module tt_um_vc32_cpu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire _14658_;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire _14727_;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire _14827_;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire _14923_;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire clknet_leaf_0_clk;
 wire \cpu.addr[10] ;
 wire \cpu.addr[11] ;
 wire \cpu.addr[12] ;
 wire \cpu.addr[13] ;
 wire \cpu.addr[14] ;
 wire \cpu.addr[15] ;
 wire \cpu.addr[1] ;
 wire \cpu.addr[2] ;
 wire \cpu.addr[3] ;
 wire \cpu.addr[4] ;
 wire \cpu.addr[5] ;
 wire \cpu.addr[6] ;
 wire \cpu.addr[7] ;
 wire \cpu.addr[8] ;
 wire \cpu.addr[9] ;
 wire \cpu.br ;
 wire \cpu.cond[0] ;
 wire \cpu.cond[1] ;
 wire \cpu.cond[2] ;
 wire \cpu.d_flush_all ;
 wire \cpu.d_rstrobe_d ;
 wire \cpu.d_wstrobe_d ;
 wire \cpu.dcache.flush_write ;
 wire \cpu.dcache.r_data[0][0] ;
 wire \cpu.dcache.r_data[0][10] ;
 wire \cpu.dcache.r_data[0][11] ;
 wire \cpu.dcache.r_data[0][12] ;
 wire \cpu.dcache.r_data[0][13] ;
 wire \cpu.dcache.r_data[0][14] ;
 wire \cpu.dcache.r_data[0][15] ;
 wire \cpu.dcache.r_data[0][16] ;
 wire \cpu.dcache.r_data[0][17] ;
 wire \cpu.dcache.r_data[0][18] ;
 wire \cpu.dcache.r_data[0][19] ;
 wire \cpu.dcache.r_data[0][1] ;
 wire \cpu.dcache.r_data[0][20] ;
 wire \cpu.dcache.r_data[0][21] ;
 wire \cpu.dcache.r_data[0][22] ;
 wire \cpu.dcache.r_data[0][23] ;
 wire \cpu.dcache.r_data[0][24] ;
 wire \cpu.dcache.r_data[0][25] ;
 wire \cpu.dcache.r_data[0][26] ;
 wire \cpu.dcache.r_data[0][27] ;
 wire \cpu.dcache.r_data[0][28] ;
 wire \cpu.dcache.r_data[0][29] ;
 wire \cpu.dcache.r_data[0][2] ;
 wire \cpu.dcache.r_data[0][30] ;
 wire \cpu.dcache.r_data[0][31] ;
 wire \cpu.dcache.r_data[0][3] ;
 wire \cpu.dcache.r_data[0][4] ;
 wire \cpu.dcache.r_data[0][5] ;
 wire \cpu.dcache.r_data[0][6] ;
 wire \cpu.dcache.r_data[0][7] ;
 wire \cpu.dcache.r_data[0][8] ;
 wire \cpu.dcache.r_data[0][9] ;
 wire \cpu.dcache.r_data[1][0] ;
 wire \cpu.dcache.r_data[1][10] ;
 wire \cpu.dcache.r_data[1][11] ;
 wire \cpu.dcache.r_data[1][12] ;
 wire \cpu.dcache.r_data[1][13] ;
 wire \cpu.dcache.r_data[1][14] ;
 wire \cpu.dcache.r_data[1][15] ;
 wire \cpu.dcache.r_data[1][16] ;
 wire \cpu.dcache.r_data[1][17] ;
 wire \cpu.dcache.r_data[1][18] ;
 wire \cpu.dcache.r_data[1][19] ;
 wire \cpu.dcache.r_data[1][1] ;
 wire \cpu.dcache.r_data[1][20] ;
 wire \cpu.dcache.r_data[1][21] ;
 wire \cpu.dcache.r_data[1][22] ;
 wire \cpu.dcache.r_data[1][23] ;
 wire \cpu.dcache.r_data[1][24] ;
 wire \cpu.dcache.r_data[1][25] ;
 wire \cpu.dcache.r_data[1][26] ;
 wire \cpu.dcache.r_data[1][27] ;
 wire \cpu.dcache.r_data[1][28] ;
 wire \cpu.dcache.r_data[1][29] ;
 wire \cpu.dcache.r_data[1][2] ;
 wire \cpu.dcache.r_data[1][30] ;
 wire \cpu.dcache.r_data[1][31] ;
 wire \cpu.dcache.r_data[1][3] ;
 wire \cpu.dcache.r_data[1][4] ;
 wire \cpu.dcache.r_data[1][5] ;
 wire \cpu.dcache.r_data[1][6] ;
 wire \cpu.dcache.r_data[1][7] ;
 wire \cpu.dcache.r_data[1][8] ;
 wire \cpu.dcache.r_data[1][9] ;
 wire \cpu.dcache.r_data[2][0] ;
 wire \cpu.dcache.r_data[2][10] ;
 wire \cpu.dcache.r_data[2][11] ;
 wire \cpu.dcache.r_data[2][12] ;
 wire \cpu.dcache.r_data[2][13] ;
 wire \cpu.dcache.r_data[2][14] ;
 wire \cpu.dcache.r_data[2][15] ;
 wire \cpu.dcache.r_data[2][16] ;
 wire \cpu.dcache.r_data[2][17] ;
 wire \cpu.dcache.r_data[2][18] ;
 wire \cpu.dcache.r_data[2][19] ;
 wire \cpu.dcache.r_data[2][1] ;
 wire \cpu.dcache.r_data[2][20] ;
 wire \cpu.dcache.r_data[2][21] ;
 wire \cpu.dcache.r_data[2][22] ;
 wire \cpu.dcache.r_data[2][23] ;
 wire \cpu.dcache.r_data[2][24] ;
 wire \cpu.dcache.r_data[2][25] ;
 wire \cpu.dcache.r_data[2][26] ;
 wire \cpu.dcache.r_data[2][27] ;
 wire \cpu.dcache.r_data[2][28] ;
 wire \cpu.dcache.r_data[2][29] ;
 wire \cpu.dcache.r_data[2][2] ;
 wire \cpu.dcache.r_data[2][30] ;
 wire \cpu.dcache.r_data[2][31] ;
 wire \cpu.dcache.r_data[2][3] ;
 wire \cpu.dcache.r_data[2][4] ;
 wire \cpu.dcache.r_data[2][5] ;
 wire \cpu.dcache.r_data[2][6] ;
 wire \cpu.dcache.r_data[2][7] ;
 wire \cpu.dcache.r_data[2][8] ;
 wire \cpu.dcache.r_data[2][9] ;
 wire \cpu.dcache.r_data[3][0] ;
 wire \cpu.dcache.r_data[3][10] ;
 wire \cpu.dcache.r_data[3][11] ;
 wire \cpu.dcache.r_data[3][12] ;
 wire \cpu.dcache.r_data[3][13] ;
 wire \cpu.dcache.r_data[3][14] ;
 wire \cpu.dcache.r_data[3][15] ;
 wire \cpu.dcache.r_data[3][16] ;
 wire \cpu.dcache.r_data[3][17] ;
 wire \cpu.dcache.r_data[3][18] ;
 wire \cpu.dcache.r_data[3][19] ;
 wire \cpu.dcache.r_data[3][1] ;
 wire \cpu.dcache.r_data[3][20] ;
 wire \cpu.dcache.r_data[3][21] ;
 wire \cpu.dcache.r_data[3][22] ;
 wire \cpu.dcache.r_data[3][23] ;
 wire \cpu.dcache.r_data[3][24] ;
 wire \cpu.dcache.r_data[3][25] ;
 wire \cpu.dcache.r_data[3][26] ;
 wire \cpu.dcache.r_data[3][27] ;
 wire \cpu.dcache.r_data[3][28] ;
 wire \cpu.dcache.r_data[3][29] ;
 wire \cpu.dcache.r_data[3][2] ;
 wire \cpu.dcache.r_data[3][30] ;
 wire \cpu.dcache.r_data[3][31] ;
 wire \cpu.dcache.r_data[3][3] ;
 wire \cpu.dcache.r_data[3][4] ;
 wire \cpu.dcache.r_data[3][5] ;
 wire \cpu.dcache.r_data[3][6] ;
 wire \cpu.dcache.r_data[3][7] ;
 wire \cpu.dcache.r_data[3][8] ;
 wire \cpu.dcache.r_data[3][9] ;
 wire \cpu.dcache.r_data[4][0] ;
 wire \cpu.dcache.r_data[4][10] ;
 wire \cpu.dcache.r_data[4][11] ;
 wire \cpu.dcache.r_data[4][12] ;
 wire \cpu.dcache.r_data[4][13] ;
 wire \cpu.dcache.r_data[4][14] ;
 wire \cpu.dcache.r_data[4][15] ;
 wire \cpu.dcache.r_data[4][16] ;
 wire \cpu.dcache.r_data[4][17] ;
 wire \cpu.dcache.r_data[4][18] ;
 wire \cpu.dcache.r_data[4][19] ;
 wire \cpu.dcache.r_data[4][1] ;
 wire \cpu.dcache.r_data[4][20] ;
 wire \cpu.dcache.r_data[4][21] ;
 wire \cpu.dcache.r_data[4][22] ;
 wire \cpu.dcache.r_data[4][23] ;
 wire \cpu.dcache.r_data[4][24] ;
 wire \cpu.dcache.r_data[4][25] ;
 wire \cpu.dcache.r_data[4][26] ;
 wire \cpu.dcache.r_data[4][27] ;
 wire \cpu.dcache.r_data[4][28] ;
 wire \cpu.dcache.r_data[4][29] ;
 wire \cpu.dcache.r_data[4][2] ;
 wire \cpu.dcache.r_data[4][30] ;
 wire \cpu.dcache.r_data[4][31] ;
 wire \cpu.dcache.r_data[4][3] ;
 wire \cpu.dcache.r_data[4][4] ;
 wire \cpu.dcache.r_data[4][5] ;
 wire \cpu.dcache.r_data[4][6] ;
 wire \cpu.dcache.r_data[4][7] ;
 wire \cpu.dcache.r_data[4][8] ;
 wire \cpu.dcache.r_data[4][9] ;
 wire \cpu.dcache.r_data[5][0] ;
 wire \cpu.dcache.r_data[5][10] ;
 wire \cpu.dcache.r_data[5][11] ;
 wire \cpu.dcache.r_data[5][12] ;
 wire \cpu.dcache.r_data[5][13] ;
 wire \cpu.dcache.r_data[5][14] ;
 wire \cpu.dcache.r_data[5][15] ;
 wire \cpu.dcache.r_data[5][16] ;
 wire \cpu.dcache.r_data[5][17] ;
 wire \cpu.dcache.r_data[5][18] ;
 wire \cpu.dcache.r_data[5][19] ;
 wire \cpu.dcache.r_data[5][1] ;
 wire \cpu.dcache.r_data[5][20] ;
 wire \cpu.dcache.r_data[5][21] ;
 wire \cpu.dcache.r_data[5][22] ;
 wire \cpu.dcache.r_data[5][23] ;
 wire \cpu.dcache.r_data[5][24] ;
 wire \cpu.dcache.r_data[5][25] ;
 wire \cpu.dcache.r_data[5][26] ;
 wire \cpu.dcache.r_data[5][27] ;
 wire \cpu.dcache.r_data[5][28] ;
 wire \cpu.dcache.r_data[5][29] ;
 wire \cpu.dcache.r_data[5][2] ;
 wire \cpu.dcache.r_data[5][30] ;
 wire \cpu.dcache.r_data[5][31] ;
 wire \cpu.dcache.r_data[5][3] ;
 wire \cpu.dcache.r_data[5][4] ;
 wire \cpu.dcache.r_data[5][5] ;
 wire \cpu.dcache.r_data[5][6] ;
 wire \cpu.dcache.r_data[5][7] ;
 wire \cpu.dcache.r_data[5][8] ;
 wire \cpu.dcache.r_data[5][9] ;
 wire \cpu.dcache.r_data[6][0] ;
 wire \cpu.dcache.r_data[6][10] ;
 wire \cpu.dcache.r_data[6][11] ;
 wire \cpu.dcache.r_data[6][12] ;
 wire \cpu.dcache.r_data[6][13] ;
 wire \cpu.dcache.r_data[6][14] ;
 wire \cpu.dcache.r_data[6][15] ;
 wire \cpu.dcache.r_data[6][16] ;
 wire \cpu.dcache.r_data[6][17] ;
 wire \cpu.dcache.r_data[6][18] ;
 wire \cpu.dcache.r_data[6][19] ;
 wire \cpu.dcache.r_data[6][1] ;
 wire \cpu.dcache.r_data[6][20] ;
 wire \cpu.dcache.r_data[6][21] ;
 wire \cpu.dcache.r_data[6][22] ;
 wire \cpu.dcache.r_data[6][23] ;
 wire \cpu.dcache.r_data[6][24] ;
 wire \cpu.dcache.r_data[6][25] ;
 wire \cpu.dcache.r_data[6][26] ;
 wire \cpu.dcache.r_data[6][27] ;
 wire \cpu.dcache.r_data[6][28] ;
 wire \cpu.dcache.r_data[6][29] ;
 wire \cpu.dcache.r_data[6][2] ;
 wire \cpu.dcache.r_data[6][30] ;
 wire \cpu.dcache.r_data[6][31] ;
 wire \cpu.dcache.r_data[6][3] ;
 wire \cpu.dcache.r_data[6][4] ;
 wire \cpu.dcache.r_data[6][5] ;
 wire \cpu.dcache.r_data[6][6] ;
 wire \cpu.dcache.r_data[6][7] ;
 wire \cpu.dcache.r_data[6][8] ;
 wire \cpu.dcache.r_data[6][9] ;
 wire \cpu.dcache.r_data[7][0] ;
 wire \cpu.dcache.r_data[7][10] ;
 wire \cpu.dcache.r_data[7][11] ;
 wire \cpu.dcache.r_data[7][12] ;
 wire \cpu.dcache.r_data[7][13] ;
 wire \cpu.dcache.r_data[7][14] ;
 wire \cpu.dcache.r_data[7][15] ;
 wire \cpu.dcache.r_data[7][16] ;
 wire \cpu.dcache.r_data[7][17] ;
 wire \cpu.dcache.r_data[7][18] ;
 wire \cpu.dcache.r_data[7][19] ;
 wire \cpu.dcache.r_data[7][1] ;
 wire \cpu.dcache.r_data[7][20] ;
 wire \cpu.dcache.r_data[7][21] ;
 wire \cpu.dcache.r_data[7][22] ;
 wire \cpu.dcache.r_data[7][23] ;
 wire \cpu.dcache.r_data[7][24] ;
 wire \cpu.dcache.r_data[7][25] ;
 wire \cpu.dcache.r_data[7][26] ;
 wire \cpu.dcache.r_data[7][27] ;
 wire \cpu.dcache.r_data[7][28] ;
 wire \cpu.dcache.r_data[7][29] ;
 wire \cpu.dcache.r_data[7][2] ;
 wire \cpu.dcache.r_data[7][30] ;
 wire \cpu.dcache.r_data[7][31] ;
 wire \cpu.dcache.r_data[7][3] ;
 wire \cpu.dcache.r_data[7][4] ;
 wire \cpu.dcache.r_data[7][5] ;
 wire \cpu.dcache.r_data[7][6] ;
 wire \cpu.dcache.r_data[7][7] ;
 wire \cpu.dcache.r_data[7][8] ;
 wire \cpu.dcache.r_data[7][9] ;
 wire \cpu.dcache.r_dirty[0] ;
 wire \cpu.dcache.r_dirty[1] ;
 wire \cpu.dcache.r_dirty[2] ;
 wire \cpu.dcache.r_dirty[3] ;
 wire \cpu.dcache.r_dirty[4] ;
 wire \cpu.dcache.r_dirty[5] ;
 wire \cpu.dcache.r_dirty[6] ;
 wire \cpu.dcache.r_dirty[7] ;
 wire \cpu.dcache.r_offset[0] ;
 wire \cpu.dcache.r_offset[1] ;
 wire \cpu.dcache.r_offset[2] ;
 wire \cpu.dcache.r_tag[0][10] ;
 wire \cpu.dcache.r_tag[0][11] ;
 wire \cpu.dcache.r_tag[0][12] ;
 wire \cpu.dcache.r_tag[0][13] ;
 wire \cpu.dcache.r_tag[0][14] ;
 wire \cpu.dcache.r_tag[0][15] ;
 wire \cpu.dcache.r_tag[0][16] ;
 wire \cpu.dcache.r_tag[0][17] ;
 wire \cpu.dcache.r_tag[0][18] ;
 wire \cpu.dcache.r_tag[0][19] ;
 wire \cpu.dcache.r_tag[0][20] ;
 wire \cpu.dcache.r_tag[0][21] ;
 wire \cpu.dcache.r_tag[0][22] ;
 wire \cpu.dcache.r_tag[0][23] ;
 wire \cpu.dcache.r_tag[0][5] ;
 wire \cpu.dcache.r_tag[0][6] ;
 wire \cpu.dcache.r_tag[0][7] ;
 wire \cpu.dcache.r_tag[0][8] ;
 wire \cpu.dcache.r_tag[0][9] ;
 wire \cpu.dcache.r_tag[1][10] ;
 wire \cpu.dcache.r_tag[1][11] ;
 wire \cpu.dcache.r_tag[1][12] ;
 wire \cpu.dcache.r_tag[1][13] ;
 wire \cpu.dcache.r_tag[1][14] ;
 wire \cpu.dcache.r_tag[1][15] ;
 wire \cpu.dcache.r_tag[1][16] ;
 wire \cpu.dcache.r_tag[1][17] ;
 wire \cpu.dcache.r_tag[1][18] ;
 wire \cpu.dcache.r_tag[1][19] ;
 wire \cpu.dcache.r_tag[1][20] ;
 wire \cpu.dcache.r_tag[1][21] ;
 wire \cpu.dcache.r_tag[1][22] ;
 wire \cpu.dcache.r_tag[1][23] ;
 wire \cpu.dcache.r_tag[1][5] ;
 wire \cpu.dcache.r_tag[1][6] ;
 wire \cpu.dcache.r_tag[1][7] ;
 wire \cpu.dcache.r_tag[1][8] ;
 wire \cpu.dcache.r_tag[1][9] ;
 wire \cpu.dcache.r_tag[2][10] ;
 wire \cpu.dcache.r_tag[2][11] ;
 wire \cpu.dcache.r_tag[2][12] ;
 wire \cpu.dcache.r_tag[2][13] ;
 wire \cpu.dcache.r_tag[2][14] ;
 wire \cpu.dcache.r_tag[2][15] ;
 wire \cpu.dcache.r_tag[2][16] ;
 wire \cpu.dcache.r_tag[2][17] ;
 wire \cpu.dcache.r_tag[2][18] ;
 wire \cpu.dcache.r_tag[2][19] ;
 wire \cpu.dcache.r_tag[2][20] ;
 wire \cpu.dcache.r_tag[2][21] ;
 wire \cpu.dcache.r_tag[2][22] ;
 wire \cpu.dcache.r_tag[2][23] ;
 wire \cpu.dcache.r_tag[2][5] ;
 wire \cpu.dcache.r_tag[2][6] ;
 wire \cpu.dcache.r_tag[2][7] ;
 wire \cpu.dcache.r_tag[2][8] ;
 wire \cpu.dcache.r_tag[2][9] ;
 wire \cpu.dcache.r_tag[3][10] ;
 wire \cpu.dcache.r_tag[3][11] ;
 wire \cpu.dcache.r_tag[3][12] ;
 wire \cpu.dcache.r_tag[3][13] ;
 wire \cpu.dcache.r_tag[3][14] ;
 wire \cpu.dcache.r_tag[3][15] ;
 wire \cpu.dcache.r_tag[3][16] ;
 wire \cpu.dcache.r_tag[3][17] ;
 wire \cpu.dcache.r_tag[3][18] ;
 wire \cpu.dcache.r_tag[3][19] ;
 wire \cpu.dcache.r_tag[3][20] ;
 wire \cpu.dcache.r_tag[3][21] ;
 wire \cpu.dcache.r_tag[3][22] ;
 wire \cpu.dcache.r_tag[3][23] ;
 wire \cpu.dcache.r_tag[3][5] ;
 wire \cpu.dcache.r_tag[3][6] ;
 wire \cpu.dcache.r_tag[3][7] ;
 wire \cpu.dcache.r_tag[3][8] ;
 wire \cpu.dcache.r_tag[3][9] ;
 wire \cpu.dcache.r_tag[4][10] ;
 wire \cpu.dcache.r_tag[4][11] ;
 wire \cpu.dcache.r_tag[4][12] ;
 wire \cpu.dcache.r_tag[4][13] ;
 wire \cpu.dcache.r_tag[4][14] ;
 wire \cpu.dcache.r_tag[4][15] ;
 wire \cpu.dcache.r_tag[4][16] ;
 wire \cpu.dcache.r_tag[4][17] ;
 wire \cpu.dcache.r_tag[4][18] ;
 wire \cpu.dcache.r_tag[4][19] ;
 wire \cpu.dcache.r_tag[4][20] ;
 wire \cpu.dcache.r_tag[4][21] ;
 wire \cpu.dcache.r_tag[4][22] ;
 wire \cpu.dcache.r_tag[4][23] ;
 wire \cpu.dcache.r_tag[4][5] ;
 wire \cpu.dcache.r_tag[4][6] ;
 wire \cpu.dcache.r_tag[4][7] ;
 wire \cpu.dcache.r_tag[4][8] ;
 wire \cpu.dcache.r_tag[4][9] ;
 wire \cpu.dcache.r_tag[5][10] ;
 wire \cpu.dcache.r_tag[5][11] ;
 wire \cpu.dcache.r_tag[5][12] ;
 wire \cpu.dcache.r_tag[5][13] ;
 wire \cpu.dcache.r_tag[5][14] ;
 wire \cpu.dcache.r_tag[5][15] ;
 wire \cpu.dcache.r_tag[5][16] ;
 wire \cpu.dcache.r_tag[5][17] ;
 wire \cpu.dcache.r_tag[5][18] ;
 wire \cpu.dcache.r_tag[5][19] ;
 wire \cpu.dcache.r_tag[5][20] ;
 wire \cpu.dcache.r_tag[5][21] ;
 wire \cpu.dcache.r_tag[5][22] ;
 wire \cpu.dcache.r_tag[5][23] ;
 wire \cpu.dcache.r_tag[5][5] ;
 wire \cpu.dcache.r_tag[5][6] ;
 wire \cpu.dcache.r_tag[5][7] ;
 wire \cpu.dcache.r_tag[5][8] ;
 wire \cpu.dcache.r_tag[5][9] ;
 wire \cpu.dcache.r_tag[6][10] ;
 wire \cpu.dcache.r_tag[6][11] ;
 wire \cpu.dcache.r_tag[6][12] ;
 wire \cpu.dcache.r_tag[6][13] ;
 wire \cpu.dcache.r_tag[6][14] ;
 wire \cpu.dcache.r_tag[6][15] ;
 wire \cpu.dcache.r_tag[6][16] ;
 wire \cpu.dcache.r_tag[6][17] ;
 wire \cpu.dcache.r_tag[6][18] ;
 wire \cpu.dcache.r_tag[6][19] ;
 wire \cpu.dcache.r_tag[6][20] ;
 wire \cpu.dcache.r_tag[6][21] ;
 wire \cpu.dcache.r_tag[6][22] ;
 wire \cpu.dcache.r_tag[6][23] ;
 wire \cpu.dcache.r_tag[6][5] ;
 wire \cpu.dcache.r_tag[6][6] ;
 wire \cpu.dcache.r_tag[6][7] ;
 wire \cpu.dcache.r_tag[6][8] ;
 wire \cpu.dcache.r_tag[6][9] ;
 wire \cpu.dcache.r_tag[7][10] ;
 wire \cpu.dcache.r_tag[7][11] ;
 wire \cpu.dcache.r_tag[7][12] ;
 wire \cpu.dcache.r_tag[7][13] ;
 wire \cpu.dcache.r_tag[7][14] ;
 wire \cpu.dcache.r_tag[7][15] ;
 wire \cpu.dcache.r_tag[7][16] ;
 wire \cpu.dcache.r_tag[7][17] ;
 wire \cpu.dcache.r_tag[7][18] ;
 wire \cpu.dcache.r_tag[7][19] ;
 wire \cpu.dcache.r_tag[7][20] ;
 wire \cpu.dcache.r_tag[7][21] ;
 wire \cpu.dcache.r_tag[7][22] ;
 wire \cpu.dcache.r_tag[7][23] ;
 wire \cpu.dcache.r_tag[7][5] ;
 wire \cpu.dcache.r_tag[7][6] ;
 wire \cpu.dcache.r_tag[7][7] ;
 wire \cpu.dcache.r_tag[7][8] ;
 wire \cpu.dcache.r_tag[7][9] ;
 wire \cpu.dcache.r_valid[0] ;
 wire \cpu.dcache.r_valid[1] ;
 wire \cpu.dcache.r_valid[2] ;
 wire \cpu.dcache.r_valid[3] ;
 wire \cpu.dcache.r_valid[4] ;
 wire \cpu.dcache.r_valid[5] ;
 wire \cpu.dcache.r_valid[6] ;
 wire \cpu.dcache.r_valid[7] ;
 wire \cpu.dcache.wdata[0] ;
 wire \cpu.dcache.wdata[10] ;
 wire \cpu.dcache.wdata[11] ;
 wire \cpu.dcache.wdata[12] ;
 wire \cpu.dcache.wdata[13] ;
 wire \cpu.dcache.wdata[14] ;
 wire \cpu.dcache.wdata[15] ;
 wire \cpu.dcache.wdata[1] ;
 wire \cpu.dcache.wdata[2] ;
 wire \cpu.dcache.wdata[3] ;
 wire \cpu.dcache.wdata[4] ;
 wire \cpu.dcache.wdata[5] ;
 wire \cpu.dcache.wdata[6] ;
 wire \cpu.dcache.wdata[7] ;
 wire \cpu.dcache.wdata[8] ;
 wire \cpu.dcache.wdata[9] ;
 wire \cpu.dec.div ;
 wire \cpu.dec.do_flush_all ;
 wire \cpu.dec.do_flush_write ;
 wire \cpu.dec.do_inv_mmu ;
 wire \cpu.dec.imm[0] ;
 wire \cpu.dec.imm[10] ;
 wire \cpu.dec.imm[11] ;
 wire \cpu.dec.imm[12] ;
 wire \cpu.dec.imm[13] ;
 wire \cpu.dec.imm[14] ;
 wire \cpu.dec.imm[15] ;
 wire \cpu.dec.imm[1] ;
 wire \cpu.dec.imm[2] ;
 wire \cpu.dec.imm[3] ;
 wire \cpu.dec.imm[4] ;
 wire \cpu.dec.imm[5] ;
 wire \cpu.dec.imm[6] ;
 wire \cpu.dec.imm[7] ;
 wire \cpu.dec.imm[8] ;
 wire \cpu.dec.imm[9] ;
 wire \cpu.dec.io ;
 wire \cpu.dec.iready ;
 wire \cpu.dec.jmp ;
 wire \cpu.dec.load ;
 wire \cpu.dec.mult ;
 wire \cpu.dec.needs_rs2 ;
 wire \cpu.dec.r_op[10] ;
 wire \cpu.dec.r_op[1] ;
 wire \cpu.dec.r_op[2] ;
 wire \cpu.dec.r_op[3] ;
 wire \cpu.dec.r_op[4] ;
 wire \cpu.dec.r_op[5] ;
 wire \cpu.dec.r_op[6] ;
 wire \cpu.dec.r_op[7] ;
 wire \cpu.dec.r_op[8] ;
 wire \cpu.dec.r_op[9] ;
 wire \cpu.dec.r_rd[0] ;
 wire \cpu.dec.r_rd[1] ;
 wire \cpu.dec.r_rd[2] ;
 wire \cpu.dec.r_rd[3] ;
 wire \cpu.dec.r_rs1[0] ;
 wire \cpu.dec.r_rs1[1] ;
 wire \cpu.dec.r_rs1[2] ;
 wire \cpu.dec.r_rs1[3] ;
 wire \cpu.dec.r_rs2[0] ;
 wire \cpu.dec.r_rs2[1] ;
 wire \cpu.dec.r_rs2[2] ;
 wire \cpu.dec.r_rs2[3] ;
 wire \cpu.dec.r_rs2_pc ;
 wire \cpu.dec.r_set_cc ;
 wire \cpu.dec.r_store ;
 wire \cpu.dec.r_swapsp ;
 wire \cpu.dec.r_sys_call ;
 wire \cpu.dec.r_trap ;
 wire \cpu.dec.supmode ;
 wire \cpu.dec.user_io ;
 wire \cpu.ex.c_div_running ;
 wire \cpu.ex.c_mult[0] ;
 wire \cpu.ex.c_mult[10] ;
 wire \cpu.ex.c_mult[11] ;
 wire \cpu.ex.c_mult[12] ;
 wire \cpu.ex.c_mult[13] ;
 wire \cpu.ex.c_mult[14] ;
 wire \cpu.ex.c_mult[15] ;
 wire \cpu.ex.c_mult[1] ;
 wire \cpu.ex.c_mult[2] ;
 wire \cpu.ex.c_mult[3] ;
 wire \cpu.ex.c_mult[4] ;
 wire \cpu.ex.c_mult[5] ;
 wire \cpu.ex.c_mult[6] ;
 wire \cpu.ex.c_mult[7] ;
 wire \cpu.ex.c_mult[8] ;
 wire \cpu.ex.c_mult[9] ;
 wire \cpu.ex.c_mult_off[0] ;
 wire \cpu.ex.c_mult_off[1] ;
 wire \cpu.ex.c_mult_off[2] ;
 wire \cpu.ex.c_mult_off[3] ;
 wire \cpu.ex.c_mult_running ;
 wire \cpu.ex.genblk3.c_supmode ;
 wire \cpu.ex.genblk3.r_mmu_d_proxy ;
 wire \cpu.ex.genblk3.r_mmu_enable ;
 wire \cpu.ex.genblk3.r_prev_supmode ;
 wire \cpu.ex.i_flush_all ;
 wire \cpu.ex.ifetch ;
 wire \cpu.ex.io_access ;
 wire \cpu.ex.mmu_read[12] ;
 wire \cpu.ex.mmu_read[13] ;
 wire \cpu.ex.mmu_read[14] ;
 wire \cpu.ex.mmu_read[15] ;
 wire \cpu.ex.mmu_read[1] ;
 wire \cpu.ex.mmu_read[2] ;
 wire \cpu.ex.mmu_read[3] ;
 wire \cpu.ex.mmu_reg_data[0] ;
 wire \cpu.ex.pc[10] ;
 wire \cpu.ex.pc[11] ;
 wire \cpu.ex.pc[12] ;
 wire \cpu.ex.pc[13] ;
 wire \cpu.ex.pc[14] ;
 wire \cpu.ex.pc[15] ;
 wire \cpu.ex.pc[1] ;
 wire \cpu.ex.pc[2] ;
 wire \cpu.ex.pc[3] ;
 wire \cpu.ex.pc[4] ;
 wire \cpu.ex.pc[5] ;
 wire \cpu.ex.pc[6] ;
 wire \cpu.ex.pc[7] ;
 wire \cpu.ex.pc[8] ;
 wire \cpu.ex.pc[9] ;
 wire \cpu.ex.r_10[0] ;
 wire \cpu.ex.r_10[10] ;
 wire \cpu.ex.r_10[11] ;
 wire \cpu.ex.r_10[12] ;
 wire \cpu.ex.r_10[13] ;
 wire \cpu.ex.r_10[14] ;
 wire \cpu.ex.r_10[15] ;
 wire \cpu.ex.r_10[1] ;
 wire \cpu.ex.r_10[2] ;
 wire \cpu.ex.r_10[3] ;
 wire \cpu.ex.r_10[4] ;
 wire \cpu.ex.r_10[5] ;
 wire \cpu.ex.r_10[6] ;
 wire \cpu.ex.r_10[7] ;
 wire \cpu.ex.r_10[8] ;
 wire \cpu.ex.r_10[9] ;
 wire \cpu.ex.r_11[0] ;
 wire \cpu.ex.r_11[10] ;
 wire \cpu.ex.r_11[11] ;
 wire \cpu.ex.r_11[12] ;
 wire \cpu.ex.r_11[13] ;
 wire \cpu.ex.r_11[14] ;
 wire \cpu.ex.r_11[15] ;
 wire \cpu.ex.r_11[1] ;
 wire \cpu.ex.r_11[2] ;
 wire \cpu.ex.r_11[3] ;
 wire \cpu.ex.r_11[4] ;
 wire \cpu.ex.r_11[5] ;
 wire \cpu.ex.r_11[6] ;
 wire \cpu.ex.r_11[7] ;
 wire \cpu.ex.r_11[8] ;
 wire \cpu.ex.r_11[9] ;
 wire \cpu.ex.r_12[0] ;
 wire \cpu.ex.r_12[10] ;
 wire \cpu.ex.r_12[11] ;
 wire \cpu.ex.r_12[12] ;
 wire \cpu.ex.r_12[13] ;
 wire \cpu.ex.r_12[14] ;
 wire \cpu.ex.r_12[15] ;
 wire \cpu.ex.r_12[1] ;
 wire \cpu.ex.r_12[2] ;
 wire \cpu.ex.r_12[3] ;
 wire \cpu.ex.r_12[4] ;
 wire \cpu.ex.r_12[5] ;
 wire \cpu.ex.r_12[6] ;
 wire \cpu.ex.r_12[7] ;
 wire \cpu.ex.r_12[8] ;
 wire \cpu.ex.r_12[9] ;
 wire \cpu.ex.r_13[0] ;
 wire \cpu.ex.r_13[10] ;
 wire \cpu.ex.r_13[11] ;
 wire \cpu.ex.r_13[12] ;
 wire \cpu.ex.r_13[13] ;
 wire \cpu.ex.r_13[14] ;
 wire \cpu.ex.r_13[15] ;
 wire \cpu.ex.r_13[1] ;
 wire \cpu.ex.r_13[2] ;
 wire \cpu.ex.r_13[3] ;
 wire \cpu.ex.r_13[4] ;
 wire \cpu.ex.r_13[5] ;
 wire \cpu.ex.r_13[6] ;
 wire \cpu.ex.r_13[7] ;
 wire \cpu.ex.r_13[8] ;
 wire \cpu.ex.r_13[9] ;
 wire \cpu.ex.r_14[0] ;
 wire \cpu.ex.r_14[10] ;
 wire \cpu.ex.r_14[11] ;
 wire \cpu.ex.r_14[12] ;
 wire \cpu.ex.r_14[13] ;
 wire \cpu.ex.r_14[14] ;
 wire \cpu.ex.r_14[15] ;
 wire \cpu.ex.r_14[1] ;
 wire \cpu.ex.r_14[2] ;
 wire \cpu.ex.r_14[3] ;
 wire \cpu.ex.r_14[4] ;
 wire \cpu.ex.r_14[5] ;
 wire \cpu.ex.r_14[6] ;
 wire \cpu.ex.r_14[7] ;
 wire \cpu.ex.r_14[8] ;
 wire \cpu.ex.r_14[9] ;
 wire \cpu.ex.r_15[0] ;
 wire \cpu.ex.r_15[10] ;
 wire \cpu.ex.r_15[11] ;
 wire \cpu.ex.r_15[12] ;
 wire \cpu.ex.r_15[13] ;
 wire \cpu.ex.r_15[14] ;
 wire \cpu.ex.r_15[15] ;
 wire \cpu.ex.r_15[1] ;
 wire \cpu.ex.r_15[2] ;
 wire \cpu.ex.r_15[3] ;
 wire \cpu.ex.r_15[4] ;
 wire \cpu.ex.r_15[5] ;
 wire \cpu.ex.r_15[6] ;
 wire \cpu.ex.r_15[7] ;
 wire \cpu.ex.r_15[8] ;
 wire \cpu.ex.r_15[9] ;
 wire \cpu.ex.r_8[0] ;
 wire \cpu.ex.r_8[10] ;
 wire \cpu.ex.r_8[11] ;
 wire \cpu.ex.r_8[12] ;
 wire \cpu.ex.r_8[13] ;
 wire \cpu.ex.r_8[14] ;
 wire \cpu.ex.r_8[15] ;
 wire \cpu.ex.r_8[1] ;
 wire \cpu.ex.r_8[2] ;
 wire \cpu.ex.r_8[3] ;
 wire \cpu.ex.r_8[4] ;
 wire \cpu.ex.r_8[5] ;
 wire \cpu.ex.r_8[6] ;
 wire \cpu.ex.r_8[7] ;
 wire \cpu.ex.r_8[8] ;
 wire \cpu.ex.r_8[9] ;
 wire \cpu.ex.r_9[0] ;
 wire \cpu.ex.r_9[10] ;
 wire \cpu.ex.r_9[11] ;
 wire \cpu.ex.r_9[12] ;
 wire \cpu.ex.r_9[13] ;
 wire \cpu.ex.r_9[14] ;
 wire \cpu.ex.r_9[15] ;
 wire \cpu.ex.r_9[1] ;
 wire \cpu.ex.r_9[2] ;
 wire \cpu.ex.r_9[3] ;
 wire \cpu.ex.r_9[4] ;
 wire \cpu.ex.r_9[5] ;
 wire \cpu.ex.r_9[6] ;
 wire \cpu.ex.r_9[7] ;
 wire \cpu.ex.r_9[8] ;
 wire \cpu.ex.r_9[9] ;
 wire \cpu.ex.r_branch_stall ;
 wire \cpu.ex.r_div_running ;
 wire \cpu.ex.r_epc[10] ;
 wire \cpu.ex.r_epc[11] ;
 wire \cpu.ex.r_epc[12] ;
 wire \cpu.ex.r_epc[13] ;
 wire \cpu.ex.r_epc[14] ;
 wire \cpu.ex.r_epc[15] ;
 wire \cpu.ex.r_epc[1] ;
 wire \cpu.ex.r_epc[2] ;
 wire \cpu.ex.r_epc[3] ;
 wire \cpu.ex.r_epc[4] ;
 wire \cpu.ex.r_epc[5] ;
 wire \cpu.ex.r_epc[6] ;
 wire \cpu.ex.r_epc[7] ;
 wire \cpu.ex.r_epc[8] ;
 wire \cpu.ex.r_epc[9] ;
 wire \cpu.ex.r_ie ;
 wire \cpu.ex.r_lr[10] ;
 wire \cpu.ex.r_lr[11] ;
 wire \cpu.ex.r_lr[12] ;
 wire \cpu.ex.r_lr[13] ;
 wire \cpu.ex.r_lr[14] ;
 wire \cpu.ex.r_lr[15] ;
 wire \cpu.ex.r_lr[1] ;
 wire \cpu.ex.r_lr[2] ;
 wire \cpu.ex.r_lr[3] ;
 wire \cpu.ex.r_lr[4] ;
 wire \cpu.ex.r_lr[5] ;
 wire \cpu.ex.r_lr[6] ;
 wire \cpu.ex.r_lr[7] ;
 wire \cpu.ex.r_lr[8] ;
 wire \cpu.ex.r_lr[9] ;
 wire \cpu.ex.r_mult[0] ;
 wire \cpu.ex.r_mult[10] ;
 wire \cpu.ex.r_mult[11] ;
 wire \cpu.ex.r_mult[12] ;
 wire \cpu.ex.r_mult[13] ;
 wire \cpu.ex.r_mult[14] ;
 wire \cpu.ex.r_mult[15] ;
 wire \cpu.ex.r_mult[16] ;
 wire \cpu.ex.r_mult[17] ;
 wire \cpu.ex.r_mult[18] ;
 wire \cpu.ex.r_mult[19] ;
 wire \cpu.ex.r_mult[1] ;
 wire \cpu.ex.r_mult[20] ;
 wire \cpu.ex.r_mult[21] ;
 wire \cpu.ex.r_mult[22] ;
 wire \cpu.ex.r_mult[23] ;
 wire \cpu.ex.r_mult[24] ;
 wire \cpu.ex.r_mult[25] ;
 wire \cpu.ex.r_mult[26] ;
 wire \cpu.ex.r_mult[27] ;
 wire \cpu.ex.r_mult[28] ;
 wire \cpu.ex.r_mult[29] ;
 wire \cpu.ex.r_mult[2] ;
 wire \cpu.ex.r_mult[30] ;
 wire \cpu.ex.r_mult[31] ;
 wire \cpu.ex.r_mult[3] ;
 wire \cpu.ex.r_mult[4] ;
 wire \cpu.ex.r_mult[5] ;
 wire \cpu.ex.r_mult[6] ;
 wire \cpu.ex.r_mult[7] ;
 wire \cpu.ex.r_mult[8] ;
 wire \cpu.ex.r_mult[9] ;
 wire \cpu.ex.r_mult_off[0] ;
 wire \cpu.ex.r_mult_off[1] ;
 wire \cpu.ex.r_mult_off[2] ;
 wire \cpu.ex.r_mult_off[3] ;
 wire \cpu.ex.r_mult_running ;
 wire \cpu.ex.r_prev_ie ;
 wire \cpu.ex.r_read_stall ;
 wire \cpu.ex.r_sp[10] ;
 wire \cpu.ex.r_sp[11] ;
 wire \cpu.ex.r_sp[12] ;
 wire \cpu.ex.r_sp[13] ;
 wire \cpu.ex.r_sp[14] ;
 wire \cpu.ex.r_sp[15] ;
 wire \cpu.ex.r_sp[1] ;
 wire \cpu.ex.r_sp[2] ;
 wire \cpu.ex.r_sp[3] ;
 wire \cpu.ex.r_sp[4] ;
 wire \cpu.ex.r_sp[5] ;
 wire \cpu.ex.r_sp[6] ;
 wire \cpu.ex.r_sp[7] ;
 wire \cpu.ex.r_sp[8] ;
 wire \cpu.ex.r_sp[9] ;
 wire \cpu.ex.r_stmp[0] ;
 wire \cpu.ex.r_stmp[10] ;
 wire \cpu.ex.r_stmp[11] ;
 wire \cpu.ex.r_stmp[12] ;
 wire \cpu.ex.r_stmp[13] ;
 wire \cpu.ex.r_stmp[14] ;
 wire \cpu.ex.r_stmp[15] ;
 wire \cpu.ex.r_stmp[1] ;
 wire \cpu.ex.r_stmp[2] ;
 wire \cpu.ex.r_stmp[3] ;
 wire \cpu.ex.r_stmp[4] ;
 wire \cpu.ex.r_stmp[5] ;
 wire \cpu.ex.r_stmp[6] ;
 wire \cpu.ex.r_stmp[7] ;
 wire \cpu.ex.r_stmp[8] ;
 wire \cpu.ex.r_stmp[9] ;
 wire \cpu.ex.r_wb_addr[0] ;
 wire \cpu.ex.r_wb_addr[1] ;
 wire \cpu.ex.r_wb_addr[2] ;
 wire \cpu.ex.r_wb_addr[3] ;
 wire \cpu.ex.r_wb_swapsp ;
 wire \cpu.ex.r_wb_valid ;
 wire \cpu.ex.r_wmask[0] ;
 wire \cpu.ex.r_wmask[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[0] ;
 wire \cpu.genblk1.mmu.r_valid_d[10] ;
 wire \cpu.genblk1.mmu.r_valid_d[11] ;
 wire \cpu.genblk1.mmu.r_valid_d[12] ;
 wire \cpu.genblk1.mmu.r_valid_d[13] ;
 wire \cpu.genblk1.mmu.r_valid_d[14] ;
 wire \cpu.genblk1.mmu.r_valid_d[15] ;
 wire \cpu.genblk1.mmu.r_valid_d[16] ;
 wire \cpu.genblk1.mmu.r_valid_d[17] ;
 wire \cpu.genblk1.mmu.r_valid_d[18] ;
 wire \cpu.genblk1.mmu.r_valid_d[19] ;
 wire \cpu.genblk1.mmu.r_valid_d[1] ;
 wire \cpu.genblk1.mmu.r_valid_d[20] ;
 wire \cpu.genblk1.mmu.r_valid_d[21] ;
 wire \cpu.genblk1.mmu.r_valid_d[22] ;
 wire \cpu.genblk1.mmu.r_valid_d[23] ;
 wire \cpu.genblk1.mmu.r_valid_d[24] ;
 wire \cpu.genblk1.mmu.r_valid_d[25] ;
 wire \cpu.genblk1.mmu.r_valid_d[26] ;
 wire \cpu.genblk1.mmu.r_valid_d[27] ;
 wire \cpu.genblk1.mmu.r_valid_d[28] ;
 wire \cpu.genblk1.mmu.r_valid_d[29] ;
 wire \cpu.genblk1.mmu.r_valid_d[2] ;
 wire \cpu.genblk1.mmu.r_valid_d[30] ;
 wire \cpu.genblk1.mmu.r_valid_d[31] ;
 wire \cpu.genblk1.mmu.r_valid_d[3] ;
 wire \cpu.genblk1.mmu.r_valid_d[4] ;
 wire \cpu.genblk1.mmu.r_valid_d[5] ;
 wire \cpu.genblk1.mmu.r_valid_d[6] ;
 wire \cpu.genblk1.mmu.r_valid_d[7] ;
 wire \cpu.genblk1.mmu.r_valid_d[8] ;
 wire \cpu.genblk1.mmu.r_valid_d[9] ;
 wire \cpu.genblk1.mmu.r_valid_i[0] ;
 wire \cpu.genblk1.mmu.r_valid_i[10] ;
 wire \cpu.genblk1.mmu.r_valid_i[11] ;
 wire \cpu.genblk1.mmu.r_valid_i[12] ;
 wire \cpu.genblk1.mmu.r_valid_i[13] ;
 wire \cpu.genblk1.mmu.r_valid_i[14] ;
 wire \cpu.genblk1.mmu.r_valid_i[15] ;
 wire \cpu.genblk1.mmu.r_valid_i[16] ;
 wire \cpu.genblk1.mmu.r_valid_i[17] ;
 wire \cpu.genblk1.mmu.r_valid_i[18] ;
 wire \cpu.genblk1.mmu.r_valid_i[19] ;
 wire \cpu.genblk1.mmu.r_valid_i[1] ;
 wire \cpu.genblk1.mmu.r_valid_i[20] ;
 wire \cpu.genblk1.mmu.r_valid_i[21] ;
 wire \cpu.genblk1.mmu.r_valid_i[22] ;
 wire \cpu.genblk1.mmu.r_valid_i[23] ;
 wire \cpu.genblk1.mmu.r_valid_i[24] ;
 wire \cpu.genblk1.mmu.r_valid_i[25] ;
 wire \cpu.genblk1.mmu.r_valid_i[26] ;
 wire \cpu.genblk1.mmu.r_valid_i[27] ;
 wire \cpu.genblk1.mmu.r_valid_i[28] ;
 wire \cpu.genblk1.mmu.r_valid_i[29] ;
 wire \cpu.genblk1.mmu.r_valid_i[2] ;
 wire \cpu.genblk1.mmu.r_valid_i[30] ;
 wire \cpu.genblk1.mmu.r_valid_i[31] ;
 wire \cpu.genblk1.mmu.r_valid_i[3] ;
 wire \cpu.genblk1.mmu.r_valid_i[4] ;
 wire \cpu.genblk1.mmu.r_valid_i[5] ;
 wire \cpu.genblk1.mmu.r_valid_i[6] ;
 wire \cpu.genblk1.mmu.r_valid_i[7] ;
 wire \cpu.genblk1.mmu.r_valid_i[8] ;
 wire \cpu.genblk1.mmu.r_valid_i[9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_d[9][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[0][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[10][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[11][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[12][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[13][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[14][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[15][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[16][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[17][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[18][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[19][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[1][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[20][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[21][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[22][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[23][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[24][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[25][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[26][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[27][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[28][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[29][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[2][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[30][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[31][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[3][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[4][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[5][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[6][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[7][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[8][9] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][0] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][10] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][11] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][1] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][2] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][3] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][4] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][5] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][6] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][7] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][8] ;
 wire \cpu.genblk1.mmu.r_vtop_i[9][9] ;
 wire \cpu.genblk1.mmu.r_writeable_d[0] ;
 wire \cpu.genblk1.mmu.r_writeable_d[10] ;
 wire \cpu.genblk1.mmu.r_writeable_d[11] ;
 wire \cpu.genblk1.mmu.r_writeable_d[12] ;
 wire \cpu.genblk1.mmu.r_writeable_d[13] ;
 wire \cpu.genblk1.mmu.r_writeable_d[14] ;
 wire \cpu.genblk1.mmu.r_writeable_d[15] ;
 wire \cpu.genblk1.mmu.r_writeable_d[16] ;
 wire \cpu.genblk1.mmu.r_writeable_d[17] ;
 wire \cpu.genblk1.mmu.r_writeable_d[18] ;
 wire \cpu.genblk1.mmu.r_writeable_d[19] ;
 wire \cpu.genblk1.mmu.r_writeable_d[1] ;
 wire \cpu.genblk1.mmu.r_writeable_d[20] ;
 wire \cpu.genblk1.mmu.r_writeable_d[21] ;
 wire \cpu.genblk1.mmu.r_writeable_d[22] ;
 wire \cpu.genblk1.mmu.r_writeable_d[23] ;
 wire \cpu.genblk1.mmu.r_writeable_d[24] ;
 wire \cpu.genblk1.mmu.r_writeable_d[25] ;
 wire \cpu.genblk1.mmu.r_writeable_d[26] ;
 wire \cpu.genblk1.mmu.r_writeable_d[27] ;
 wire \cpu.genblk1.mmu.r_writeable_d[28] ;
 wire \cpu.genblk1.mmu.r_writeable_d[29] ;
 wire \cpu.genblk1.mmu.r_writeable_d[2] ;
 wire \cpu.genblk1.mmu.r_writeable_d[30] ;
 wire \cpu.genblk1.mmu.r_writeable_d[31] ;
 wire \cpu.genblk1.mmu.r_writeable_d[3] ;
 wire \cpu.genblk1.mmu.r_writeable_d[4] ;
 wire \cpu.genblk1.mmu.r_writeable_d[5] ;
 wire \cpu.genblk1.mmu.r_writeable_d[6] ;
 wire \cpu.genblk1.mmu.r_writeable_d[7] ;
 wire \cpu.genblk1.mmu.r_writeable_d[8] ;
 wire \cpu.genblk1.mmu.r_writeable_d[9] ;
 wire \cpu.gpio.genblk1[3].srcs_o[0] ;
 wire \cpu.gpio.genblk1[3].srcs_o[11] ;
 wire \cpu.gpio.genblk1[3].srcs_o[1] ;
 wire \cpu.gpio.genblk1[3].srcs_o[2] ;
 wire \cpu.gpio.genblk1[3].srcs_o[3] ;
 wire \cpu.gpio.genblk1[3].srcs_o[4] ;
 wire \cpu.gpio.genblk1[3].srcs_o[5] ;
 wire \cpu.gpio.genblk1[3].srcs_o[6] ;
 wire \cpu.gpio.genblk1[3].srcs_o[7] ;
 wire \cpu.gpio.genblk1[3].srcs_o[8] ;
 wire \cpu.gpio.genblk1[4].srcs_o[0] ;
 wire \cpu.gpio.genblk1[5].srcs_o[0] ;
 wire \cpu.gpio.genblk1[6].srcs_o[0] ;
 wire \cpu.gpio.genblk1[7].srcs_o[0] ;
 wire \cpu.gpio.genblk2[4].srcs_io[0] ;
 wire \cpu.gpio.genblk2[5].srcs_io[0] ;
 wire \cpu.gpio.genblk2[6].srcs_io[0] ;
 wire \cpu.gpio.genblk2[7].srcs_io[0] ;
 wire \cpu.gpio.r_enable_in[0] ;
 wire \cpu.gpio.r_enable_in[1] ;
 wire \cpu.gpio.r_enable_in[2] ;
 wire \cpu.gpio.r_enable_in[3] ;
 wire \cpu.gpio.r_enable_in[4] ;
 wire \cpu.gpio.r_enable_in[5] ;
 wire \cpu.gpio.r_enable_in[6] ;
 wire \cpu.gpio.r_enable_in[7] ;
 wire \cpu.gpio.r_enable_io[4] ;
 wire \cpu.gpio.r_enable_io[5] ;
 wire \cpu.gpio.r_enable_io[6] ;
 wire \cpu.gpio.r_enable_io[7] ;
 wire \cpu.gpio.r_spi_miso_src[0][0] ;
 wire \cpu.gpio.r_spi_miso_src[0][1] ;
 wire \cpu.gpio.r_spi_miso_src[0][2] ;
 wire \cpu.gpio.r_spi_miso_src[0][3] ;
 wire \cpu.gpio.r_spi_miso_src[1][0] ;
 wire \cpu.gpio.r_spi_miso_src[1][1] ;
 wire \cpu.gpio.r_spi_miso_src[1][2] ;
 wire \cpu.gpio.r_spi_miso_src[1][3] ;
 wire \cpu.gpio.r_src_io[4][0] ;
 wire \cpu.gpio.r_src_io[4][1] ;
 wire \cpu.gpio.r_src_io[4][2] ;
 wire \cpu.gpio.r_src_io[4][3] ;
 wire \cpu.gpio.r_src_io[5][0] ;
 wire \cpu.gpio.r_src_io[5][1] ;
 wire \cpu.gpio.r_src_io[5][2] ;
 wire \cpu.gpio.r_src_io[5][3] ;
 wire \cpu.gpio.r_src_io[6][0] ;
 wire \cpu.gpio.r_src_io[6][1] ;
 wire \cpu.gpio.r_src_io[6][2] ;
 wire \cpu.gpio.r_src_io[6][3] ;
 wire \cpu.gpio.r_src_io[7][0] ;
 wire \cpu.gpio.r_src_io[7][1] ;
 wire \cpu.gpio.r_src_io[7][2] ;
 wire \cpu.gpio.r_src_io[7][3] ;
 wire \cpu.gpio.r_src_o[3][0] ;
 wire \cpu.gpio.r_src_o[3][1] ;
 wire \cpu.gpio.r_src_o[3][2] ;
 wire \cpu.gpio.r_src_o[3][3] ;
 wire \cpu.gpio.r_src_o[4][0] ;
 wire \cpu.gpio.r_src_o[4][1] ;
 wire \cpu.gpio.r_src_o[4][2] ;
 wire \cpu.gpio.r_src_o[4][3] ;
 wire \cpu.gpio.r_src_o[5][0] ;
 wire \cpu.gpio.r_src_o[5][1] ;
 wire \cpu.gpio.r_src_o[5][2] ;
 wire \cpu.gpio.r_src_o[5][3] ;
 wire \cpu.gpio.r_src_o[6][0] ;
 wire \cpu.gpio.r_src_o[6][1] ;
 wire \cpu.gpio.r_src_o[6][2] ;
 wire \cpu.gpio.r_src_o[6][3] ;
 wire \cpu.gpio.r_src_o[7][0] ;
 wire \cpu.gpio.r_src_o[7][1] ;
 wire \cpu.gpio.r_src_o[7][2] ;
 wire \cpu.gpio.r_src_o[7][3] ;
 wire \cpu.gpio.r_uart_rx_src[0] ;
 wire \cpu.gpio.r_uart_rx_src[1] ;
 wire \cpu.gpio.r_uart_rx_src[2] ;
 wire \cpu.gpio.uart_rx ;
 wire \cpu.i_wstrobe_d ;
 wire \cpu.icache.r_data[0][0] ;
 wire \cpu.icache.r_data[0][10] ;
 wire \cpu.icache.r_data[0][11] ;
 wire \cpu.icache.r_data[0][12] ;
 wire \cpu.icache.r_data[0][13] ;
 wire \cpu.icache.r_data[0][14] ;
 wire \cpu.icache.r_data[0][15] ;
 wire \cpu.icache.r_data[0][16] ;
 wire \cpu.icache.r_data[0][17] ;
 wire \cpu.icache.r_data[0][18] ;
 wire \cpu.icache.r_data[0][19] ;
 wire \cpu.icache.r_data[0][1] ;
 wire \cpu.icache.r_data[0][20] ;
 wire \cpu.icache.r_data[0][21] ;
 wire \cpu.icache.r_data[0][22] ;
 wire \cpu.icache.r_data[0][23] ;
 wire \cpu.icache.r_data[0][24] ;
 wire \cpu.icache.r_data[0][25] ;
 wire \cpu.icache.r_data[0][26] ;
 wire \cpu.icache.r_data[0][27] ;
 wire \cpu.icache.r_data[0][28] ;
 wire \cpu.icache.r_data[0][29] ;
 wire \cpu.icache.r_data[0][2] ;
 wire \cpu.icache.r_data[0][30] ;
 wire \cpu.icache.r_data[0][31] ;
 wire \cpu.icache.r_data[0][3] ;
 wire \cpu.icache.r_data[0][4] ;
 wire \cpu.icache.r_data[0][5] ;
 wire \cpu.icache.r_data[0][6] ;
 wire \cpu.icache.r_data[0][7] ;
 wire \cpu.icache.r_data[0][8] ;
 wire \cpu.icache.r_data[0][9] ;
 wire \cpu.icache.r_data[1][0] ;
 wire \cpu.icache.r_data[1][10] ;
 wire \cpu.icache.r_data[1][11] ;
 wire \cpu.icache.r_data[1][12] ;
 wire \cpu.icache.r_data[1][13] ;
 wire \cpu.icache.r_data[1][14] ;
 wire \cpu.icache.r_data[1][15] ;
 wire \cpu.icache.r_data[1][16] ;
 wire \cpu.icache.r_data[1][17] ;
 wire \cpu.icache.r_data[1][18] ;
 wire \cpu.icache.r_data[1][19] ;
 wire \cpu.icache.r_data[1][1] ;
 wire \cpu.icache.r_data[1][20] ;
 wire \cpu.icache.r_data[1][21] ;
 wire \cpu.icache.r_data[1][22] ;
 wire \cpu.icache.r_data[1][23] ;
 wire \cpu.icache.r_data[1][24] ;
 wire \cpu.icache.r_data[1][25] ;
 wire \cpu.icache.r_data[1][26] ;
 wire \cpu.icache.r_data[1][27] ;
 wire \cpu.icache.r_data[1][28] ;
 wire \cpu.icache.r_data[1][29] ;
 wire \cpu.icache.r_data[1][2] ;
 wire \cpu.icache.r_data[1][30] ;
 wire \cpu.icache.r_data[1][31] ;
 wire \cpu.icache.r_data[1][3] ;
 wire \cpu.icache.r_data[1][4] ;
 wire \cpu.icache.r_data[1][5] ;
 wire \cpu.icache.r_data[1][6] ;
 wire \cpu.icache.r_data[1][7] ;
 wire \cpu.icache.r_data[1][8] ;
 wire \cpu.icache.r_data[1][9] ;
 wire \cpu.icache.r_data[2][0] ;
 wire \cpu.icache.r_data[2][10] ;
 wire \cpu.icache.r_data[2][11] ;
 wire \cpu.icache.r_data[2][12] ;
 wire \cpu.icache.r_data[2][13] ;
 wire \cpu.icache.r_data[2][14] ;
 wire \cpu.icache.r_data[2][15] ;
 wire \cpu.icache.r_data[2][16] ;
 wire \cpu.icache.r_data[2][17] ;
 wire \cpu.icache.r_data[2][18] ;
 wire \cpu.icache.r_data[2][19] ;
 wire \cpu.icache.r_data[2][1] ;
 wire \cpu.icache.r_data[2][20] ;
 wire \cpu.icache.r_data[2][21] ;
 wire \cpu.icache.r_data[2][22] ;
 wire \cpu.icache.r_data[2][23] ;
 wire \cpu.icache.r_data[2][24] ;
 wire \cpu.icache.r_data[2][25] ;
 wire \cpu.icache.r_data[2][26] ;
 wire \cpu.icache.r_data[2][27] ;
 wire \cpu.icache.r_data[2][28] ;
 wire \cpu.icache.r_data[2][29] ;
 wire \cpu.icache.r_data[2][2] ;
 wire \cpu.icache.r_data[2][30] ;
 wire \cpu.icache.r_data[2][31] ;
 wire \cpu.icache.r_data[2][3] ;
 wire \cpu.icache.r_data[2][4] ;
 wire \cpu.icache.r_data[2][5] ;
 wire \cpu.icache.r_data[2][6] ;
 wire \cpu.icache.r_data[2][7] ;
 wire \cpu.icache.r_data[2][8] ;
 wire \cpu.icache.r_data[2][9] ;
 wire \cpu.icache.r_data[3][0] ;
 wire \cpu.icache.r_data[3][10] ;
 wire \cpu.icache.r_data[3][11] ;
 wire \cpu.icache.r_data[3][12] ;
 wire \cpu.icache.r_data[3][13] ;
 wire \cpu.icache.r_data[3][14] ;
 wire \cpu.icache.r_data[3][15] ;
 wire \cpu.icache.r_data[3][16] ;
 wire \cpu.icache.r_data[3][17] ;
 wire \cpu.icache.r_data[3][18] ;
 wire \cpu.icache.r_data[3][19] ;
 wire \cpu.icache.r_data[3][1] ;
 wire \cpu.icache.r_data[3][20] ;
 wire \cpu.icache.r_data[3][21] ;
 wire \cpu.icache.r_data[3][22] ;
 wire \cpu.icache.r_data[3][23] ;
 wire \cpu.icache.r_data[3][24] ;
 wire \cpu.icache.r_data[3][25] ;
 wire \cpu.icache.r_data[3][26] ;
 wire \cpu.icache.r_data[3][27] ;
 wire \cpu.icache.r_data[3][28] ;
 wire \cpu.icache.r_data[3][29] ;
 wire \cpu.icache.r_data[3][2] ;
 wire \cpu.icache.r_data[3][30] ;
 wire \cpu.icache.r_data[3][31] ;
 wire \cpu.icache.r_data[3][3] ;
 wire \cpu.icache.r_data[3][4] ;
 wire \cpu.icache.r_data[3][5] ;
 wire \cpu.icache.r_data[3][6] ;
 wire \cpu.icache.r_data[3][7] ;
 wire \cpu.icache.r_data[3][8] ;
 wire \cpu.icache.r_data[3][9] ;
 wire \cpu.icache.r_data[4][0] ;
 wire \cpu.icache.r_data[4][10] ;
 wire \cpu.icache.r_data[4][11] ;
 wire \cpu.icache.r_data[4][12] ;
 wire \cpu.icache.r_data[4][13] ;
 wire \cpu.icache.r_data[4][14] ;
 wire \cpu.icache.r_data[4][15] ;
 wire \cpu.icache.r_data[4][16] ;
 wire \cpu.icache.r_data[4][17] ;
 wire \cpu.icache.r_data[4][18] ;
 wire \cpu.icache.r_data[4][19] ;
 wire \cpu.icache.r_data[4][1] ;
 wire \cpu.icache.r_data[4][20] ;
 wire \cpu.icache.r_data[4][21] ;
 wire \cpu.icache.r_data[4][22] ;
 wire \cpu.icache.r_data[4][23] ;
 wire \cpu.icache.r_data[4][24] ;
 wire \cpu.icache.r_data[4][25] ;
 wire \cpu.icache.r_data[4][26] ;
 wire \cpu.icache.r_data[4][27] ;
 wire \cpu.icache.r_data[4][28] ;
 wire \cpu.icache.r_data[4][29] ;
 wire \cpu.icache.r_data[4][2] ;
 wire \cpu.icache.r_data[4][30] ;
 wire \cpu.icache.r_data[4][31] ;
 wire \cpu.icache.r_data[4][3] ;
 wire \cpu.icache.r_data[4][4] ;
 wire \cpu.icache.r_data[4][5] ;
 wire \cpu.icache.r_data[4][6] ;
 wire \cpu.icache.r_data[4][7] ;
 wire \cpu.icache.r_data[4][8] ;
 wire \cpu.icache.r_data[4][9] ;
 wire \cpu.icache.r_data[5][0] ;
 wire \cpu.icache.r_data[5][10] ;
 wire \cpu.icache.r_data[5][11] ;
 wire \cpu.icache.r_data[5][12] ;
 wire \cpu.icache.r_data[5][13] ;
 wire \cpu.icache.r_data[5][14] ;
 wire \cpu.icache.r_data[5][15] ;
 wire \cpu.icache.r_data[5][16] ;
 wire \cpu.icache.r_data[5][17] ;
 wire \cpu.icache.r_data[5][18] ;
 wire \cpu.icache.r_data[5][19] ;
 wire \cpu.icache.r_data[5][1] ;
 wire \cpu.icache.r_data[5][20] ;
 wire \cpu.icache.r_data[5][21] ;
 wire \cpu.icache.r_data[5][22] ;
 wire \cpu.icache.r_data[5][23] ;
 wire \cpu.icache.r_data[5][24] ;
 wire \cpu.icache.r_data[5][25] ;
 wire \cpu.icache.r_data[5][26] ;
 wire \cpu.icache.r_data[5][27] ;
 wire \cpu.icache.r_data[5][28] ;
 wire \cpu.icache.r_data[5][29] ;
 wire \cpu.icache.r_data[5][2] ;
 wire \cpu.icache.r_data[5][30] ;
 wire \cpu.icache.r_data[5][31] ;
 wire \cpu.icache.r_data[5][3] ;
 wire \cpu.icache.r_data[5][4] ;
 wire \cpu.icache.r_data[5][5] ;
 wire \cpu.icache.r_data[5][6] ;
 wire \cpu.icache.r_data[5][7] ;
 wire \cpu.icache.r_data[5][8] ;
 wire \cpu.icache.r_data[5][9] ;
 wire \cpu.icache.r_data[6][0] ;
 wire \cpu.icache.r_data[6][10] ;
 wire \cpu.icache.r_data[6][11] ;
 wire \cpu.icache.r_data[6][12] ;
 wire \cpu.icache.r_data[6][13] ;
 wire \cpu.icache.r_data[6][14] ;
 wire \cpu.icache.r_data[6][15] ;
 wire \cpu.icache.r_data[6][16] ;
 wire \cpu.icache.r_data[6][17] ;
 wire \cpu.icache.r_data[6][18] ;
 wire \cpu.icache.r_data[6][19] ;
 wire \cpu.icache.r_data[6][1] ;
 wire \cpu.icache.r_data[6][20] ;
 wire \cpu.icache.r_data[6][21] ;
 wire \cpu.icache.r_data[6][22] ;
 wire \cpu.icache.r_data[6][23] ;
 wire \cpu.icache.r_data[6][24] ;
 wire \cpu.icache.r_data[6][25] ;
 wire \cpu.icache.r_data[6][26] ;
 wire \cpu.icache.r_data[6][27] ;
 wire \cpu.icache.r_data[6][28] ;
 wire \cpu.icache.r_data[6][29] ;
 wire \cpu.icache.r_data[6][2] ;
 wire \cpu.icache.r_data[6][30] ;
 wire \cpu.icache.r_data[6][31] ;
 wire \cpu.icache.r_data[6][3] ;
 wire \cpu.icache.r_data[6][4] ;
 wire \cpu.icache.r_data[6][5] ;
 wire \cpu.icache.r_data[6][6] ;
 wire \cpu.icache.r_data[6][7] ;
 wire \cpu.icache.r_data[6][8] ;
 wire \cpu.icache.r_data[6][9] ;
 wire \cpu.icache.r_data[7][0] ;
 wire \cpu.icache.r_data[7][10] ;
 wire \cpu.icache.r_data[7][11] ;
 wire \cpu.icache.r_data[7][12] ;
 wire \cpu.icache.r_data[7][13] ;
 wire \cpu.icache.r_data[7][14] ;
 wire \cpu.icache.r_data[7][15] ;
 wire \cpu.icache.r_data[7][16] ;
 wire \cpu.icache.r_data[7][17] ;
 wire \cpu.icache.r_data[7][18] ;
 wire \cpu.icache.r_data[7][19] ;
 wire \cpu.icache.r_data[7][1] ;
 wire \cpu.icache.r_data[7][20] ;
 wire \cpu.icache.r_data[7][21] ;
 wire \cpu.icache.r_data[7][22] ;
 wire \cpu.icache.r_data[7][23] ;
 wire \cpu.icache.r_data[7][24] ;
 wire \cpu.icache.r_data[7][25] ;
 wire \cpu.icache.r_data[7][26] ;
 wire \cpu.icache.r_data[7][27] ;
 wire \cpu.icache.r_data[7][28] ;
 wire \cpu.icache.r_data[7][29] ;
 wire \cpu.icache.r_data[7][2] ;
 wire \cpu.icache.r_data[7][30] ;
 wire \cpu.icache.r_data[7][31] ;
 wire \cpu.icache.r_data[7][3] ;
 wire \cpu.icache.r_data[7][4] ;
 wire \cpu.icache.r_data[7][5] ;
 wire \cpu.icache.r_data[7][6] ;
 wire \cpu.icache.r_data[7][7] ;
 wire \cpu.icache.r_data[7][8] ;
 wire \cpu.icache.r_data[7][9] ;
 wire \cpu.icache.r_offset[0] ;
 wire \cpu.icache.r_offset[1] ;
 wire \cpu.icache.r_offset[2] ;
 wire \cpu.icache.r_tag[0][10] ;
 wire \cpu.icache.r_tag[0][11] ;
 wire \cpu.icache.r_tag[0][12] ;
 wire \cpu.icache.r_tag[0][13] ;
 wire \cpu.icache.r_tag[0][14] ;
 wire \cpu.icache.r_tag[0][15] ;
 wire \cpu.icache.r_tag[0][16] ;
 wire \cpu.icache.r_tag[0][17] ;
 wire \cpu.icache.r_tag[0][18] ;
 wire \cpu.icache.r_tag[0][19] ;
 wire \cpu.icache.r_tag[0][20] ;
 wire \cpu.icache.r_tag[0][21] ;
 wire \cpu.icache.r_tag[0][22] ;
 wire \cpu.icache.r_tag[0][23] ;
 wire \cpu.icache.r_tag[0][5] ;
 wire \cpu.icache.r_tag[0][6] ;
 wire \cpu.icache.r_tag[0][7] ;
 wire \cpu.icache.r_tag[0][8] ;
 wire \cpu.icache.r_tag[0][9] ;
 wire \cpu.icache.r_tag[1][10] ;
 wire \cpu.icache.r_tag[1][11] ;
 wire \cpu.icache.r_tag[1][12] ;
 wire \cpu.icache.r_tag[1][13] ;
 wire \cpu.icache.r_tag[1][14] ;
 wire \cpu.icache.r_tag[1][15] ;
 wire \cpu.icache.r_tag[1][16] ;
 wire \cpu.icache.r_tag[1][17] ;
 wire \cpu.icache.r_tag[1][18] ;
 wire \cpu.icache.r_tag[1][19] ;
 wire \cpu.icache.r_tag[1][20] ;
 wire \cpu.icache.r_tag[1][21] ;
 wire \cpu.icache.r_tag[1][22] ;
 wire \cpu.icache.r_tag[1][23] ;
 wire \cpu.icache.r_tag[1][5] ;
 wire \cpu.icache.r_tag[1][6] ;
 wire \cpu.icache.r_tag[1][7] ;
 wire \cpu.icache.r_tag[1][8] ;
 wire \cpu.icache.r_tag[1][9] ;
 wire \cpu.icache.r_tag[2][10] ;
 wire \cpu.icache.r_tag[2][11] ;
 wire \cpu.icache.r_tag[2][12] ;
 wire \cpu.icache.r_tag[2][13] ;
 wire \cpu.icache.r_tag[2][14] ;
 wire \cpu.icache.r_tag[2][15] ;
 wire \cpu.icache.r_tag[2][16] ;
 wire \cpu.icache.r_tag[2][17] ;
 wire \cpu.icache.r_tag[2][18] ;
 wire \cpu.icache.r_tag[2][19] ;
 wire \cpu.icache.r_tag[2][20] ;
 wire \cpu.icache.r_tag[2][21] ;
 wire \cpu.icache.r_tag[2][22] ;
 wire \cpu.icache.r_tag[2][23] ;
 wire \cpu.icache.r_tag[2][5] ;
 wire \cpu.icache.r_tag[2][6] ;
 wire \cpu.icache.r_tag[2][7] ;
 wire \cpu.icache.r_tag[2][8] ;
 wire \cpu.icache.r_tag[2][9] ;
 wire \cpu.icache.r_tag[3][10] ;
 wire \cpu.icache.r_tag[3][11] ;
 wire \cpu.icache.r_tag[3][12] ;
 wire \cpu.icache.r_tag[3][13] ;
 wire \cpu.icache.r_tag[3][14] ;
 wire \cpu.icache.r_tag[3][15] ;
 wire \cpu.icache.r_tag[3][16] ;
 wire \cpu.icache.r_tag[3][17] ;
 wire \cpu.icache.r_tag[3][18] ;
 wire \cpu.icache.r_tag[3][19] ;
 wire \cpu.icache.r_tag[3][20] ;
 wire \cpu.icache.r_tag[3][21] ;
 wire \cpu.icache.r_tag[3][22] ;
 wire \cpu.icache.r_tag[3][23] ;
 wire \cpu.icache.r_tag[3][5] ;
 wire \cpu.icache.r_tag[3][6] ;
 wire \cpu.icache.r_tag[3][7] ;
 wire \cpu.icache.r_tag[3][8] ;
 wire \cpu.icache.r_tag[3][9] ;
 wire \cpu.icache.r_tag[4][10] ;
 wire \cpu.icache.r_tag[4][11] ;
 wire \cpu.icache.r_tag[4][12] ;
 wire \cpu.icache.r_tag[4][13] ;
 wire \cpu.icache.r_tag[4][14] ;
 wire \cpu.icache.r_tag[4][15] ;
 wire \cpu.icache.r_tag[4][16] ;
 wire \cpu.icache.r_tag[4][17] ;
 wire \cpu.icache.r_tag[4][18] ;
 wire \cpu.icache.r_tag[4][19] ;
 wire \cpu.icache.r_tag[4][20] ;
 wire \cpu.icache.r_tag[4][21] ;
 wire \cpu.icache.r_tag[4][22] ;
 wire \cpu.icache.r_tag[4][23] ;
 wire \cpu.icache.r_tag[4][5] ;
 wire \cpu.icache.r_tag[4][6] ;
 wire \cpu.icache.r_tag[4][7] ;
 wire \cpu.icache.r_tag[4][8] ;
 wire \cpu.icache.r_tag[4][9] ;
 wire \cpu.icache.r_tag[5][10] ;
 wire \cpu.icache.r_tag[5][11] ;
 wire \cpu.icache.r_tag[5][12] ;
 wire \cpu.icache.r_tag[5][13] ;
 wire \cpu.icache.r_tag[5][14] ;
 wire \cpu.icache.r_tag[5][15] ;
 wire \cpu.icache.r_tag[5][16] ;
 wire \cpu.icache.r_tag[5][17] ;
 wire \cpu.icache.r_tag[5][18] ;
 wire \cpu.icache.r_tag[5][19] ;
 wire \cpu.icache.r_tag[5][20] ;
 wire \cpu.icache.r_tag[5][21] ;
 wire \cpu.icache.r_tag[5][22] ;
 wire \cpu.icache.r_tag[5][23] ;
 wire \cpu.icache.r_tag[5][5] ;
 wire \cpu.icache.r_tag[5][6] ;
 wire \cpu.icache.r_tag[5][7] ;
 wire \cpu.icache.r_tag[5][8] ;
 wire \cpu.icache.r_tag[5][9] ;
 wire \cpu.icache.r_tag[6][10] ;
 wire \cpu.icache.r_tag[6][11] ;
 wire \cpu.icache.r_tag[6][12] ;
 wire \cpu.icache.r_tag[6][13] ;
 wire \cpu.icache.r_tag[6][14] ;
 wire \cpu.icache.r_tag[6][15] ;
 wire \cpu.icache.r_tag[6][16] ;
 wire \cpu.icache.r_tag[6][17] ;
 wire \cpu.icache.r_tag[6][18] ;
 wire \cpu.icache.r_tag[6][19] ;
 wire \cpu.icache.r_tag[6][20] ;
 wire \cpu.icache.r_tag[6][21] ;
 wire \cpu.icache.r_tag[6][22] ;
 wire \cpu.icache.r_tag[6][23] ;
 wire \cpu.icache.r_tag[6][5] ;
 wire \cpu.icache.r_tag[6][6] ;
 wire \cpu.icache.r_tag[6][7] ;
 wire \cpu.icache.r_tag[6][8] ;
 wire \cpu.icache.r_tag[6][9] ;
 wire \cpu.icache.r_tag[7][10] ;
 wire \cpu.icache.r_tag[7][11] ;
 wire \cpu.icache.r_tag[7][12] ;
 wire \cpu.icache.r_tag[7][13] ;
 wire \cpu.icache.r_tag[7][14] ;
 wire \cpu.icache.r_tag[7][15] ;
 wire \cpu.icache.r_tag[7][16] ;
 wire \cpu.icache.r_tag[7][17] ;
 wire \cpu.icache.r_tag[7][18] ;
 wire \cpu.icache.r_tag[7][19] ;
 wire \cpu.icache.r_tag[7][20] ;
 wire \cpu.icache.r_tag[7][21] ;
 wire \cpu.icache.r_tag[7][22] ;
 wire \cpu.icache.r_tag[7][23] ;
 wire \cpu.icache.r_tag[7][5] ;
 wire \cpu.icache.r_tag[7][6] ;
 wire \cpu.icache.r_tag[7][7] ;
 wire \cpu.icache.r_tag[7][8] ;
 wire \cpu.icache.r_tag[7][9] ;
 wire \cpu.icache.r_valid[0] ;
 wire \cpu.icache.r_valid[1] ;
 wire \cpu.icache.r_valid[2] ;
 wire \cpu.icache.r_valid[3] ;
 wire \cpu.icache.r_valid[4] ;
 wire \cpu.icache.r_valid[5] ;
 wire \cpu.icache.r_valid[6] ;
 wire \cpu.icache.r_valid[7] ;
 wire \cpu.intr.r_clock ;
 wire \cpu.intr.r_clock_cmp[0] ;
 wire \cpu.intr.r_clock_cmp[10] ;
 wire \cpu.intr.r_clock_cmp[11] ;
 wire \cpu.intr.r_clock_cmp[12] ;
 wire \cpu.intr.r_clock_cmp[13] ;
 wire \cpu.intr.r_clock_cmp[14] ;
 wire \cpu.intr.r_clock_cmp[15] ;
 wire \cpu.intr.r_clock_cmp[16] ;
 wire \cpu.intr.r_clock_cmp[17] ;
 wire \cpu.intr.r_clock_cmp[18] ;
 wire \cpu.intr.r_clock_cmp[19] ;
 wire \cpu.intr.r_clock_cmp[1] ;
 wire \cpu.intr.r_clock_cmp[20] ;
 wire \cpu.intr.r_clock_cmp[21] ;
 wire \cpu.intr.r_clock_cmp[22] ;
 wire \cpu.intr.r_clock_cmp[23] ;
 wire \cpu.intr.r_clock_cmp[24] ;
 wire \cpu.intr.r_clock_cmp[25] ;
 wire \cpu.intr.r_clock_cmp[26] ;
 wire \cpu.intr.r_clock_cmp[27] ;
 wire \cpu.intr.r_clock_cmp[28] ;
 wire \cpu.intr.r_clock_cmp[29] ;
 wire \cpu.intr.r_clock_cmp[2] ;
 wire \cpu.intr.r_clock_cmp[30] ;
 wire \cpu.intr.r_clock_cmp[31] ;
 wire \cpu.intr.r_clock_cmp[3] ;
 wire \cpu.intr.r_clock_cmp[4] ;
 wire \cpu.intr.r_clock_cmp[5] ;
 wire \cpu.intr.r_clock_cmp[6] ;
 wire \cpu.intr.r_clock_cmp[7] ;
 wire \cpu.intr.r_clock_cmp[8] ;
 wire \cpu.intr.r_clock_cmp[9] ;
 wire \cpu.intr.r_clock_count[0] ;
 wire \cpu.intr.r_clock_count[10] ;
 wire \cpu.intr.r_clock_count[11] ;
 wire \cpu.intr.r_clock_count[12] ;
 wire \cpu.intr.r_clock_count[13] ;
 wire \cpu.intr.r_clock_count[14] ;
 wire \cpu.intr.r_clock_count[15] ;
 wire \cpu.intr.r_clock_count[16] ;
 wire \cpu.intr.r_clock_count[17] ;
 wire \cpu.intr.r_clock_count[18] ;
 wire \cpu.intr.r_clock_count[19] ;
 wire \cpu.intr.r_clock_count[1] ;
 wire \cpu.intr.r_clock_count[20] ;
 wire \cpu.intr.r_clock_count[21] ;
 wire \cpu.intr.r_clock_count[22] ;
 wire \cpu.intr.r_clock_count[23] ;
 wire \cpu.intr.r_clock_count[24] ;
 wire \cpu.intr.r_clock_count[25] ;
 wire \cpu.intr.r_clock_count[26] ;
 wire \cpu.intr.r_clock_count[27] ;
 wire \cpu.intr.r_clock_count[28] ;
 wire \cpu.intr.r_clock_count[29] ;
 wire \cpu.intr.r_clock_count[2] ;
 wire \cpu.intr.r_clock_count[30] ;
 wire \cpu.intr.r_clock_count[31] ;
 wire \cpu.intr.r_clock_count[3] ;
 wire \cpu.intr.r_clock_count[4] ;
 wire \cpu.intr.r_clock_count[5] ;
 wire \cpu.intr.r_clock_count[6] ;
 wire \cpu.intr.r_clock_count[7] ;
 wire \cpu.intr.r_clock_count[8] ;
 wire \cpu.intr.r_clock_count[9] ;
 wire \cpu.intr.r_enable[0] ;
 wire \cpu.intr.r_enable[1] ;
 wire \cpu.intr.r_enable[2] ;
 wire \cpu.intr.r_enable[3] ;
 wire \cpu.intr.r_enable[4] ;
 wire \cpu.intr.r_enable[5] ;
 wire \cpu.intr.r_swi ;
 wire \cpu.intr.r_timer ;
 wire \cpu.intr.r_timer_count[0] ;
 wire \cpu.intr.r_timer_count[10] ;
 wire \cpu.intr.r_timer_count[11] ;
 wire \cpu.intr.r_timer_count[12] ;
 wire \cpu.intr.r_timer_count[13] ;
 wire \cpu.intr.r_timer_count[14] ;
 wire \cpu.intr.r_timer_count[15] ;
 wire \cpu.intr.r_timer_count[16] ;
 wire \cpu.intr.r_timer_count[17] ;
 wire \cpu.intr.r_timer_count[18] ;
 wire \cpu.intr.r_timer_count[19] ;
 wire \cpu.intr.r_timer_count[1] ;
 wire \cpu.intr.r_timer_count[20] ;
 wire \cpu.intr.r_timer_count[21] ;
 wire \cpu.intr.r_timer_count[22] ;
 wire \cpu.intr.r_timer_count[23] ;
 wire \cpu.intr.r_timer_count[2] ;
 wire \cpu.intr.r_timer_count[3] ;
 wire \cpu.intr.r_timer_count[4] ;
 wire \cpu.intr.r_timer_count[5] ;
 wire \cpu.intr.r_timer_count[6] ;
 wire \cpu.intr.r_timer_count[7] ;
 wire \cpu.intr.r_timer_count[8] ;
 wire \cpu.intr.r_timer_count[9] ;
 wire \cpu.intr.r_timer_reload[0] ;
 wire \cpu.intr.r_timer_reload[10] ;
 wire \cpu.intr.r_timer_reload[11] ;
 wire \cpu.intr.r_timer_reload[12] ;
 wire \cpu.intr.r_timer_reload[13] ;
 wire \cpu.intr.r_timer_reload[14] ;
 wire \cpu.intr.r_timer_reload[15] ;
 wire \cpu.intr.r_timer_reload[16] ;
 wire \cpu.intr.r_timer_reload[17] ;
 wire \cpu.intr.r_timer_reload[18] ;
 wire \cpu.intr.r_timer_reload[19] ;
 wire \cpu.intr.r_timer_reload[1] ;
 wire \cpu.intr.r_timer_reload[20] ;
 wire \cpu.intr.r_timer_reload[21] ;
 wire \cpu.intr.r_timer_reload[22] ;
 wire \cpu.intr.r_timer_reload[23] ;
 wire \cpu.intr.r_timer_reload[2] ;
 wire \cpu.intr.r_timer_reload[3] ;
 wire \cpu.intr.r_timer_reload[4] ;
 wire \cpu.intr.r_timer_reload[5] ;
 wire \cpu.intr.r_timer_reload[6] ;
 wire \cpu.intr.r_timer_reload[7] ;
 wire \cpu.intr.r_timer_reload[8] ;
 wire \cpu.intr.r_timer_reload[9] ;
 wire \cpu.intr.spi_intr ;
 wire \cpu.qspi.c_rstrobe_d ;
 wire \cpu.qspi.c_wstrobe_d ;
 wire \cpu.qspi.c_wstrobe_i ;
 wire \cpu.qspi.r_count[0] ;
 wire \cpu.qspi.r_count[1] ;
 wire \cpu.qspi.r_count[2] ;
 wire \cpu.qspi.r_count[3] ;
 wire \cpu.qspi.r_count[4] ;
 wire \cpu.qspi.r_ind ;
 wire \cpu.qspi.r_mask[0] ;
 wire \cpu.qspi.r_mask[1] ;
 wire \cpu.qspi.r_mask[2] ;
 wire \cpu.qspi.r_quad[0] ;
 wire \cpu.qspi.r_quad[1] ;
 wire \cpu.qspi.r_quad[2] ;
 wire \cpu.qspi.r_read_delay[0][0] ;
 wire \cpu.qspi.r_read_delay[0][1] ;
 wire \cpu.qspi.r_read_delay[0][2] ;
 wire \cpu.qspi.r_read_delay[0][3] ;
 wire \cpu.qspi.r_read_delay[1][0] ;
 wire \cpu.qspi.r_read_delay[1][1] ;
 wire \cpu.qspi.r_read_delay[1][2] ;
 wire \cpu.qspi.r_read_delay[1][3] ;
 wire \cpu.qspi.r_read_delay[2][0] ;
 wire \cpu.qspi.r_read_delay[2][1] ;
 wire \cpu.qspi.r_read_delay[2][2] ;
 wire \cpu.qspi.r_read_delay[2][3] ;
 wire \cpu.qspi.r_rom_mode[0] ;
 wire \cpu.qspi.r_rom_mode[1] ;
 wire \cpu.qspi.r_state[0] ;
 wire \cpu.qspi.r_state[10] ;
 wire \cpu.qspi.r_state[11] ;
 wire \cpu.qspi.r_state[12] ;
 wire \cpu.qspi.r_state[13] ;
 wire \cpu.qspi.r_state[14] ;
 wire \cpu.qspi.r_state[15] ;
 wire \cpu.qspi.r_state[16] ;
 wire \cpu.qspi.r_state[17] ;
 wire \cpu.qspi.r_state[1] ;
 wire \cpu.qspi.r_state[2] ;
 wire \cpu.qspi.r_state[3] ;
 wire \cpu.qspi.r_state[4] ;
 wire \cpu.qspi.r_state[5] ;
 wire \cpu.qspi.r_state[6] ;
 wire \cpu.qspi.r_state[7] ;
 wire \cpu.qspi.r_state[8] ;
 wire \cpu.qspi.r_state[9] ;
 wire \cpu.r_clk_invert ;
 wire \cpu.spi.r_bits[0] ;
 wire \cpu.spi.r_bits[1] ;
 wire \cpu.spi.r_bits[2] ;
 wire \cpu.spi.r_clk_count[0][0] ;
 wire \cpu.spi.r_clk_count[0][1] ;
 wire \cpu.spi.r_clk_count[0][2] ;
 wire \cpu.spi.r_clk_count[0][3] ;
 wire \cpu.spi.r_clk_count[0][4] ;
 wire \cpu.spi.r_clk_count[0][5] ;
 wire \cpu.spi.r_clk_count[0][6] ;
 wire \cpu.spi.r_clk_count[0][7] ;
 wire \cpu.spi.r_clk_count[1][0] ;
 wire \cpu.spi.r_clk_count[1][1] ;
 wire \cpu.spi.r_clk_count[1][2] ;
 wire \cpu.spi.r_clk_count[1][3] ;
 wire \cpu.spi.r_clk_count[1][4] ;
 wire \cpu.spi.r_clk_count[1][5] ;
 wire \cpu.spi.r_clk_count[1][6] ;
 wire \cpu.spi.r_clk_count[1][7] ;
 wire \cpu.spi.r_clk_count[2][0] ;
 wire \cpu.spi.r_clk_count[2][1] ;
 wire \cpu.spi.r_clk_count[2][2] ;
 wire \cpu.spi.r_clk_count[2][3] ;
 wire \cpu.spi.r_clk_count[2][4] ;
 wire \cpu.spi.r_clk_count[2][5] ;
 wire \cpu.spi.r_clk_count[2][6] ;
 wire \cpu.spi.r_clk_count[2][7] ;
 wire \cpu.spi.r_count[0] ;
 wire \cpu.spi.r_count[1] ;
 wire \cpu.spi.r_count[2] ;
 wire \cpu.spi.r_count[3] ;
 wire \cpu.spi.r_count[4] ;
 wire \cpu.spi.r_count[5] ;
 wire \cpu.spi.r_count[6] ;
 wire \cpu.spi.r_count[7] ;
 wire \cpu.spi.r_in[0] ;
 wire \cpu.spi.r_in[1] ;
 wire \cpu.spi.r_in[2] ;
 wire \cpu.spi.r_in[3] ;
 wire \cpu.spi.r_in[4] ;
 wire \cpu.spi.r_in[5] ;
 wire \cpu.spi.r_in[6] ;
 wire \cpu.spi.r_in[7] ;
 wire \cpu.spi.r_mode[0][0] ;
 wire \cpu.spi.r_mode[0][1] ;
 wire \cpu.spi.r_mode[1][0] ;
 wire \cpu.spi.r_mode[1][1] ;
 wire \cpu.spi.r_mode[2][0] ;
 wire \cpu.spi.r_mode[2][1] ;
 wire \cpu.spi.r_out[0] ;
 wire \cpu.spi.r_out[1] ;
 wire \cpu.spi.r_out[2] ;
 wire \cpu.spi.r_out[3] ;
 wire \cpu.spi.r_out[4] ;
 wire \cpu.spi.r_out[5] ;
 wire \cpu.spi.r_out[6] ;
 wire \cpu.spi.r_out[7] ;
 wire \cpu.spi.r_ready ;
 wire \cpu.spi.r_searching ;
 wire \cpu.spi.r_sel[0] ;
 wire \cpu.spi.r_sel[1] ;
 wire \cpu.spi.r_src[0] ;
 wire \cpu.spi.r_src[1] ;
 wire \cpu.spi.r_src[2] ;
 wire \cpu.spi.r_state[0] ;
 wire \cpu.spi.r_state[1] ;
 wire \cpu.spi.r_state[2] ;
 wire \cpu.spi.r_state[3] ;
 wire \cpu.spi.r_state[4] ;
 wire \cpu.spi.r_state[5] ;
 wire \cpu.spi.r_state[6] ;
 wire \cpu.spi.r_timeout[0] ;
 wire \cpu.spi.r_timeout[1] ;
 wire \cpu.spi.r_timeout[2] ;
 wire \cpu.spi.r_timeout[3] ;
 wire \cpu.spi.r_timeout[4] ;
 wire \cpu.spi.r_timeout[5] ;
 wire \cpu.spi.r_timeout[6] ;
 wire \cpu.spi.r_timeout[7] ;
 wire \cpu.spi.r_timeout_count[0] ;
 wire \cpu.spi.r_timeout_count[1] ;
 wire \cpu.spi.r_timeout_count[2] ;
 wire \cpu.spi.r_timeout_count[3] ;
 wire \cpu.spi.r_timeout_count[4] ;
 wire \cpu.spi.r_timeout_count[5] ;
 wire \cpu.spi.r_timeout_count[6] ;
 wire \cpu.spi.r_timeout_count[7] ;
 wire \cpu.uart.r_div[0] ;
 wire \cpu.uart.r_div[10] ;
 wire \cpu.uart.r_div[11] ;
 wire \cpu.uart.r_div[1] ;
 wire \cpu.uart.r_div[2] ;
 wire \cpu.uart.r_div[3] ;
 wire \cpu.uart.r_div[4] ;
 wire \cpu.uart.r_div[5] ;
 wire \cpu.uart.r_div[6] ;
 wire \cpu.uart.r_div[7] ;
 wire \cpu.uart.r_div[8] ;
 wire \cpu.uart.r_div[9] ;
 wire \cpu.uart.r_div_value[0] ;
 wire \cpu.uart.r_div_value[10] ;
 wire \cpu.uart.r_div_value[11] ;
 wire \cpu.uart.r_div_value[1] ;
 wire \cpu.uart.r_div_value[2] ;
 wire \cpu.uart.r_div_value[3] ;
 wire \cpu.uart.r_div_value[4] ;
 wire \cpu.uart.r_div_value[5] ;
 wire \cpu.uart.r_div_value[6] ;
 wire \cpu.uart.r_div_value[7] ;
 wire \cpu.uart.r_div_value[8] ;
 wire \cpu.uart.r_div_value[9] ;
 wire \cpu.uart.r_ib[0] ;
 wire \cpu.uart.r_ib[1] ;
 wire \cpu.uart.r_ib[2] ;
 wire \cpu.uart.r_ib[3] ;
 wire \cpu.uart.r_ib[4] ;
 wire \cpu.uart.r_ib[5] ;
 wire \cpu.uart.r_ib[6] ;
 wire \cpu.uart.r_in[0] ;
 wire \cpu.uart.r_in[1] ;
 wire \cpu.uart.r_in[2] ;
 wire \cpu.uart.r_in[3] ;
 wire \cpu.uart.r_in[4] ;
 wire \cpu.uart.r_in[5] ;
 wire \cpu.uart.r_in[6] ;
 wire \cpu.uart.r_in[7] ;
 wire \cpu.uart.r_out[0] ;
 wire \cpu.uart.r_out[1] ;
 wire \cpu.uart.r_out[2] ;
 wire \cpu.uart.r_out[3] ;
 wire \cpu.uart.r_out[4] ;
 wire \cpu.uart.r_out[5] ;
 wire \cpu.uart.r_out[6] ;
 wire \cpu.uart.r_out[7] ;
 wire \cpu.uart.r_r ;
 wire \cpu.uart.r_r_int ;
 wire \cpu.uart.r_r_invert ;
 wire \cpu.uart.r_rcnt[0] ;
 wire \cpu.uart.r_rcnt[1] ;
 wire \cpu.uart.r_rstate[0] ;
 wire \cpu.uart.r_rstate[1] ;
 wire \cpu.uart.r_rstate[2] ;
 wire \cpu.uart.r_rstate[3] ;
 wire \cpu.uart.r_x_int ;
 wire \cpu.uart.r_x_invert ;
 wire \cpu.uart.r_xcnt[0] ;
 wire \cpu.uart.r_xcnt[1] ;
 wire \cpu.uart.r_xstate[0] ;
 wire \cpu.uart.r_xstate[1] ;
 wire \cpu.uart.r_xstate[2] ;
 wire \cpu.uart.r_xstate[3] ;
 wire r_reset;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net2418;
 wire net2419;
 wire net2420;
 wire net2421;
 wire net2422;
 wire net2423;
 wire net2424;
 wire net2425;
 wire net2426;
 wire net2427;
 wire net2428;
 wire net2429;
 wire net2430;
 wire net2431;
 wire net2432;
 wire net2433;
 wire net2434;
 wire net2435;
 wire net2436;
 wire net2437;
 wire net2438;
 wire net2439;
 wire net2440;
 wire net2441;
 wire net2442;
 wire net2443;
 wire net2444;
 wire net2445;
 wire net2446;
 wire net2447;
 wire net2448;
 wire net2449;
 wire net2450;
 wire net2451;
 wire net2452;
 wire net2453;
 wire net2454;
 wire net2455;
 wire net2456;
 wire net2457;
 wire net2458;
 wire net2459;
 wire net2460;
 wire net2461;
 wire net2462;
 wire net2463;
 wire net2464;
 wire net2465;
 wire net2466;
 wire net2467;
 wire net2468;
 wire net2469;
 wire net2470;
 wire net2471;
 wire net2472;
 wire net2473;
 wire net2474;
 wire net2475;
 wire net2476;
 wire net2477;
 wire net2478;
 wire net2479;
 wire net2480;
 wire net2481;
 wire net2482;
 wire net2483;
 wire net2484;
 wire net2485;
 wire net2486;
 wire net2487;
 wire net2488;
 wire net2489;
 wire net2490;
 wire net2491;
 wire net2492;
 wire net2493;
 wire net2494;
 wire net2495;
 wire net2496;
 wire net2497;
 wire net2498;
 wire net2499;
 wire net2500;
 wire net2501;
 wire net2502;
 wire net2503;
 wire net2504;
 wire net2505;
 wire net2506;
 wire net2507;
 wire net2508;
 wire net2509;
 wire net2510;
 wire net2511;
 wire net2512;
 wire net2513;
 wire net2514;
 wire net2515;
 wire net2516;
 wire net2517;
 wire net2518;
 wire net2519;
 wire net2520;
 wire net2521;
 wire net2522;
 wire net2523;
 wire net2524;
 wire net2525;
 wire net2526;
 wire net2527;
 wire net2528;
 wire net2529;
 wire net2530;
 wire net2531;
 wire net2532;
 wire net2533;
 wire net2534;
 wire net2535;
 wire net2536;
 wire net2537;
 wire net2538;
 wire net2539;
 wire net2540;
 wire net2541;
 wire net2542;
 wire net2543;
 wire net2544;
 wire net2545;
 wire net2546;
 wire net2547;
 wire net2548;
 wire net2549;
 wire net2550;
 wire net2551;
 wire net2552;
 wire net2553;
 wire net2554;
 wire net2555;
 wire net2556;
 wire net2557;
 wire net2558;
 wire net2559;
 wire net2560;
 wire net2561;
 wire net2562;
 wire net2563;
 wire net2564;
 wire net2565;
 wire net2566;
 wire net2567;
 wire net2568;
 wire net2569;
 wire net2570;
 wire net2571;
 wire net2572;
 wire net2573;
 wire net2574;
 wire net2575;
 wire net2576;
 wire net2577;
 wire net2578;
 wire net2579;
 wire net2580;
 wire net2581;
 wire net2582;
 wire net2583;
 wire net2584;
 wire net2585;
 wire net2586;
 wire net2587;
 wire net2588;
 wire net2589;
 wire net2590;
 wire net2591;
 wire net2592;
 wire net2593;
 wire net2594;
 wire net2595;
 wire net2596;
 wire net2597;
 wire net2598;
 wire net2599;
 wire net2600;
 wire net2601;
 wire net2602;
 wire net2603;
 wire net2604;
 wire net2605;
 wire net2606;
 wire net2607;
 wire net2608;
 wire net2609;
 wire net2610;
 wire net2611;
 wire net2612;
 wire net2613;
 wire net2614;
 wire net2615;
 wire net2616;
 wire net2617;
 wire net2618;
 wire net2619;
 wire net2620;
 wire net2621;
 wire net2622;
 wire net2623;
 wire net2624;
 wire net2625;
 wire net2626;
 wire net2627;
 wire net2628;
 wire net2629;
 wire net2630;
 wire net2631;
 wire net2632;
 wire net2633;
 wire net2634;
 wire net2635;
 wire net2636;
 wire net2637;
 wire net2638;
 wire net2639;
 wire net2640;
 wire net2641;
 wire net2642;
 wire net2643;
 wire net2644;
 wire net2645;
 wire net2646;
 wire net2647;
 wire net2648;
 wire net2649;
 wire net2650;
 wire net2651;
 wire net2652;
 wire net2653;
 wire net2654;
 wire net2655;
 wire net2656;
 wire net2657;
 wire net2658;
 wire net2659;
 wire net2660;
 wire net2661;
 wire net2662;
 wire net2663;
 wire net2664;
 wire net2665;
 wire net2666;
 wire net2667;
 wire net2668;
 wire net2669;
 wire net2670;
 wire net2671;
 wire net2672;
 wire net2673;
 wire net2674;
 wire net2675;
 wire net2676;
 wire net2677;
 wire net2678;
 wire net2679;
 wire net2680;
 wire net2681;
 wire net2682;
 wire net2683;
 wire net2684;
 wire net2685;
 wire net2686;
 wire net2687;
 wire net2688;
 wire net2689;
 wire net2690;
 wire net2691;
 wire net2692;
 wire net2693;
 wire net2694;
 wire net2695;
 wire net2696;
 wire net2697;
 wire net2698;
 wire net2699;
 wire net2700;
 wire net2701;
 wire net2702;
 wire net2703;
 wire net2704;
 wire net2705;
 wire net2706;
 wire net2707;
 wire net2708;
 wire net2709;
 wire net2710;
 wire net2711;
 wire net2712;
 wire net2713;
 wire net2714;
 wire net2715;
 wire net2716;
 wire net2717;
 wire net2718;
 wire net2719;
 wire net2720;
 wire net2721;
 wire net2722;
 wire net2723;
 wire net2724;
 wire net2725;
 wire net2726;
 wire net2727;
 wire net2728;
 wire net2729;
 wire net2730;
 wire net2731;
 wire net2732;
 wire net2733;
 wire net2734;
 wire net2735;
 wire net2736;
 wire net2737;
 wire net2738;
 wire net2739;
 wire net2740;
 wire net2741;
 wire net2742;
 wire net2743;
 wire net2744;
 wire net2745;
 wire net2746;
 wire net2747;
 wire net2748;
 wire net2749;
 wire net2750;
 wire net2751;
 wire net2752;
 wire net2753;
 wire net2754;
 wire net2755;
 wire net2756;
 wire net2757;
 wire net2758;
 wire net2759;
 wire net2760;
 wire net2761;
 wire net2762;
 wire net2763;
 wire net2764;
 wire net2765;
 wire net2766;
 wire net2767;
 wire net2768;
 wire net2769;
 wire net2770;
 wire net2771;
 wire net2772;
 wire net2773;
 wire net2774;
 wire net2775;
 wire net2776;
 wire net2777;
 wire net2778;
 wire net2779;
 wire net2780;
 wire net2781;
 wire net2782;
 wire net2783;
 wire net2784;
 wire net2785;
 wire net2786;
 wire net2787;
 wire net2788;
 wire net2789;
 wire net2790;
 wire net2791;
 wire net2792;
 wire net2793;
 wire net2794;
 wire net2795;
 wire net2796;
 wire net2797;
 wire net2798;
 wire net2799;
 wire net2800;
 wire net2801;
 wire net2802;
 wire net2803;
 wire net2804;
 wire net2805;
 wire net2806;
 wire net2807;
 wire net2808;
 wire net2809;
 wire net2810;
 wire net2811;
 wire net2812;
 wire net2813;
 wire net2814;
 wire net2815;
 wire net2816;
 wire net2817;
 wire net2818;
 wire net2819;
 wire net2820;
 wire net2821;
 wire net2822;
 wire net2823;
 wire net2824;
 wire net2825;
 wire net2826;
 wire net2827;
 wire net2828;
 wire net2829;
 wire net2830;
 wire net2831;
 wire net2832;
 wire net2833;
 wire net2834;
 wire net2835;
 wire net2836;
 wire net2837;
 wire net2838;
 wire net2839;
 wire net2840;
 wire net2841;
 wire net2842;
 wire net2843;
 wire net2844;
 wire net2845;
 wire net2846;
 wire net2847;
 wire net2848;
 wire net2849;
 wire net2850;
 wire net2851;
 wire net2852;
 wire net2853;
 wire net2854;
 wire net2855;
 wire net2856;
 wire net2857;
 wire net2858;
 wire net2859;
 wire net2860;
 wire net2861;
 wire net2862;
 wire net2863;
 wire net2864;
 wire net2865;
 wire net2866;
 wire net2867;
 wire net2868;
 wire net2869;
 wire net2870;
 wire net2871;
 wire net2872;
 wire net2873;
 wire net2874;
 wire net2875;
 wire net2876;
 wire net2877;
 wire net2878;
 wire net2879;
 wire net2880;
 wire net2881;
 wire net2882;
 wire net2883;
 wire net2884;
 wire net2885;
 wire net2886;
 wire net2887;
 wire net2888;
 wire net2889;
 wire net2890;
 wire net2891;
 wire net2892;
 wire net2893;
 wire net2894;
 wire net2895;
 wire net2896;
 wire net2897;
 wire net2898;
 wire net2899;
 wire net2900;
 wire net2901;
 wire net2902;
 wire net2903;
 wire net2904;
 wire net2905;
 wire net2906;
 wire net2907;
 wire net2908;
 wire net2909;
 wire net2910;
 wire net2911;
 wire net2912;
 wire net2913;
 wire net2914;
 wire net2915;
 wire net2916;
 wire net2917;
 wire net2918;
 wire net2919;
 wire net2920;
 wire net2921;
 wire net2922;
 wire net2923;
 wire net2924;
 wire net2925;
 wire net2926;
 wire net2927;
 wire net2928;
 wire net2929;
 wire net2930;
 wire net2931;
 wire net2932;
 wire net2933;
 wire net2934;
 wire net2935;
 wire net2936;
 wire net2937;
 wire net2938;
 wire net2939;
 wire net2940;
 wire net2941;
 wire net2942;
 wire net2943;
 wire net2944;
 wire net2945;
 wire net2946;
 wire net2947;
 wire net2948;
 wire net2949;
 wire net2950;
 wire net2951;
 wire net2952;
 wire net2953;
 wire net2954;
 wire net2955;
 wire net2956;
 wire net2957;
 wire net2958;
 wire net2959;
 wire net2960;
 wire net2961;
 wire net2962;
 wire net2963;
 wire net2964;
 wire net2965;
 wire net2966;
 wire net2967;
 wire net2968;
 wire net2969;
 wire net2970;
 wire net2971;
 wire net2972;
 wire net2973;
 wire net2974;
 wire net2975;
 wire net2976;
 wire net2977;
 wire net2978;
 wire net2979;
 wire net2980;
 wire net2981;
 wire net2982;
 wire net2983;
 wire net2984;
 wire net2985;
 wire net2986;
 wire net2987;
 wire net2988;
 wire net2989;
 wire net2990;
 wire net2991;
 wire net2992;
 wire net2993;
 wire net2994;
 wire net2995;
 wire net2996;
 wire net2997;
 wire net2998;
 wire net2999;
 wire net3000;
 wire net3001;
 wire net3002;
 wire net3003;
 wire net3004;
 wire net3005;
 wire net3006;
 wire net3007;
 wire net3008;
 wire net3009;
 wire net3010;
 wire net3011;
 wire net3012;
 wire net3013;
 wire net3014;
 wire net3015;
 wire net3016;
 wire net3017;
 wire net3018;
 wire net3019;
 wire net3020;
 wire net3021;
 wire net3022;
 wire net3023;
 wire net3024;
 wire net3025;
 wire net3026;
 wire net3027;
 wire net3028;
 wire net3029;
 wire net3030;
 wire net3031;
 wire net3032;
 wire net3033;
 wire net3034;
 wire net3035;
 wire net3036;
 wire net3037;
 wire net3038;
 wire net3039;
 wire net3040;
 wire net3041;
 wire net3042;
 wire net3043;
 wire net3044;
 wire net3045;
 wire net3046;
 wire net3047;
 wire net3048;
 wire net3049;
 wire net3050;
 wire net3051;
 wire net3052;
 wire net3053;
 wire net3054;
 wire net3055;
 wire net3056;
 wire net3057;
 wire net3058;
 wire net3059;
 wire net3060;
 wire net3061;
 wire net3062;
 wire net3063;
 wire net3064;
 wire net3065;
 wire net3066;
 wire net3067;
 wire net3068;
 wire net3069;
 wire net3070;
 wire net3071;
 wire net3072;
 wire net3073;
 wire net3074;
 wire net3075;
 wire net3076;
 wire net3077;
 wire net3078;
 wire net3079;
 wire net3080;
 wire net3081;
 wire net3082;
 wire net3083;
 wire net3084;
 wire net3085;
 wire net3086;
 wire net3087;
 wire net3088;
 wire net3089;
 wire net3090;
 wire net3091;
 wire net3092;
 wire net3093;
 wire net3094;
 wire net3095;
 wire net3096;
 wire net3097;
 wire net3098;
 wire net3099;
 wire net3100;
 wire net3101;
 wire net3102;
 wire net3103;
 wire net3104;
 wire net3105;
 wire net3106;
 wire net3107;
 wire net3108;
 wire net3109;
 wire net3110;
 wire net3111;
 wire net3112;
 wire net3113;
 wire net3114;
 wire net3115;
 wire net3116;
 wire net3117;
 wire net3118;
 wire net3119;
 wire net3120;
 wire net3121;
 wire net3122;
 wire net3123;
 wire net3124;
 wire net3125;
 wire net3126;
 wire net3127;
 wire net3128;
 wire net3129;
 wire net3130;
 wire net3131;
 wire net3132;
 wire net3133;
 wire net3134;
 wire net3135;
 wire net3136;
 wire net3137;
 wire net3138;
 wire net3139;
 wire net3140;
 wire net3141;
 wire net3142;
 wire net3143;
 wire net3144;
 wire net3145;
 wire net3146;
 wire net3147;
 wire net3148;
 wire net3149;
 wire net3150;
 wire net3151;
 wire net3152;
 wire net3153;
 wire net3154;
 wire net3155;
 wire net3156;
 wire net3157;
 wire net3158;
 wire net3159;
 wire net3160;
 wire net3161;
 wire net3162;
 wire net3163;
 wire net3164;
 wire net3165;
 wire net3166;
 wire net3167;
 wire net3168;
 wire net3169;
 wire net3170;
 wire net3171;
 wire net3172;
 wire net3173;
 wire net3174;
 wire net3175;
 wire net3176;
 wire net3177;
 wire net3178;
 wire net3179;
 wire net3180;
 wire net3181;
 wire net3182;
 wire net3183;
 wire net3184;
 wire net3185;
 wire net3186;
 wire net3187;
 wire net3188;
 wire net3189;
 wire net3190;
 wire net3191;
 wire net3192;
 wire net3193;
 wire net3194;
 wire net3195;
 wire net3196;
 wire net3197;
 wire net3198;
 wire net3199;
 wire net3200;
 wire net3201;
 wire net3202;
 wire net3203;
 wire net3204;
 wire net3205;
 wire net3206;
 wire net3207;
 wire net3208;
 wire net3209;
 wire net3210;
 wire net3211;
 wire net3212;
 wire net3213;
 wire net3214;
 wire net3215;
 wire net3216;
 wire net3217;
 wire net3218;
 wire net3219;
 wire net3220;
 wire net3221;
 wire net3222;
 wire net3223;
 wire net3224;
 wire net3225;
 wire net3226;
 wire net3227;
 wire net3228;
 wire net3229;
 wire net3230;
 wire net3231;
 wire net3232;
 wire net3233;
 wire net3234;
 wire net3235;
 wire net3236;
 wire net3237;
 wire net3238;
 wire net3239;
 wire net3240;
 wire net3241;
 wire net3242;
 wire net3243;
 wire net3244;
 wire net3245;
 wire net3246;
 wire net3247;
 wire net3248;
 wire net3249;
 wire net3250;
 wire net3251;
 wire net3252;
 wire net3253;
 wire net3254;
 wire net3255;
 wire net3256;
 wire net3257;
 wire net3258;
 wire net3259;
 wire net3260;
 wire net3261;
 wire net3262;
 wire net3263;
 wire net3264;
 wire net3265;
 wire net3266;
 wire net3267;
 wire net3268;
 wire net3269;
 wire net3270;
 wire net3271;
 wire net3272;
 wire net3273;
 wire net3274;
 wire net3275;
 wire net3276;
 wire net3277;
 wire net3278;
 wire net3279;
 wire net3280;
 wire net3281;
 wire net3282;
 wire net3283;
 wire net3284;
 wire net3285;
 wire net3286;
 wire net3287;
 wire net3288;
 wire net3289;
 wire net3290;
 wire net3291;
 wire net3292;
 wire net3293;
 wire net3294;
 wire net3295;
 wire net3296;
 wire net3297;
 wire net3298;
 wire net3299;
 wire net3300;
 wire net3301;
 wire net3302;
 wire net3303;
 wire net3304;
 wire net3305;
 wire net3306;
 wire net3307;
 wire net3308;
 wire net3309;
 wire net3310;
 wire net3311;
 wire net3312;
 wire net3313;
 wire net3314;
 wire net3315;
 wire net3316;
 wire net3317;
 wire net3318;
 wire net3319;
 wire net3320;
 wire net3321;
 wire net3322;
 wire net3323;
 wire net3324;
 wire net3325;
 wire net3326;
 wire net3327;
 wire net3328;
 wire net3329;
 wire net3330;
 wire net3331;
 wire net3332;
 wire net3333;
 wire net3334;
 wire net3335;
 wire net3336;
 wire net3337;
 wire net3338;
 wire net3339;
 wire net3340;
 wire net3341;
 wire net3342;
 wire net3343;
 wire net3344;
 wire net3345;
 wire net3346;
 wire net3347;
 wire net3348;
 wire net3349;
 wire net3350;
 wire net3351;
 wire net3352;
 wire net3353;
 wire net3354;
 wire net3355;
 wire net3356;
 wire net3357;
 wire net3358;
 wire net3359;
 wire net3360;
 wire net3361;
 wire net3362;
 wire net3363;
 wire net3364;
 wire net3365;
 wire net3366;
 wire net3367;
 wire net3368;
 wire net3369;
 wire net3370;
 wire net3371;
 wire net3372;
 wire net3373;
 wire net3374;
 wire net3375;
 wire net3376;
 wire net3377;
 wire net3378;
 wire net3379;
 wire net3380;
 wire net3381;
 wire net3382;
 wire net3383;
 wire net3384;
 wire net3385;
 wire net3386;
 wire net3387;
 wire net3388;
 wire net3389;
 wire net3390;
 wire net3391;
 wire net3392;
 wire net3393;
 wire net3394;
 wire net3395;
 wire net3396;
 wire net3397;
 wire net3398;
 wire net3399;
 wire net3400;
 wire net3401;
 wire net3402;
 wire net3403;
 wire net3404;
 wire net3405;
 wire net3406;
 wire net3407;
 wire net3408;
 wire net3409;
 wire net3410;
 wire net3411;
 wire net3412;
 wire net3413;
 wire net3414;
 wire net3415;
 wire net3416;
 wire net3417;
 wire net3418;
 wire net3419;
 wire net3420;
 wire net3421;
 wire net3422;
 wire net3423;
 wire net3424;
 wire net3425;
 wire net3426;
 wire net3427;
 wire net3428;
 wire net3429;
 wire net3430;
 wire net3431;
 wire net3432;
 wire net3433;
 wire net3434;
 wire net3435;
 wire net3436;
 wire net3437;
 wire net3438;
 wire net3439;
 wire net3440;
 wire net3441;
 wire net3442;
 wire net3443;
 wire net3444;
 wire net3445;
 wire net3446;
 wire net3447;
 wire net3448;
 wire net3449;
 wire net3450;
 wire net3451;
 wire net3452;
 wire net3453;
 wire net3454;
 wire net3455;
 wire net3456;
 wire net3457;
 wire net3458;
 wire net3459;
 wire net3460;
 wire net3461;
 wire net3462;
 wire net3463;
 wire net3464;
 wire net3465;
 wire net3466;
 wire net3467;
 wire net3468;
 wire net3469;
 wire net3470;
 wire net3471;
 wire net3472;
 wire net3473;
 wire net3474;
 wire net3475;
 wire net3476;
 wire net3477;
 wire net3478;
 wire net3479;
 wire net3480;
 wire net3481;
 wire net3482;
 wire net3483;
 wire net3484;
 wire net3485;
 wire net3486;
 wire net3487;
 wire net3488;
 wire net3489;
 wire net3490;
 wire net3491;
 wire net3492;
 wire net3493;
 wire net3494;
 wire net3495;
 wire net3496;
 wire net3497;
 wire net3498;
 wire net3499;
 wire net3500;
 wire net3501;
 wire net3502;
 wire net3503;
 wire net3504;
 wire net3505;
 wire net3506;
 wire net3507;
 wire net3508;
 wire net3509;
 wire net3510;
 wire net3511;
 wire net3512;
 wire net3513;
 wire net3514;
 wire net3515;
 wire net3516;
 wire net3517;
 wire net3518;
 wire net3519;
 wire net3520;
 wire net3521;
 wire net3522;
 wire net3523;
 wire net3524;
 wire net3525;
 wire net3526;
 wire net3527;
 wire net3528;
 wire net3529;
 wire net3530;
 wire net3531;
 wire net3532;
 wire net3533;
 wire net3534;
 wire net3535;
 wire net3536;
 wire net3537;
 wire net3538;
 wire net3539;
 wire net3540;
 wire net3541;
 wire net3542;
 wire net3543;
 wire net3544;
 wire net3545;
 wire net3546;
 wire net3547;
 wire net3548;
 wire net3549;
 wire net3550;
 wire net3551;
 wire net3552;
 wire net3553;
 wire net3554;
 wire net3555;
 wire net3556;
 wire net3557;
 wire net3558;
 wire net3559;
 wire net3560;
 wire net3561;
 wire net3562;
 wire net3563;
 wire net3564;
 wire net3565;
 wire net3566;
 wire net3567;
 wire net3568;
 wire net3569;
 wire net3570;
 wire net3571;
 wire net3572;
 wire net3573;
 wire net3574;
 wire net3575;
 wire net3576;
 wire net3577;
 wire net3578;
 wire net3579;
 wire net3580;
 wire net3581;
 wire net3582;
 wire net3583;
 wire net3584;
 wire net3585;
 wire net3586;
 wire net3587;
 wire net3588;
 wire net3589;
 wire net3590;
 wire net3591;
 wire net3592;
 wire net3593;
 wire net3594;
 wire net3595;
 wire net3596;
 wire net3597;
 wire net3598;
 wire net3599;
 wire net3600;
 wire net3601;
 wire net3602;
 wire net3603;
 wire net3604;
 wire net3605;
 wire net3606;
 wire net3607;
 wire net3608;
 wire net3609;
 wire net3610;
 wire net3611;
 wire net3612;
 wire net3613;
 wire net3614;
 wire net3615;
 wire net3616;
 wire net3617;
 wire net3618;
 wire net3619;
 wire net3620;
 wire net3621;
 wire net3622;
 wire net3623;
 wire net3624;
 wire net3625;
 wire net3626;
 wire net3627;
 wire net3628;
 wire net3629;
 wire net3630;
 wire net3631;
 wire net3632;
 wire net3633;
 wire net3634;
 wire net3635;
 wire net3636;
 wire net3637;
 wire net3638;
 wire net3639;
 wire net3640;
 wire net3641;
 wire net3642;
 wire net3643;
 wire net3644;
 wire net3645;
 wire net3646;
 wire net3647;
 wire net3648;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_2 _15019_ (.A(\cpu.dec.r_op[6] ),
    .X(_08242_));
 sg13g2_buf_1 _15020_ (.A(_08242_),
    .X(_08243_));
 sg13g2_buf_1 _15021_ (.A(net1091),
    .X(_08244_));
 sg13g2_buf_1 _15022_ (.A(_00187_),
    .X(_08245_));
 sg13g2_buf_8 _15023_ (.A(\cpu.addr[13] ),
    .X(_08246_));
 sg13g2_buf_8 _15024_ (.A(\cpu.addr[15] ),
    .X(_08247_));
 sg13g2_nor2b_1 _15025_ (.A(_08246_),
    .B_N(_08247_),
    .Y(_08248_));
 sg13g2_buf_16 _15026_ (.X(_08249_),
    .A(\cpu.addr[12] ));
 sg13g2_buf_8 _15027_ (.A(\cpu.addr[14] ),
    .X(_08250_));
 sg13g2_buf_8 _15028_ (.A(_08250_),
    .X(_08251_));
 sg13g2_mux4_1 _15029_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .S1(net1090),
    .X(_08252_));
 sg13g2_and2_1 _15030_ (.A(_08248_),
    .B(_08252_),
    .X(_08253_));
 sg13g2_buf_8 _15031_ (.A(_08250_),
    .X(_08254_));
 sg13g2_nand2_1 _15032_ (.Y(_08255_),
    .A(_08254_),
    .B(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_nand2b_1 _15033_ (.Y(_08256_),
    .B(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A_N(_08251_));
 sg13g2_buf_8 _15034_ (.A(_08249_),
    .X(_08257_));
 sg13g2_nand3b_1 _15035_ (.B(_08246_),
    .C(_08247_),
    .Y(_08258_),
    .A_N(net1088));
 sg13g2_a21oi_1 _15036_ (.A1(_08255_),
    .A2(_08256_),
    .Y(_08259_),
    .B1(_08258_));
 sg13g2_buf_8 _15037_ (.A(_08246_),
    .X(_08260_));
 sg13g2_and2_1 _15038_ (.A(_08249_),
    .B(_08247_),
    .X(_08261_));
 sg13g2_buf_1 _15039_ (.A(_08261_),
    .X(_08262_));
 sg13g2_mux2_1 _15040_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .S(net1090),
    .X(_08263_));
 sg13g2_and3_1 _15041_ (.X(_08264_),
    .A(_08260_),
    .B(_08262_),
    .C(_08263_));
 sg13g2_buf_2 _15042_ (.A(_00191_),
    .X(_08265_));
 sg13g2_inv_1 _15043_ (.Y(_08266_),
    .A(_08265_));
 sg13g2_buf_2 _15044_ (.A(\cpu.ex.r_wmask[1] ),
    .X(_08267_));
 sg13g2_buf_8 _15045_ (.A(\cpu.ex.r_wmask[0] ),
    .X(_08268_));
 sg13g2_or2_1 _15046_ (.X(_08269_),
    .B(_08268_),
    .A(_08267_));
 sg13g2_buf_1 _15047_ (.A(\cpu.ex.io_access ),
    .X(_08270_));
 sg13g2_buf_8 _15048_ (.A(\cpu.ex.genblk3.r_mmu_enable ),
    .X(_08271_));
 sg13g2_nor2b_1 _15049_ (.A(net1166),
    .B_N(net1165),
    .Y(_08272_));
 sg13g2_buf_8 _15050_ (.A(\cpu.ex.ifetch ),
    .X(_08273_));
 sg13g2_buf_2 _15051_ (.A(\cpu.ex.genblk3.r_mmu_d_proxy ),
    .X(_08274_));
 sg13g2_nand2b_1 _15052_ (.Y(_08275_),
    .B(_08274_),
    .A_N(net1164));
 sg13g2_nand4_1 _15053_ (.B(_08269_),
    .C(_08272_),
    .A(_08266_),
    .Y(_08276_),
    .D(_08275_));
 sg13g2_nor4_1 _15054_ (.A(_08253_),
    .B(_08259_),
    .C(_08264_),
    .D(_08276_),
    .Y(_08277_));
 sg13g2_buf_1 _15055_ (.A(_08247_),
    .X(_08278_));
 sg13g2_mux4_1 _15056_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .S1(net1090),
    .X(_08279_));
 sg13g2_mux4_1 _15057_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .S1(net1090),
    .X(_08280_));
 sg13g2_mux2_1 _15058_ (.A0(_08279_),
    .A1(_08280_),
    .S(net1087),
    .X(_08281_));
 sg13g2_nand2b_1 _15059_ (.Y(_08282_),
    .B(_08281_),
    .A_N(net1086));
 sg13g2_mux4_1 _15060_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .S1(net1090),
    .X(_08283_));
 sg13g2_nand2_1 _15061_ (.Y(_08284_),
    .A(_08248_),
    .B(_08283_));
 sg13g2_mux2_1 _15062_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .S(net1090),
    .X(_08285_));
 sg13g2_nand2b_1 _15063_ (.Y(_08286_),
    .B(_08285_),
    .A_N(_08258_));
 sg13g2_mux2_1 _15064_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .S(net1090),
    .X(_08287_));
 sg13g2_nand3_1 _15065_ (.B(_08262_),
    .C(_08287_),
    .A(net1087),
    .Y(_08288_));
 sg13g2_inv_1 _15066_ (.Y(_08289_),
    .A(_08267_));
 sg13g2_inv_1 _15067_ (.Y(_08290_),
    .A(_08268_));
 sg13g2_nand2b_1 _15068_ (.Y(_08291_),
    .B(net1165),
    .A_N(net1166));
 sg13g2_a221oi_1 _15069_ (.B2(_08275_),
    .C1(_08291_),
    .B1(_08266_),
    .A1(_08289_),
    .Y(_08292_),
    .A2(_08290_));
 sg13g2_and4_1 _15070_ (.A(_08284_),
    .B(_08286_),
    .C(_08288_),
    .D(_08292_),
    .X(_08293_));
 sg13g2_mux4_1 _15071_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .S1(_08251_),
    .X(_08294_));
 sg13g2_mux4_1 _15072_ (.S0(_08249_),
    .A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A2(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A3(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .S1(net1090),
    .X(_08295_));
 sg13g2_mux2_1 _15073_ (.A0(_08294_),
    .A1(_08295_),
    .S(_08260_),
    .X(_08296_));
 sg13g2_nand2b_1 _15074_ (.Y(_08297_),
    .B(_08296_),
    .A_N(net1086));
 sg13g2_a22oi_1 _15075_ (.Y(_08298_),
    .B1(_08293_),
    .B2(_08297_),
    .A2(_08282_),
    .A1(_08277_));
 sg13g2_buf_8 _15076_ (.A(_08298_),
    .X(_08299_));
 sg13g2_buf_8 _15077_ (.A(_08299_),
    .X(_08300_));
 sg13g2_buf_8 _15078_ (.A(\cpu.dec.supmode ),
    .X(_08301_));
 sg13g2_buf_1 _15079_ (.A(\cpu.ex.pc[15] ),
    .X(_08302_));
 sg13g2_nor2b_1 _15080_ (.A(net1163),
    .B_N(_08302_),
    .Y(_08303_));
 sg13g2_buf_8 _15081_ (.A(\cpu.ex.pc[14] ),
    .X(_08304_));
 sg13g2_mux2_1 _15082_ (.A0(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[12] ),
    .S(_08304_),
    .X(_08305_));
 sg13g2_mux2_1 _15083_ (.A0(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[13] ),
    .S(_08304_),
    .X(_08306_));
 sg13g2_mux2_1 _15084_ (.A0(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[14] ),
    .S(_08304_),
    .X(_08307_));
 sg13g2_mux2_1 _15085_ (.A0(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[15] ),
    .S(_08304_),
    .X(_08308_));
 sg13g2_buf_8 _15086_ (.A(\cpu.ex.pc[12] ),
    .X(_08309_));
 sg13g2_buf_8 _15087_ (.A(\cpu.ex.pc[13] ),
    .X(_08310_));
 sg13g2_buf_1 _15088_ (.A(_08310_),
    .X(_08311_));
 sg13g2_mux4_1 _15089_ (.S0(_08309_),
    .A0(_08305_),
    .A1(_08306_),
    .A2(_08307_),
    .A3(_08308_),
    .S1(net1085),
    .X(_08312_));
 sg13g2_buf_2 _15090_ (.A(_08302_),
    .X(_08313_));
 sg13g2_and2_1 _15091_ (.A(_08313_),
    .B(net1163),
    .X(_08314_));
 sg13g2_buf_8 _15092_ (.A(_08304_),
    .X(_08315_));
 sg13g2_mux2_1 _15093_ (.A0(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[28] ),
    .S(net1083),
    .X(_08316_));
 sg13g2_mux2_1 _15094_ (.A0(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[29] ),
    .S(net1083),
    .X(_08317_));
 sg13g2_mux2_1 _15095_ (.A0(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[30] ),
    .S(_08304_),
    .X(_08318_));
 sg13g2_mux2_1 _15096_ (.A0(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[31] ),
    .S(net1083),
    .X(_08319_));
 sg13g2_mux4_1 _15097_ (.S0(_08309_),
    .A0(_08316_),
    .A1(_08317_),
    .A2(_08318_),
    .A3(_08319_),
    .S1(net1085),
    .X(_08320_));
 sg13g2_a22oi_1 _15098_ (.Y(_08321_),
    .B1(_08314_),
    .B2(_08320_),
    .A2(_08312_),
    .A1(_08303_));
 sg13g2_nand2b_1 _15099_ (.Y(_08322_),
    .B(_08310_),
    .A_N(_08309_));
 sg13g2_mux2_1 _15100_ (.A0(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[6] ),
    .S(net1083),
    .X(_08323_));
 sg13g2_nor2_1 _15101_ (.A(_08322_),
    .B(_08323_),
    .Y(_08324_));
 sg13g2_nand2b_1 _15102_ (.Y(_08325_),
    .B(_08309_),
    .A_N(_08310_));
 sg13g2_mux2_1 _15103_ (.A0(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[5] ),
    .S(_08304_),
    .X(_08326_));
 sg13g2_nor2_1 _15104_ (.A(_08302_),
    .B(net1163),
    .Y(_08327_));
 sg13g2_o21ai_1 _15105_ (.B1(_08327_),
    .Y(_08328_),
    .A1(_08325_),
    .A2(_08326_));
 sg13g2_nand2_1 _15106_ (.Y(_08329_),
    .A(_08309_),
    .B(_08310_));
 sg13g2_mux2_1 _15107_ (.A0(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[7] ),
    .S(_08315_),
    .X(_08330_));
 sg13g2_nor2_1 _15108_ (.A(_08329_),
    .B(_08330_),
    .Y(_08331_));
 sg13g2_buf_1 _15109_ (.A(_08309_),
    .X(_08332_));
 sg13g2_mux2_1 _15110_ (.A0(\cpu.genblk1.mmu.r_valid_i[0] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[4] ),
    .S(net1083),
    .X(_08333_));
 sg13g2_nor3_1 _15111_ (.A(_08332_),
    .B(_08311_),
    .C(_08333_),
    .Y(_08334_));
 sg13g2_or4_1 _15112_ (.A(_08324_),
    .B(_08328_),
    .C(_08331_),
    .D(_08334_),
    .X(_08335_));
 sg13g2_inv_2 _15113_ (.Y(_08336_),
    .A(net1165));
 sg13g2_inv_2 _15114_ (.Y(_08337_),
    .A(_08273_));
 sg13g2_buf_8 _15115_ (.A(_08337_),
    .X(_08338_));
 sg13g2_nor2_1 _15116_ (.A(_08336_),
    .B(_08338_),
    .Y(_08339_));
 sg13g2_mux2_1 _15117_ (.A0(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[22] ),
    .S(net1083),
    .X(_08340_));
 sg13g2_nor2_1 _15118_ (.A(_08322_),
    .B(_08340_),
    .Y(_08341_));
 sg13g2_mux2_1 _15119_ (.A0(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[21] ),
    .S(_08304_),
    .X(_08342_));
 sg13g2_nor2b_1 _15120_ (.A(_08302_),
    .B_N(net1163),
    .Y(_08343_));
 sg13g2_o21ai_1 _15121_ (.B1(_08343_),
    .Y(_08344_),
    .A1(_08325_),
    .A2(_08342_));
 sg13g2_mux2_1 _15122_ (.A0(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[23] ),
    .S(net1083),
    .X(_08345_));
 sg13g2_nor2_1 _15123_ (.A(_08329_),
    .B(_08345_),
    .Y(_08346_));
 sg13g2_mux2_1 _15124_ (.A0(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A1(\cpu.genblk1.mmu.r_valid_i[20] ),
    .S(net1083),
    .X(_08347_));
 sg13g2_nor3_1 _15125_ (.A(_08332_),
    .B(_08311_),
    .C(_08347_),
    .Y(_08348_));
 sg13g2_or4_1 _15126_ (.A(_08341_),
    .B(_08344_),
    .C(_08346_),
    .D(_08348_),
    .X(_08349_));
 sg13g2_nand4_1 _15127_ (.B(_08335_),
    .C(_08339_),
    .A(_08321_),
    .Y(_08350_),
    .D(_08349_));
 sg13g2_buf_8 _15128_ (.A(_08350_),
    .X(_08351_));
 sg13g2_buf_1 _15129_ (.A(\cpu.ex.r_read_stall ),
    .X(_08352_));
 sg13g2_inv_1 _15130_ (.Y(_08353_),
    .A(_08352_));
 sg13g2_nor2_1 _15131_ (.A(_08267_),
    .B(_08268_),
    .Y(_08354_));
 sg13g2_buf_2 _15132_ (.A(_08354_),
    .X(_08355_));
 sg13g2_nand3_1 _15133_ (.B(_08353_),
    .C(_08355_),
    .A(_08245_),
    .Y(_08356_));
 sg13g2_buf_1 _15134_ (.A(_08356_),
    .X(_08357_));
 sg13g2_nor2b_1 _15135_ (.A(_08351_),
    .B_N(_08357_),
    .Y(_08358_));
 sg13g2_buf_8 _15136_ (.A(_08358_),
    .X(_08359_));
 sg13g2_buf_8 _15137_ (.A(net1087),
    .X(_08360_));
 sg13g2_a21oi_1 _15138_ (.A1(_08338_),
    .A2(_08274_),
    .Y(_08361_),
    .B1(_08265_));
 sg13g2_mux4_1 _15139_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[23] ),
    .S1(net1089),
    .X(_08362_));
 sg13g2_mux4_1 _15140_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[31] ),
    .S1(net1089),
    .X(_08363_));
 sg13g2_mux2_1 _15141_ (.A0(_08362_),
    .A1(_08363_),
    .S(_08247_),
    .X(_08364_));
 sg13g2_nand3_1 _15142_ (.B(_08361_),
    .C(_08364_),
    .A(net949),
    .Y(_08365_));
 sg13g2_buf_8 _15143_ (.A(net1089),
    .X(_08366_));
 sg13g2_nand2_1 _15144_ (.Y(_08367_),
    .A(_08266_),
    .B(_08275_));
 sg13g2_buf_8 _15145_ (.A(_08367_),
    .X(_08368_));
 sg13g2_mux4_1 _15146_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[7] ),
    .S1(_08246_),
    .X(_08369_));
 sg13g2_mux4_1 _15147_ (.S0(net1088),
    .A0(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A3(\cpu.genblk1.mmu.r_valid_d[15] ),
    .S1(_08246_),
    .X(_08370_));
 sg13g2_mux2_1 _15148_ (.A0(_08369_),
    .A1(_08370_),
    .S(_08247_),
    .X(_08371_));
 sg13g2_nand3_1 _15149_ (.B(_08368_),
    .C(_08371_),
    .A(net948),
    .Y(_08372_));
 sg13g2_and2_1 _15150_ (.A(_08365_),
    .B(_08372_),
    .X(_08373_));
 sg13g2_buf_1 _15151_ (.A(\cpu.cond[0] ),
    .X(_08374_));
 sg13g2_inv_2 _15152_ (.Y(_08375_),
    .A(_08374_));
 sg13g2_buf_1 _15153_ (.A(\cpu.ex.mmu_reg_data[0] ),
    .X(_08376_));
 sg13g2_buf_1 _15154_ (.A(_00196_),
    .X(_08377_));
 sg13g2_buf_8 _15155_ (.A(_08352_),
    .X(_08378_));
 sg13g2_nand2_1 _15156_ (.Y(_08379_),
    .A(net1162),
    .B(net1081));
 sg13g2_o21ai_1 _15157_ (.B1(_08379_),
    .Y(_08380_),
    .A1(net1162),
    .A2(net1161));
 sg13g2_nand2_1 _15158_ (.Y(_08381_),
    .A(net1161),
    .B(_08353_));
 sg13g2_o21ai_1 _15159_ (.B1(_08381_),
    .Y(_08382_),
    .A1(_08375_),
    .A2(_08380_));
 sg13g2_buf_2 _15160_ (.A(_08382_),
    .X(_08383_));
 sg13g2_nand3_1 _15161_ (.B(_00195_),
    .C(_08357_),
    .A(net1165),
    .Y(_08384_));
 sg13g2_nand2_1 _15162_ (.Y(_08385_),
    .A(_08269_),
    .B(_08272_));
 sg13g2_o21ai_1 _15163_ (.B1(_08385_),
    .Y(_08386_),
    .A1(_08383_),
    .A2(_08384_));
 sg13g2_nor2_1 _15164_ (.A(net1088),
    .B(net1086),
    .Y(_08387_));
 sg13g2_nand2b_1 _15165_ (.Y(_08388_),
    .B(\cpu.genblk1.mmu.r_valid_d[0] ),
    .A_N(net1087));
 sg13g2_nand2_1 _15166_ (.Y(_08389_),
    .A(\cpu.genblk1.mmu.r_valid_d[2] ),
    .B(net1087));
 sg13g2_nand3_1 _15167_ (.B(_08388_),
    .C(_08389_),
    .A(_08387_),
    .Y(_08390_));
 sg13g2_nand2b_1 _15168_ (.Y(_08391_),
    .B(_08246_),
    .A_N(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_o21ai_1 _15169_ (.B1(_08391_),
    .Y(_08392_),
    .A1(net1087),
    .A2(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_nor2b_1 _15170_ (.A(_08247_),
    .B_N(net1088),
    .Y(_08393_));
 sg13g2_nand2b_1 _15171_ (.Y(_08394_),
    .B(net1087),
    .A_N(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_o21ai_1 _15172_ (.B1(_08394_),
    .Y(_08395_),
    .A1(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(net1087));
 sg13g2_a22oi_1 _15173_ (.Y(_08396_),
    .B1(_08393_),
    .B2(_08395_),
    .A2(_08392_),
    .A1(_08262_));
 sg13g2_nand2b_1 _15174_ (.Y(_08397_),
    .B(_08247_),
    .A_N(net1088));
 sg13g2_mux2_1 _15175_ (.A0(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[10] ),
    .S(_08246_),
    .X(_08398_));
 sg13g2_nor2_1 _15176_ (.A(_08397_),
    .B(_08398_),
    .Y(_08399_));
 sg13g2_nor3_1 _15177_ (.A(net948),
    .B(_08361_),
    .C(_08399_),
    .Y(_08400_));
 sg13g2_nand3_1 _15178_ (.B(_08396_),
    .C(_08400_),
    .A(_08390_),
    .Y(_08401_));
 sg13g2_nand2b_1 _15179_ (.Y(_08402_),
    .B(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A_N(net1089));
 sg13g2_nand2_1 _15180_ (.Y(_08403_),
    .A(net948),
    .B(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_nand3_1 _15181_ (.B(_08402_),
    .C(_08403_),
    .A(_08387_),
    .Y(_08404_));
 sg13g2_nand2b_1 _15182_ (.Y(_08405_),
    .B(net1089),
    .A_N(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_o21ai_1 _15183_ (.B1(_08405_),
    .Y(_08406_),
    .A1(net1089),
    .A2(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_nand2b_1 _15184_ (.Y(_08407_),
    .B(net1089),
    .A_N(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_o21ai_1 _15185_ (.B1(_08407_),
    .Y(_08408_),
    .A1(_08254_),
    .A2(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_a22oi_1 _15186_ (.Y(_08409_),
    .B1(_08408_),
    .B2(_08393_),
    .A2(_08406_),
    .A1(_08262_));
 sg13g2_mux2_1 _15187_ (.A0(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A1(\cpu.genblk1.mmu.r_valid_d[28] ),
    .S(net1089),
    .X(_08410_));
 sg13g2_nor2_1 _15188_ (.A(_08397_),
    .B(_08410_),
    .Y(_08411_));
 sg13g2_nor3_1 _15189_ (.A(net949),
    .B(_08368_),
    .C(_08411_),
    .Y(_08412_));
 sg13g2_nand3_1 _15190_ (.B(_08409_),
    .C(_08412_),
    .A(_08404_),
    .Y(_08413_));
 sg13g2_and4_1 _15191_ (.A(_08373_),
    .B(_08386_),
    .C(_08401_),
    .D(_08413_),
    .X(_08414_));
 sg13g2_buf_2 _15192_ (.A(_08414_),
    .X(_08415_));
 sg13g2_nor2_1 _15193_ (.A(_08359_),
    .B(_08415_),
    .Y(_08416_));
 sg13g2_buf_1 _15194_ (.A(_08416_),
    .X(_08417_));
 sg13g2_nand2_1 _15195_ (.Y(_08418_),
    .A(net498),
    .B(net358));
 sg13g2_buf_2 _15196_ (.A(_08418_),
    .X(_08419_));
 sg13g2_nor2_1 _15197_ (.A(_08245_),
    .B(_08419_),
    .Y(_08420_));
 sg13g2_buf_1 _15198_ (.A(net1085),
    .X(_08421_));
 sg13g2_buf_1 _15199_ (.A(net947),
    .X(_08422_));
 sg13g2_buf_2 _15200_ (.A(_08422_),
    .X(_08423_));
 sg13g2_buf_1 _15201_ (.A(_08271_),
    .X(_08424_));
 sg13g2_buf_4 _15202_ (.X(_08425_),
    .A(net1082));
 sg13g2_buf_2 _15203_ (.A(_08425_),
    .X(_08426_));
 sg13g2_buf_1 _15204_ (.A(net947),
    .X(_08427_));
 sg13g2_mux4_1 _15205_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .S1(net836),
    .X(_08428_));
 sg13g2_mux4_1 _15206_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .S1(net836),
    .X(_08429_));
 sg13g2_buf_2 _15207_ (.A(_08425_),
    .X(_08430_));
 sg13g2_buf_1 _15208_ (.A(net947),
    .X(_08431_));
 sg13g2_mux4_1 _15209_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .S1(net834),
    .X(_08432_));
 sg13g2_mux4_1 _15210_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .S1(net834),
    .X(_08433_));
 sg13g2_buf_2 _15211_ (.A(_08315_),
    .X(_08434_));
 sg13g2_mux4_1 _15212_ (.S0(net946),
    .A0(_08428_),
    .A1(_08429_),
    .A2(_08432_),
    .A3(_08433_),
    .S1(net1084),
    .X(_08435_));
 sg13g2_nand2_1 _15213_ (.Y(_08436_),
    .A(net1163),
    .B(_08435_));
 sg13g2_inv_1 _15214_ (.Y(_08437_),
    .A(net1163));
 sg13g2_buf_1 _15215_ (.A(_08437_),
    .X(_08438_));
 sg13g2_mux4_1 _15216_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .S1(net836),
    .X(_08439_));
 sg13g2_mux4_1 _15217_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .S1(net836),
    .X(_08440_));
 sg13g2_mux4_1 _15218_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .S1(net834),
    .X(_08441_));
 sg13g2_mux4_1 _15219_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .S1(net834),
    .X(_08442_));
 sg13g2_mux4_1 _15220_ (.S0(net946),
    .A0(_08439_),
    .A1(_08440_),
    .A2(_08441_),
    .A3(_08442_),
    .S1(net1084),
    .X(_08443_));
 sg13g2_nand2_1 _15221_ (.Y(_08444_),
    .A(net945),
    .B(_08443_));
 sg13g2_nand3_1 _15222_ (.B(_08436_),
    .C(_08444_),
    .A(net1080),
    .Y(_08445_));
 sg13g2_o21ai_1 _15223_ (.B1(_08445_),
    .Y(_08446_),
    .A1(net735),
    .A2(net1080));
 sg13g2_buf_1 _15224_ (.A(_08446_),
    .X(_08447_));
 sg13g2_buf_2 _15225_ (.A(_00188_),
    .X(_08448_));
 sg13g2_buf_1 _15226_ (.A(_08448_),
    .X(_08449_));
 sg13g2_buf_1 _15227_ (.A(\cpu.ex.pc[2] ),
    .X(_08450_));
 sg13g2_buf_2 _15228_ (.A(\cpu.ex.pc[4] ),
    .X(_08451_));
 sg13g2_buf_1 _15229_ (.A(\cpu.ex.pc[3] ),
    .X(_08452_));
 sg13g2_nor2b_1 _15230_ (.A(net1159),
    .B_N(net1158),
    .Y(_08453_));
 sg13g2_nand2b_1 _15231_ (.Y(_08454_),
    .B(net1159),
    .A_N(net1158));
 sg13g2_o21ai_1 _15232_ (.B1(_08454_),
    .Y(_08455_),
    .A1(net1160),
    .A2(_08453_));
 sg13g2_nand2_1 _15233_ (.Y(_08456_),
    .A(net1079),
    .B(_08455_));
 sg13g2_buf_1 _15234_ (.A(_08456_),
    .X(_08457_));
 sg13g2_buf_1 _15235_ (.A(net734),
    .X(_08458_));
 sg13g2_buf_1 _15236_ (.A(_08458_),
    .X(_08459_));
 sg13g2_buf_1 _15237_ (.A(net734),
    .X(_08460_));
 sg13g2_buf_1 _15238_ (.A(_08460_),
    .X(_08461_));
 sg13g2_buf_1 _15239_ (.A(net1158),
    .X(_08462_));
 sg13g2_buf_2 _15240_ (.A(net1078),
    .X(_08463_));
 sg13g2_buf_1 _15241_ (.A(_08463_),
    .X(_08464_));
 sg13g2_buf_2 _15242_ (.A(net1079),
    .X(_08465_));
 sg13g2_mux2_1 _15243_ (.A0(\cpu.icache.r_tag[7][13] ),
    .A1(\cpu.icache.r_tag[3][13] ),
    .S(net943),
    .X(_08466_));
 sg13g2_nor2_1 _15244_ (.A(net1078),
    .B(_08449_),
    .Y(_08467_));
 sg13g2_buf_1 _15245_ (.A(_08467_),
    .X(_08468_));
 sg13g2_a22oi_1 _15246_ (.Y(_08469_),
    .B1(net832),
    .B2(\cpu.icache.r_tag[5][13] ),
    .A2(_08466_),
    .A1(net833));
 sg13g2_buf_2 _15247_ (.A(net1160),
    .X(_08470_));
 sg13g2_buf_2 _15248_ (.A(net1077),
    .X(_08471_));
 sg13g2_buf_1 _15249_ (.A(net942),
    .X(_08472_));
 sg13g2_nand2b_1 _15250_ (.Y(_08473_),
    .B(net831),
    .A_N(_08469_));
 sg13g2_inv_1 _15251_ (.Y(_08474_),
    .A(net1160));
 sg13g2_buf_2 _15252_ (.A(_08474_),
    .X(_08475_));
 sg13g2_nor3_1 _15253_ (.A(net941),
    .B(net1158),
    .C(net1159),
    .Y(_08476_));
 sg13g2_buf_2 _15254_ (.A(_08476_),
    .X(_08477_));
 sg13g2_buf_1 _15255_ (.A(_08477_),
    .X(_08478_));
 sg13g2_buf_1 _15256_ (.A(net657),
    .X(_08479_));
 sg13g2_nor2_1 _15257_ (.A(net1160),
    .B(_08448_),
    .Y(_08480_));
 sg13g2_buf_1 _15258_ (.A(_08480_),
    .X(_08481_));
 sg13g2_buf_1 _15259_ (.A(net940),
    .X(_08482_));
 sg13g2_mux2_1 _15260_ (.A0(\cpu.icache.r_tag[4][13] ),
    .A1(\cpu.icache.r_tag[6][13] ),
    .S(net833),
    .X(_08483_));
 sg13g2_a22oi_1 _15261_ (.Y(_08484_),
    .B1(net830),
    .B2(_08483_),
    .A2(net577),
    .A1(\cpu.icache.r_tag[1][13] ));
 sg13g2_and2_1 _15262_ (.A(net941),
    .B(_08453_),
    .X(_08485_));
 sg13g2_buf_2 _15263_ (.A(_08485_),
    .X(_08486_));
 sg13g2_buf_1 _15264_ (.A(_08486_),
    .X(_08487_));
 sg13g2_buf_1 _15265_ (.A(_08487_),
    .X(_08488_));
 sg13g2_nand2_1 _15266_ (.Y(_08489_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(net576));
 sg13g2_nand4_1 _15267_ (.B(_08473_),
    .C(_08484_),
    .A(net578),
    .Y(_08490_),
    .D(_08489_));
 sg13g2_o21ai_1 _15268_ (.B1(_08490_),
    .Y(_08491_),
    .A1(\cpu.icache.r_tag[0][13] ),
    .A2(net579));
 sg13g2_xnor2_1 _15269_ (.Y(_08492_),
    .A(net400),
    .B(_08491_));
 sg13g2_buf_2 _15270_ (.A(_08425_),
    .X(_08493_));
 sg13g2_buf_2 _15271_ (.A(net829),
    .X(_08494_));
 sg13g2_mux4_1 _15272_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .S1(net834),
    .X(_08495_));
 sg13g2_mux4_1 _15273_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .S1(net836),
    .X(_08496_));
 sg13g2_mux4_1 _15274_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .S1(net834),
    .X(_08497_));
 sg13g2_mux4_1 _15275_ (.S0(net835),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .S1(net834),
    .X(_08498_));
 sg13g2_mux4_1 _15276_ (.S0(net946),
    .A0(_08495_),
    .A1(_08496_),
    .A2(_08497_),
    .A3(_08498_),
    .S1(net1084),
    .X(_08499_));
 sg13g2_nand2_1 _15277_ (.Y(_08500_),
    .A(net1163),
    .B(_08499_));
 sg13g2_mux4_1 _15278_ (.S0(_08430_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .S1(net834),
    .X(_08501_));
 sg13g2_mux4_1 _15279_ (.S0(_08430_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .S1(_08431_),
    .X(_08502_));
 sg13g2_buf_4 _15280_ (.X(_08503_),
    .A(_08425_));
 sg13g2_buf_2 _15281_ (.A(net947),
    .X(_08504_));
 sg13g2_mux4_1 _15282_ (.S0(_08503_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .S1(_08504_),
    .X(_08505_));
 sg13g2_mux4_1 _15283_ (.S0(_08503_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .S1(_08431_),
    .X(_08506_));
 sg13g2_mux4_1 _15284_ (.S0(net946),
    .A0(_08501_),
    .A1(_08502_),
    .A2(_08505_),
    .A3(_08506_),
    .S1(net1084),
    .X(_08507_));
 sg13g2_nand2_1 _15285_ (.Y(_08508_),
    .A(net945),
    .B(_08507_));
 sg13g2_nand3_1 _15286_ (.B(_08500_),
    .C(_08508_),
    .A(net1080),
    .Y(_08509_));
 sg13g2_o21ai_1 _15287_ (.B1(_08509_),
    .Y(_08510_),
    .A1(net733),
    .A2(net1080));
 sg13g2_buf_1 _15288_ (.A(_08510_),
    .X(_08511_));
 sg13g2_buf_1 _15289_ (.A(_08460_),
    .X(_08512_));
 sg13g2_buf_1 _15290_ (.A(_08477_),
    .X(_08513_));
 sg13g2_buf_1 _15291_ (.A(net655),
    .X(_08514_));
 sg13g2_buf_2 _15292_ (.A(net944),
    .X(_08515_));
 sg13g2_mux2_1 _15293_ (.A0(\cpu.icache.r_tag[4][12] ),
    .A1(\cpu.icache.r_tag[6][12] ),
    .S(net828),
    .X(_08516_));
 sg13g2_a22oi_1 _15294_ (.Y(_08517_),
    .B1(net830),
    .B2(_08516_),
    .A2(net574),
    .A1(\cpu.icache.r_tag[1][12] ));
 sg13g2_buf_1 _15295_ (.A(_08486_),
    .X(_08518_));
 sg13g2_buf_1 _15296_ (.A(net654),
    .X(_08519_));
 sg13g2_buf_1 _15297_ (.A(net943),
    .X(_08520_));
 sg13g2_nand2_1 _15298_ (.Y(_08521_),
    .A(net1160),
    .B(net1158));
 sg13g2_buf_2 _15299_ (.A(_08521_),
    .X(_08522_));
 sg13g2_nor2_1 _15300_ (.A(net827),
    .B(_08522_),
    .Y(_08523_));
 sg13g2_a22oi_1 _15301_ (.Y(_08524_),
    .B1(_08523_),
    .B2(\cpu.icache.r_tag[7][12] ),
    .A2(net573),
    .A1(\cpu.icache.r_tag[2][12] ));
 sg13g2_inv_1 _15302_ (.Y(_08525_),
    .A(_08448_));
 sg13g2_nor2_1 _15303_ (.A(net1076),
    .B(_08522_),
    .Y(_08526_));
 sg13g2_buf_1 _15304_ (.A(_08526_),
    .X(_08527_));
 sg13g2_buf_1 _15305_ (.A(_08527_),
    .X(_08528_));
 sg13g2_buf_2 _15306_ (.A(net653),
    .X(_08529_));
 sg13g2_nor3_1 _15307_ (.A(net941),
    .B(net1158),
    .C(_08448_),
    .Y(_08530_));
 sg13g2_buf_2 _15308_ (.A(_08530_),
    .X(_08531_));
 sg13g2_buf_2 _15309_ (.A(_08531_),
    .X(_08532_));
 sg13g2_buf_2 _15310_ (.A(net652),
    .X(_08533_));
 sg13g2_a22oi_1 _15311_ (.Y(_08534_),
    .B1(net571),
    .B2(\cpu.icache.r_tag[5][12] ),
    .A2(net572),
    .A1(\cpu.icache.r_tag[3][12] ));
 sg13g2_nand4_1 _15312_ (.B(_08517_),
    .C(_08524_),
    .A(net575),
    .Y(_08535_),
    .D(_08534_));
 sg13g2_o21ai_1 _15313_ (.B1(_08535_),
    .Y(_08536_),
    .A1(\cpu.icache.r_tag[0][12] ),
    .A2(net579));
 sg13g2_xnor2_1 _15314_ (.Y(_08537_),
    .A(net399),
    .B(_08536_));
 sg13g2_nand2_1 _15315_ (.Y(_08538_),
    .A(_08492_),
    .B(_08537_));
 sg13g2_inv_1 _15316_ (.Y(_08539_),
    .A(_08538_));
 sg13g2_buf_2 _15317_ (.A(_00190_),
    .X(_08540_));
 sg13g2_buf_1 _15318_ (.A(_08540_),
    .X(_08541_));
 sg13g2_buf_2 _15319_ (.A(_08503_),
    .X(_08542_));
 sg13g2_buf_1 _15320_ (.A(_08504_),
    .X(_08543_));
 sg13g2_mux4_1 _15321_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S1(net731),
    .X(_08544_));
 sg13g2_buf_2 _15322_ (.A(_08503_),
    .X(_08545_));
 sg13g2_mux4_1 _15323_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S1(net731),
    .X(_08546_));
 sg13g2_buf_1 _15324_ (.A(_08504_),
    .X(_08547_));
 sg13g2_mux4_1 _15325_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S1(net729),
    .X(_08548_));
 sg13g2_mux4_1 _15326_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S1(net729),
    .X(_08549_));
 sg13g2_buf_2 _15327_ (.A(net946),
    .X(_08550_));
 sg13g2_buf_1 _15328_ (.A(_08313_),
    .X(_08551_));
 sg13g2_mux4_1 _15329_ (.S0(net826),
    .A0(_08544_),
    .A1(_08546_),
    .A2(_08548_),
    .A3(_08549_),
    .S1(net939),
    .X(_08552_));
 sg13g2_mux4_1 _15330_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S1(net729),
    .X(_08553_));
 sg13g2_mux4_1 _15331_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S1(net729),
    .X(_08554_));
 sg13g2_buf_2 _15332_ (.A(_08503_),
    .X(_08555_));
 sg13g2_buf_1 _15333_ (.A(_08504_),
    .X(_08556_));
 sg13g2_mux4_1 _15334_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S1(net727),
    .X(_08557_));
 sg13g2_mux4_1 _15335_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S1(net727),
    .X(_08558_));
 sg13g2_mux4_1 _15336_ (.S0(net826),
    .A0(_08553_),
    .A1(_08554_),
    .A2(_08557_),
    .A3(_08558_),
    .S1(net939),
    .X(_08559_));
 sg13g2_buf_1 _15337_ (.A(net945),
    .X(_08560_));
 sg13g2_mux2_1 _15338_ (.A0(_08552_),
    .A1(_08559_),
    .S(net825),
    .X(_08561_));
 sg13g2_nand2b_1 _15339_ (.Y(_08562_),
    .B(_08561_),
    .A_N(_08541_));
 sg13g2_buf_1 _15340_ (.A(_08562_),
    .X(_08563_));
 sg13g2_a22oi_1 _15341_ (.Y(_08564_),
    .B1(net573),
    .B2(\cpu.icache.r_tag[2][21] ),
    .A2(net574),
    .A1(\cpu.icache.r_tag[1][21] ));
 sg13g2_and2_1 _15342_ (.A(net1078),
    .B(net940),
    .X(_08565_));
 sg13g2_buf_2 _15343_ (.A(_08565_),
    .X(_08566_));
 sg13g2_buf_2 _15344_ (.A(_08566_),
    .X(_08567_));
 sg13g2_a22oi_1 _15345_ (.Y(_08568_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][21] ),
    .A2(net572),
    .A1(\cpu.icache.r_tag[3][21] ));
 sg13g2_buf_1 _15346_ (.A(_08449_),
    .X(_08569_));
 sg13g2_buf_1 _15347_ (.A(net938),
    .X(_08570_));
 sg13g2_nor2_1 _15348_ (.A(net1160),
    .B(net1158),
    .Y(_08571_));
 sg13g2_buf_2 _15349_ (.A(_08571_),
    .X(_08572_));
 sg13g2_mux2_1 _15350_ (.A0(\cpu.icache.r_tag[5][21] ),
    .A1(\cpu.icache.r_tag[7][21] ),
    .S(net944),
    .X(_08573_));
 sg13g2_a22oi_1 _15351_ (.Y(_08574_),
    .B1(_08573_),
    .B2(net942),
    .A2(_08572_),
    .A1(\cpu.icache.r_tag[4][21] ));
 sg13g2_or2_1 _15352_ (.X(_08575_),
    .B(_08574_),
    .A(net824));
 sg13g2_nand3_1 _15353_ (.B(_08568_),
    .C(_08575_),
    .A(_08564_),
    .Y(_08576_));
 sg13g2_mux2_1 _15354_ (.A0(\cpu.icache.r_tag[0][21] ),
    .A1(_08576_),
    .S(net578),
    .X(_08577_));
 sg13g2_xnor2_1 _15355_ (.Y(_08578_),
    .A(net398),
    .B(_08577_));
 sg13g2_mux4_1 _15356_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S1(net729),
    .X(_08579_));
 sg13g2_mux4_1 _15357_ (.S0(_08542_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S1(net729),
    .X(_08580_));
 sg13g2_mux4_1 _15358_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S1(net727),
    .X(_08581_));
 sg13g2_mux4_1 _15359_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S1(net727),
    .X(_08582_));
 sg13g2_mux4_1 _15360_ (.S0(net826),
    .A0(_08579_),
    .A1(_08580_),
    .A2(_08581_),
    .A3(_08582_),
    .S1(net939),
    .X(_08583_));
 sg13g2_mux4_1 _15361_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S1(net727),
    .X(_08584_));
 sg13g2_mux4_1 _15362_ (.S0(_08555_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S1(net727),
    .X(_08585_));
 sg13g2_mux4_1 _15363_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S1(_08556_),
    .X(_08586_));
 sg13g2_mux4_1 _15364_ (.S0(_08555_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S1(_08556_),
    .X(_08587_));
 sg13g2_mux4_1 _15365_ (.S0(_08550_),
    .A0(_08584_),
    .A1(_08585_),
    .A2(_08586_),
    .A3(_08587_),
    .S1(_08551_),
    .X(_08588_));
 sg13g2_mux2_1 _15366_ (.A0(_08583_),
    .A1(_08588_),
    .S(_08438_),
    .X(_08589_));
 sg13g2_nand2b_1 _15367_ (.Y(_08590_),
    .B(_08589_),
    .A_N(net1075));
 sg13g2_buf_1 _15368_ (.A(_08590_),
    .X(_08591_));
 sg13g2_nor3_2 _15369_ (.A(_08450_),
    .B(_08462_),
    .C(net1079),
    .Y(_08592_));
 sg13g2_buf_1 _15370_ (.A(_08592_),
    .X(_08593_));
 sg13g2_buf_1 _15371_ (.A(net823),
    .X(_08594_));
 sg13g2_mux2_1 _15372_ (.A0(\cpu.icache.r_tag[7][22] ),
    .A1(\cpu.icache.r_tag[3][22] ),
    .S(net827),
    .X(_08595_));
 sg13g2_and2_1 _15373_ (.A(net1160),
    .B(net1158),
    .X(_08596_));
 sg13g2_buf_2 _15374_ (.A(_08596_),
    .X(_08597_));
 sg13g2_buf_1 _15375_ (.A(_08597_),
    .X(_08598_));
 sg13g2_a22oi_1 _15376_ (.Y(_08599_),
    .B1(_08595_),
    .B2(net822),
    .A2(net726),
    .A1(\cpu.icache.r_tag[4][22] ));
 sg13g2_a22oi_1 _15377_ (.Y(_08600_),
    .B1(net573),
    .B2(\cpu.icache.r_tag[2][22] ),
    .A2(net574),
    .A1(\cpu.icache.r_tag[1][22] ));
 sg13g2_a22oi_1 _15378_ (.Y(_08601_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][22] ),
    .A2(net652),
    .A1(\cpu.icache.r_tag[5][22] ));
 sg13g2_nand4_1 _15379_ (.B(_08599_),
    .C(_08600_),
    .A(net575),
    .Y(_08602_),
    .D(_08601_));
 sg13g2_o21ai_1 _15380_ (.B1(_08602_),
    .Y(_08603_),
    .A1(\cpu.icache.r_tag[0][22] ),
    .A2(net579));
 sg13g2_xor2_1 _15381_ (.B(_08603_),
    .A(net397),
    .X(_08604_));
 sg13g2_buf_2 _15382_ (.A(_08503_),
    .X(_08605_));
 sg13g2_buf_1 _15383_ (.A(_08504_),
    .X(_08606_));
 sg13g2_mux4_1 _15384_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .S1(net724),
    .X(_08607_));
 sg13g2_mux4_1 _15385_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .S1(net724),
    .X(_08608_));
 sg13g2_mux4_1 _15386_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .S1(net731),
    .X(_08609_));
 sg13g2_mux4_1 _15387_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .S1(net724),
    .X(_08610_));
 sg13g2_mux4_1 _15388_ (.S0(net826),
    .A0(_08607_),
    .A1(_08608_),
    .A2(_08609_),
    .A3(_08610_),
    .S1(net939),
    .X(_08611_));
 sg13g2_mux4_1 _15389_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .S1(net724),
    .X(_08612_));
 sg13g2_mux4_1 _15390_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .S1(net724),
    .X(_08613_));
 sg13g2_mux4_1 _15391_ (.S0(_08545_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .S1(_08543_),
    .X(_08614_));
 sg13g2_mux4_1 _15392_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .S1(_08543_),
    .X(_08615_));
 sg13g2_mux4_1 _15393_ (.S0(_08550_),
    .A0(_08612_),
    .A1(_08613_),
    .A2(_08614_),
    .A3(_08615_),
    .S1(_08551_),
    .X(_08616_));
 sg13g2_mux2_1 _15394_ (.A0(_08611_),
    .A1(_08616_),
    .S(net825),
    .X(_08617_));
 sg13g2_nand2b_1 _15395_ (.Y(_08618_),
    .B(_08617_),
    .A_N(net1075));
 sg13g2_buf_2 _15396_ (.A(_08618_),
    .X(_08619_));
 sg13g2_buf_1 _15397_ (.A(net651),
    .X(_08620_));
 sg13g2_a22oi_1 _15398_ (.Y(_08621_),
    .B1(net570),
    .B2(\cpu.icache.r_tag[6][16] ),
    .A2(net577),
    .A1(\cpu.icache.r_tag[1][16] ));
 sg13g2_a22oi_1 _15399_ (.Y(_08622_),
    .B1(net726),
    .B2(\cpu.icache.r_tag[4][16] ),
    .A2(net576),
    .A1(\cpu.icache.r_tag[2][16] ));
 sg13g2_mux2_1 _15400_ (.A0(\cpu.icache.r_tag[7][16] ),
    .A1(\cpu.icache.r_tag[3][16] ),
    .S(net938),
    .X(_08623_));
 sg13g2_buf_1 _15401_ (.A(net828),
    .X(_08624_));
 sg13g2_a22oi_1 _15402_ (.Y(_08625_),
    .B1(_08623_),
    .B2(net723),
    .A2(net832),
    .A1(\cpu.icache.r_tag[5][16] ));
 sg13g2_nand2b_1 _15403_ (.Y(_08626_),
    .B(net831),
    .A_N(_08625_));
 sg13g2_nand4_1 _15404_ (.B(_08621_),
    .C(_08622_),
    .A(net578),
    .Y(_08627_),
    .D(_08626_));
 sg13g2_o21ai_1 _15405_ (.B1(_08627_),
    .Y(_08628_),
    .A1(\cpu.icache.r_tag[0][16] ),
    .A2(net579));
 sg13g2_xor2_1 _15406_ (.B(_08628_),
    .A(_08619_),
    .X(_08629_));
 sg13g2_buf_1 _15407_ (.A(_08504_),
    .X(_08630_));
 sg13g2_mux4_1 _15408_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .S1(net722),
    .X(_08631_));
 sg13g2_buf_2 _15409_ (.A(_08503_),
    .X(_08632_));
 sg13g2_mux4_1 _15410_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .S1(net722),
    .X(_08633_));
 sg13g2_mux4_1 _15411_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .S1(net724),
    .X(_08634_));
 sg13g2_mux4_1 _15412_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .S1(net724),
    .X(_08635_));
 sg13g2_buf_1 _15413_ (.A(_08434_),
    .X(_08636_));
 sg13g2_buf_1 _15414_ (.A(net1084),
    .X(_08637_));
 sg13g2_mux4_1 _15415_ (.S0(net821),
    .A0(_08631_),
    .A1(_08633_),
    .A2(_08634_),
    .A3(_08635_),
    .S1(net937),
    .X(_08638_));
 sg13g2_mux4_1 _15416_ (.S0(net725),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .S1(net724),
    .X(_08639_));
 sg13g2_mux4_1 _15417_ (.S0(_08605_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .S1(_08606_),
    .X(_08640_));
 sg13g2_mux4_1 _15418_ (.S0(_08545_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .S1(net731),
    .X(_08641_));
 sg13g2_mux4_1 _15419_ (.S0(_08605_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .S1(_08606_),
    .X(_08642_));
 sg13g2_mux4_1 _15420_ (.S0(net826),
    .A0(_08639_),
    .A1(_08640_),
    .A2(_08641_),
    .A3(_08642_),
    .S1(net937),
    .X(_08643_));
 sg13g2_mux2_1 _15421_ (.A0(_08638_),
    .A1(_08643_),
    .S(net825),
    .X(_08644_));
 sg13g2_nand2b_1 _15422_ (.Y(_08645_),
    .B(_08644_),
    .A_N(net1075));
 sg13g2_buf_2 _15423_ (.A(_08645_),
    .X(_08646_));
 sg13g2_mux2_1 _15424_ (.A0(\cpu.icache.r_tag[7][17] ),
    .A1(\cpu.icache.r_tag[3][17] ),
    .S(net938),
    .X(_08647_));
 sg13g2_a22oi_1 _15425_ (.Y(_08648_),
    .B1(_08647_),
    .B2(net723),
    .A2(net832),
    .A1(\cpu.icache.r_tag[5][17] ));
 sg13g2_nand2b_1 _15426_ (.Y(_08649_),
    .B(net831),
    .A_N(_08648_));
 sg13g2_mux2_1 _15427_ (.A0(\cpu.icache.r_tag[4][17] ),
    .A1(\cpu.icache.r_tag[6][17] ),
    .S(net833),
    .X(_08650_));
 sg13g2_a22oi_1 _15428_ (.Y(_08651_),
    .B1(net830),
    .B2(_08650_),
    .A2(net577),
    .A1(\cpu.icache.r_tag[1][17] ));
 sg13g2_nand2_1 _15429_ (.Y(_08652_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net576));
 sg13g2_nand4_1 _15430_ (.B(_08649_),
    .C(_08651_),
    .A(net578),
    .Y(_08653_),
    .D(_08652_));
 sg13g2_o21ai_1 _15431_ (.B1(_08653_),
    .Y(_08654_),
    .A1(\cpu.icache.r_tag[0][17] ),
    .A2(net579));
 sg13g2_xor2_1 _15432_ (.B(_08654_),
    .A(net395),
    .X(_08655_));
 sg13g2_nor4_1 _15433_ (.A(_08578_),
    .B(_08604_),
    .C(_08629_),
    .D(_08655_),
    .Y(_08656_));
 sg13g2_mux4_1 _15434_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S1(net727),
    .X(_08657_));
 sg13g2_mux4_1 _15435_ (.S0(net728),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S1(net727),
    .X(_08658_));
 sg13g2_mux4_1 _15436_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S1(net838),
    .X(_08659_));
 sg13g2_mux4_1 _15437_ (.S0(_08493_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S1(_08422_),
    .X(_08660_));
 sg13g2_mux4_1 _15438_ (.S0(net945),
    .A0(_08657_),
    .A1(_08658_),
    .A2(_08659_),
    .A3(_08660_),
    .S1(net939),
    .X(_08661_));
 sg13g2_nand2b_1 _15439_ (.Y(_08662_),
    .B(net1080),
    .A_N(_08661_));
 sg13g2_mux4_1 _15440_ (.S0(net733),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S1(net735),
    .X(_08663_));
 sg13g2_mux4_1 _15441_ (.S0(net733),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S1(net735),
    .X(_08664_));
 sg13g2_mux4_1 _15442_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S1(net735),
    .X(_08665_));
 sg13g2_mux4_1 _15443_ (.S0(net733),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S1(net735),
    .X(_08666_));
 sg13g2_mux4_1 _15444_ (.S0(net945),
    .A0(_08663_),
    .A1(_08664_),
    .A2(_08665_),
    .A3(_08666_),
    .S1(net937),
    .X(_08667_));
 sg13g2_nor2_1 _15445_ (.A(net821),
    .B(_08336_),
    .Y(_08668_));
 sg13g2_a22oi_1 _15446_ (.Y(_08669_),
    .B1(_08667_),
    .B2(_08668_),
    .A2(_08662_),
    .A1(net821));
 sg13g2_buf_2 _15447_ (.A(_08669_),
    .X(_08670_));
 sg13g2_mux2_1 _15448_ (.A0(\cpu.icache.r_tag[7][14] ),
    .A1(\cpu.icache.r_tag[3][14] ),
    .S(net943),
    .X(_08671_));
 sg13g2_a22oi_1 _15449_ (.Y(_08672_),
    .B1(_08671_),
    .B2(net833),
    .A2(net832),
    .A1(\cpu.icache.r_tag[5][14] ));
 sg13g2_nand2b_1 _15450_ (.Y(_08673_),
    .B(net831),
    .A_N(_08672_));
 sg13g2_mux2_1 _15451_ (.A0(\cpu.icache.r_tag[4][14] ),
    .A1(\cpu.icache.r_tag[6][14] ),
    .S(net828),
    .X(_08674_));
 sg13g2_a22oi_1 _15452_ (.Y(_08675_),
    .B1(net830),
    .B2(_08674_),
    .A2(net574),
    .A1(\cpu.icache.r_tag[1][14] ));
 sg13g2_nand2_1 _15453_ (.Y(_08676_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(net576));
 sg13g2_nand4_1 _15454_ (.B(_08673_),
    .C(_08675_),
    .A(net575),
    .Y(_08677_),
    .D(_08676_));
 sg13g2_o21ai_1 _15455_ (.B1(_08677_),
    .Y(_08678_),
    .A1(\cpu.icache.r_tag[0][14] ),
    .A2(net579));
 sg13g2_xor2_1 _15456_ (.B(_08678_),
    .A(net394),
    .X(_08679_));
 sg13g2_mux4_1 _15457_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S1(net731),
    .X(_08680_));
 sg13g2_mux4_1 _15458_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S1(net731),
    .X(_08681_));
 sg13g2_mux4_1 _15459_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S1(net729),
    .X(_08682_));
 sg13g2_mux4_1 _15460_ (.S0(_08542_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S1(net729),
    .X(_08683_));
 sg13g2_mux4_1 _15461_ (.S0(net826),
    .A0(_08680_),
    .A1(_08681_),
    .A2(_08682_),
    .A3(_08683_),
    .S1(net939),
    .X(_08684_));
 sg13g2_mux4_1 _15462_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S1(net731),
    .X(_08685_));
 sg13g2_mux4_1 _15463_ (.S0(net730),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S1(net731),
    .X(_08686_));
 sg13g2_mux4_1 _15464_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S1(_08547_),
    .X(_08687_));
 sg13g2_mux4_1 _15465_ (.S0(net732),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S1(_08547_),
    .X(_08688_));
 sg13g2_mux4_1 _15466_ (.S0(net826),
    .A0(_08685_),
    .A1(_08686_),
    .A2(_08687_),
    .A3(_08688_),
    .S1(net939),
    .X(_08689_));
 sg13g2_mux2_1 _15467_ (.A0(_08684_),
    .A1(_08689_),
    .S(net825),
    .X(_08690_));
 sg13g2_nand2b_1 _15468_ (.Y(_08691_),
    .B(_08690_),
    .A_N(_08541_));
 sg13g2_buf_1 _15469_ (.A(_08691_),
    .X(_08692_));
 sg13g2_mux2_1 _15470_ (.A0(\cpu.icache.r_tag[7][20] ),
    .A1(\cpu.icache.r_tag[3][20] ),
    .S(net827),
    .X(_08693_));
 sg13g2_a22oi_1 _15471_ (.Y(_08694_),
    .B1(_08693_),
    .B2(net822),
    .A2(net726),
    .A1(\cpu.icache.r_tag[4][20] ));
 sg13g2_a22oi_1 _15472_ (.Y(_08695_),
    .B1(net576),
    .B2(\cpu.icache.r_tag[2][20] ),
    .A2(net577),
    .A1(\cpu.icache.r_tag[1][20] ));
 sg13g2_a22oi_1 _15473_ (.Y(_08696_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][20] ),
    .A2(net652),
    .A1(\cpu.icache.r_tag[5][20] ));
 sg13g2_nand4_1 _15474_ (.B(_08694_),
    .C(_08695_),
    .A(net578),
    .Y(_08697_),
    .D(_08696_));
 sg13g2_o21ai_1 _15475_ (.B1(_08697_),
    .Y(_08698_),
    .A1(\cpu.icache.r_tag[0][20] ),
    .A2(net579));
 sg13g2_xor2_1 _15476_ (.B(_08698_),
    .A(net393),
    .X(_08699_));
 sg13g2_mux4_1 _15477_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S1(net722),
    .X(_08700_));
 sg13g2_mux4_1 _15478_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S1(net722),
    .X(_08701_));
 sg13g2_mux4_1 _15479_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S1(net722),
    .X(_08702_));
 sg13g2_mux4_1 _15480_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S1(net722),
    .X(_08703_));
 sg13g2_mux4_1 _15481_ (.S0(net821),
    .A0(_08700_),
    .A1(_08701_),
    .A2(_08702_),
    .A3(_08703_),
    .S1(net937),
    .X(_08704_));
 sg13g2_mux4_1 _15482_ (.S0(_08632_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S1(net722),
    .X(_08705_));
 sg13g2_mux4_1 _15483_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S1(net722),
    .X(_08706_));
 sg13g2_mux4_1 _15484_ (.S0(_08632_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S1(_08630_),
    .X(_08707_));
 sg13g2_mux4_1 _15485_ (.S0(net721),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S1(_08630_),
    .X(_08708_));
 sg13g2_mux4_1 _15486_ (.S0(net821),
    .A0(_08705_),
    .A1(_08706_),
    .A2(_08707_),
    .A3(_08708_),
    .S1(net937),
    .X(_08709_));
 sg13g2_mux2_1 _15487_ (.A0(_08704_),
    .A1(_08709_),
    .S(net825),
    .X(_08710_));
 sg13g2_nand2b_1 _15488_ (.Y(_08711_),
    .B(_08710_),
    .A_N(net1075));
 sg13g2_buf_2 _15489_ (.A(_08711_),
    .X(_08712_));
 sg13g2_buf_1 _15490_ (.A(net575),
    .X(_08713_));
 sg13g2_a22oi_1 _15491_ (.Y(_08714_),
    .B1(net576),
    .B2(\cpu.icache.r_tag[2][19] ),
    .A2(net577),
    .A1(\cpu.icache.r_tag[1][19] ));
 sg13g2_mux4_1 _15492_ (.S0(net942),
    .A0(\cpu.icache.r_tag[4][19] ),
    .A1(\cpu.icache.r_tag[5][19] ),
    .A2(\cpu.icache.r_tag[6][19] ),
    .A3(\cpu.icache.r_tag[7][19] ),
    .S1(net833),
    .X(_08715_));
 sg13g2_a22oi_1 _15493_ (.Y(_08716_),
    .B1(_08715_),
    .B2(net1076),
    .A2(net572),
    .A1(\cpu.icache.r_tag[3][19] ));
 sg13g2_nand3_1 _15494_ (.B(_08714_),
    .C(_08716_),
    .A(net578),
    .Y(_08717_));
 sg13g2_o21ai_1 _15495_ (.B1(_08717_),
    .Y(_08718_),
    .A1(\cpu.icache.r_tag[0][19] ),
    .A2(_08713_));
 sg13g2_xor2_1 _15496_ (.B(_08718_),
    .A(net392),
    .X(_08719_));
 sg13g2_mux4_1 _15497_ (.S0(_08425_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .S1(_08504_),
    .X(_08720_));
 sg13g2_mux4_1 _15498_ (.S0(_08503_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .S1(_08504_),
    .X(_08721_));
 sg13g2_mux4_1 _15499_ (.S0(_08425_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .S1(_08421_),
    .X(_08722_));
 sg13g2_mux4_1 _15500_ (.S0(_08425_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .S1(net947),
    .X(_08723_));
 sg13g2_mux4_1 _15501_ (.S0(net945),
    .A0(_08720_),
    .A1(_08721_),
    .A2(_08722_),
    .A3(_08723_),
    .S1(net946),
    .X(_08724_));
 sg13g2_nand2b_1 _15502_ (.Y(_08725_),
    .B(net1080),
    .A_N(_08724_));
 sg13g2_mux4_1 _15503_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .S1(net838),
    .X(_08726_));
 sg13g2_mux4_1 _15504_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .S1(net838),
    .X(_08727_));
 sg13g2_mux4_1 _15505_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .S1(net838),
    .X(_08728_));
 sg13g2_mux4_1 _15506_ (.S0(_08493_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .S1(net838),
    .X(_08729_));
 sg13g2_mux4_1 _15507_ (.S0(_08438_),
    .A0(_08726_),
    .A1(_08727_),
    .A2(_08728_),
    .A3(_08729_),
    .S1(net821),
    .X(_08730_));
 sg13g2_nor2_1 _15508_ (.A(net937),
    .B(_08336_),
    .Y(_08731_));
 sg13g2_a22oi_1 _15509_ (.Y(_08732_),
    .B1(_08730_),
    .B2(_08731_),
    .A2(_08725_),
    .A1(net937));
 sg13g2_buf_1 _15510_ (.A(_08732_),
    .X(_08733_));
 sg13g2_and2_1 _15511_ (.A(net1079),
    .B(_08455_),
    .X(_08734_));
 sg13g2_buf_1 _15512_ (.A(_08734_),
    .X(_08735_));
 sg13g2_buf_1 _15513_ (.A(_08735_),
    .X(_08736_));
 sg13g2_mux2_1 _15514_ (.A0(\cpu.icache.r_tag[7][15] ),
    .A1(\cpu.icache.r_tag[3][15] ),
    .S(net1079),
    .X(_08737_));
 sg13g2_a22oi_1 _15515_ (.Y(_08738_),
    .B1(_08737_),
    .B2(net828),
    .A2(_08467_),
    .A1(\cpu.icache.r_tag[5][15] ));
 sg13g2_nand2b_1 _15516_ (.Y(_08739_),
    .B(net942),
    .A_N(_08738_));
 sg13g2_a22oi_1 _15517_ (.Y(_08740_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][15] ),
    .A2(net656),
    .A1(\cpu.icache.r_tag[2][15] ));
 sg13g2_a22oi_1 _15518_ (.Y(_08741_),
    .B1(net823),
    .B2(\cpu.icache.r_tag[4][15] ),
    .A2(net655),
    .A1(\cpu.icache.r_tag[1][15] ));
 sg13g2_nand3_1 _15519_ (.B(_08740_),
    .C(_08741_),
    .A(_08739_),
    .Y(_08742_));
 sg13g2_a21oi_1 _15520_ (.A1(\cpu.icache.r_tag[0][15] ),
    .A2(_08736_),
    .Y(_08743_),
    .B1(_08742_));
 sg13g2_xor2_1 _15521_ (.B(_08743_),
    .A(net448),
    .X(_08744_));
 sg13g2_mux4_1 _15522_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S1(net838),
    .X(_08745_));
 sg13g2_mux4_1 _15523_ (.S0(net829),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S1(net838),
    .X(_08746_));
 sg13g2_mux4_1 _15524_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S1(net836),
    .X(_08747_));
 sg13g2_mux4_1 _15525_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S1(net836),
    .X(_08748_));
 sg13g2_mux4_1 _15526_ (.S0(net826),
    .A0(_08745_),
    .A1(_08746_),
    .A2(_08747_),
    .A3(_08748_),
    .S1(net939),
    .X(_08749_));
 sg13g2_mux4_1 _15527_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S1(net836),
    .X(_08750_));
 sg13g2_mux4_1 _15528_ (.S0(net837),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S1(net838),
    .X(_08751_));
 sg13g2_mux4_1 _15529_ (.S0(_08426_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S1(_08427_),
    .X(_08752_));
 sg13g2_mux4_1 _15530_ (.S0(_08426_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S1(_08427_),
    .X(_08753_));
 sg13g2_mux4_1 _15531_ (.S0(_08434_),
    .A0(_08750_),
    .A1(_08751_),
    .A2(_08752_),
    .A3(_08753_),
    .S1(net1084),
    .X(_08754_));
 sg13g2_mux2_1 _15532_ (.A0(_08749_),
    .A1(_08754_),
    .S(net945),
    .X(_08755_));
 sg13g2_nand2b_1 _15533_ (.Y(_08756_),
    .B(_08755_),
    .A_N(net1075));
 sg13g2_buf_1 _15534_ (.A(_08756_),
    .X(_08757_));
 sg13g2_and2_1 _15535_ (.A(\cpu.icache.r_tag[6][18] ),
    .B(_08566_),
    .X(_08758_));
 sg13g2_a221oi_1 _15536_ (.B2(\cpu.icache.r_tag[5][18] ),
    .C1(_08758_),
    .B1(net652),
    .A1(\cpu.icache.r_tag[3][18] ),
    .Y(_08759_),
    .A2(net653));
 sg13g2_a22oi_1 _15537_ (.Y(_08760_),
    .B1(_08523_),
    .B2(\cpu.icache.r_tag[7][18] ),
    .A2(net573),
    .A1(\cpu.icache.r_tag[2][18] ));
 sg13g2_a22oi_1 _15538_ (.Y(_08761_),
    .B1(net823),
    .B2(\cpu.icache.r_tag[4][18] ),
    .A2(net574),
    .A1(\cpu.icache.r_tag[1][18] ));
 sg13g2_nand4_1 _15539_ (.B(_08759_),
    .C(_08760_),
    .A(net659),
    .Y(_08762_),
    .D(_08761_));
 sg13g2_o21ai_1 _15540_ (.B1(_08762_),
    .Y(_08763_),
    .A1(\cpu.icache.r_tag[0][18] ),
    .A2(net578));
 sg13g2_xnor2_1 _15541_ (.Y(_08764_),
    .A(net447),
    .B(_08763_));
 sg13g2_mux4_1 _15542_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S1(net947),
    .X(_08765_));
 sg13g2_mux4_1 _15543_ (.S0(_08425_),
    .A0(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S1(net947),
    .X(_08766_));
 sg13g2_mux4_1 _15544_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S1(net1085),
    .X(_08767_));
 sg13g2_mux4_1 _15545_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S1(net1085),
    .X(_08768_));
 sg13g2_mux4_1 _15546_ (.S0(net946),
    .A0(_08765_),
    .A1(_08766_),
    .A2(_08767_),
    .A3(_08768_),
    .S1(net1084),
    .X(_08769_));
 sg13g2_mux4_1 _15547_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S1(net1085),
    .X(_08770_));
 sg13g2_mux4_1 _15548_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S1(net947),
    .X(_08771_));
 sg13g2_mux4_1 _15549_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S1(net1085),
    .X(_08772_));
 sg13g2_mux4_1 _15550_ (.S0(net1082),
    .A0(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S1(net1085),
    .X(_08773_));
 sg13g2_mux4_1 _15551_ (.S0(net946),
    .A0(_08770_),
    .A1(_08771_),
    .A2(_08772_),
    .A3(_08773_),
    .S1(net1084),
    .X(_08774_));
 sg13g2_mux2_1 _15552_ (.A0(_08769_),
    .A1(_08774_),
    .S(net945),
    .X(_08775_));
 sg13g2_nand2b_1 _15553_ (.Y(_08776_),
    .B(_08775_),
    .A_N(net1075));
 sg13g2_buf_1 _15554_ (.A(_08776_),
    .X(_08777_));
 sg13g2_a22oi_1 _15555_ (.Y(_08778_),
    .B1(net823),
    .B2(\cpu.icache.r_tag[4][23] ),
    .A2(_08531_),
    .A1(\cpu.icache.r_tag[5][23] ));
 sg13g2_a22oi_1 _15556_ (.Y(_08779_),
    .B1(_08566_),
    .B2(\cpu.icache.r_tag[6][23] ),
    .A2(net655),
    .A1(\cpu.icache.r_tag[1][23] ));
 sg13g2_mux2_1 _15557_ (.A0(\cpu.icache.r_tag[7][23] ),
    .A1(\cpu.icache.r_tag[3][23] ),
    .S(net943),
    .X(_08780_));
 sg13g2_a22oi_1 _15558_ (.Y(_08781_),
    .B1(net822),
    .B2(_08780_),
    .A2(net654),
    .A1(\cpu.icache.r_tag[2][23] ));
 sg13g2_nand4_1 _15559_ (.B(_08778_),
    .C(_08779_),
    .A(net658),
    .Y(_08782_),
    .D(_08781_));
 sg13g2_o21ai_1 _15560_ (.B1(_08782_),
    .Y(_08783_),
    .A1(\cpu.icache.r_tag[0][23] ),
    .A2(net659));
 sg13g2_xor2_1 _15561_ (.B(_08783_),
    .A(net496),
    .X(_08784_));
 sg13g2_buf_1 _15562_ (.A(\cpu.ex.pc[7] ),
    .X(_08785_));
 sg13g2_a22oi_1 _15563_ (.Y(_08786_),
    .B1(net652),
    .B2(\cpu.icache.r_tag[5][7] ),
    .A2(net656),
    .A1(\cpu.icache.r_tag[2][7] ));
 sg13g2_a22oi_1 _15564_ (.Y(_08787_),
    .B1(net653),
    .B2(\cpu.icache.r_tag[3][7] ),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][7] ));
 sg13g2_buf_1 _15565_ (.A(net1078),
    .X(_08788_));
 sg13g2_mux2_1 _15566_ (.A0(\cpu.icache.r_tag[4][7] ),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(net936),
    .X(_08789_));
 sg13g2_a22oi_1 _15567_ (.Y(_08790_),
    .B1(_08789_),
    .B2(net941),
    .A2(_08597_),
    .A1(\cpu.icache.r_tag[7][7] ));
 sg13g2_or2_1 _15568_ (.X(_08791_),
    .B(_08790_),
    .A(net827));
 sg13g2_nand3_1 _15569_ (.B(_08787_),
    .C(_08791_),
    .A(_08786_),
    .Y(_08792_));
 sg13g2_mux2_1 _15570_ (.A0(\cpu.icache.r_tag[0][7] ),
    .A1(_08792_),
    .S(net659),
    .X(_08793_));
 sg13g2_xnor2_1 _15571_ (.Y(_08794_),
    .A(_08785_),
    .B(_08793_));
 sg13g2_inv_1 _15572_ (.Y(_08795_),
    .A(\cpu.ex.pc[8] ));
 sg13g2_a22oi_1 _15573_ (.Y(_08796_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][8] ),
    .A2(net656),
    .A1(\cpu.icache.r_tag[2][8] ));
 sg13g2_a22oi_1 _15574_ (.Y(_08797_),
    .B1(net653),
    .B2(\cpu.icache.r_tag[3][8] ),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][8] ));
 sg13g2_mux2_1 _15575_ (.A0(\cpu.icache.r_tag[5][8] ),
    .A1(\cpu.icache.r_tag[7][8] ),
    .S(net936),
    .X(_08798_));
 sg13g2_a22oi_1 _15576_ (.Y(_08799_),
    .B1(_08798_),
    .B2(net1077),
    .A2(_08572_),
    .A1(\cpu.icache.r_tag[4][8] ));
 sg13g2_or2_1 _15577_ (.X(_08800_),
    .B(_08799_),
    .A(net827));
 sg13g2_nand4_1 _15578_ (.B(_08796_),
    .C(_08797_),
    .A(net658),
    .Y(_08801_),
    .D(_08800_));
 sg13g2_o21ai_1 _15579_ (.B1(_08801_),
    .Y(_08802_),
    .A1(\cpu.icache.r_tag[0][8] ),
    .A2(net575));
 sg13g2_xnor2_1 _15580_ (.Y(_08803_),
    .A(_08795_),
    .B(_08802_));
 sg13g2_buf_2 _15581_ (.A(\cpu.ex.pc[5] ),
    .X(_08804_));
 sg13g2_mux2_1 _15582_ (.A0(\cpu.icache.r_tag[7][5] ),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net943),
    .X(_08805_));
 sg13g2_a22oi_1 _15583_ (.Y(_08806_),
    .B1(_08805_),
    .B2(net828),
    .A2(net832),
    .A1(\cpu.icache.r_tag[5][5] ));
 sg13g2_nand2b_1 _15584_ (.Y(_08807_),
    .B(net942),
    .A_N(_08806_));
 sg13g2_mux2_1 _15585_ (.A0(\cpu.icache.r_tag[4][5] ),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net944),
    .X(_08808_));
 sg13g2_a22oi_1 _15586_ (.Y(_08809_),
    .B1(net940),
    .B2(_08808_),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][5] ));
 sg13g2_nand2_1 _15587_ (.Y(_08810_),
    .A(\cpu.icache.r_tag[2][5] ),
    .B(net573));
 sg13g2_nand4_1 _15588_ (.B(_08807_),
    .C(_08809_),
    .A(net659),
    .Y(_08811_),
    .D(_08810_));
 sg13g2_o21ai_1 _15589_ (.B1(_08811_),
    .Y(_08812_),
    .A1(\cpu.icache.r_tag[0][5] ),
    .A2(net575));
 sg13g2_xor2_1 _15590_ (.B(_08812_),
    .A(_08804_),
    .X(_08813_));
 sg13g2_buf_1 _15591_ (.A(_08624_),
    .X(_08814_));
 sg13g2_mux4_1 _15592_ (.S0(net831),
    .A0(\cpu.icache.r_valid[0] ),
    .A1(\cpu.icache.r_valid[1] ),
    .A2(\cpu.icache.r_valid[2] ),
    .A3(\cpu.icache.r_valid[3] ),
    .S1(net649),
    .X(_08815_));
 sg13g2_mux4_1 _15593_ (.S0(net831),
    .A0(\cpu.icache.r_valid[4] ),
    .A1(\cpu.icache.r_valid[5] ),
    .A2(\cpu.icache.r_valid[6] ),
    .A3(\cpu.icache.r_valid[7] ),
    .S1(net723),
    .X(_08816_));
 sg13g2_mux2_1 _15594_ (.A0(_08815_),
    .A1(_08816_),
    .S(_08451_),
    .X(_08817_));
 sg13g2_nand4_1 _15595_ (.B(_08803_),
    .C(_08813_),
    .A(_08794_),
    .Y(_08818_),
    .D(_08817_));
 sg13g2_buf_1 _15596_ (.A(\cpu.ex.pc[6] ),
    .X(_08819_));
 sg13g2_mux2_1 _15597_ (.A0(\cpu.icache.r_tag[7][6] ),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net1079),
    .X(_08820_));
 sg13g2_a22oi_1 _15598_ (.Y(_08821_),
    .B1(_08820_),
    .B2(net828),
    .A2(_08467_),
    .A1(\cpu.icache.r_tag[5][6] ));
 sg13g2_nand2b_1 _15599_ (.Y(_08822_),
    .B(net942),
    .A_N(_08821_));
 sg13g2_mux2_1 _15600_ (.A0(\cpu.icache.r_tag[4][6] ),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net944),
    .X(_08823_));
 sg13g2_a22oi_1 _15601_ (.Y(_08824_),
    .B1(net940),
    .B2(_08823_),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][6] ));
 sg13g2_nand2_1 _15602_ (.Y(_08825_),
    .A(\cpu.icache.r_tag[2][6] ),
    .B(net656));
 sg13g2_nand4_1 _15603_ (.B(_08822_),
    .C(_08824_),
    .A(net658),
    .Y(_08826_),
    .D(_08825_));
 sg13g2_o21ai_1 _15604_ (.B1(_08826_),
    .Y(_08827_),
    .A1(\cpu.icache.r_tag[0][6] ),
    .A2(net575));
 sg13g2_xor2_1 _15605_ (.B(_08827_),
    .A(_08819_),
    .X(_08828_));
 sg13g2_buf_1 _15606_ (.A(\cpu.ex.pc[10] ),
    .X(_08829_));
 sg13g2_mux2_1 _15607_ (.A0(\cpu.icache.r_tag[7][10] ),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(net943),
    .X(_08830_));
 sg13g2_a22oi_1 _15608_ (.Y(_08831_),
    .B1(_08830_),
    .B2(net822),
    .A2(net823),
    .A1(\cpu.icache.r_tag[4][10] ));
 sg13g2_a22oi_1 _15609_ (.Y(_08832_),
    .B1(net652),
    .B2(\cpu.icache.r_tag[5][10] ),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][10] ));
 sg13g2_a22oi_1 _15610_ (.Y(_08833_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][10] ),
    .A2(net654),
    .A1(\cpu.icache.r_tag[2][10] ));
 sg13g2_nand4_1 _15611_ (.B(_08831_),
    .C(_08832_),
    .A(net658),
    .Y(_08834_),
    .D(_08833_));
 sg13g2_o21ai_1 _15612_ (.B1(_08834_),
    .Y(_08835_),
    .A1(\cpu.icache.r_tag[0][10] ),
    .A2(net659));
 sg13g2_xor2_1 _15613_ (.B(_08835_),
    .A(_08829_),
    .X(_08836_));
 sg13g2_buf_1 _15614_ (.A(\cpu.ex.pc[11] ),
    .X(_08837_));
 sg13g2_mux2_1 _15615_ (.A0(\cpu.icache.r_tag[7][11] ),
    .A1(\cpu.icache.r_tag[3][11] ),
    .S(net943),
    .X(_08838_));
 sg13g2_a22oi_1 _15616_ (.Y(_08839_),
    .B1(_08838_),
    .B2(net822),
    .A2(net823),
    .A1(\cpu.icache.r_tag[4][11] ));
 sg13g2_a22oi_1 _15617_ (.Y(_08840_),
    .B1(net652),
    .B2(\cpu.icache.r_tag[5][11] ),
    .A2(net656),
    .A1(\cpu.icache.r_tag[2][11] ));
 sg13g2_a22oi_1 _15618_ (.Y(_08841_),
    .B1(net651),
    .B2(\cpu.icache.r_tag[6][11] ),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][11] ));
 sg13g2_nand3_1 _15619_ (.B(_08840_),
    .C(_08841_),
    .A(_08839_),
    .Y(_08842_));
 sg13g2_mux2_1 _15620_ (.A0(\cpu.icache.r_tag[0][11] ),
    .A1(_08842_),
    .S(net659),
    .X(_08843_));
 sg13g2_xnor2_1 _15621_ (.Y(_08844_),
    .A(_08837_),
    .B(_08843_));
 sg13g2_buf_1 _15622_ (.A(\cpu.ex.pc[9] ),
    .X(_08845_));
 sg13g2_a22oi_1 _15623_ (.Y(_08846_),
    .B1(net652),
    .B2(\cpu.icache.r_tag[5][9] ),
    .A2(net657),
    .A1(\cpu.icache.r_tag[1][9] ));
 sg13g2_a22oi_1 _15624_ (.Y(_08847_),
    .B1(net823),
    .B2(\cpu.icache.r_tag[4][9] ),
    .A2(net656),
    .A1(\cpu.icache.r_tag[2][9] ));
 sg13g2_mux2_1 _15625_ (.A0(\cpu.icache.r_tag[7][9] ),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(net1079),
    .X(_08848_));
 sg13g2_a22oi_1 _15626_ (.Y(_08849_),
    .B1(_08848_),
    .B2(net1077),
    .A2(net940),
    .A1(\cpu.icache.r_tag[6][9] ));
 sg13g2_nand2b_1 _15627_ (.Y(_08850_),
    .B(net833),
    .A_N(_08849_));
 sg13g2_nand4_1 _15628_ (.B(_08846_),
    .C(_08847_),
    .A(net659),
    .Y(_08851_),
    .D(_08850_));
 sg13g2_o21ai_1 _15629_ (.B1(_08851_),
    .Y(_08852_),
    .A1(\cpu.icache.r_tag[0][9] ),
    .A2(net575));
 sg13g2_xor2_1 _15630_ (.B(_08852_),
    .A(_08845_),
    .X(_08853_));
 sg13g2_nand4_1 _15631_ (.B(_08836_),
    .C(_08844_),
    .A(_08828_),
    .Y(_08854_),
    .D(_08853_));
 sg13g2_nor3_1 _15632_ (.A(_08784_),
    .B(_08818_),
    .C(_08854_),
    .Y(_08855_));
 sg13g2_nand3b_1 _15633_ (.B(_08764_),
    .C(_08855_),
    .Y(_08856_),
    .A_N(_08744_));
 sg13g2_nor4_1 _15634_ (.A(_08679_),
    .B(_08699_),
    .C(_08719_),
    .D(_08856_),
    .Y(_08857_));
 sg13g2_nand4_1 _15635_ (.B(_08539_),
    .C(_08656_),
    .A(_08420_),
    .Y(_08858_),
    .D(_08857_));
 sg13g2_buf_1 _15636_ (.A(_08858_),
    .X(_08859_));
 sg13g2_buf_1 _15637_ (.A(_08859_),
    .X(_08860_));
 sg13g2_buf_1 _15638_ (.A(net114),
    .X(_08861_));
 sg13g2_buf_1 _15639_ (.A(\cpu.ex.pc[1] ),
    .X(_08862_));
 sg13g2_buf_1 _15640_ (.A(_08862_),
    .X(_08863_));
 sg13g2_nor2_2 _15641_ (.A(net941),
    .B(net1078),
    .Y(_08864_));
 sg13g2_mux2_1 _15642_ (.A0(\cpu.icache.r_data[4][5] ),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(net936),
    .X(_08865_));
 sg13g2_buf_2 _15643_ (.A(net941),
    .X(_08866_));
 sg13g2_a22oi_1 _15644_ (.Y(_08867_),
    .B1(_08865_),
    .B2(net820),
    .A2(_08864_),
    .A1(\cpu.icache.r_data[5][5] ));
 sg13g2_nand2_1 _15645_ (.Y(_08868_),
    .A(_08465_),
    .B(\cpu.icache.r_data[3][5] ));
 sg13g2_nand2_1 _15646_ (.Y(_08869_),
    .A(net1076),
    .B(\cpu.icache.r_data[7][5] ));
 sg13g2_a21oi_1 _15647_ (.A1(_08868_),
    .A2(_08869_),
    .Y(_08870_),
    .B1(_08522_));
 sg13g2_a221oi_1 _15648_ (.B2(\cpu.icache.r_data[2][5] ),
    .C1(_08870_),
    .B1(net654),
    .A1(\cpu.icache.r_data[1][5] ),
    .Y(_08871_),
    .A2(net655));
 sg13g2_o21ai_1 _15649_ (.B1(_08871_),
    .Y(_08872_),
    .A1(net824),
    .A2(_08867_));
 sg13g2_nand2_1 _15650_ (.Y(_08873_),
    .A(_00207_),
    .B(net720));
 sg13g2_o21ai_1 _15651_ (.B1(_08873_),
    .Y(_08874_),
    .A1(net650),
    .A2(_08872_));
 sg13g2_nor2_1 _15652_ (.A(_00208_),
    .B(net658),
    .Y(_08875_));
 sg13g2_mux2_1 _15653_ (.A0(\cpu.icache.r_data[4][21] ),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(net936),
    .X(_08876_));
 sg13g2_a22oi_1 _15654_ (.Y(_08877_),
    .B1(_08876_),
    .B2(_08475_),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][21] ));
 sg13g2_or2_1 _15655_ (.X(_08878_),
    .B(_08877_),
    .A(_08520_));
 sg13g2_a22oi_1 _15656_ (.Y(_08879_),
    .B1(net653),
    .B2(\cpu.icache.r_data[3][21] ),
    .A2(net654),
    .A1(\cpu.icache.r_data[2][21] ));
 sg13g2_a22oi_1 _15657_ (.Y(_08880_),
    .B1(_08532_),
    .B2(\cpu.icache.r_data[5][21] ),
    .A2(net655),
    .A1(\cpu.icache.r_data[1][21] ));
 sg13g2_nand3_1 _15658_ (.B(_08879_),
    .C(_08880_),
    .A(_08878_),
    .Y(_08881_));
 sg13g2_o21ai_1 _15659_ (.B1(net1074),
    .Y(_08882_),
    .A1(_08875_),
    .A2(_08881_));
 sg13g2_o21ai_1 _15660_ (.B1(_08882_),
    .Y(_08883_),
    .A1(net1074),
    .A2(_08874_));
 sg13g2_buf_2 _15661_ (.A(_08883_),
    .X(_08884_));
 sg13g2_inv_1 _15662_ (.Y(_08885_),
    .A(_08884_));
 sg13g2_buf_1 _15663_ (.A(_08863_),
    .X(_08886_));
 sg13g2_nor2_1 _15664_ (.A(_00210_),
    .B(net658),
    .Y(_08887_));
 sg13g2_buf_1 _15665_ (.A(_08520_),
    .X(_08888_));
 sg13g2_mux2_1 _15666_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(\cpu.icache.r_data[7][22] ),
    .S(net944),
    .X(_08889_));
 sg13g2_nor2b_1 _15667_ (.A(net1160),
    .B_N(_08462_),
    .Y(_08890_));
 sg13g2_buf_2 _15668_ (.A(_08890_),
    .X(_08891_));
 sg13g2_a22oi_1 _15669_ (.Y(_08892_),
    .B1(_08891_),
    .B2(\cpu.icache.r_data[6][22] ),
    .A2(_08889_),
    .A1(net942));
 sg13g2_nor2_1 _15670_ (.A(_08888_),
    .B(_08892_),
    .Y(_08893_));
 sg13g2_a22oi_1 _15671_ (.Y(_08894_),
    .B1(net823),
    .B2(\cpu.icache.r_data[4][22] ),
    .A2(net653),
    .A1(\cpu.icache.r_data[3][22] ));
 sg13g2_a22oi_1 _15672_ (.Y(_08895_),
    .B1(net656),
    .B2(\cpu.icache.r_data[2][22] ),
    .A2(_08478_),
    .A1(\cpu.icache.r_data[1][22] ));
 sg13g2_nand2_1 _15673_ (.Y(_08896_),
    .A(_08894_),
    .B(_08895_));
 sg13g2_nor3_1 _15674_ (.A(_08887_),
    .B(_08893_),
    .C(_08896_),
    .Y(_08897_));
 sg13g2_nand2_1 _15675_ (.Y(_08898_),
    .A(_00209_),
    .B(net720));
 sg13g2_a22oi_1 _15676_ (.Y(_08899_),
    .B1(_08532_),
    .B2(\cpu.icache.r_data[5][6] ),
    .A2(_08478_),
    .A1(\cpu.icache.r_data[1][6] ));
 sg13g2_a22oi_1 _15677_ (.Y(_08900_),
    .B1(net653),
    .B2(\cpu.icache.r_data[3][6] ),
    .A2(_08487_),
    .A1(\cpu.icache.r_data[2][6] ));
 sg13g2_mux2_1 _15678_ (.A0(\cpu.icache.r_data[4][6] ),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(net936),
    .X(_08901_));
 sg13g2_a22oi_1 _15679_ (.Y(_08902_),
    .B1(_08901_),
    .B2(_08866_),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][6] ));
 sg13g2_or2_1 _15680_ (.X(_08903_),
    .B(_08902_),
    .A(net827));
 sg13g2_nand4_1 _15681_ (.B(_08899_),
    .C(_08900_),
    .A(net658),
    .Y(_08904_),
    .D(_08903_));
 sg13g2_a21oi_1 _15682_ (.A1(_08898_),
    .A2(_08904_),
    .Y(_08905_),
    .B1(_08863_));
 sg13g2_a21oi_1 _15683_ (.A1(net935),
    .A2(_08897_),
    .Y(_08906_),
    .B1(_08905_));
 sg13g2_buf_1 _15684_ (.A(_08906_),
    .X(_08907_));
 sg13g2_inv_1 _15685_ (.Y(_08908_),
    .A(net357));
 sg13g2_nand2_1 _15686_ (.Y(_08909_),
    .A(_08885_),
    .B(_08908_));
 sg13g2_nor2_1 _15687_ (.A(_00206_),
    .B(net578),
    .Y(_08910_));
 sg13g2_mux2_1 _15688_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(\cpu.icache.r_data[7][31] ),
    .S(net723),
    .X(_08911_));
 sg13g2_buf_1 _15689_ (.A(_08472_),
    .X(_08912_));
 sg13g2_a22oi_1 _15690_ (.Y(_08913_),
    .B1(_08911_),
    .B2(net718),
    .A2(_08891_),
    .A1(\cpu.icache.r_data[6][31] ));
 sg13g2_nor2_1 _15691_ (.A(net719),
    .B(_08913_),
    .Y(_08914_));
 sg13g2_buf_1 _15692_ (.A(net574),
    .X(_08915_));
 sg13g2_buf_1 _15693_ (.A(net573),
    .X(_08916_));
 sg13g2_a22oi_1 _15694_ (.Y(_08917_),
    .B1(net494),
    .B2(\cpu.icache.r_data[2][31] ),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][31] ));
 sg13g2_a22oi_1 _15695_ (.Y(_08918_),
    .B1(net726),
    .B2(\cpu.icache.r_data[4][31] ),
    .A2(net572),
    .A1(\cpu.icache.r_data[3][31] ));
 sg13g2_nand2_1 _15696_ (.Y(_08919_),
    .A(_08917_),
    .B(_08918_));
 sg13g2_nor3_1 _15697_ (.A(_08910_),
    .B(_08914_),
    .C(_08919_),
    .Y(_08920_));
 sg13g2_nand2_1 _15698_ (.Y(_08921_),
    .A(_00205_),
    .B(net650));
 sg13g2_mux2_1 _15699_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_08569_),
    .X(_08922_));
 sg13g2_a22oi_1 _15700_ (.Y(_08923_),
    .B1(_08922_),
    .B2(net723),
    .A2(net832),
    .A1(\cpu.icache.r_data[5][15] ));
 sg13g2_nand2b_1 _15701_ (.Y(_08924_),
    .B(net718),
    .A_N(_08923_));
 sg13g2_mux2_1 _15702_ (.A0(\cpu.icache.r_data[4][15] ),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(net833),
    .X(_08925_));
 sg13g2_a22oi_1 _15703_ (.Y(_08926_),
    .B1(net830),
    .B2(_08925_),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][15] ));
 sg13g2_nand2_1 _15704_ (.Y(_08927_),
    .A(\cpu.icache.r_data[2][15] ),
    .B(net576));
 sg13g2_nand4_1 _15705_ (.B(_08924_),
    .C(_08926_),
    .A(_08459_),
    .Y(_08928_),
    .D(_08927_));
 sg13g2_a21oi_1 _15706_ (.A1(_08921_),
    .A2(_08928_),
    .Y(_08929_),
    .B1(net935));
 sg13g2_a21o_1 _15707_ (.A2(_08920_),
    .A1(net935),
    .B1(_08929_),
    .X(_08930_));
 sg13g2_buf_1 _15708_ (.A(_08930_),
    .X(_08931_));
 sg13g2_mux2_1 _15709_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(net938),
    .X(_08932_));
 sg13g2_a22oi_1 _15710_ (.Y(_08933_),
    .B1(_08932_),
    .B2(net723),
    .A2(net832),
    .A1(\cpu.icache.r_data[5][29] ));
 sg13g2_nand2b_1 _15711_ (.Y(_08934_),
    .B(net831),
    .A_N(_08933_));
 sg13g2_a22oi_1 _15712_ (.Y(_08935_),
    .B1(_08567_),
    .B2(\cpu.icache.r_data[6][29] ),
    .A2(net573),
    .A1(\cpu.icache.r_data[2][29] ));
 sg13g2_a22oi_1 _15713_ (.Y(_08936_),
    .B1(net726),
    .B2(\cpu.icache.r_data[4][29] ),
    .A2(net577),
    .A1(\cpu.icache.r_data[1][29] ));
 sg13g2_nand3_1 _15714_ (.B(_08935_),
    .C(_08936_),
    .A(_08934_),
    .Y(_08937_));
 sg13g2_a21oi_1 _15715_ (.A1(\cpu.icache.r_data[0][29] ),
    .A2(net650),
    .Y(_08938_),
    .B1(_08937_));
 sg13g2_nand2b_1 _15716_ (.Y(_08939_),
    .B(net650),
    .A_N(\cpu.icache.r_data[0][13] ));
 sg13g2_a22oi_1 _15717_ (.Y(_08940_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][13] ),
    .A2(net577),
    .A1(\cpu.icache.r_data[1][13] ));
 sg13g2_a22oi_1 _15718_ (.Y(_08941_),
    .B1(net572),
    .B2(\cpu.icache.r_data[3][13] ),
    .A2(net573),
    .A1(\cpu.icache.r_data[2][13] ));
 sg13g2_mux2_1 _15719_ (.A0(\cpu.icache.r_data[4][13] ),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(net944),
    .X(_08942_));
 sg13g2_a22oi_1 _15720_ (.Y(_08943_),
    .B1(_08942_),
    .B2(net820),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][13] ));
 sg13g2_or2_1 _15721_ (.X(_08944_),
    .B(_08943_),
    .A(net719));
 sg13g2_nand4_1 _15722_ (.B(_08940_),
    .C(_08941_),
    .A(_08512_),
    .Y(_08945_),
    .D(_08944_));
 sg13g2_a21oi_1 _15723_ (.A1(_08939_),
    .A2(_08945_),
    .Y(_08946_),
    .B1(_08886_));
 sg13g2_a21oi_1 _15724_ (.A1(net935),
    .A2(_08938_),
    .Y(_08947_),
    .B1(_08946_));
 sg13g2_buf_2 _15725_ (.A(_08947_),
    .X(_08948_));
 sg13g2_mux2_1 _15726_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(net938),
    .X(_08949_));
 sg13g2_a22oi_1 _15727_ (.Y(_08950_),
    .B1(_08949_),
    .B2(net723),
    .A2(net832),
    .A1(\cpu.icache.r_data[5][30] ));
 sg13g2_inv_1 _15728_ (.Y(_08951_),
    .A(_08950_));
 sg13g2_mux2_1 _15729_ (.A0(\cpu.icache.r_data[4][30] ),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_08515_),
    .X(_08952_));
 sg13g2_a22oi_1 _15730_ (.Y(_08953_),
    .B1(net940),
    .B2(_08952_),
    .A2(net574),
    .A1(\cpu.icache.r_data[1][30] ));
 sg13g2_inv_1 _15731_ (.Y(_08954_),
    .A(_08953_));
 sg13g2_a221oi_1 _15732_ (.B2(net718),
    .C1(_08954_),
    .B1(_08951_),
    .A1(\cpu.icache.r_data[2][30] ),
    .Y(_08955_),
    .A2(net576));
 sg13g2_o21ai_1 _15733_ (.B1(_08955_),
    .Y(_08956_),
    .A1(_00204_),
    .A2(net579));
 sg13g2_inv_1 _15734_ (.Y(_08957_),
    .A(_08862_));
 sg13g2_buf_1 _15735_ (.A(_08957_),
    .X(_08958_));
 sg13g2_nand2_1 _15736_ (.Y(_08959_),
    .A(_00203_),
    .B(net650));
 sg13g2_mux2_1 _15737_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_08465_),
    .X(_08960_));
 sg13g2_a22oi_1 _15738_ (.Y(_08961_),
    .B1(_08960_),
    .B2(_08624_),
    .A2(_08468_),
    .A1(\cpu.icache.r_data[5][14] ));
 sg13g2_nand2b_1 _15739_ (.Y(_08962_),
    .B(_08472_),
    .A_N(_08961_));
 sg13g2_mux2_1 _15740_ (.A0(\cpu.icache.r_data[4][14] ),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(net833),
    .X(_08963_));
 sg13g2_a22oi_1 _15741_ (.Y(_08964_),
    .B1(net830),
    .B2(_08963_),
    .A2(net577),
    .A1(\cpu.icache.r_data[1][14] ));
 sg13g2_nand2_1 _15742_ (.Y(_08965_),
    .A(\cpu.icache.r_data[2][14] ),
    .B(_08488_));
 sg13g2_nand4_1 _15743_ (.B(_08962_),
    .C(_08964_),
    .A(_08461_),
    .Y(_08966_),
    .D(_08965_));
 sg13g2_and3_1 _15744_ (.X(_08967_),
    .A(net934),
    .B(_08959_),
    .C(_08966_));
 sg13g2_a21o_1 _15745_ (.A2(_08956_),
    .A1(net935),
    .B1(_08967_),
    .X(_08968_));
 sg13g2_buf_1 _15746_ (.A(_08968_),
    .X(_08969_));
 sg13g2_nor3_1 _15747_ (.A(_08931_),
    .B(_08948_),
    .C(net263),
    .Y(_08970_));
 sg13g2_buf_2 _15748_ (.A(_08970_),
    .X(_08971_));
 sg13g2_buf_1 _15749_ (.A(_08886_),
    .X(_08972_));
 sg13g2_nand2_1 _15750_ (.Y(_08973_),
    .A(\cpu.icache.r_data[0][16] ),
    .B(net650));
 sg13g2_mux2_1 _15751_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(net719),
    .X(_08974_));
 sg13g2_a22oi_1 _15752_ (.Y(_08975_),
    .B1(_08974_),
    .B2(net649),
    .A2(_08468_),
    .A1(\cpu.icache.r_data[5][16] ));
 sg13g2_nand2b_1 _15753_ (.Y(_08976_),
    .B(net718),
    .A_N(_08975_));
 sg13g2_nand2_1 _15754_ (.Y(_08977_),
    .A(\cpu.icache.r_data[2][16] ),
    .B(_08916_));
 sg13g2_mux2_1 _15755_ (.A0(\cpu.icache.r_data[4][16] ),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(net649),
    .X(_08978_));
 sg13g2_a22oi_1 _15756_ (.Y(_08979_),
    .B1(_08482_),
    .B2(_08978_),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][16] ));
 sg13g2_nand4_1 _15757_ (.B(_08976_),
    .C(_08977_),
    .A(_08973_),
    .Y(_08980_),
    .D(_08979_));
 sg13g2_mux2_1 _15758_ (.A0(\cpu.icache.r_data[4][0] ),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_08464_),
    .X(_08981_));
 sg13g2_a22oi_1 _15759_ (.Y(_08982_),
    .B1(_08981_),
    .B2(net820),
    .A2(_08864_),
    .A1(\cpu.icache.r_data[5][0] ));
 sg13g2_mux2_1 _15760_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(net824),
    .X(_08983_));
 sg13g2_a22oi_1 _15761_ (.Y(_08984_),
    .B1(net822),
    .B2(_08983_),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[1][0] ));
 sg13g2_o21ai_1 _15762_ (.B1(_08984_),
    .Y(_08985_),
    .A1(net719),
    .A2(_08982_));
 sg13g2_a21oi_1 _15763_ (.A1(\cpu.icache.r_data[2][0] ),
    .A2(net494),
    .Y(_08986_),
    .B1(_08985_));
 sg13g2_nand2_1 _15764_ (.Y(_08987_),
    .A(net497),
    .B(_08986_));
 sg13g2_o21ai_1 _15765_ (.B1(_08987_),
    .Y(_08988_),
    .A1(\cpu.icache.r_data[0][0] ),
    .A2(net497));
 sg13g2_nor2_1 _15766_ (.A(net819),
    .B(_08988_),
    .Y(_08989_));
 sg13g2_a21oi_1 _15767_ (.A1(net819),
    .A2(_08980_),
    .Y(_08990_),
    .B1(_08989_));
 sg13g2_buf_1 _15768_ (.A(_08990_),
    .X(_08991_));
 sg13g2_mux2_1 _15769_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(net824),
    .X(_08992_));
 sg13g2_a22oi_1 _15770_ (.Y(_08993_),
    .B1(_08992_),
    .B2(net831),
    .A2(_08482_),
    .A1(\cpu.icache.r_data[6][17] ));
 sg13g2_nand2b_1 _15771_ (.Y(_08994_),
    .B(net649),
    .A_N(_08993_));
 sg13g2_a22oi_1 _15772_ (.Y(_08995_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][17] ),
    .A2(net494),
    .A1(\cpu.icache.r_data[2][17] ));
 sg13g2_a22oi_1 _15773_ (.Y(_08996_),
    .B1(net726),
    .B2(\cpu.icache.r_data[4][17] ),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][17] ));
 sg13g2_nand3_1 _15774_ (.B(_08995_),
    .C(_08996_),
    .A(_08994_),
    .Y(_08997_));
 sg13g2_a21oi_1 _15775_ (.A1(\cpu.icache.r_data[0][17] ),
    .A2(net650),
    .Y(_08998_),
    .B1(_08997_));
 sg13g2_a22oi_1 _15776_ (.Y(_08999_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][1] ),
    .A2(_08915_),
    .A1(\cpu.icache.r_data[1][1] ));
 sg13g2_a22oi_1 _15777_ (.Y(_09000_),
    .B1(net572),
    .B2(\cpu.icache.r_data[3][1] ),
    .A2(net494),
    .A1(\cpu.icache.r_data[2][1] ));
 sg13g2_mux2_1 _15778_ (.A0(\cpu.icache.r_data[4][1] ),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_08515_),
    .X(_09001_));
 sg13g2_a22oi_1 _15779_ (.Y(_09002_),
    .B1(_09001_),
    .B2(net820),
    .A2(_08598_),
    .A1(\cpu.icache.r_data[7][1] ));
 sg13g2_or2_1 _15780_ (.X(_09003_),
    .B(_09002_),
    .A(net719));
 sg13g2_nand4_1 _15781_ (.B(_08999_),
    .C(_09000_),
    .A(_08459_),
    .Y(_09004_),
    .D(_09003_));
 sg13g2_o21ai_1 _15782_ (.B1(_09004_),
    .Y(_09005_),
    .A1(\cpu.icache.r_data[0][1] ),
    .A2(_08713_));
 sg13g2_mux2_1 _15783_ (.A0(_08998_),
    .A1(_09005_),
    .S(net934),
    .X(_09006_));
 sg13g2_buf_1 _15784_ (.A(_09006_),
    .X(_09007_));
 sg13g2_inv_1 _15785_ (.Y(_09008_),
    .A(_09007_));
 sg13g2_buf_1 _15786_ (.A(_09008_),
    .X(_09009_));
 sg13g2_nor2_1 _15787_ (.A(_08991_),
    .B(net210),
    .Y(_09010_));
 sg13g2_buf_1 _15788_ (.A(_09010_),
    .X(_09011_));
 sg13g2_nand2_1 _15789_ (.Y(_09012_),
    .A(_08971_),
    .B(_09011_));
 sg13g2_buf_1 _15790_ (.A(_09012_),
    .X(_09013_));
 sg13g2_nand2b_1 _15791_ (.Y(_09014_),
    .B(net720),
    .A_N(_00202_));
 sg13g2_mux2_1 _15792_ (.A0(\cpu.icache.r_data[5][27] ),
    .A1(\cpu.icache.r_data[7][27] ),
    .S(net1078),
    .X(_09015_));
 sg13g2_a22oi_1 _15793_ (.Y(_09016_),
    .B1(_09015_),
    .B2(net1077),
    .A2(_08572_),
    .A1(\cpu.icache.r_data[4][27] ));
 sg13g2_or2_1 _15794_ (.X(_09017_),
    .B(_09016_),
    .A(net938));
 sg13g2_a22oi_1 _15795_ (.Y(_09018_),
    .B1(_08566_),
    .B2(\cpu.icache.r_data[6][27] ),
    .A2(net654),
    .A1(\cpu.icache.r_data[2][27] ));
 sg13g2_a22oi_1 _15796_ (.Y(_09019_),
    .B1(net653),
    .B2(\cpu.icache.r_data[3][27] ),
    .A2(net655),
    .A1(\cpu.icache.r_data[1][27] ));
 sg13g2_nand4_1 _15797_ (.B(_09017_),
    .C(_09018_),
    .A(_09014_),
    .Y(_09020_),
    .D(_09019_));
 sg13g2_mux2_1 _15798_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(net1078),
    .X(_09021_));
 sg13g2_a22oi_1 _15799_ (.Y(_09022_),
    .B1(_09021_),
    .B2(net941),
    .A2(_08864_),
    .A1(\cpu.icache.r_data[5][11] ));
 sg13g2_nand2_1 _15800_ (.Y(_09023_),
    .A(_08448_),
    .B(\cpu.icache.r_data[3][11] ));
 sg13g2_nand2_1 _15801_ (.Y(_09024_),
    .A(net1076),
    .B(\cpu.icache.r_data[7][11] ));
 sg13g2_a21oi_1 _15802_ (.A1(_09023_),
    .A2(_09024_),
    .Y(_09025_),
    .B1(_08522_));
 sg13g2_a221oi_1 _15803_ (.B2(\cpu.icache.r_data[2][11] ),
    .C1(_09025_),
    .B1(_08486_),
    .A1(\cpu.icache.r_data[1][11] ),
    .Y(_09026_),
    .A2(_08477_));
 sg13g2_o21ai_1 _15804_ (.B1(_09026_),
    .Y(_09027_),
    .A1(net938),
    .A2(_09022_));
 sg13g2_nand2_1 _15805_ (.Y(_09028_),
    .A(_00201_),
    .B(net720));
 sg13g2_o21ai_1 _15806_ (.B1(_09028_),
    .Y(_09029_),
    .A1(net720),
    .A2(_09027_));
 sg13g2_nor2_1 _15807_ (.A(_08862_),
    .B(_09029_),
    .Y(_09030_));
 sg13g2_a21oi_1 _15808_ (.A1(net1074),
    .A2(_09020_),
    .Y(_09031_),
    .B1(_09030_));
 sg13g2_buf_1 _15809_ (.A(_09031_),
    .X(_09032_));
 sg13g2_nor2_1 _15810_ (.A(_00200_),
    .B(net734),
    .Y(_09033_));
 sg13g2_mux2_1 _15811_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(\cpu.icache.r_data[7][26] ),
    .S(_08788_),
    .X(_09034_));
 sg13g2_a22oi_1 _15812_ (.Y(_09035_),
    .B1(_09034_),
    .B2(net1077),
    .A2(_08572_),
    .A1(\cpu.icache.r_data[4][26] ));
 sg13g2_nor2_1 _15813_ (.A(net827),
    .B(_09035_),
    .Y(_09036_));
 sg13g2_a22oi_1 _15814_ (.Y(_09037_),
    .B1(net654),
    .B2(\cpu.icache.r_data[2][26] ),
    .A2(net655),
    .A1(\cpu.icache.r_data[1][26] ));
 sg13g2_a22oi_1 _15815_ (.Y(_09038_),
    .B1(_08566_),
    .B2(\cpu.icache.r_data[6][26] ),
    .A2(_08527_),
    .A1(\cpu.icache.r_data[3][26] ));
 sg13g2_nand2_1 _15816_ (.Y(_09039_),
    .A(_09037_),
    .B(_09038_));
 sg13g2_nor4_1 _15817_ (.A(_08957_),
    .B(_09033_),
    .C(_09036_),
    .D(_09039_),
    .Y(_09040_));
 sg13g2_nand2_1 _15818_ (.Y(_09041_),
    .A(_00199_),
    .B(net720));
 sg13g2_a22oi_1 _15819_ (.Y(_09042_),
    .B1(_08531_),
    .B2(\cpu.icache.r_data[5][10] ),
    .A2(_08477_),
    .A1(\cpu.icache.r_data[1][10] ));
 sg13g2_a22oi_1 _15820_ (.Y(_09043_),
    .B1(_08592_),
    .B2(\cpu.icache.r_data[4][10] ),
    .A2(_08486_),
    .A1(\cpu.icache.r_data[2][10] ));
 sg13g2_mux2_1 _15821_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(\cpu.icache.r_data[3][10] ),
    .S(_08448_),
    .X(_09044_));
 sg13g2_a22oi_1 _15822_ (.Y(_09045_),
    .B1(_09044_),
    .B2(net1077),
    .A2(net940),
    .A1(\cpu.icache.r_data[6][10] ));
 sg13g2_nand2b_1 _15823_ (.Y(_09046_),
    .B(_08463_),
    .A_N(_09045_));
 sg13g2_nand4_1 _15824_ (.B(_09042_),
    .C(_09043_),
    .A(net734),
    .Y(_09047_),
    .D(_09046_));
 sg13g2_a21oi_1 _15825_ (.A1(_09041_),
    .A2(_09047_),
    .Y(_09048_),
    .B1(net1074));
 sg13g2_or2_1 _15826_ (.X(_09049_),
    .B(_09048_),
    .A(_09040_));
 sg13g2_buf_1 _15827_ (.A(_09049_),
    .X(_09050_));
 sg13g2_nor2_1 _15828_ (.A(_09032_),
    .B(net355),
    .Y(_09051_));
 sg13g2_inv_1 _15829_ (.Y(_09052_),
    .A(_09051_));
 sg13g2_nor4_1 _15830_ (.A(net114),
    .B(_08909_),
    .C(_09013_),
    .D(_09052_),
    .Y(_09053_));
 sg13g2_a21o_1 _15831_ (.A2(net95),
    .A1(_08244_),
    .B1(_09053_),
    .X(_00017_));
 sg13g2_buf_1 _15832_ (.A(\cpu.dec.r_op[4] ),
    .X(_09054_));
 sg13g2_buf_1 _15833_ (.A(_09054_),
    .X(_09055_));
 sg13g2_buf_1 _15834_ (.A(_08859_),
    .X(_09056_));
 sg13g2_a22oi_1 _15835_ (.Y(_09057_),
    .B1(_08566_),
    .B2(\cpu.icache.r_data[6][12] ),
    .A2(_08486_),
    .A1(\cpu.icache.r_data[2][12] ));
 sg13g2_a22oi_1 _15836_ (.Y(_09058_),
    .B1(_08527_),
    .B2(\cpu.icache.r_data[3][12] ),
    .A2(_08477_),
    .A1(\cpu.icache.r_data[1][12] ));
 sg13g2_mux2_1 _15837_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(\cpu.icache.r_data[7][12] ),
    .S(_08452_),
    .X(_09059_));
 sg13g2_a22oi_1 _15838_ (.Y(_09060_),
    .B1(_09059_),
    .B2(net1077),
    .A2(_08572_),
    .A1(\cpu.icache.r_data[4][12] ));
 sg13g2_or2_1 _15839_ (.X(_09061_),
    .B(_09060_),
    .A(net943));
 sg13g2_and4_1 _15840_ (.A(_08457_),
    .B(_09057_),
    .C(_09058_),
    .D(_09061_),
    .X(_09062_));
 sg13g2_a21oi_1 _15841_ (.A1(_00211_),
    .A2(net720),
    .Y(_09063_),
    .B1(_09062_));
 sg13g2_nor2_1 _15842_ (.A(_00212_),
    .B(_08457_),
    .Y(_09064_));
 sg13g2_mux2_1 _15843_ (.A0(\cpu.icache.r_data[4][28] ),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_08788_),
    .X(_09065_));
 sg13g2_a22oi_1 _15844_ (.Y(_09066_),
    .B1(_09065_),
    .B2(_08475_),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][28] ));
 sg13g2_nor2_1 _15845_ (.A(net827),
    .B(_09066_),
    .Y(_09067_));
 sg13g2_a22oi_1 _15846_ (.Y(_09068_),
    .B1(_08486_),
    .B2(\cpu.icache.r_data[2][28] ),
    .A2(_08477_),
    .A1(\cpu.icache.r_data[1][28] ));
 sg13g2_a22oi_1 _15847_ (.Y(_09069_),
    .B1(_08531_),
    .B2(\cpu.icache.r_data[5][28] ),
    .A2(_08527_),
    .A1(\cpu.icache.r_data[3][28] ));
 sg13g2_nand2_1 _15848_ (.Y(_09070_),
    .A(_09068_),
    .B(_09069_));
 sg13g2_or4_1 _15849_ (.A(_08957_),
    .B(_09064_),
    .C(_09067_),
    .D(_09070_),
    .X(_09071_));
 sg13g2_o21ai_1 _15850_ (.B1(_09071_),
    .Y(_09072_),
    .A1(net1074),
    .A2(_09063_));
 sg13g2_buf_1 _15851_ (.A(_09072_),
    .X(_09073_));
 sg13g2_buf_1 _15852_ (.A(_09073_),
    .X(_09074_));
 sg13g2_buf_1 _15853_ (.A(_09007_),
    .X(_09075_));
 sg13g2_nor2_1 _15854_ (.A(_08991_),
    .B(_09075_),
    .Y(_09076_));
 sg13g2_buf_2 _15855_ (.A(_09076_),
    .X(_09077_));
 sg13g2_nand3_1 _15856_ (.B(_09051_),
    .C(_09077_),
    .A(_08971_),
    .Y(_09078_));
 sg13g2_buf_1 _15857_ (.A(_09078_),
    .X(_09079_));
 sg13g2_or2_1 _15858_ (.X(_09080_),
    .B(_09079_),
    .A(_08909_));
 sg13g2_nor3_1 _15859_ (.A(net113),
    .B(net354),
    .C(_09080_),
    .Y(_09081_));
 sg13g2_a21o_1 _15860_ (.A2(net95),
    .A1(_09055_),
    .B1(_09081_),
    .X(_00015_));
 sg13g2_buf_1 _15861_ (.A(\cpu.dec.r_op[5] ),
    .X(_09082_));
 sg13g2_inv_1 _15862_ (.Y(_09083_),
    .A(_09032_));
 sg13g2_nor4_1 _15863_ (.A(net114),
    .B(_09013_),
    .C(_09083_),
    .D(net355),
    .Y(_09084_));
 sg13g2_a21o_1 _15864_ (.A2(net95),
    .A1(_09082_),
    .B1(_09084_),
    .X(_00016_));
 sg13g2_buf_1 _15865_ (.A(\cpu.dec.r_op[7] ),
    .X(_09085_));
 sg13g2_nand2_1 _15866_ (.Y(_09086_),
    .A(_08884_),
    .B(net357));
 sg13g2_nor3_1 _15867_ (.A(net113),
    .B(_09079_),
    .C(_09086_),
    .Y(_09087_));
 sg13g2_a21o_1 _15868_ (.A2(net95),
    .A1(_09085_),
    .B1(_09087_),
    .X(_00018_));
 sg13g2_nand2_1 _15869_ (.Y(_09088_),
    .A(_09051_),
    .B(net354));
 sg13g2_buf_1 _15870_ (.A(_08884_),
    .X(_09089_));
 sg13g2_nand2_1 _15871_ (.Y(_09090_),
    .A(_09089_),
    .B(_08908_));
 sg13g2_nor3_1 _15872_ (.A(_09013_),
    .B(_09088_),
    .C(_09090_),
    .Y(_09091_));
 sg13g2_buf_2 _15873_ (.A(\cpu.dec.r_op[3] ),
    .X(_09092_));
 sg13g2_buf_1 _15874_ (.A(_09092_),
    .X(_09093_));
 sg13g2_buf_1 _15875_ (.A(net114),
    .X(_09094_));
 sg13g2_mux2_1 _15876_ (.A0(_09091_),
    .A1(_09093_),
    .S(net94),
    .X(_00014_));
 sg13g2_buf_1 _15877_ (.A(net114),
    .X(_09095_));
 sg13g2_buf_1 _15878_ (.A(_08971_),
    .X(_09096_));
 sg13g2_nand2_1 _15879_ (.Y(_09097_),
    .A(_09083_),
    .B(net355));
 sg13g2_o21ai_1 _15880_ (.B1(_09097_),
    .Y(_09098_),
    .A1(_09086_),
    .A2(_09088_));
 sg13g2_nand3_1 _15881_ (.B(_09011_),
    .C(_09098_),
    .A(_09096_),
    .Y(_09099_));
 sg13g2_buf_1 _15882_ (.A(\cpu.dec.r_op[2] ),
    .X(_09100_));
 sg13g2_buf_1 _15883_ (.A(_08859_),
    .X(_09101_));
 sg13g2_nand2_1 _15884_ (.Y(_09102_),
    .A(_09100_),
    .B(_09101_));
 sg13g2_o21ai_1 _15885_ (.B1(_09102_),
    .Y(_00013_),
    .A1(_09095_),
    .A2(_09099_));
 sg13g2_nor2b_1 _15886_ (.A(r_reset),
    .B_N(net1),
    .Y(_09103_));
 sg13g2_buf_1 _15887_ (.A(_09103_),
    .X(_09104_));
 sg13g2_buf_1 _15888_ (.A(net1071),
    .X(_09105_));
 sg13g2_buf_1 _15889_ (.A(net933),
    .X(_09106_));
 sg13g2_buf_2 _15890_ (.A(net818),
    .X(_09107_));
 sg13g2_inv_2 _15891_ (.Y(_09108_),
    .A(_08299_));
 sg13g2_nor3_2 _15892_ (.A(_09108_),
    .B(_08359_),
    .C(_08415_),
    .Y(_09109_));
 sg13g2_buf_2 _15893_ (.A(\cpu.dec.r_trap ),
    .X(_09110_));
 sg13g2_nand2_1 _15894_ (.Y(_09111_),
    .A(\cpu.intr.r_clock ),
    .B(\cpu.intr.r_enable[1] ));
 sg13g2_buf_2 _15895_ (.A(\cpu.intr.r_timer ),
    .X(_09112_));
 sg13g2_nand2_1 _15896_ (.Y(_09113_),
    .A(_09112_),
    .B(\cpu.intr.r_enable[2] ));
 sg13g2_buf_1 _15897_ (.A(\cpu.uart.r_x_int ),
    .X(_09114_));
 sg13g2_buf_1 _15898_ (.A(\cpu.uart.r_r_int ),
    .X(_09115_));
 sg13g2_buf_1 _15899_ (.A(\cpu.intr.r_enable[0] ),
    .X(_09116_));
 sg13g2_o21ai_1 _15900_ (.B1(_09116_),
    .Y(_09117_),
    .A1(_09114_),
    .A2(_09115_));
 sg13g2_buf_1 _15901_ (.A(\cpu.intr.r_swi ),
    .X(_09118_));
 sg13g2_buf_2 _15902_ (.A(\cpu.intr.spi_intr ),
    .X(_09119_));
 sg13g2_buf_2 _15903_ (.A(\cpu.intr.r_enable[5] ),
    .X(_09120_));
 sg13g2_a22oi_1 _15904_ (.Y(_09121_),
    .B1(_09119_),
    .B2(_09120_),
    .A2(_09118_),
    .A1(\cpu.intr.r_enable[3] ));
 sg13g2_and4_1 _15905_ (.A(_09111_),
    .B(_09113_),
    .C(_09117_),
    .D(_09121_),
    .X(_09122_));
 sg13g2_buf_8 _15906_ (.A(_09122_),
    .X(_09123_));
 sg13g2_inv_1 _15907_ (.Y(_09124_),
    .A(_09123_));
 sg13g2_buf_1 _15908_ (.A(\cpu.gpio.r_enable_in[1] ),
    .X(_09125_));
 sg13g2_buf_2 _15909_ (.A(ui_in[1]),
    .X(_09126_));
 sg13g2_buf_1 _15910_ (.A(\cpu.gpio.r_enable_in[5] ),
    .X(_09127_));
 sg13g2_buf_2 _15911_ (.A(ui_in[5]),
    .X(_09128_));
 sg13g2_a22oi_1 _15912_ (.Y(_09129_),
    .B1(_09127_),
    .B2(_09128_),
    .A2(_09126_),
    .A1(_09125_));
 sg13g2_buf_1 _15913_ (.A(\cpu.gpio.r_enable_io[6] ),
    .X(_09130_));
 sg13g2_buf_1 _15914_ (.A(uio_in[6]),
    .X(_09131_));
 sg13g2_buf_2 _15915_ (.A(uio_in[7]),
    .X(_09132_));
 sg13g2_a22oi_1 _15916_ (.Y(_09133_),
    .B1(\cpu.gpio.r_enable_io[7] ),
    .B2(_09132_),
    .A2(_09131_),
    .A1(_09130_));
 sg13g2_and2_1 _15917_ (.A(_09129_),
    .B(_09133_),
    .X(_09134_));
 sg13g2_buf_1 _15918_ (.A(_09134_),
    .X(_09135_));
 sg13g2_buf_1 _15919_ (.A(\cpu.gpio.r_enable_in[2] ),
    .X(_09136_));
 sg13g2_buf_1 _15920_ (.A(ui_in[2]),
    .X(_09137_));
 sg13g2_buf_2 _15921_ (.A(\cpu.gpio.r_enable_in[7] ),
    .X(_09138_));
 sg13g2_buf_2 _15922_ (.A(ui_in[7]),
    .X(_09139_));
 sg13g2_a22oi_1 _15923_ (.Y(_09140_),
    .B1(_09138_),
    .B2(_09139_),
    .A2(_09137_),
    .A1(_09136_));
 sg13g2_buf_1 _15924_ (.A(uio_in[4]),
    .X(_09141_));
 sg13g2_buf_1 _15925_ (.A(uio_in[5]),
    .X(_09142_));
 sg13g2_a22oi_1 _15926_ (.Y(_09143_),
    .B1(\cpu.gpio.r_enable_io[5] ),
    .B2(_09142_),
    .A2(_09141_),
    .A1(\cpu.gpio.r_enable_io[4] ));
 sg13g2_buf_1 _15927_ (.A(\cpu.gpio.r_enable_in[3] ),
    .X(_09144_));
 sg13g2_buf_8 _15928_ (.A(ui_in[3]),
    .X(_09145_));
 sg13g2_buf_1 _15929_ (.A(\cpu.gpio.r_enable_in[4] ),
    .X(_09146_));
 sg13g2_buf_2 _15930_ (.A(ui_in[4]),
    .X(_09147_));
 sg13g2_a22oi_1 _15931_ (.Y(_09148_),
    .B1(_09146_),
    .B2(_09147_),
    .A2(_09145_),
    .A1(_09144_));
 sg13g2_buf_8 _15932_ (.A(ui_in[0]),
    .X(_09149_));
 sg13g2_buf_1 _15933_ (.A(\cpu.gpio.r_enable_in[6] ),
    .X(_09150_));
 sg13g2_buf_2 _15934_ (.A(ui_in[6]),
    .X(_09151_));
 sg13g2_a22oi_1 _15935_ (.Y(_09152_),
    .B1(_09150_),
    .B2(_09151_),
    .A2(_09149_),
    .A1(\cpu.gpio.r_enable_in[0] ));
 sg13g2_and4_1 _15936_ (.A(_09140_),
    .B(_09143_),
    .C(_09148_),
    .D(_09152_),
    .X(_09153_));
 sg13g2_buf_1 _15937_ (.A(_09153_),
    .X(_09154_));
 sg13g2_buf_1 _15938_ (.A(\cpu.intr.r_enable[4] ),
    .X(_09155_));
 sg13g2_inv_1 _15939_ (.Y(_09156_),
    .A(_09155_));
 sg13g2_a21oi_1 _15940_ (.A1(_09135_),
    .A2(_09154_),
    .Y(_09157_),
    .B1(_09156_));
 sg13g2_buf_2 _15941_ (.A(\cpu.ex.r_ie ),
    .X(_09158_));
 sg13g2_o21ai_1 _15942_ (.B1(_09158_),
    .Y(_09159_),
    .A1(_09124_),
    .A2(_09157_));
 sg13g2_buf_1 _15943_ (.A(_09159_),
    .X(_09160_));
 sg13g2_nor2_1 _15944_ (.A(_08437_),
    .B(_09160_),
    .Y(_09161_));
 sg13g2_nor2_2 _15945_ (.A(_09110_),
    .B(_09161_),
    .Y(_09162_));
 sg13g2_nand2_2 _15946_ (.Y(_09163_),
    .A(_09109_),
    .B(_09162_));
 sg13g2_buf_2 _15947_ (.A(\cpu.addr[6] ),
    .X(_09164_));
 sg13g2_buf_4 _15948_ (.X(_09165_),
    .A(\cpu.addr[8] ));
 sg13g2_buf_1 _15949_ (.A(\cpu.addr[7] ),
    .X(_09166_));
 sg13g2_inv_2 _15950_ (.Y(_09167_),
    .A(net1154));
 sg13g2_nor2_1 _15951_ (.A(_09165_),
    .B(_09167_),
    .Y(_09168_));
 sg13g2_and2_1 _15952_ (.A(_09164_),
    .B(_09168_),
    .X(_09169_));
 sg13g2_buf_1 _15953_ (.A(_09169_),
    .X(_09170_));
 sg13g2_buf_1 _15954_ (.A(_00215_),
    .X(_09171_));
 sg13g2_buf_1 _15955_ (.A(\cpu.addr[2] ),
    .X(_09172_));
 sg13g2_buf_1 _15956_ (.A(_09172_),
    .X(_09173_));
 sg13g2_buf_1 _15957_ (.A(_09173_),
    .X(_09174_));
 sg13g2_buf_2 _15958_ (.A(net932),
    .X(_09175_));
 sg13g2_buf_1 _15959_ (.A(net817),
    .X(_09176_));
 sg13g2_buf_2 _15960_ (.A(\cpu.addr[1] ),
    .X(_09177_));
 sg13g2_buf_1 _15961_ (.A(_09177_),
    .X(_09178_));
 sg13g2_buf_1 _15962_ (.A(net1069),
    .X(_09179_));
 sg13g2_nor2_1 _15963_ (.A(net716),
    .B(net931),
    .Y(_09180_));
 sg13g2_buf_2 _15964_ (.A(_09180_),
    .X(_09181_));
 sg13g2_and2_1 _15965_ (.A(_09171_),
    .B(_09181_),
    .X(_09182_));
 sg13g2_buf_1 _15966_ (.A(_09182_),
    .X(_09183_));
 sg13g2_nand2_1 _15967_ (.Y(_09184_),
    .A(_09170_),
    .B(_09183_));
 sg13g2_nor4_2 _15968_ (.A(_00195_),
    .B(_08383_),
    .C(_09163_),
    .Y(_09185_),
    .D(_09184_));
 sg13g2_buf_2 _15969_ (.A(\cpu.addr[3] ),
    .X(_09186_));
 sg13g2_buf_2 _15970_ (.A(_09186_),
    .X(_09187_));
 sg13g2_buf_8 _15971_ (.A(net1068),
    .X(_09188_));
 sg13g2_buf_8 _15972_ (.A(net930),
    .X(_09189_));
 sg13g2_buf_2 _15973_ (.A(net816),
    .X(_09190_));
 sg13g2_buf_1 _15974_ (.A(net715),
    .X(_09191_));
 sg13g2_buf_1 _15975_ (.A(net648),
    .X(_09192_));
 sg13g2_buf_1 _15976_ (.A(net569),
    .X(_09193_));
 sg13g2_inv_1 _15977_ (.Y(_09194_),
    .A(net1166));
 sg13g2_nor3_2 _15978_ (.A(net1067),
    .B(_08355_),
    .C(_09163_),
    .Y(_09195_));
 sg13g2_and2_1 _15979_ (.A(_09170_),
    .B(_09195_),
    .X(_09196_));
 sg13g2_buf_1 _15980_ (.A(_09196_),
    .X(_09197_));
 sg13g2_nor2b_1 _15981_ (.A(net493),
    .B_N(_09197_),
    .Y(_09198_));
 sg13g2_buf_1 _15982_ (.A(_09198_),
    .X(_09199_));
 sg13g2_buf_1 _15983_ (.A(\cpu.spi.r_state[1] ),
    .X(_09200_));
 sg13g2_nand2b_1 _15984_ (.Y(_09201_),
    .B(net1152),
    .A_N(_09199_));
 sg13g2_buf_2 _15985_ (.A(_09201_),
    .X(_09202_));
 sg13g2_buf_1 _15986_ (.A(\cpu.spi.r_state[6] ),
    .X(_09203_));
 sg13g2_buf_1 _15987_ (.A(\cpu.spi.r_bits[0] ),
    .X(_09204_));
 sg13g2_buf_1 _15988_ (.A(\cpu.spi.r_bits[1] ),
    .X(_09205_));
 sg13g2_nor3_1 _15989_ (.A(_09204_),
    .B(_09205_),
    .C(\cpu.spi.r_bits[2] ),
    .Y(_09206_));
 sg13g2_nor3_2 _15990_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .C(\cpu.spi.r_timeout_count[2] ),
    .Y(_09207_));
 sg13g2_nor2b_1 _15991_ (.A(\cpu.spi.r_timeout_count[3] ),
    .B_N(_09207_),
    .Y(_09208_));
 sg13g2_nand2b_1 _15992_ (.Y(_09209_),
    .B(_09208_),
    .A_N(\cpu.spi.r_timeout_count[4] ));
 sg13g2_nor2_1 _15993_ (.A(\cpu.spi.r_timeout_count[5] ),
    .B(_09209_),
    .Y(_09210_));
 sg13g2_nand2b_1 _15994_ (.Y(_09211_),
    .B(_09210_),
    .A_N(\cpu.spi.r_timeout_count[6] ));
 sg13g2_buf_1 _15995_ (.A(_09211_),
    .X(_09212_));
 sg13g2_o21ai_1 _15996_ (.B1(\cpu.spi.r_searching ),
    .Y(_09213_),
    .A1(\cpu.spi.r_timeout_count[7] ),
    .A2(_09212_));
 sg13g2_nand2_1 _15997_ (.Y(_09214_),
    .A(_09206_),
    .B(_09213_));
 sg13g2_buf_1 _15998_ (.A(\cpu.spi.r_in[3] ),
    .X(_09215_));
 sg13g2_buf_1 _15999_ (.A(\cpu.spi.r_in[1] ),
    .X(_09216_));
 sg13g2_buf_1 _16000_ (.A(\cpu.spi.r_in[0] ),
    .X(_09217_));
 sg13g2_nand2_1 _16001_ (.Y(_09218_),
    .A(_09216_),
    .B(_09217_));
 sg13g2_nand3_1 _16002_ (.B(\cpu.spi.r_in[7] ),
    .C(_09218_),
    .A(_09215_),
    .Y(_09219_));
 sg13g2_buf_1 _16003_ (.A(\cpu.spi.r_in[2] ),
    .X(_09220_));
 sg13g2_buf_1 _16004_ (.A(\cpu.spi.r_in[5] ),
    .X(_09221_));
 sg13g2_buf_1 _16005_ (.A(\cpu.spi.r_in[4] ),
    .X(_09222_));
 sg13g2_buf_1 _16006_ (.A(\cpu.spi.r_in[6] ),
    .X(_09223_));
 sg13g2_nand4_1 _16007_ (.B(_09221_),
    .C(_09222_),
    .A(_09220_),
    .Y(_09224_),
    .D(_09223_));
 sg13g2_nor2_1 _16008_ (.A(_09219_),
    .B(_09224_),
    .Y(_09225_));
 sg13g2_o21ai_1 _16009_ (.B1(\cpu.spi.r_searching ),
    .Y(_09226_),
    .A1(_00214_),
    .A2(_09225_));
 sg13g2_nand2_2 _16010_ (.Y(_09227_),
    .A(_09214_),
    .B(_09226_));
 sg13g2_buf_1 _16011_ (.A(\cpu.spi.r_count[7] ),
    .X(_09228_));
 sg13g2_buf_1 _16012_ (.A(\cpu.spi.r_count[2] ),
    .X(_09229_));
 sg13g2_buf_1 _16013_ (.A(\cpu.spi.r_count[0] ),
    .X(_09230_));
 sg13g2_or2_1 _16014_ (.X(_09231_),
    .B(\cpu.spi.r_count[1] ),
    .A(_09230_));
 sg13g2_buf_1 _16015_ (.A(_09231_),
    .X(_09232_));
 sg13g2_nor3_1 _16016_ (.A(_09229_),
    .B(\cpu.spi.r_count[3] ),
    .C(_09232_),
    .Y(_09233_));
 sg13g2_nor2b_1 _16017_ (.A(\cpu.spi.r_count[4] ),
    .B_N(_09233_),
    .Y(_09234_));
 sg13g2_nor2b_1 _16018_ (.A(\cpu.spi.r_count[5] ),
    .B_N(_09234_),
    .Y(_09235_));
 sg13g2_nor2b_1 _16019_ (.A(\cpu.spi.r_count[6] ),
    .B_N(_09235_),
    .Y(_09236_));
 sg13g2_buf_1 _16020_ (.A(_09236_),
    .X(_09237_));
 sg13g2_nor2b_1 _16021_ (.A(_09228_),
    .B_N(_09237_),
    .Y(_09238_));
 sg13g2_buf_1 _16022_ (.A(_09238_),
    .X(_09239_));
 sg13g2_buf_1 _16023_ (.A(_09239_),
    .X(_09240_));
 sg13g2_nand3_1 _16024_ (.B(_09227_),
    .C(net353),
    .A(net1151),
    .Y(_09241_));
 sg13g2_o21ai_1 _16025_ (.B1(_09241_),
    .Y(_09242_),
    .A1(_09185_),
    .A2(_09202_));
 sg13g2_and2_1 _16026_ (.A(net717),
    .B(_09242_),
    .X(_00030_));
 sg13g2_buf_1 _16027_ (.A(net1152),
    .X(_09243_));
 sg13g2_buf_1 _16028_ (.A(_09199_),
    .X(_09244_));
 sg13g2_buf_1 _16029_ (.A(net157),
    .X(_09245_));
 sg13g2_a21oi_1 _16030_ (.A1(_09243_),
    .A2(_09245_),
    .Y(_09246_),
    .B1(\cpu.spi.r_state[5] ));
 sg13g2_buf_1 _16031_ (.A(\cpu.spi.r_state[4] ),
    .X(_09247_));
 sg13g2_nand2b_1 _16032_ (.Y(_09248_),
    .B(_09237_),
    .A_N(_09228_));
 sg13g2_buf_2 _16033_ (.A(_09248_),
    .X(_09249_));
 sg13g2_buf_1 _16034_ (.A(_09249_),
    .X(_09250_));
 sg13g2_inv_2 _16035_ (.Y(_09251_),
    .A(net1151));
 sg13g2_nor2_1 _16036_ (.A(_09251_),
    .B(_09227_),
    .Y(_09252_));
 sg13g2_nor3_1 _16037_ (.A(net1150),
    .B(net352),
    .C(_09252_),
    .Y(_09253_));
 sg13g2_buf_2 _16038_ (.A(\cpu.spi.r_state[2] ),
    .X(_09254_));
 sg13g2_o21ai_1 _16039_ (.B1(net818),
    .Y(_09255_),
    .A1(_09254_),
    .A2(net353));
 sg13g2_a21oi_1 _16040_ (.A1(_09246_),
    .A2(_09253_),
    .Y(_00031_),
    .B1(_09255_));
 sg13g2_nand2b_1 _16041_ (.Y(_09256_),
    .B(net1),
    .A_N(r_reset));
 sg13g2_buf_1 _16042_ (.A(_09256_),
    .X(_09257_));
 sg13g2_buf_1 _16043_ (.A(_09257_),
    .X(_09258_));
 sg13g2_buf_1 _16044_ (.A(net929),
    .X(_09259_));
 sg13g2_buf_1 _16045_ (.A(_09259_),
    .X(_09260_));
 sg13g2_inv_1 _16046_ (.Y(_09261_),
    .A(net1152));
 sg13g2_nor2_1 _16047_ (.A(_09261_),
    .B(_09199_),
    .Y(_09262_));
 sg13g2_buf_1 _16048_ (.A(\cpu.spi.r_state[3] ),
    .X(_09263_));
 sg13g2_a21oi_1 _16049_ (.A1(_09185_),
    .A2(_09262_),
    .Y(_09264_),
    .B1(_09263_));
 sg13g2_nor3_1 _16050_ (.A(net714),
    .B(_09240_),
    .C(_09264_),
    .Y(_00032_));
 sg13g2_buf_2 _16051_ (.A(\cpu.spi.r_state[0] ),
    .X(_09265_));
 sg13g2_nand4_1 _16052_ (.B(net933),
    .C(_09183_),
    .A(_09265_),
    .Y(_09266_),
    .D(_09197_));
 sg13g2_buf_1 _16053_ (.A(_09266_),
    .X(_09267_));
 sg13g2_nand3_1 _16054_ (.B(net818),
    .C(_09250_),
    .A(net1150),
    .Y(_09268_));
 sg13g2_nand2_1 _16055_ (.Y(_00033_),
    .A(_09267_),
    .B(_09268_));
 sg13g2_nor3_1 _16056_ (.A(net714),
    .B(_09240_),
    .C(_09246_),
    .Y(_00034_));
 sg13g2_buf_1 _16057_ (.A(_09260_),
    .X(_09269_));
 sg13g2_nor2_1 _16058_ (.A(_09251_),
    .B(net353),
    .Y(_09270_));
 sg13g2_a21oi_1 _16059_ (.A1(_09254_),
    .A2(net353),
    .Y(_09271_),
    .B1(_09270_));
 sg13g2_nor2_1 _16060_ (.A(net647),
    .B(_09271_),
    .Y(_00035_));
 sg13g2_buf_1 _16061_ (.A(\cpu.ex.r_div_running ),
    .X(_09272_));
 sg13g2_buf_1 _16062_ (.A(\cpu.ex.r_mult_off[1] ),
    .X(_09273_));
 sg13g2_buf_1 _16063_ (.A(\cpu.ex.r_mult_off[2] ),
    .X(_09274_));
 sg13g2_buf_1 _16064_ (.A(\cpu.ex.r_mult_off[3] ),
    .X(_09275_));
 sg13g2_buf_1 _16065_ (.A(\cpu.ex.r_mult_off[0] ),
    .X(_09276_));
 sg13g2_buf_1 _16066_ (.A(\cpu.dec.div ),
    .X(_09277_));
 sg13g2_buf_1 _16067_ (.A(\cpu.dec.mult ),
    .X(_09278_));
 sg13g2_nand3b_1 _16068_ (.B(\cpu.dec.iready ),
    .C(_00197_),
    .Y(_09279_),
    .A_N(\cpu.ex.r_branch_stall ));
 sg13g2_buf_2 _16069_ (.A(_09279_),
    .X(_09280_));
 sg13g2_nor2_1 _16070_ (.A(_09257_),
    .B(_09280_),
    .Y(_09281_));
 sg13g2_o21ai_1 _16071_ (.B1(_09281_),
    .Y(_09282_),
    .A1(_09277_),
    .A2(_09278_));
 sg13g2_buf_1 _16072_ (.A(_09282_),
    .X(_09283_));
 sg13g2_buf_1 _16073_ (.A(_09283_),
    .X(_09284_));
 sg13g2_and2_1 _16074_ (.A(_09276_),
    .B(net646),
    .X(_09285_));
 sg13g2_buf_2 _16075_ (.A(_09285_),
    .X(_09286_));
 sg13g2_inv_1 _16076_ (.Y(\cpu.ex.c_mult_off[0] ),
    .A(_09286_));
 sg13g2_nor4_2 _16077_ (.A(_09273_),
    .B(_09274_),
    .C(_09275_),
    .Y(_09287_),
    .D(\cpu.ex.c_mult_off[0] ));
 sg13g2_buf_1 _16078_ (.A(_09281_),
    .X(_09288_));
 sg13g2_and2_1 _16079_ (.A(_09277_),
    .B(net814),
    .X(_09289_));
 sg13g2_buf_1 _16080_ (.A(_09289_),
    .X(_09290_));
 sg13g2_buf_1 _16081_ (.A(_09290_),
    .X(_09291_));
 sg13g2_o21ai_1 _16082_ (.B1(net1071),
    .Y(_09292_),
    .A1(_09272_),
    .A2(_09291_));
 sg13g2_a21oi_1 _16083_ (.A1(_09272_),
    .A2(_09287_),
    .Y(\cpu.ex.c_div_running ),
    .B1(_09292_));
 sg13g2_buf_2 _16084_ (.A(\cpu.ex.r_mult_running ),
    .X(_09293_));
 sg13g2_inv_2 _16085_ (.Y(_09294_),
    .A(_09293_));
 sg13g2_nand2_1 _16086_ (.Y(_09295_),
    .A(_09278_),
    .B(_09288_));
 sg13g2_buf_1 _16087_ (.A(_09295_),
    .X(_09296_));
 sg13g2_nand2_1 _16088_ (.Y(_09297_),
    .A(_09294_),
    .B(_09296_));
 sg13g2_buf_1 _16089_ (.A(_09297_),
    .X(_09298_));
 sg13g2_nand2_1 _16090_ (.Y(_09299_),
    .A(net1071),
    .B(net492));
 sg13g2_a21oi_1 _16091_ (.A1(_09293_),
    .A2(_09287_),
    .Y(\cpu.ex.c_mult_running ),
    .B1(_09299_));
 sg13g2_inv_1 _16092_ (.Y(_09300_),
    .A(_09265_));
 sg13g2_a21oi_1 _16093_ (.A1(_09183_),
    .A2(_09197_),
    .Y(_09301_),
    .B1(_09300_));
 sg13g2_nor2_1 _16094_ (.A(net929),
    .B(_09301_),
    .Y(_09302_));
 sg13g2_o21ai_1 _16095_ (.B1(_09302_),
    .Y(_00029_),
    .A1(net352),
    .A2(_09264_));
 sg13g2_buf_2 _16096_ (.A(\cpu.dcache.flush_write ),
    .X(_09303_));
 sg13g2_buf_1 _16097_ (.A(_08361_),
    .X(_09304_));
 sg13g2_buf_8 _16098_ (.A(_08257_),
    .X(_09305_));
 sg13g2_buf_8 _16099_ (.A(_09305_),
    .X(_09306_));
 sg13g2_buf_2 _16100_ (.A(_09306_),
    .X(_09307_));
 sg13g2_buf_1 _16101_ (.A(net949),
    .X(_09308_));
 sg13g2_buf_2 _16102_ (.A(_09308_),
    .X(_09309_));
 sg13g2_mux4_1 _16103_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .S1(net711),
    .X(_09310_));
 sg13g2_mux4_1 _16104_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .S1(net711),
    .X(_09311_));
 sg13g2_buf_8 _16105_ (.A(_09305_),
    .X(_09312_));
 sg13g2_buf_2 _16106_ (.A(net811),
    .X(_09313_));
 sg13g2_buf_1 _16107_ (.A(_08360_),
    .X(_09314_));
 sg13g2_buf_2 _16108_ (.A(_09314_),
    .X(_09315_));
 sg13g2_mux4_1 _16109_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .S1(net709),
    .X(_09316_));
 sg13g2_mux4_1 _16110_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .S1(net709),
    .X(_09317_));
 sg13g2_buf_2 _16111_ (.A(net948),
    .X(_09318_));
 sg13g2_buf_2 _16112_ (.A(net1086),
    .X(_09319_));
 sg13g2_buf_1 _16113_ (.A(_09319_),
    .X(_09320_));
 sg13g2_mux4_1 _16114_ (.S0(net809),
    .A0(_09310_),
    .A1(_09311_),
    .A2(_09316_),
    .A3(_09317_),
    .S1(net808),
    .X(_09321_));
 sg13g2_nand2_1 _16115_ (.Y(_09322_),
    .A(net713),
    .B(_09321_));
 sg13g2_buf_1 _16116_ (.A(_08368_),
    .X(_09323_));
 sg13g2_mux4_1 _16117_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .S1(net709),
    .X(_09324_));
 sg13g2_mux4_1 _16118_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .S1(net709),
    .X(_09325_));
 sg13g2_mux4_1 _16119_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .S1(net709),
    .X(_09326_));
 sg13g2_mux4_1 _16120_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .S1(net709),
    .X(_09327_));
 sg13g2_mux4_1 _16121_ (.S0(net809),
    .A0(_09324_),
    .A1(_09325_),
    .A2(_09326_),
    .A3(_09327_),
    .S1(net808),
    .X(_09328_));
 sg13g2_nand2_1 _16122_ (.Y(_09329_),
    .A(net708),
    .B(_09328_));
 sg13g2_a21oi_2 _16123_ (.B1(_08540_),
    .Y(_09330_),
    .A2(_09329_),
    .A1(_09322_));
 sg13g2_buf_1 _16124_ (.A(_09330_),
    .X(_09331_));
 sg13g2_inv_1 _16125_ (.Y(_09332_),
    .A(_00240_));
 sg13g2_buf_8 _16126_ (.A(\cpu.addr[4] ),
    .X(_09333_));
 sg13g2_or2_1 _16127_ (.X(_09334_),
    .B(_09186_),
    .A(_09333_));
 sg13g2_buf_2 _16128_ (.A(_09334_),
    .X(_09335_));
 sg13g2_buf_1 _16129_ (.A(_00220_),
    .X(_09336_));
 sg13g2_and2_1 _16130_ (.A(net1153),
    .B(_09336_),
    .X(_09337_));
 sg13g2_buf_1 _16131_ (.A(_09337_),
    .X(_09338_));
 sg13g2_nor2_1 _16132_ (.A(_09335_),
    .B(_09338_),
    .Y(_09339_));
 sg13g2_buf_1 _16133_ (.A(_09339_),
    .X(_09340_));
 sg13g2_nand2_1 _16134_ (.Y(_09341_),
    .A(net1153),
    .B(_09333_));
 sg13g2_nor2_1 _16135_ (.A(net930),
    .B(_09341_),
    .Y(_09342_));
 sg13g2_buf_1 _16136_ (.A(_09342_),
    .X(_09343_));
 sg13g2_a22oi_1 _16137_ (.Y(_09344_),
    .B1(net706),
    .B2(\cpu.dcache.r_tag[5][17] ),
    .A2(net707),
    .A1(_09332_));
 sg13g2_nor2b_1 _16138_ (.A(net1153),
    .B_N(_09333_),
    .Y(_09345_));
 sg13g2_buf_2 _16139_ (.A(_09345_),
    .X(_09346_));
 sg13g2_and2_1 _16140_ (.A(net1068),
    .B(_09346_),
    .X(_09347_));
 sg13g2_buf_2 _16141_ (.A(_09347_),
    .X(_09348_));
 sg13g2_buf_1 _16142_ (.A(_09348_),
    .X(_09349_));
 sg13g2_buf_1 _16143_ (.A(_09336_),
    .X(_09350_));
 sg13g2_nor2b_1 _16144_ (.A(_09186_),
    .B_N(net1065),
    .Y(_09351_));
 sg13g2_and2_1 _16145_ (.A(net1153),
    .B(_09351_),
    .X(_09352_));
 sg13g2_buf_8 _16146_ (.A(_09352_),
    .X(_09353_));
 sg13g2_buf_1 _16147_ (.A(net705),
    .X(_09354_));
 sg13g2_a22oi_1 _16148_ (.Y(_09355_),
    .B1(net643),
    .B2(\cpu.dcache.r_tag[1][17] ),
    .A2(net644),
    .A1(\cpu.dcache.r_tag[6][17] ));
 sg13g2_and2_1 _16149_ (.A(_09186_),
    .B(_09336_),
    .X(_09356_));
 sg13g2_buf_2 _16150_ (.A(_09356_),
    .X(_09357_));
 sg13g2_and2_1 _16151_ (.A(net1070),
    .B(_09357_),
    .X(_09358_));
 sg13g2_buf_2 _16152_ (.A(_09358_),
    .X(_09359_));
 sg13g2_buf_1 _16153_ (.A(_09359_),
    .X(_09360_));
 sg13g2_nor2b_1 _16154_ (.A(net1068),
    .B_N(_09346_),
    .Y(_09361_));
 sg13g2_buf_1 _16155_ (.A(_09361_),
    .X(_09362_));
 sg13g2_a22oi_1 _16156_ (.Y(_09363_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[4][17] ),
    .A2(net642),
    .A1(\cpu.dcache.r_tag[3][17] ));
 sg13g2_and3_1 _16157_ (.X(_09364_),
    .A(net1153),
    .B(_09333_),
    .C(_09187_));
 sg13g2_buf_1 _16158_ (.A(_09364_),
    .X(_09365_));
 sg13g2_buf_2 _16159_ (.A(_09365_),
    .X(_09366_));
 sg13g2_inv_1 _16160_ (.Y(_09367_),
    .A(net1153));
 sg13g2_and2_1 _16161_ (.A(_09367_),
    .B(_09357_),
    .X(_09368_));
 sg13g2_buf_2 _16162_ (.A(_09368_),
    .X(_09369_));
 sg13g2_buf_1 _16163_ (.A(_09369_),
    .X(_09370_));
 sg13g2_a22oi_1 _16164_ (.Y(_09371_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][17] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[7][17] ));
 sg13g2_nand4_1 _16165_ (.B(_09355_),
    .C(_09363_),
    .A(_09344_),
    .Y(_09372_),
    .D(_09371_));
 sg13g2_xor2_1 _16166_ (.B(_09372_),
    .A(net391),
    .X(_09373_));
 sg13g2_mux4_1 _16167_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .S1(net711),
    .X(_09374_));
 sg13g2_mux4_1 _16168_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .S1(net711),
    .X(_09375_));
 sg13g2_mux4_1 _16169_ (.S0(_09313_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .S1(_09315_),
    .X(_09376_));
 sg13g2_mux4_1 _16170_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .S1(net709),
    .X(_09377_));
 sg13g2_mux4_1 _16171_ (.S0(net809),
    .A0(_09374_),
    .A1(_09375_),
    .A2(_09376_),
    .A3(_09377_),
    .S1(_09320_),
    .X(_09378_));
 sg13g2_nand2_1 _16172_ (.Y(_09379_),
    .A(net713),
    .B(_09378_));
 sg13g2_mux4_1 _16173_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .S1(net711),
    .X(_09380_));
 sg13g2_mux4_1 _16174_ (.S0(_09307_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .S1(_09309_),
    .X(_09381_));
 sg13g2_mux4_1 _16175_ (.S0(net710),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .S1(net709),
    .X(_09382_));
 sg13g2_mux4_1 _16176_ (.S0(_09313_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .S1(_09315_),
    .X(_09383_));
 sg13g2_mux4_1 _16177_ (.S0(net809),
    .A0(_09380_),
    .A1(_09381_),
    .A2(_09382_),
    .A3(_09383_),
    .S1(net808),
    .X(_09384_));
 sg13g2_nand2_1 _16178_ (.Y(_09385_),
    .A(net708),
    .B(_09384_));
 sg13g2_a21oi_2 _16179_ (.B1(net1075),
    .Y(_09386_),
    .A2(_09385_),
    .A1(_09379_));
 sg13g2_buf_1 _16180_ (.A(_09386_),
    .X(_09387_));
 sg13g2_inv_1 _16181_ (.Y(_09388_),
    .A(_00239_));
 sg13g2_a22oi_1 _16182_ (.Y(_09389_),
    .B1(net706),
    .B2(\cpu.dcache.r_tag[5][16] ),
    .A2(net707),
    .A1(_09388_));
 sg13g2_buf_1 _16183_ (.A(net704),
    .X(_09390_));
 sg13g2_a22oi_1 _16184_ (.Y(_09391_),
    .B1(_09390_),
    .B2(\cpu.dcache.r_tag[4][16] ),
    .A2(net705),
    .A1(\cpu.dcache.r_tag[1][16] ));
 sg13g2_a22oi_1 _16185_ (.Y(_09392_),
    .B1(net642),
    .B2(\cpu.dcache.r_tag[3][16] ),
    .A2(net644),
    .A1(\cpu.dcache.r_tag[6][16] ));
 sg13g2_a22oi_1 _16186_ (.Y(_09393_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][16] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[7][16] ));
 sg13g2_nand4_1 _16187_ (.B(_09391_),
    .C(_09392_),
    .A(_09389_),
    .Y(_09394_),
    .D(_09393_));
 sg13g2_xor2_1 _16188_ (.B(_09394_),
    .A(net390),
    .X(_09395_));
 sg13g2_buf_8 _16189_ (.A(_09305_),
    .X(_09396_));
 sg13g2_buf_2 _16190_ (.A(_09396_),
    .X(_09397_));
 sg13g2_buf_2 _16191_ (.A(net812),
    .X(_09398_));
 sg13g2_mux4_1 _16192_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .S1(net701),
    .X(_09399_));
 sg13g2_mux4_1 _16193_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .S1(net701),
    .X(_09400_));
 sg13g2_mux4_1 _16194_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .S1(net711),
    .X(_09401_));
 sg13g2_mux4_1 _16195_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .S1(net711),
    .X(_09402_));
 sg13g2_mux4_1 _16196_ (.S0(net809),
    .A0(_09399_),
    .A1(_09400_),
    .A2(_09401_),
    .A3(_09402_),
    .S1(_09320_),
    .X(_09403_));
 sg13g2_nand2_1 _16197_ (.Y(_09404_),
    .A(net713),
    .B(_09403_));
 sg13g2_mux4_1 _16198_ (.S0(_09397_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .S1(_09398_),
    .X(_09405_));
 sg13g2_mux4_1 _16199_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .S1(net701),
    .X(_09406_));
 sg13g2_mux4_1 _16200_ (.S0(_09307_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .S1(_09309_),
    .X(_09407_));
 sg13g2_mux4_1 _16201_ (.S0(net712),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .S1(net711),
    .X(_09408_));
 sg13g2_mux4_1 _16202_ (.S0(net809),
    .A0(_09405_),
    .A1(_09406_),
    .A2(_09407_),
    .A3(_09408_),
    .S1(net808),
    .X(_09409_));
 sg13g2_nand2_1 _16203_ (.Y(_09410_),
    .A(net708),
    .B(_09409_));
 sg13g2_a21oi_2 _16204_ (.B1(net1075),
    .Y(_09411_),
    .A2(_09410_),
    .A1(_09404_));
 sg13g2_buf_1 _16205_ (.A(_09411_),
    .X(_09412_));
 sg13g2_inv_1 _16206_ (.Y(_09413_),
    .A(_00242_));
 sg13g2_buf_2 _16207_ (.A(net706),
    .X(_09414_));
 sg13g2_a22oi_1 _16208_ (.Y(_09415_),
    .B1(_09414_),
    .B2(\cpu.dcache.r_tag[5][19] ),
    .A2(net707),
    .A1(_09413_));
 sg13g2_a22oi_1 _16209_ (.Y(_09416_),
    .B1(_09390_),
    .B2(\cpu.dcache.r_tag[4][19] ),
    .A2(net643),
    .A1(\cpu.dcache.r_tag[1][19] ));
 sg13g2_a22oi_1 _16210_ (.Y(_09417_),
    .B1(net642),
    .B2(\cpu.dcache.r_tag[3][19] ),
    .A2(net644),
    .A1(\cpu.dcache.r_tag[6][19] ));
 sg13g2_a22oi_1 _16211_ (.Y(_09418_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][19] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[7][19] ));
 sg13g2_nand4_1 _16212_ (.B(_09416_),
    .C(_09417_),
    .A(_09415_),
    .Y(_09419_),
    .D(_09418_));
 sg13g2_xor2_1 _16213_ (.B(_09419_),
    .A(_09412_),
    .X(_09420_));
 sg13g2_nor3_1 _16214_ (.A(_09373_),
    .B(_09395_),
    .C(_09420_),
    .Y(_09421_));
 sg13g2_mux4_1 _16215_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .S1(net701),
    .X(_09422_));
 sg13g2_mux4_1 _16216_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .S1(net701),
    .X(_09423_));
 sg13g2_mux4_1 _16217_ (.S0(net702),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .S1(net701),
    .X(_09424_));
 sg13g2_mux4_1 _16218_ (.S0(_09397_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .S1(_09398_),
    .X(_09425_));
 sg13g2_mux4_1 _16219_ (.S0(_09318_),
    .A0(_09422_),
    .A1(_09423_),
    .A2(_09424_),
    .A3(_09425_),
    .S1(net808),
    .X(_09426_));
 sg13g2_buf_1 _16220_ (.A(_08257_),
    .X(_09427_));
 sg13g2_buf_2 _16221_ (.A(net927),
    .X(_09428_));
 sg13g2_buf_8 _16222_ (.A(net949),
    .X(_09429_));
 sg13g2_buf_1 _16223_ (.A(net805),
    .X(_09430_));
 sg13g2_mux4_1 _16224_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .S1(net700),
    .X(_09431_));
 sg13g2_mux4_1 _16225_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .S1(net700),
    .X(_09432_));
 sg13g2_mux4_1 _16226_ (.S0(_09428_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .S1(_09430_),
    .X(_09433_));
 sg13g2_mux4_1 _16227_ (.S0(_09428_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .S1(_09430_),
    .X(_09434_));
 sg13g2_buf_2 _16228_ (.A(net948),
    .X(_09435_));
 sg13g2_mux4_1 _16229_ (.S0(net804),
    .A0(_09431_),
    .A1(_09432_),
    .A2(_09433_),
    .A3(_09434_),
    .S1(_09319_),
    .X(_09436_));
 sg13g2_and2_1 _16230_ (.A(_09304_),
    .B(_09436_),
    .X(_09437_));
 sg13g2_a21oi_1 _16231_ (.A1(net708),
    .A2(_09426_),
    .Y(_09438_),
    .B1(_09437_));
 sg13g2_nor2_1 _16232_ (.A(net1080),
    .B(net702),
    .Y(_09439_));
 sg13g2_a21oi_2 _16233_ (.B1(_09439_),
    .Y(_09440_),
    .A2(_09438_),
    .A1(net1080));
 sg13g2_buf_1 _16234_ (.A(_09440_),
    .X(_09441_));
 sg13g2_nor2_1 _16235_ (.A(_09333_),
    .B(net1068),
    .Y(_09442_));
 sg13g2_buf_1 _16236_ (.A(_09442_),
    .X(_09443_));
 sg13g2_a22oi_1 _16237_ (.Y(_09444_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[7][12] ),
    .A2(net642),
    .A1(\cpu.dcache.r_tag[3][12] ));
 sg13g2_a22oi_1 _16238_ (.Y(_09445_),
    .B1(_09349_),
    .B2(\cpu.dcache.r_tag[6][12] ),
    .A2(net706),
    .A1(\cpu.dcache.r_tag[5][12] ));
 sg13g2_a22oi_1 _16239_ (.Y(_09446_),
    .B1(_09369_),
    .B2(\cpu.dcache.r_tag[2][12] ),
    .A2(net704),
    .A1(\cpu.dcache.r_tag[4][12] ));
 sg13g2_nand3_1 _16240_ (.B(_09445_),
    .C(_09446_),
    .A(_09444_),
    .Y(_09447_));
 sg13g2_nand2_1 _16241_ (.Y(_09448_),
    .A(_00235_),
    .B(_09443_));
 sg13g2_o21ai_1 _16242_ (.B1(_09448_),
    .Y(_09449_),
    .A1(_09443_),
    .A2(_09447_));
 sg13g2_o21ai_1 _16243_ (.B1(net643),
    .Y(_09450_),
    .A1(\cpu.dcache.r_tag[1][12] ),
    .A2(_09447_));
 sg13g2_o21ai_1 _16244_ (.B1(_09450_),
    .Y(_09451_),
    .A1(net643),
    .A2(_09449_));
 sg13g2_xnor2_1 _16245_ (.Y(_09452_),
    .A(_09441_),
    .B(_09451_));
 sg13g2_buf_1 _16246_ (.A(_09333_),
    .X(_09453_));
 sg13g2_inv_2 _16247_ (.Y(_09454_),
    .A(net1064));
 sg13g2_buf_1 _16248_ (.A(_09367_),
    .X(_09455_));
 sg13g2_mux2_1 _16249_ (.A0(\cpu.dcache.r_tag[4][13] ),
    .A1(\cpu.dcache.r_tag[6][13] ),
    .S(_09189_),
    .X(_09456_));
 sg13g2_and2_1 _16250_ (.A(net932),
    .B(net816),
    .X(_09457_));
 sg13g2_a22oi_1 _16251_ (.Y(_09458_),
    .B1(_09457_),
    .B2(\cpu.dcache.r_tag[7][13] ),
    .A2(_09456_),
    .A1(net926));
 sg13g2_nand2b_1 _16252_ (.Y(_09459_),
    .B(_09443_),
    .A_N(_09338_));
 sg13g2_buf_2 _16253_ (.A(_09459_),
    .X(_09460_));
 sg13g2_a22oi_1 _16254_ (.Y(_09461_),
    .B1(net705),
    .B2(\cpu.dcache.r_tag[1][13] ),
    .A2(net706),
    .A1(\cpu.dcache.r_tag[5][13] ));
 sg13g2_o21ai_1 _16255_ (.B1(_09461_),
    .Y(_09462_),
    .A1(_00236_),
    .A2(_09460_));
 sg13g2_a221oi_1 _16256_ (.B2(\cpu.dcache.r_tag[2][13] ),
    .C1(_09462_),
    .B1(net641),
    .A1(\cpu.dcache.r_tag[3][13] ),
    .Y(_09463_),
    .A2(net642));
 sg13g2_o21ai_1 _16257_ (.B1(_09463_),
    .Y(_09464_),
    .A1(_09454_),
    .A2(_09458_));
 sg13g2_mux4_1 _16258_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .S1(_09308_),
    .X(_09465_));
 sg13g2_mux4_1 _16259_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .S1(net812),
    .X(_09466_));
 sg13g2_mux4_1 _16260_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .S1(net812),
    .X(_09467_));
 sg13g2_mux4_1 _16261_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .S1(net812),
    .X(_09468_));
 sg13g2_mux4_1 _16262_ (.S0(net804),
    .A0(_09465_),
    .A1(_09466_),
    .A2(_09467_),
    .A3(_09468_),
    .S1(net928),
    .X(_09469_));
 sg13g2_mux4_1 _16263_ (.S0(_09305_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .S1(net949),
    .X(_09470_));
 sg13g2_mux4_1 _16264_ (.S0(_09305_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .S1(_09429_),
    .X(_09471_));
 sg13g2_mux4_1 _16265_ (.S0(_09305_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .S1(net949),
    .X(_09472_));
 sg13g2_mux4_1 _16266_ (.S0(_09305_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .S1(net949),
    .X(_09473_));
 sg13g2_mux4_1 _16267_ (.S0(net948),
    .A0(_09470_),
    .A1(_09471_),
    .A2(_09472_),
    .A3(_09473_),
    .S1(net1086),
    .X(_09474_));
 sg13g2_and2_1 _16268_ (.A(_09304_),
    .B(_09474_),
    .X(_09475_));
 sg13g2_a21oi_1 _16269_ (.A1(_09323_),
    .A2(_09469_),
    .Y(_09476_),
    .B1(_09475_));
 sg13g2_nor2_1 _16270_ (.A(net1165),
    .B(net701),
    .Y(_09477_));
 sg13g2_a21oi_2 _16271_ (.B1(_09477_),
    .Y(_09478_),
    .A2(_09476_),
    .A1(_08424_));
 sg13g2_buf_1 _16272_ (.A(_09478_),
    .X(_09479_));
 sg13g2_xor2_1 _16273_ (.B(_09479_),
    .A(_09464_),
    .X(_09480_));
 sg13g2_nand2_1 _16274_ (.Y(_09481_),
    .A(net932),
    .B(_09351_));
 sg13g2_buf_1 _16275_ (.A(_09481_),
    .X(_09482_));
 sg13g2_a22oi_1 _16276_ (.Y(_09483_),
    .B1(_09359_),
    .B2(\cpu.dcache.r_tag[3][10] ),
    .A2(_09342_),
    .A1(\cpu.dcache.r_tag[5][10] ));
 sg13g2_a22oi_1 _16277_ (.Y(_09484_),
    .B1(_09361_),
    .B2(\cpu.dcache.r_tag[4][10] ),
    .A2(_09348_),
    .A1(\cpu.dcache.r_tag[6][10] ));
 sg13g2_a22oi_1 _16278_ (.Y(_09485_),
    .B1(_09369_),
    .B2(\cpu.dcache.r_tag[2][10] ),
    .A2(_09365_),
    .A1(\cpu.dcache.r_tag[7][10] ));
 sg13g2_and3_1 _16279_ (.X(_09486_),
    .A(_09483_),
    .B(_09484_),
    .C(_09485_));
 sg13g2_mux2_1 _16280_ (.A0(_00232_),
    .A1(_09486_),
    .S(_09335_),
    .X(_09487_));
 sg13g2_nor2_1 _16281_ (.A(\cpu.dcache.r_tag[1][10] ),
    .B(net699),
    .Y(_09488_));
 sg13g2_a22oi_1 _16282_ (.Y(_09489_),
    .B1(_09488_),
    .B2(_09486_),
    .A2(_09487_),
    .A1(net699));
 sg13g2_xnor2_1 _16283_ (.Y(_09490_),
    .A(_00231_),
    .B(_09489_));
 sg13g2_a22oi_1 _16284_ (.Y(_09491_),
    .B1(_09369_),
    .B2(\cpu.dcache.r_tag[2][6] ),
    .A2(_09365_),
    .A1(\cpu.dcache.r_tag[7][6] ));
 sg13g2_a22oi_1 _16285_ (.Y(_09492_),
    .B1(_09348_),
    .B2(\cpu.dcache.r_tag[6][6] ),
    .A2(_09342_),
    .A1(\cpu.dcache.r_tag[5][6] ));
 sg13g2_a22oi_1 _16286_ (.Y(_09493_),
    .B1(_09362_),
    .B2(\cpu.dcache.r_tag[4][6] ),
    .A2(_09359_),
    .A1(\cpu.dcache.r_tag[3][6] ));
 sg13g2_and3_1 _16287_ (.X(_09494_),
    .A(_09491_),
    .B(_09492_),
    .C(_09493_));
 sg13g2_mux2_1 _16288_ (.A0(_00224_),
    .A1(_09494_),
    .S(_09335_),
    .X(_09495_));
 sg13g2_nor2_1 _16289_ (.A(\cpu.dcache.r_tag[1][6] ),
    .B(_09482_),
    .Y(_09496_));
 sg13g2_a22oi_1 _16290_ (.Y(_09497_),
    .B1(_09496_),
    .B2(_09494_),
    .A2(_09495_),
    .A1(_09482_));
 sg13g2_xnor2_1 _16291_ (.Y(_09498_),
    .A(_00223_),
    .B(_09497_));
 sg13g2_mux2_1 _16292_ (.A0(\cpu.dcache.r_tag[4][11] ),
    .A1(\cpu.dcache.r_tag[6][11] ),
    .S(net930),
    .X(_09499_));
 sg13g2_buf_1 _16293_ (.A(net1064),
    .X(_09500_));
 sg13g2_a22oi_1 _16294_ (.Y(_09501_),
    .B1(_09499_),
    .B2(_09500_),
    .A2(_09357_),
    .A1(\cpu.dcache.r_tag[2][11] ));
 sg13g2_mux2_1 _16295_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(\cpu.dcache.r_tag[7][11] ),
    .S(net930),
    .X(_09502_));
 sg13g2_a221oi_1 _16296_ (.B2(_09453_),
    .C1(_09455_),
    .B1(_09502_),
    .A1(\cpu.dcache.r_tag[3][11] ),
    .Y(_09503_),
    .A2(_09357_));
 sg13g2_a21oi_1 _16297_ (.A1(net926),
    .A2(_09501_),
    .Y(_09504_),
    .B1(_09503_));
 sg13g2_nor2_1 _16298_ (.A(\cpu.dcache.r_tag[1][11] ),
    .B(_09504_),
    .Y(_09505_));
 sg13g2_nor2_1 _16299_ (.A(_00234_),
    .B(_09335_),
    .Y(_09506_));
 sg13g2_nor3_1 _16300_ (.A(_09354_),
    .B(_09506_),
    .C(_09504_),
    .Y(_09507_));
 sg13g2_a21o_1 _16301_ (.A2(_09505_),
    .A1(_09354_),
    .B1(_09507_),
    .X(_09508_));
 sg13g2_xor2_1 _16302_ (.B(_09508_),
    .A(_00233_),
    .X(_09509_));
 sg13g2_nor4_1 _16303_ (.A(_09480_),
    .B(_09490_),
    .C(_09498_),
    .D(_09509_),
    .Y(_09510_));
 sg13g2_inv_1 _16304_ (.Y(_09511_),
    .A(net1065));
 sg13g2_mux2_1 _16305_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(\cpu.dcache.r_tag[3][14] ),
    .S(net930),
    .X(_09512_));
 sg13g2_nor2b_1 _16306_ (.A(net932),
    .B_N(net930),
    .Y(_09513_));
 sg13g2_a22oi_1 _16307_ (.Y(_09514_),
    .B1(_09513_),
    .B2(\cpu.dcache.r_tag[2][14] ),
    .A2(_09512_),
    .A1(net932));
 sg13g2_nor2_1 _16308_ (.A(_09511_),
    .B(_09514_),
    .Y(_09515_));
 sg13g2_mux2_1 _16309_ (.A0(\cpu.dcache.r_tag[4][14] ),
    .A1(\cpu.dcache.r_tag[6][14] ),
    .S(net930),
    .X(_09516_));
 sg13g2_nor2_2 _16310_ (.A(_09367_),
    .B(net816),
    .Y(_09517_));
 sg13g2_a22oi_1 _16311_ (.Y(_09518_),
    .B1(_09517_),
    .B2(\cpu.dcache.r_tag[5][14] ),
    .A2(_09516_),
    .A1(net926));
 sg13g2_nor2_1 _16312_ (.A(_09454_),
    .B(_09518_),
    .Y(_09519_));
 sg13g2_nand2_1 _16313_ (.Y(_09520_),
    .A(\cpu.dcache.r_tag[7][14] ),
    .B(_09365_));
 sg13g2_o21ai_1 _16314_ (.B1(_09520_),
    .Y(_09521_),
    .A1(_00237_),
    .A2(_09460_));
 sg13g2_nor3_1 _16315_ (.A(_09515_),
    .B(_09519_),
    .C(_09521_),
    .Y(_09522_));
 sg13g2_buf_1 _16316_ (.A(net809),
    .X(_09523_));
 sg13g2_mux4_1 _16317_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .S1(_09429_),
    .X(_09524_));
 sg13g2_buf_8 _16318_ (.A(_09305_),
    .X(_09525_));
 sg13g2_buf_8 _16319_ (.A(net949),
    .X(_09526_));
 sg13g2_mux4_1 _16320_ (.S0(_09525_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .S1(_09526_),
    .X(_09527_));
 sg13g2_mux4_1 _16321_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .S1(net805),
    .X(_09528_));
 sg13g2_mux4_1 _16322_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .S1(net805),
    .X(_09529_));
 sg13g2_mux4_1 _16323_ (.S0(_08368_),
    .A0(_09524_),
    .A1(_09527_),
    .A2(_09528_),
    .A3(_09529_),
    .S1(net1086),
    .X(_09530_));
 sg13g2_nand2_1 _16324_ (.Y(_09531_),
    .A(_08271_),
    .B(_09530_));
 sg13g2_mux4_1 _16325_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .S1(net802),
    .X(_09532_));
 sg13g2_mux4_1 _16326_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .S1(net802),
    .X(_09533_));
 sg13g2_mux4_1 _16327_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .S1(net805),
    .X(_09534_));
 sg13g2_mux4_1 _16328_ (.S0(_09427_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .S1(net805),
    .X(_09535_));
 sg13g2_mux4_1 _16329_ (.S0(_08368_),
    .A0(_09532_),
    .A1(_09533_),
    .A2(_09534_),
    .A3(_09535_),
    .S1(_08278_),
    .X(_09536_));
 sg13g2_o21ai_1 _16330_ (.B1(_09318_),
    .Y(_09537_),
    .A1(_08336_),
    .A2(_09536_));
 sg13g2_o21ai_1 _16331_ (.B1(_09537_),
    .Y(_09538_),
    .A1(net698),
    .A2(_09531_));
 sg13g2_buf_1 _16332_ (.A(_09538_),
    .X(_09539_));
 sg13g2_xor2_1 _16333_ (.B(_09539_),
    .A(_09522_),
    .X(_09540_));
 sg13g2_inv_1 _16334_ (.Y(_09541_),
    .A(_00225_));
 sg13g2_nand3b_1 _16335_ (.B(\cpu.dcache.r_tag[4][7] ),
    .C(net1064),
    .Y(_09542_),
    .A_N(net1068));
 sg13g2_nand4_1 _16336_ (.B(net1068),
    .C(net1065),
    .A(net1070),
    .Y(_09543_),
    .D(\cpu.dcache.r_tag[3][7] ));
 sg13g2_o21ai_1 _16337_ (.B1(_09543_),
    .Y(_09544_),
    .A1(net1070),
    .A2(_09542_));
 sg13g2_inv_1 _16338_ (.Y(_09545_),
    .A(\cpu.dcache.r_tag[5][7] ));
 sg13g2_nand3b_1 _16339_ (.B(_09333_),
    .C(_09172_),
    .Y(_09546_),
    .A_N(_09186_));
 sg13g2_buf_1 _16340_ (.A(_09546_),
    .X(_09547_));
 sg13g2_nand4_1 _16341_ (.B(net1064),
    .C(net1068),
    .A(net1070),
    .Y(_09548_),
    .D(\cpu.dcache.r_tag[7][7] ));
 sg13g2_o21ai_1 _16342_ (.B1(_09548_),
    .Y(_09549_),
    .A1(_09545_),
    .A2(_09547_));
 sg13g2_inv_1 _16343_ (.Y(_09550_),
    .A(\cpu.dcache.r_tag[2][7] ));
 sg13g2_nand3b_1 _16344_ (.B(net1068),
    .C(net1065),
    .Y(_09551_),
    .A_N(net1153));
 sg13g2_buf_1 _16345_ (.A(_09551_),
    .X(_09552_));
 sg13g2_nor2_1 _16346_ (.A(_09550_),
    .B(_09552_),
    .Y(_09553_));
 sg13g2_inv_1 _16347_ (.Y(_09554_),
    .A(\cpu.dcache.r_tag[6][7] ));
 sg13g2_nand3b_1 _16348_ (.B(_09333_),
    .C(_09186_),
    .Y(_09555_),
    .A_N(net1153));
 sg13g2_buf_2 _16349_ (.A(_09555_),
    .X(_09556_));
 sg13g2_nor2_1 _16350_ (.A(_09554_),
    .B(_09556_),
    .Y(_09557_));
 sg13g2_nor4_1 _16351_ (.A(_09544_),
    .B(_09549_),
    .C(_09553_),
    .D(_09557_),
    .Y(_09558_));
 sg13g2_mux2_1 _16352_ (.A0(_00226_),
    .A1(_09558_),
    .S(_09335_),
    .X(_09559_));
 sg13g2_nor2_1 _16353_ (.A(\cpu.dcache.r_tag[1][7] ),
    .B(_09481_),
    .Y(_09560_));
 sg13g2_a22oi_1 _16354_ (.Y(_09561_),
    .B1(_09560_),
    .B2(_09558_),
    .A2(_09559_),
    .A1(_09481_));
 sg13g2_xnor2_1 _16355_ (.Y(_09562_),
    .A(_09541_),
    .B(_09561_));
 sg13g2_buf_1 _16356_ (.A(_00221_),
    .X(_09563_));
 sg13g2_inv_2 _16357_ (.Y(_09564_),
    .A(_09563_));
 sg13g2_mux2_1 _16358_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(\cpu.dcache.r_tag[7][5] ),
    .S(_09188_),
    .X(_09565_));
 sg13g2_a22oi_1 _16359_ (.Y(_09566_),
    .B1(_09565_),
    .B2(_09453_),
    .A2(_09357_),
    .A1(\cpu.dcache.r_tag[3][5] ));
 sg13g2_nand2b_1 _16360_ (.Y(_09567_),
    .B(net932),
    .A_N(_09566_));
 sg13g2_and2_1 _16361_ (.A(net1064),
    .B(_09187_),
    .X(_09568_));
 sg13g2_and3_1 _16362_ (.X(_09569_),
    .A(_09367_),
    .B(\cpu.dcache.r_tag[6][5] ),
    .C(_09568_));
 sg13g2_a221oi_1 _16363_ (.B2(\cpu.dcache.r_tag[4][5] ),
    .C1(_09569_),
    .B1(net704),
    .A1(\cpu.dcache.r_tag[1][5] ),
    .Y(_09570_),
    .A2(net705));
 sg13g2_nand2b_1 _16364_ (.Y(_09571_),
    .B(net707),
    .A_N(_00222_));
 sg13g2_nand3_1 _16365_ (.B(\cpu.dcache.r_tag[2][5] ),
    .C(_09357_),
    .A(net926),
    .Y(_09572_));
 sg13g2_and4_1 _16366_ (.A(_09567_),
    .B(_09570_),
    .C(_09571_),
    .D(_09572_),
    .X(_09573_));
 sg13g2_xnor2_1 _16367_ (.Y(_09574_),
    .A(_09564_),
    .B(_09573_));
 sg13g2_inv_1 _16368_ (.Y(_09575_),
    .A(_00228_));
 sg13g2_a22oi_1 _16369_ (.Y(_09576_),
    .B1(net706),
    .B2(\cpu.dcache.r_tag[5][8] ),
    .A2(_09339_),
    .A1(_09575_));
 sg13g2_a22oi_1 _16370_ (.Y(_09577_),
    .B1(\cpu.dcache.r_tag[3][8] ),
    .B2(net1065),
    .A2(\cpu.dcache.r_tag[7][8] ),
    .A1(net1064));
 sg13g2_a221oi_1 _16371_ (.B2(net1065),
    .C1(net1070),
    .B1(\cpu.dcache.r_tag[2][8] ),
    .A1(net1064),
    .Y(_09578_),
    .A2(\cpu.dcache.r_tag[6][8] ));
 sg13g2_a21oi_1 _16372_ (.A1(net932),
    .A2(_09577_),
    .Y(_09579_),
    .B1(_09578_));
 sg13g2_nand2_1 _16373_ (.Y(_09580_),
    .A(net816),
    .B(_09579_));
 sg13g2_a22oi_1 _16374_ (.Y(_09581_),
    .B1(_09346_),
    .B2(\cpu.dcache.r_tag[4][8] ),
    .A2(_09338_),
    .A1(\cpu.dcache.r_tag[1][8] ));
 sg13g2_or2_1 _16375_ (.X(_09582_),
    .B(_09581_),
    .A(net816));
 sg13g2_nand3_1 _16376_ (.B(_09580_),
    .C(_09582_),
    .A(_09576_),
    .Y(_09583_));
 sg13g2_xnor2_1 _16377_ (.Y(_09584_),
    .A(_00227_),
    .B(_09583_));
 sg13g2_a22oi_1 _16378_ (.Y(_09585_),
    .B1(\cpu.dcache.r_tag[2][9] ),
    .B2(_09350_),
    .A2(\cpu.dcache.r_tag[6][9] ),
    .A1(net1064));
 sg13g2_nand3_1 _16379_ (.B(_09350_),
    .C(\cpu.dcache.r_tag[3][9] ),
    .A(net1070),
    .Y(_09586_));
 sg13g2_o21ai_1 _16380_ (.B1(_09586_),
    .Y(_09587_),
    .A1(_09174_),
    .A2(_09585_));
 sg13g2_nand2_1 _16381_ (.Y(_09588_),
    .A(net816),
    .B(_09587_));
 sg13g2_inv_1 _16382_ (.Y(_09589_),
    .A(_00230_));
 sg13g2_a22oi_1 _16383_ (.Y(_09590_),
    .B1(net705),
    .B2(\cpu.dcache.r_tag[1][9] ),
    .A2(net707),
    .A1(_09589_));
 sg13g2_mux2_1 _16384_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(\cpu.dcache.r_tag[7][9] ),
    .S(_09188_),
    .X(_09591_));
 sg13g2_nor2_1 _16385_ (.A(net1070),
    .B(net930),
    .Y(_09592_));
 sg13g2_a22oi_1 _16386_ (.Y(_09593_),
    .B1(_09592_),
    .B2(\cpu.dcache.r_tag[4][9] ),
    .A2(_09591_),
    .A1(net1070));
 sg13g2_nand2b_1 _16387_ (.Y(_09594_),
    .B(net925),
    .A_N(_09593_));
 sg13g2_and3_1 _16388_ (.X(_09595_),
    .A(_09588_),
    .B(_09590_),
    .C(_09594_));
 sg13g2_xor2_1 _16389_ (.B(_09595_),
    .A(_00229_),
    .X(_09596_));
 sg13g2_nor3_1 _16390_ (.A(_09574_),
    .B(_09584_),
    .C(_09596_),
    .Y(_09597_));
 sg13g2_nand3_1 _16391_ (.B(_09562_),
    .C(_09597_),
    .A(_09540_),
    .Y(_09598_));
 sg13g2_buf_2 _16392_ (.A(net927),
    .X(_09599_));
 sg13g2_buf_1 _16393_ (.A(net805),
    .X(_09600_));
 sg13g2_mux4_1 _16394_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .S1(net697),
    .X(_09601_));
 sg13g2_mux4_1 _16395_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .S1(net700),
    .X(_09602_));
 sg13g2_mux4_1 _16396_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .S1(net697),
    .X(_09603_));
 sg13g2_mux4_1 _16397_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .S1(net697),
    .X(_09604_));
 sg13g2_mux4_1 _16398_ (.S0(net804),
    .A0(_09601_),
    .A1(_09602_),
    .A2(_09603_),
    .A3(_09604_),
    .S1(net928),
    .X(_09605_));
 sg13g2_nand2_1 _16399_ (.Y(_09606_),
    .A(net713),
    .B(_09605_));
 sg13g2_mux4_1 _16400_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .S1(net697),
    .X(_09607_));
 sg13g2_mux4_1 _16401_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .S1(net697),
    .X(_09608_));
 sg13g2_mux4_1 _16402_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .S1(net697),
    .X(_09609_));
 sg13g2_mux4_1 _16403_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .S1(net697),
    .X(_09610_));
 sg13g2_mux4_1 _16404_ (.S0(net804),
    .A0(_09607_),
    .A1(_09608_),
    .A2(_09609_),
    .A3(_09610_),
    .S1(net928),
    .X(_09611_));
 sg13g2_nand2_1 _16405_ (.Y(_09612_),
    .A(net708),
    .B(_09611_));
 sg13g2_a21oi_2 _16406_ (.B1(_08540_),
    .Y(_09613_),
    .A2(_09612_),
    .A1(_09606_));
 sg13g2_buf_2 _16407_ (.A(_09613_),
    .X(_09614_));
 sg13g2_inv_1 _16408_ (.Y(_09615_),
    .A(_00243_));
 sg13g2_a22oi_1 _16409_ (.Y(_09616_),
    .B1(net706),
    .B2(\cpu.dcache.r_tag[5][23] ),
    .A2(net707),
    .A1(_09615_));
 sg13g2_a22oi_1 _16410_ (.Y(_09617_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[4][23] ),
    .A2(net705),
    .A1(\cpu.dcache.r_tag[1][23] ));
 sg13g2_a22oi_1 _16411_ (.Y(_09618_),
    .B1(net642),
    .B2(\cpu.dcache.r_tag[3][23] ),
    .A2(net644),
    .A1(\cpu.dcache.r_tag[6][23] ));
 sg13g2_a22oi_1 _16412_ (.Y(_09619_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][23] ),
    .A2(net703),
    .A1(\cpu.dcache.r_tag[7][23] ));
 sg13g2_nand4_1 _16413_ (.B(_09617_),
    .C(_09618_),
    .A(_09616_),
    .Y(_09620_),
    .D(_09619_));
 sg13g2_xor2_1 _16414_ (.B(_09620_),
    .A(_09614_),
    .X(_09621_));
 sg13g2_mux4_1 _16415_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .S1(net700),
    .X(_09622_));
 sg13g2_mux4_1 _16416_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .S1(net700),
    .X(_09623_));
 sg13g2_mux4_1 _16417_ (.S0(net801),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .S1(net697),
    .X(_09624_));
 sg13g2_mux4_1 _16418_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .S1(net700),
    .X(_09625_));
 sg13g2_mux4_1 _16419_ (.S0(net804),
    .A0(_09622_),
    .A1(_09623_),
    .A2(_09624_),
    .A3(_09625_),
    .S1(net928),
    .X(_09626_));
 sg13g2_nand2_1 _16420_ (.Y(_09627_),
    .A(net713),
    .B(_09626_));
 sg13g2_mux4_1 _16421_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .S1(net700),
    .X(_09628_));
 sg13g2_mux4_1 _16422_ (.S0(net806),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .S1(net700),
    .X(_09629_));
 sg13g2_mux4_1 _16423_ (.S0(_09599_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .S1(_09600_),
    .X(_09630_));
 sg13g2_mux4_1 _16424_ (.S0(_09599_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .S1(_09600_),
    .X(_09631_));
 sg13g2_mux4_1 _16425_ (.S0(net804),
    .A0(_09628_),
    .A1(_09629_),
    .A2(_09630_),
    .A3(_09631_),
    .S1(net928),
    .X(_09632_));
 sg13g2_nand2_1 _16426_ (.Y(_09633_),
    .A(net708),
    .B(_09632_));
 sg13g2_a21oi_2 _16427_ (.B1(_08540_),
    .Y(_09634_),
    .A2(_09633_),
    .A1(_09627_));
 sg13g2_buf_1 _16428_ (.A(_09634_),
    .X(_09635_));
 sg13g2_mux2_1 _16429_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(\cpu.dcache.r_tag[7][21] ),
    .S(net816),
    .X(_09636_));
 sg13g2_nand2b_1 _16430_ (.Y(_09637_),
    .B(_09636_),
    .A_N(_09341_));
 sg13g2_mux2_1 _16431_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(\cpu.dcache.r_tag[3][21] ),
    .S(net816),
    .X(_09638_));
 sg13g2_mux2_1 _16432_ (.A0(\cpu.dcache.r_tag[4][21] ),
    .A1(\cpu.dcache.r_tag[6][21] ),
    .S(_09189_),
    .X(_09639_));
 sg13g2_a22oi_1 _16433_ (.Y(_09640_),
    .B1(_09639_),
    .B2(_09346_),
    .A2(_09638_),
    .A1(_09338_));
 sg13g2_buf_1 _16434_ (.A(net707),
    .X(_09641_));
 sg13g2_a22oi_1 _16435_ (.Y(_09642_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][21] ),
    .A2(_09641_),
    .A1(\cpu.dcache.r_tag[0][21] ));
 sg13g2_nand3_1 _16436_ (.B(_09640_),
    .C(_09642_),
    .A(_09637_),
    .Y(_09643_));
 sg13g2_xor2_1 _16437_ (.B(_09643_),
    .A(net387),
    .X(_09644_));
 sg13g2_mux4_1 _16438_ (.S0(_09396_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .S1(net812),
    .X(_09645_));
 sg13g2_mux4_1 _16439_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .S1(net812),
    .X(_09646_));
 sg13g2_mux4_1 _16440_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .S1(net810),
    .X(_09647_));
 sg13g2_mux4_1 _16441_ (.S0(_09306_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .S1(_09314_),
    .X(_09648_));
 sg13g2_mux4_1 _16442_ (.S0(net804),
    .A0(_09645_),
    .A1(_09646_),
    .A2(_09647_),
    .A3(_09648_),
    .S1(net928),
    .X(_09649_));
 sg13g2_nand2_1 _16443_ (.Y(_09650_),
    .A(net713),
    .B(_09649_));
 sg13g2_mux4_1 _16444_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .S1(net812),
    .X(_09651_));
 sg13g2_mux4_1 _16445_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .S1(net812),
    .X(_09652_));
 sg13g2_mux4_1 _16446_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .S1(net810),
    .X(_09653_));
 sg13g2_mux4_1 _16447_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .S1(net810),
    .X(_09654_));
 sg13g2_mux4_1 _16448_ (.S0(net804),
    .A0(_09651_),
    .A1(_09652_),
    .A2(_09653_),
    .A3(_09654_),
    .S1(net928),
    .X(_09655_));
 sg13g2_nand2_1 _16449_ (.Y(_09656_),
    .A(_09323_),
    .B(_09655_));
 sg13g2_a21oi_2 _16450_ (.B1(_08540_),
    .Y(_09657_),
    .A2(_09656_),
    .A1(_09650_));
 sg13g2_buf_1 _16451_ (.A(_09657_),
    .X(_09658_));
 sg13g2_inv_1 _16452_ (.Y(_09659_),
    .A(_00241_));
 sg13g2_a22oi_1 _16453_ (.Y(_09660_),
    .B1(net641),
    .B2(\cpu.dcache.r_tag[2][18] ),
    .A2(net707),
    .A1(_09659_));
 sg13g2_a22oi_1 _16454_ (.Y(_09661_),
    .B1(net705),
    .B2(\cpu.dcache.r_tag[1][18] ),
    .A2(_09349_),
    .A1(\cpu.dcache.r_tag[6][18] ));
 sg13g2_a22oi_1 _16455_ (.Y(_09662_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[7][18] ),
    .A2(net706),
    .A1(\cpu.dcache.r_tag[5][18] ));
 sg13g2_a22oi_1 _16456_ (.Y(_09663_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[4][18] ),
    .A2(net642),
    .A1(\cpu.dcache.r_tag[3][18] ));
 sg13g2_nand4_1 _16457_ (.B(_09661_),
    .C(_09662_),
    .A(_09660_),
    .Y(_09664_),
    .D(_09663_));
 sg13g2_xnor2_1 _16458_ (.Y(_09665_),
    .A(net445),
    .B(_09664_));
 sg13g2_mux4_1 _16459_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .S1(net810),
    .X(_09666_));
 sg13g2_mux4_1 _16460_ (.S0(net807),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .S1(net810),
    .X(_09667_));
 sg13g2_buf_1 _16461_ (.A(_08360_),
    .X(_09668_));
 sg13g2_mux4_1 _16462_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .S1(net800),
    .X(_09669_));
 sg13g2_mux4_1 _16463_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .S1(net800),
    .X(_09670_));
 sg13g2_mux4_1 _16464_ (.S0(net948),
    .A0(_09666_),
    .A1(_09667_),
    .A2(_09669_),
    .A3(_09670_),
    .S1(net928),
    .X(_09671_));
 sg13g2_nand2_1 _16465_ (.Y(_09672_),
    .A(net713),
    .B(_09671_));
 sg13g2_mux4_1 _16466_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .S1(net810),
    .X(_09673_));
 sg13g2_mux4_1 _16467_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .S1(net810),
    .X(_09674_));
 sg13g2_mux4_1 _16468_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .S1(net800),
    .X(_09675_));
 sg13g2_mux4_1 _16469_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .S1(net800),
    .X(_09676_));
 sg13g2_mux4_1 _16470_ (.S0(net948),
    .A0(_09673_),
    .A1(_09674_),
    .A2(_09675_),
    .A3(_09676_),
    .S1(net1086),
    .X(_09677_));
 sg13g2_nand2_1 _16471_ (.Y(_09678_),
    .A(net708),
    .B(_09677_));
 sg13g2_a21oi_2 _16472_ (.B1(_08540_),
    .Y(_09679_),
    .A2(_09678_),
    .A1(_09672_));
 sg13g2_buf_1 _16473_ (.A(_09679_),
    .X(_09680_));
 sg13g2_a22oi_1 _16474_ (.Y(_09681_),
    .B1(_09370_),
    .B2(\cpu.dcache.r_tag[2][20] ),
    .A2(_09340_),
    .A1(\cpu.dcache.r_tag[0][20] ));
 sg13g2_a22oi_1 _16475_ (.Y(_09682_),
    .B1(net644),
    .B2(\cpu.dcache.r_tag[6][20] ),
    .A2(_09343_),
    .A1(\cpu.dcache.r_tag[5][20] ));
 sg13g2_a22oi_1 _16476_ (.Y(_09683_),
    .B1(net703),
    .B2(\cpu.dcache.r_tag[7][20] ),
    .A2(_09360_),
    .A1(\cpu.dcache.r_tag[3][20] ));
 sg13g2_a22oi_1 _16477_ (.Y(_09684_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[4][20] ),
    .A2(_09353_),
    .A1(\cpu.dcache.r_tag[1][20] ));
 sg13g2_nand4_1 _16478_ (.B(_09682_),
    .C(_09683_),
    .A(_09681_),
    .Y(_09685_),
    .D(_09684_));
 sg13g2_xnor2_1 _16479_ (.Y(_09686_),
    .A(net444),
    .B(_09685_));
 sg13g2_mux4_1 _16480_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .S1(_09668_),
    .X(_09687_));
 sg13g2_mux4_1 _16481_ (.S0(net813),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .S1(net810),
    .X(_09688_));
 sg13g2_mux4_1 _16482_ (.S0(_09312_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .S1(net800),
    .X(_09689_));
 sg13g2_mux4_1 _16483_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .S1(net800),
    .X(_09690_));
 sg13g2_mux4_1 _16484_ (.S0(_08366_),
    .A0(_09687_),
    .A1(_09688_),
    .A2(_09689_),
    .A3(_09690_),
    .S1(_08278_),
    .X(_09691_));
 sg13g2_nand2_1 _16485_ (.Y(_09692_),
    .A(net713),
    .B(_09691_));
 sg13g2_mux4_1 _16486_ (.S0(_09312_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .S1(_09668_),
    .X(_09693_));
 sg13g2_mux4_1 _16487_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .S1(net800),
    .X(_09694_));
 sg13g2_mux4_1 _16488_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .S1(net802),
    .X(_09695_));
 sg13g2_mux4_1 _16489_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .S1(net802),
    .X(_09696_));
 sg13g2_mux4_1 _16490_ (.S0(_08366_),
    .A0(_09693_),
    .A1(_09694_),
    .A2(_09695_),
    .A3(_09696_),
    .S1(net1086),
    .X(_09697_));
 sg13g2_nand2_1 _16491_ (.Y(_09698_),
    .A(_08368_),
    .B(_09697_));
 sg13g2_a21oi_2 _16492_ (.B1(_08540_),
    .Y(_09699_),
    .A2(_09698_),
    .A1(_09692_));
 sg13g2_buf_1 _16493_ (.A(_09699_),
    .X(_09700_));
 sg13g2_nand2_1 _16494_ (.Y(_09701_),
    .A(\cpu.dcache.r_tag[6][22] ),
    .B(_09348_));
 sg13g2_a22oi_1 _16495_ (.Y(_09702_),
    .B1(_09369_),
    .B2(\cpu.dcache.r_tag[2][22] ),
    .A2(_09362_),
    .A1(\cpu.dcache.r_tag[4][22] ));
 sg13g2_a22oi_1 _16496_ (.Y(_09703_),
    .B1(_09366_),
    .B2(\cpu.dcache.r_tag[7][22] ),
    .A2(_09359_),
    .A1(\cpu.dcache.r_tag[3][22] ));
 sg13g2_a22oi_1 _16497_ (.Y(_09704_),
    .B1(_09353_),
    .B2(\cpu.dcache.r_tag[1][22] ),
    .A2(_09342_),
    .A1(\cpu.dcache.r_tag[5][22] ));
 sg13g2_nand4_1 _16498_ (.B(_09702_),
    .C(_09703_),
    .A(_09701_),
    .Y(_09705_),
    .D(_09704_));
 sg13g2_mux2_1 _16499_ (.A0(\cpu.dcache.r_tag[0][22] ),
    .A1(_09705_),
    .S(_09460_),
    .X(_09706_));
 sg13g2_xnor2_1 _16500_ (.Y(_09707_),
    .A(_09700_),
    .B(_09706_));
 sg13g2_inv_1 _16501_ (.Y(_09708_),
    .A(_00238_));
 sg13g2_a22oi_1 _16502_ (.Y(_09709_),
    .B1(_09370_),
    .B2(\cpu.dcache.r_tag[2][15] ),
    .A2(_09340_),
    .A1(_09708_));
 sg13g2_a22oi_1 _16503_ (.Y(_09710_),
    .B1(net705),
    .B2(\cpu.dcache.r_tag[1][15] ),
    .A2(_09348_),
    .A1(\cpu.dcache.r_tag[6][15] ));
 sg13g2_a22oi_1 _16504_ (.Y(_09711_),
    .B1(_09366_),
    .B2(\cpu.dcache.r_tag[7][15] ),
    .A2(_09343_),
    .A1(\cpu.dcache.r_tag[5][15] ));
 sg13g2_a22oi_1 _16505_ (.Y(_09712_),
    .B1(net704),
    .B2(\cpu.dcache.r_tag[4][15] ),
    .A2(net642),
    .A1(\cpu.dcache.r_tag[3][15] ));
 sg13g2_nand4_1 _16506_ (.B(_09710_),
    .C(_09711_),
    .A(_09709_),
    .Y(_09713_),
    .D(_09712_));
 sg13g2_mux4_1 _16507_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .S1(net802),
    .X(_09714_));
 sg13g2_mux4_1 _16508_ (.S0(_09525_),
    .A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .S1(_09526_),
    .X(_09715_));
 sg13g2_mux4_1 _16509_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .S1(net805),
    .X(_09716_));
 sg13g2_mux4_1 _16510_ (.S0(net927),
    .A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .S1(net805),
    .X(_09717_));
 sg13g2_mux4_1 _16511_ (.S0(_08368_),
    .A0(_09714_),
    .A1(_09715_),
    .A2(_09716_),
    .A3(_09717_),
    .S1(_09435_),
    .X(_09718_));
 sg13g2_nand2_1 _16512_ (.Y(_09719_),
    .A(net1165),
    .B(_09718_));
 sg13g2_mux4_1 _16513_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .S1(net802),
    .X(_09720_));
 sg13g2_mux4_1 _16514_ (.S0(net811),
    .A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .S1(net800),
    .X(_09721_));
 sg13g2_mux4_1 _16515_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .S1(net802),
    .X(_09722_));
 sg13g2_mux4_1 _16516_ (.S0(net803),
    .A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A2(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A3(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .S1(net802),
    .X(_09723_));
 sg13g2_mux4_1 _16517_ (.S0(_08368_),
    .A0(_09720_),
    .A1(_09721_),
    .A2(_09722_),
    .A3(_09723_),
    .S1(_09435_),
    .X(_09724_));
 sg13g2_o21ai_1 _16518_ (.B1(net808),
    .Y(_09725_),
    .A1(_08336_),
    .A2(_09724_));
 sg13g2_o21ai_1 _16519_ (.B1(_09725_),
    .Y(_09726_),
    .A1(net808),
    .A2(_09719_));
 sg13g2_buf_1 _16520_ (.A(_09726_),
    .X(_09727_));
 sg13g2_xnor2_1 _16521_ (.Y(_09728_),
    .A(_09713_),
    .B(net442));
 sg13g2_nand4_1 _16522_ (.B(_09686_),
    .C(_09707_),
    .A(_09665_),
    .Y(_09729_),
    .D(_09728_));
 sg13g2_nor4_1 _16523_ (.A(_09598_),
    .B(_09621_),
    .C(_09644_),
    .D(_09729_),
    .Y(_09730_));
 sg13g2_nand4_1 _16524_ (.B(_09452_),
    .C(_09510_),
    .A(_09421_),
    .Y(_09731_),
    .D(_09730_));
 sg13g2_mux4_1 _16525_ (.S0(_09175_),
    .A0(\cpu.dcache.r_valid[4] ),
    .A1(\cpu.dcache.r_valid[5] ),
    .A2(\cpu.dcache.r_valid[6] ),
    .A3(\cpu.dcache.r_valid[7] ),
    .S1(net715),
    .X(_09732_));
 sg13g2_mux4_1 _16526_ (.S0(net932),
    .A0(\cpu.dcache.r_valid[0] ),
    .A1(\cpu.dcache.r_valid[1] ),
    .A2(\cpu.dcache.r_valid[2] ),
    .A3(\cpu.dcache.r_valid[3] ),
    .S1(net715),
    .X(_09733_));
 sg13g2_mux2_1 _16527_ (.A0(_09732_),
    .A1(_09733_),
    .S(_09454_),
    .X(_09734_));
 sg13g2_mux4_1 _16528_ (.S0(net817),
    .A0(\cpu.dcache.r_dirty[4] ),
    .A1(\cpu.dcache.r_dirty[5] ),
    .A2(\cpu.dcache.r_dirty[6] ),
    .A3(\cpu.dcache.r_dirty[7] ),
    .S1(net715),
    .X(_09735_));
 sg13g2_mux4_1 _16529_ (.S0(_09175_),
    .A0(\cpu.dcache.r_dirty[0] ),
    .A1(\cpu.dcache.r_dirty[1] ),
    .A2(\cpu.dcache.r_dirty[2] ),
    .A3(\cpu.dcache.r_dirty[3] ),
    .S1(net715),
    .X(_09736_));
 sg13g2_mux2_1 _16530_ (.A0(_09735_),
    .A1(_09736_),
    .S(_09454_),
    .X(_09737_));
 sg13g2_and4_1 _16531_ (.A(_09109_),
    .B(_09162_),
    .C(_09734_),
    .D(_09737_),
    .X(_09738_));
 sg13g2_o21ai_1 _16532_ (.B1(_09738_),
    .Y(_09739_),
    .A1(_09303_),
    .A2(_09731_));
 sg13g2_buf_1 _16533_ (.A(_09739_),
    .X(_09740_));
 sg13g2_inv_1 _16534_ (.Y(_09741_),
    .A(_09740_));
 sg13g2_nor2b_1 _16535_ (.A(_09731_),
    .B_N(_09734_),
    .Y(_09742_));
 sg13g2_nor3_1 _16536_ (.A(_09303_),
    .B(_09738_),
    .C(_09742_),
    .Y(_09743_));
 sg13g2_buf_1 _16537_ (.A(_09743_),
    .X(_09744_));
 sg13g2_buf_1 _16538_ (.A(_09109_),
    .X(_09745_));
 sg13g2_nand3_1 _16539_ (.B(net350),
    .C(_09162_),
    .A(net1067),
    .Y(_09746_));
 sg13g2_buf_1 _16540_ (.A(_09746_),
    .X(_09747_));
 sg13g2_a21oi_1 _16541_ (.A1(_08355_),
    .A2(_08383_),
    .Y(_09748_),
    .B1(_09747_));
 sg13g2_o21ai_1 _16542_ (.B1(_09748_),
    .Y(_09749_),
    .A1(_09741_),
    .A2(_09744_));
 sg13g2_or2_1 _16543_ (.X(_09750_),
    .B(_08744_),
    .A(_08784_));
 sg13g2_nand4_1 _16544_ (.B(_08828_),
    .C(_08803_),
    .A(_08794_),
    .Y(_09751_),
    .D(_08836_));
 sg13g2_nand4_1 _16545_ (.B(_08844_),
    .C(_08817_),
    .A(_08813_),
    .Y(_09752_),
    .D(_08853_));
 sg13g2_nor4_1 _16546_ (.A(_09750_),
    .B(_08578_),
    .C(_09751_),
    .D(_09752_),
    .Y(_09753_));
 sg13g2_inv_1 _16547_ (.Y(_09754_),
    .A(_08764_));
 sg13g2_nor4_1 _16548_ (.A(_08604_),
    .B(_08679_),
    .C(_08699_),
    .D(_09754_),
    .Y(_09755_));
 sg13g2_nor3_1 _16549_ (.A(_08629_),
    .B(_08655_),
    .C(_08719_),
    .Y(_09756_));
 sg13g2_nand4_1 _16550_ (.B(_09753_),
    .C(_09755_),
    .A(_08539_),
    .Y(_09757_),
    .D(_09756_));
 sg13g2_nand2_1 _16551_ (.Y(_09758_),
    .A(net1164),
    .B(_09757_));
 sg13g2_nand3_1 _16552_ (.B(_09749_),
    .C(_09758_),
    .A(\cpu.qspi.r_state[17] ),
    .Y(_09759_));
 sg13g2_buf_1 _16553_ (.A(_09759_),
    .X(_09760_));
 sg13g2_buf_1 _16554_ (.A(\cpu.qspi.r_state[7] ),
    .X(_09761_));
 sg13g2_buf_2 _16555_ (.A(\cpu.qspi.r_ind ),
    .X(_09762_));
 sg13g2_buf_1 _16556_ (.A(\cpu.qspi.r_count[0] ),
    .X(_09763_));
 sg13g2_buf_2 _16557_ (.A(\cpu.qspi.r_count[1] ),
    .X(_09764_));
 sg13g2_buf_1 _16558_ (.A(\cpu.qspi.r_count[2] ),
    .X(_09765_));
 sg13g2_nor4_2 _16559_ (.A(_09763_),
    .B(_09764_),
    .C(\cpu.qspi.r_count[3] ),
    .Y(_09766_),
    .D(_09765_));
 sg13g2_and2_1 _16560_ (.A(_00244_),
    .B(_09766_),
    .X(_09767_));
 sg13g2_buf_1 _16561_ (.A(_09767_),
    .X(_09768_));
 sg13g2_buf_1 _16562_ (.A(\cpu.qspi.r_state[2] ),
    .X(_09769_));
 sg13g2_buf_1 _16563_ (.A(\cpu.qspi.r_state[1] ),
    .X(_09770_));
 sg13g2_a221oi_1 _16564_ (.B2(_09769_),
    .C1(_09770_),
    .B1(_09768_),
    .A1(_09761_),
    .Y(_09771_),
    .A2(_09762_));
 sg13g2_buf_2 _16565_ (.A(net815),
    .X(_09772_));
 sg13g2_buf_1 _16566_ (.A(_09772_),
    .X(_09773_));
 sg13g2_a21oi_1 _16567_ (.A1(_09760_),
    .A2(_09771_),
    .Y(_00026_),
    .B1(_09773_));
 sg13g2_buf_1 _16568_ (.A(\cpu.qspi.r_state[16] ),
    .X(_09774_));
 sg13g2_nand2_1 _16569_ (.Y(_09775_),
    .A(_00244_),
    .B(_09766_));
 sg13g2_buf_1 _16570_ (.A(_09775_),
    .X(_09776_));
 sg13g2_nor2_1 _16571_ (.A(net1164),
    .B(_09740_),
    .Y(_09777_));
 sg13g2_buf_8 _16572_ (.A(_09777_),
    .X(_09778_));
 sg13g2_buf_2 _16573_ (.A(\cpu.qspi.r_state[8] ),
    .X(_09779_));
 sg13g2_a22oi_1 _16574_ (.Y(_09780_),
    .B1(_09778_),
    .B2(_09779_),
    .A2(net799),
    .A1(net1149));
 sg13g2_nor2_1 _16575_ (.A(_09269_),
    .B(_09780_),
    .Y(_00025_));
 sg13g2_buf_1 _16576_ (.A(\cpu.qspi.r_state[4] ),
    .X(_09781_));
 sg13g2_buf_1 _16577_ (.A(\cpu.qspi.r_state[9] ),
    .X(_09782_));
 sg13g2_a21oi_1 _16578_ (.A1(_09781_),
    .A2(_09768_),
    .Y(_09783_),
    .B1(_09782_));
 sg13g2_nor2_1 _16579_ (.A(net647),
    .B(_09783_),
    .Y(_00022_));
 sg13g2_buf_1 _16580_ (.A(_00270_),
    .X(_09784_));
 sg13g2_buf_1 _16581_ (.A(\cpu.qspi.r_state[12] ),
    .X(_09785_));
 sg13g2_nand2_1 _16582_ (.Y(_09786_),
    .A(_09785_),
    .B(net799));
 sg13g2_a21oi_1 _16583_ (.A1(_09784_),
    .A2(_09786_),
    .Y(_00023_),
    .B1(_09773_));
 sg13g2_buf_1 _16584_ (.A(\cpu.qspi.r_rom_mode[1] ),
    .X(_09787_));
 sg13g2_buf_1 _16585_ (.A(\cpu.qspi.r_rom_mode[0] ),
    .X(_09788_));
 sg13g2_inv_1 _16586_ (.Y(_09789_),
    .A(_09614_));
 sg13g2_or2_1 _16587_ (.X(_09790_),
    .B(_08777_),
    .A(net950));
 sg13g2_o21ai_1 _16588_ (.B1(_09790_),
    .Y(_09791_),
    .A1(net1164),
    .A2(_09789_));
 sg13g2_nor2_1 _16589_ (.A(_09788_),
    .B(_09791_),
    .Y(_09792_));
 sg13g2_a21oi_1 _16590_ (.A1(_09788_),
    .A2(_09778_),
    .Y(_09793_),
    .B1(_09792_));
 sg13g2_and2_1 _16591_ (.A(_09787_),
    .B(_09793_),
    .X(_09794_));
 sg13g2_buf_8 _16592_ (.A(_09794_),
    .X(_09795_));
 sg13g2_inv_1 _16593_ (.Y(_09796_),
    .A(_09791_));
 sg13g2_nor3_1 _16594_ (.A(_09788_),
    .B(_09787_),
    .C(_09796_),
    .Y(_09797_));
 sg13g2_buf_2 _16595_ (.A(_09797_),
    .X(_09798_));
 sg13g2_nor2_1 _16596_ (.A(_09798_),
    .B(_09795_),
    .Y(_09799_));
 sg13g2_buf_2 _16597_ (.A(_09799_),
    .X(_09800_));
 sg13g2_and2_1 _16598_ (.A(\cpu.qspi.r_quad[2] ),
    .B(_09798_),
    .X(_09801_));
 sg13g2_a221oi_1 _16599_ (.B2(\cpu.qspi.r_quad[0] ),
    .C1(_09801_),
    .B1(_09800_),
    .A1(\cpu.qspi.r_quad[1] ),
    .Y(_09802_),
    .A2(_09795_));
 sg13g2_buf_2 _16600_ (.A(_09802_),
    .X(_09803_));
 sg13g2_inv_1 _16601_ (.Y(_09804_),
    .A(\cpu.qspi.r_state[17] ));
 sg13g2_a21oi_1 _16602_ (.A1(_09749_),
    .A2(_09758_),
    .Y(_09805_),
    .B1(_09804_));
 sg13g2_a22oi_1 _16603_ (.Y(_09806_),
    .B1(_09803_),
    .B2(_09805_),
    .A2(net799),
    .A1(_09781_));
 sg13g2_nor2_1 _16604_ (.A(net647),
    .B(_09806_),
    .Y(_00028_));
 sg13g2_buf_1 _16605_ (.A(\cpu.qspi.r_state[14] ),
    .X(_09807_));
 sg13g2_and2_1 _16606_ (.A(_09769_),
    .B(_09775_),
    .X(_09808_));
 sg13g2_buf_1 _16607_ (.A(_09808_),
    .X(_09809_));
 sg13g2_a21oi_1 _16608_ (.A1(_09807_),
    .A2(_09768_),
    .Y(_09810_),
    .B1(_09809_));
 sg13g2_nor2_1 _16609_ (.A(net647),
    .B(_09810_),
    .Y(_00027_));
 sg13g2_inv_1 _16610_ (.Y(_09811_),
    .A(_09761_));
 sg13g2_buf_1 _16611_ (.A(net818),
    .X(_09812_));
 sg13g2_o21ai_1 _16612_ (.B1(net696),
    .Y(_00021_),
    .A1(_09811_),
    .A2(_09762_));
 sg13g2_buf_2 _16613_ (.A(\cpu.dec.r_op[1] ),
    .X(_09813_));
 sg13g2_nor4_1 _16614_ (.A(net114),
    .B(net304),
    .C(_08908_),
    .D(_09079_),
    .Y(_09814_));
 sg13g2_a21o_1 _16615_ (.A2(_08861_),
    .A1(_09813_),
    .B1(_09814_),
    .X(_00012_));
 sg13g2_buf_1 _16616_ (.A(\cpu.dec.r_op[10] ),
    .X(_09815_));
 sg13g2_nand2_1 _16617_ (.Y(_09816_),
    .A(net356),
    .B(net355));
 sg13g2_nor3_1 _16618_ (.A(net113),
    .B(_09013_),
    .C(_09816_),
    .Y(_09817_));
 sg13g2_a21o_1 _16619_ (.A2(_08861_),
    .A1(_09815_),
    .B1(_09817_),
    .X(_00011_));
 sg13g2_buf_1 _16620_ (.A(\cpu.dec.r_op[9] ),
    .X(_09818_));
 sg13g2_buf_1 _16621_ (.A(net1145),
    .X(_09819_));
 sg13g2_buf_1 _16622_ (.A(net114),
    .X(_09820_));
 sg13g2_inv_1 _16623_ (.Y(_09821_),
    .A(_08931_));
 sg13g2_nor2_1 _16624_ (.A(_08948_),
    .B(_08969_),
    .Y(_09822_));
 sg13g2_buf_2 _16625_ (.A(_09822_),
    .X(_09823_));
 sg13g2_nand2_1 _16626_ (.Y(_09824_),
    .A(_09821_),
    .B(_09823_));
 sg13g2_buf_1 _16627_ (.A(_09824_),
    .X(_09825_));
 sg13g2_buf_1 _16628_ (.A(_08991_),
    .X(_09826_));
 sg13g2_buf_1 _16629_ (.A(net236),
    .X(_09827_));
 sg13g2_nor3_1 _16630_ (.A(_09089_),
    .B(_08908_),
    .C(_09088_),
    .Y(_09828_));
 sg13g2_nor2_1 _16631_ (.A(_09827_),
    .B(_09097_),
    .Y(_09829_));
 sg13g2_a21oi_1 _16632_ (.A1(_09827_),
    .A2(_09828_),
    .Y(_09830_),
    .B1(_09829_));
 sg13g2_nor4_1 _16633_ (.A(_08860_),
    .B(net156),
    .C(net186),
    .D(_09830_),
    .Y(_09831_));
 sg13g2_a21o_1 _16634_ (.A2(net92),
    .A1(net1063),
    .B1(_09831_),
    .X(_00020_));
 sg13g2_buf_2 _16635_ (.A(\cpu.qspi.r_state[5] ),
    .X(_09832_));
 sg13g2_a21oi_1 _16636_ (.A1(net1147),
    .A2(net799),
    .Y(_09833_),
    .B1(_09832_));
 sg13g2_nor2_1 _16637_ (.A(_09269_),
    .B(_09833_),
    .Y(_00024_));
 sg13g2_inv_1 _16638_ (.Y(_09834_),
    .A(_08948_));
 sg13g2_nand2_1 _16639_ (.Y(_09835_),
    .A(_08931_),
    .B(_09834_));
 sg13g2_buf_1 _16640_ (.A(_09835_),
    .X(_09836_));
 sg13g2_nor2_1 _16641_ (.A(net263),
    .B(_09836_),
    .Y(_09837_));
 sg13g2_buf_1 _16642_ (.A(_09837_),
    .X(_09838_));
 sg13g2_a21o_1 _16643_ (.A2(_08980_),
    .A1(net819),
    .B1(_08989_),
    .X(_09839_));
 sg13g2_buf_1 _16644_ (.A(_09839_),
    .X(_09840_));
 sg13g2_nor2_1 _16645_ (.A(_09840_),
    .B(net236),
    .Y(_09841_));
 sg13g2_buf_1 _16646_ (.A(_09841_),
    .X(_09842_));
 sg13g2_nand2_1 _16647_ (.Y(_09843_),
    .A(net155),
    .B(_09842_));
 sg13g2_buf_2 _16648_ (.A(\cpu.dec.r_op[8] ),
    .X(_09844_));
 sg13g2_buf_1 _16649_ (.A(_09844_),
    .X(_09845_));
 sg13g2_nand2_1 _16650_ (.Y(_09846_),
    .A(net1062),
    .B(net112));
 sg13g2_o21ai_1 _16651_ (.B1(_09846_),
    .Y(_00019_),
    .A1(net93),
    .A2(_09843_));
 sg13g2_buf_1 _16652_ (.A(\cpu.uart.r_div[11] ),
    .X(_09847_));
 sg13g2_nor3_1 _16653_ (.A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ),
    .C(\cpu.uart.r_div[2] ),
    .Y(_09848_));
 sg13g2_nor2b_1 _16654_ (.A(\cpu.uart.r_div[3] ),
    .B_N(_09848_),
    .Y(_09849_));
 sg13g2_nor2b_1 _16655_ (.A(\cpu.uart.r_div[4] ),
    .B_N(_09849_),
    .Y(_09850_));
 sg13g2_nor2b_1 _16656_ (.A(\cpu.uart.r_div[5] ),
    .B_N(_09850_),
    .Y(_09851_));
 sg13g2_nor2b_1 _16657_ (.A(\cpu.uart.r_div[6] ),
    .B_N(_09851_),
    .Y(_09852_));
 sg13g2_nand2b_1 _16658_ (.Y(_09853_),
    .B(_09852_),
    .A_N(\cpu.uart.r_div[7] ));
 sg13g2_nor2_1 _16659_ (.A(\cpu.uart.r_div[8] ),
    .B(_09853_),
    .Y(_09854_));
 sg13g2_nand2b_1 _16660_ (.Y(_09855_),
    .B(_09854_),
    .A_N(\cpu.uart.r_div[9] ));
 sg13g2_buf_1 _16661_ (.A(_09855_),
    .X(_09856_));
 sg13g2_nor3_2 _16662_ (.A(_09847_),
    .B(\cpu.uart.r_div[10] ),
    .C(_09856_),
    .Y(_09857_));
 sg13g2_buf_1 _16663_ (.A(_09857_),
    .X(_09858_));
 sg13g2_nor2_1 _16664_ (.A(net929),
    .B(net349),
    .Y(_09859_));
 sg13g2_buf_1 _16665_ (.A(_09859_),
    .X(_09860_));
 sg13g2_buf_1 _16666_ (.A(net262),
    .X(_09861_));
 sg13g2_mux2_1 _16667_ (.A0(\cpu.uart.r_div_value[0] ),
    .A1(_00272_),
    .S(_09861_),
    .X(_00079_));
 sg13g2_xnor2_1 _16668_ (.Y(_09862_),
    .A(\cpu.uart.r_div[0] ),
    .B(\cpu.uart.r_div[1] ));
 sg13g2_mux2_1 _16669_ (.A0(\cpu.uart.r_div_value[1] ),
    .A1(_09862_),
    .S(net235),
    .X(_00082_));
 sg13g2_o21ai_1 _16670_ (.B1(\cpu.uart.r_div[2] ),
    .Y(_09863_),
    .A1(\cpu.uart.r_div[0] ),
    .A2(\cpu.uart.r_div[1] ));
 sg13g2_nor2b_1 _16671_ (.A(_09848_),
    .B_N(_09863_),
    .Y(_09864_));
 sg13g2_nor2_1 _16672_ (.A(\cpu.uart.r_div_value[2] ),
    .B(net262),
    .Y(_09865_));
 sg13g2_a21oi_1 _16673_ (.A1(_09861_),
    .A2(_09864_),
    .Y(_00083_),
    .B1(_09865_));
 sg13g2_xnor2_1 _16674_ (.Y(_09866_),
    .A(\cpu.uart.r_div[3] ),
    .B(_09848_));
 sg13g2_nor2_1 _16675_ (.A(\cpu.uart.r_div_value[3] ),
    .B(_09860_),
    .Y(_09867_));
 sg13g2_a21oi_1 _16676_ (.A1(net235),
    .A2(_09866_),
    .Y(_00084_),
    .B1(_09867_));
 sg13g2_xnor2_1 _16677_ (.Y(_09868_),
    .A(\cpu.uart.r_div[4] ),
    .B(_09849_));
 sg13g2_nor2_1 _16678_ (.A(\cpu.uart.r_div_value[4] ),
    .B(net262),
    .Y(_09869_));
 sg13g2_a21oi_1 _16679_ (.A1(net235),
    .A2(_09868_),
    .Y(_00085_),
    .B1(_09869_));
 sg13g2_xnor2_1 _16680_ (.Y(_09870_),
    .A(\cpu.uart.r_div[5] ),
    .B(_09850_));
 sg13g2_nor2_1 _16681_ (.A(\cpu.uart.r_div_value[5] ),
    .B(net262),
    .Y(_09871_));
 sg13g2_a21oi_1 _16682_ (.A1(net235),
    .A2(_09870_),
    .Y(_00086_),
    .B1(_09871_));
 sg13g2_xnor2_1 _16683_ (.Y(_09872_),
    .A(\cpu.uart.r_div[6] ),
    .B(_09851_));
 sg13g2_nor2_1 _16684_ (.A(\cpu.uart.r_div_value[6] ),
    .B(net262),
    .Y(_09873_));
 sg13g2_a21oi_1 _16685_ (.A1(net235),
    .A2(_09872_),
    .Y(_00087_),
    .B1(_09873_));
 sg13g2_xnor2_1 _16686_ (.Y(_09874_),
    .A(\cpu.uart.r_div[7] ),
    .B(_09852_));
 sg13g2_nor2_1 _16687_ (.A(\cpu.uart.r_div_value[7] ),
    .B(net262),
    .Y(_09875_));
 sg13g2_a21oi_1 _16688_ (.A1(net235),
    .A2(_09874_),
    .Y(_00088_),
    .B1(_09875_));
 sg13g2_xor2_1 _16689_ (.B(_09853_),
    .A(\cpu.uart.r_div[8] ),
    .X(_09876_));
 sg13g2_nor2_1 _16690_ (.A(\cpu.uart.r_div_value[8] ),
    .B(net262),
    .Y(_09877_));
 sg13g2_a21oi_1 _16691_ (.A1(net235),
    .A2(_09876_),
    .Y(_00089_),
    .B1(_09877_));
 sg13g2_xnor2_1 _16692_ (.Y(_09878_),
    .A(\cpu.uart.r_div[9] ),
    .B(_09854_));
 sg13g2_nor2_1 _16693_ (.A(\cpu.uart.r_div_value[9] ),
    .B(net262),
    .Y(_09879_));
 sg13g2_a21oi_1 _16694_ (.A1(net235),
    .A2(_09878_),
    .Y(_00090_),
    .B1(_09879_));
 sg13g2_inv_1 _16695_ (.Y(_09880_),
    .A(\cpu.uart.r_div_value[10] ));
 sg13g2_nand2_1 _16696_ (.Y(_09881_),
    .A(net933),
    .B(_09856_));
 sg13g2_o21ai_1 _16697_ (.B1(_09881_),
    .Y(_09882_),
    .A1(_09847_),
    .A2(\cpu.uart.r_div_value[10] ));
 sg13g2_inv_1 _16698_ (.Y(_09883_),
    .A(\cpu.uart.r_div[10] ));
 sg13g2_nor3_1 _16699_ (.A(_09883_),
    .B(net815),
    .C(_09856_),
    .Y(_09884_));
 sg13g2_a221oi_1 _16700_ (.B2(_09883_),
    .C1(_09884_),
    .B1(_09882_),
    .A1(_09880_),
    .Y(_00080_),
    .A2(net714));
 sg13g2_nor2_1 _16701_ (.A(\cpu.uart.r_div[10] ),
    .B(_09856_),
    .Y(_09885_));
 sg13g2_nand2_1 _16702_ (.Y(_09886_),
    .A(_09847_),
    .B(net818));
 sg13g2_o21ai_1 _16703_ (.B1(\cpu.uart.r_div_value[11] ),
    .Y(_09887_),
    .A1(net815),
    .A2(net349));
 sg13g2_o21ai_1 _16704_ (.B1(_09887_),
    .Y(_00081_),
    .A1(_09885_),
    .A2(_09886_));
 sg13g2_inv_2 _16705_ (.Y(_09888_),
    .A(_09177_));
 sg13g2_buf_1 _16706_ (.A(_09888_),
    .X(_09889_));
 sg13g2_buf_1 _16707_ (.A(net923),
    .X(_09890_));
 sg13g2_nand3_1 _16708_ (.B(net925),
    .C(_09192_),
    .A(_09176_),
    .Y(_09891_));
 sg13g2_buf_2 _16709_ (.A(_09891_),
    .X(_09892_));
 sg13g2_buf_2 _16710_ (.A(\cpu.addr[5] ),
    .X(_09893_));
 sg13g2_buf_1 _16711_ (.A(_09893_),
    .X(_09894_));
 sg13g2_nor3_1 _16712_ (.A(_09894_),
    .B(_09165_),
    .C(net1154),
    .Y(_09895_));
 sg13g2_and2_1 _16713_ (.A(_09164_),
    .B(_09895_),
    .X(_09896_));
 sg13g2_buf_1 _16714_ (.A(_09896_),
    .X(_09897_));
 sg13g2_nand2_1 _16715_ (.Y(_09898_),
    .A(_09195_),
    .B(_09897_));
 sg13g2_nor3_1 _16716_ (.A(net798),
    .B(_09892_),
    .C(_09898_),
    .Y(_09899_));
 sg13g2_buf_1 _16717_ (.A(_09899_),
    .X(_09900_));
 sg13g2_buf_1 _16718_ (.A(\cpu.intr.r_timer_count[19] ),
    .X(_09901_));
 sg13g2_buf_1 _16719_ (.A(\cpu.intr.r_timer_count[18] ),
    .X(_09902_));
 sg13g2_buf_1 _16720_ (.A(\cpu.intr.r_timer_count[17] ),
    .X(_09903_));
 sg13g2_buf_1 _16721_ (.A(\cpu.intr.r_timer_count[16] ),
    .X(_09904_));
 sg13g2_buf_1 _16722_ (.A(\cpu.intr.r_timer_count[10] ),
    .X(_09905_));
 sg13g2_buf_1 _16723_ (.A(\cpu.intr.r_timer_count[7] ),
    .X(_09906_));
 sg13g2_buf_1 _16724_ (.A(\cpu.intr.r_timer_count[1] ),
    .X(_09907_));
 sg13g2_nor3_1 _16725_ (.A(_09907_),
    .B(\cpu.intr.r_timer_count[0] ),
    .C(\cpu.intr.r_timer_count[2] ),
    .Y(_09908_));
 sg13g2_nor2b_1 _16726_ (.A(\cpu.intr.r_timer_count[3] ),
    .B_N(_09908_),
    .Y(_09909_));
 sg13g2_nor2b_1 _16727_ (.A(\cpu.intr.r_timer_count[4] ),
    .B_N(_09909_),
    .Y(_09910_));
 sg13g2_nor2b_1 _16728_ (.A(\cpu.intr.r_timer_count[5] ),
    .B_N(_09910_),
    .Y(_09911_));
 sg13g2_nand2b_1 _16729_ (.Y(_09912_),
    .B(_09911_),
    .A_N(\cpu.intr.r_timer_count[6] ));
 sg13g2_nor3_1 _16730_ (.A(_09906_),
    .B(\cpu.intr.r_timer_count[8] ),
    .C(_09912_),
    .Y(_09913_));
 sg13g2_nand2b_1 _16731_ (.Y(_09914_),
    .B(_09913_),
    .A_N(\cpu.intr.r_timer_count[9] ));
 sg13g2_nor3_1 _16732_ (.A(\cpu.intr.r_timer_count[11] ),
    .B(_09905_),
    .C(_09914_),
    .Y(_09915_));
 sg13g2_nor2b_1 _16733_ (.A(\cpu.intr.r_timer_count[12] ),
    .B_N(_09915_),
    .Y(_09916_));
 sg13g2_nor2b_1 _16734_ (.A(\cpu.intr.r_timer_count[13] ),
    .B_N(_09916_),
    .Y(_09917_));
 sg13g2_nor2b_1 _16735_ (.A(\cpu.intr.r_timer_count[14] ),
    .B_N(_09917_),
    .Y(_09918_));
 sg13g2_nand2b_2 _16736_ (.Y(_09919_),
    .B(_09918_),
    .A_N(\cpu.intr.r_timer_count[15] ));
 sg13g2_nor3_2 _16737_ (.A(_09903_),
    .B(_09904_),
    .C(_09919_),
    .Y(_09920_));
 sg13g2_nand2b_1 _16738_ (.Y(_09921_),
    .B(_09920_),
    .A_N(_09902_));
 sg13g2_or2_1 _16739_ (.X(_09922_),
    .B(_09921_),
    .A(_09901_));
 sg13g2_buf_1 _16740_ (.A(_09922_),
    .X(_09923_));
 sg13g2_buf_1 _16741_ (.A(\cpu.intr.r_timer_count[21] ),
    .X(_09924_));
 sg13g2_buf_2 _16742_ (.A(\cpu.intr.r_timer_count[20] ),
    .X(_09925_));
 sg13g2_buf_1 _16743_ (.A(\cpu.intr.r_timer_count[23] ),
    .X(_09926_));
 sg13g2_buf_1 _16744_ (.A(\cpu.intr.r_timer_count[22] ),
    .X(_09927_));
 sg13g2_nor4_2 _16745_ (.A(_09924_),
    .B(_09925_),
    .C(_09926_),
    .Y(_09928_),
    .D(_09927_));
 sg13g2_nand2b_1 _16746_ (.Y(_09929_),
    .B(_09928_),
    .A_N(_09923_));
 sg13g2_buf_2 _16747_ (.A(_09929_),
    .X(_09930_));
 sg13g2_nor2b_1 _16748_ (.A(_09900_),
    .B_N(_09930_),
    .Y(_09931_));
 sg13g2_buf_1 _16749_ (.A(_09931_),
    .X(_09932_));
 sg13g2_buf_1 _16750_ (.A(_09932_),
    .X(_09933_));
 sg13g2_mux2_1 _16751_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(_00278_),
    .S(net65),
    .X(_00055_));
 sg13g2_xnor2_1 _16752_ (.Y(_09934_),
    .A(_09907_),
    .B(\cpu.intr.r_timer_count[0] ));
 sg13g2_mux2_1 _16753_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(_09934_),
    .S(net65),
    .X(_00066_));
 sg13g2_buf_1 _16754_ (.A(_09932_),
    .X(_09935_));
 sg13g2_o21ai_1 _16755_ (.B1(\cpu.intr.r_timer_count[2] ),
    .Y(_09936_),
    .A1(_09907_),
    .A2(\cpu.intr.r_timer_count[0] ));
 sg13g2_nor2b_1 _16756_ (.A(_09908_),
    .B_N(_09936_),
    .Y(_09937_));
 sg13g2_nor2_1 _16757_ (.A(\cpu.intr.r_timer_reload[2] ),
    .B(net65),
    .Y(_09938_));
 sg13g2_a21oi_1 _16758_ (.A1(net64),
    .A2(_09937_),
    .Y(_00071_),
    .B1(_09938_));
 sg13g2_xnor2_1 _16759_ (.Y(_09939_),
    .A(\cpu.intr.r_timer_count[3] ),
    .B(_09908_));
 sg13g2_nor2_1 _16760_ (.A(\cpu.intr.r_timer_reload[3] ),
    .B(net65),
    .Y(_09940_));
 sg13g2_a21oi_1 _16761_ (.A1(net64),
    .A2(_09939_),
    .Y(_00072_),
    .B1(_09940_));
 sg13g2_xnor2_1 _16762_ (.Y(_09941_),
    .A(\cpu.intr.r_timer_count[4] ),
    .B(_09909_));
 sg13g2_nor2_1 _16763_ (.A(\cpu.intr.r_timer_reload[4] ),
    .B(net65),
    .Y(_09942_));
 sg13g2_a21oi_1 _16764_ (.A1(net64),
    .A2(_09941_),
    .Y(_00073_),
    .B1(_09942_));
 sg13g2_xnor2_1 _16765_ (.Y(_09943_),
    .A(\cpu.intr.r_timer_count[5] ),
    .B(_09910_));
 sg13g2_nor2_1 _16766_ (.A(\cpu.intr.r_timer_reload[5] ),
    .B(net65),
    .Y(_09944_));
 sg13g2_a21oi_1 _16767_ (.A1(net64),
    .A2(_09943_),
    .Y(_00074_),
    .B1(_09944_));
 sg13g2_xnor2_1 _16768_ (.Y(_09945_),
    .A(\cpu.intr.r_timer_count[6] ),
    .B(_09911_));
 sg13g2_buf_1 _16769_ (.A(_09932_),
    .X(_09946_));
 sg13g2_nor2_1 _16770_ (.A(\cpu.intr.r_timer_reload[6] ),
    .B(net63),
    .Y(_09947_));
 sg13g2_a21oi_1 _16771_ (.A1(_09935_),
    .A2(_09945_),
    .Y(_00075_),
    .B1(_09947_));
 sg13g2_xor2_1 _16772_ (.B(_09912_),
    .A(_09906_),
    .X(_09948_));
 sg13g2_nor2_1 _16773_ (.A(\cpu.intr.r_timer_reload[7] ),
    .B(net63),
    .Y(_09949_));
 sg13g2_a21oi_1 _16774_ (.A1(_09935_),
    .A2(_09948_),
    .Y(_00076_),
    .B1(_09949_));
 sg13g2_nor2_1 _16775_ (.A(_09906_),
    .B(_09912_),
    .Y(_09950_));
 sg13g2_xnor2_1 _16776_ (.Y(_09951_),
    .A(\cpu.intr.r_timer_count[8] ),
    .B(_09950_));
 sg13g2_nor2_1 _16777_ (.A(\cpu.intr.r_timer_reload[8] ),
    .B(net63),
    .Y(_09952_));
 sg13g2_a21oi_1 _16778_ (.A1(net64),
    .A2(_09951_),
    .Y(_00077_),
    .B1(_09952_));
 sg13g2_xnor2_1 _16779_ (.Y(_09953_),
    .A(\cpu.intr.r_timer_count[9] ),
    .B(_09913_));
 sg13g2_nor2_1 _16780_ (.A(\cpu.intr.r_timer_reload[9] ),
    .B(_09946_),
    .Y(_09954_));
 sg13g2_a21oi_1 _16781_ (.A1(net64),
    .A2(_09953_),
    .Y(_00078_),
    .B1(_09954_));
 sg13g2_xor2_1 _16782_ (.B(_09914_),
    .A(_09905_),
    .X(_09955_));
 sg13g2_nor2_1 _16783_ (.A(\cpu.intr.r_timer_reload[10] ),
    .B(net63),
    .Y(_09956_));
 sg13g2_a21oi_1 _16784_ (.A1(net64),
    .A2(_09955_),
    .Y(_00056_),
    .B1(_09956_));
 sg13g2_o21ai_1 _16785_ (.B1(\cpu.intr.r_timer_count[11] ),
    .Y(_09957_),
    .A1(_09905_),
    .A2(_09914_));
 sg13g2_nor2b_1 _16786_ (.A(_09915_),
    .B_N(_09957_),
    .Y(_09958_));
 sg13g2_nor2_1 _16787_ (.A(\cpu.intr.r_timer_reload[11] ),
    .B(net63),
    .Y(_09959_));
 sg13g2_a21oi_1 _16788_ (.A1(net64),
    .A2(_09958_),
    .Y(_00057_),
    .B1(_09959_));
 sg13g2_xnor2_1 _16789_ (.Y(_09960_),
    .A(\cpu.intr.r_timer_count[12] ),
    .B(_09915_));
 sg13g2_nor2_1 _16790_ (.A(\cpu.intr.r_timer_reload[12] ),
    .B(net63),
    .Y(_09961_));
 sg13g2_a21oi_1 _16791_ (.A1(net65),
    .A2(_09960_),
    .Y(_00058_),
    .B1(_09961_));
 sg13g2_xnor2_1 _16792_ (.Y(_09962_),
    .A(\cpu.intr.r_timer_count[13] ),
    .B(_09916_));
 sg13g2_nor2_1 _16793_ (.A(\cpu.intr.r_timer_reload[13] ),
    .B(_09946_),
    .Y(_09963_));
 sg13g2_a21oi_1 _16794_ (.A1(net65),
    .A2(_09962_),
    .Y(_00059_),
    .B1(_09963_));
 sg13g2_xnor2_1 _16795_ (.Y(_09964_),
    .A(\cpu.intr.r_timer_count[14] ),
    .B(_09917_));
 sg13g2_nor2_1 _16796_ (.A(\cpu.intr.r_timer_reload[14] ),
    .B(net63),
    .Y(_09965_));
 sg13g2_a21oi_1 _16797_ (.A1(_09933_),
    .A2(_09964_),
    .Y(_00060_),
    .B1(_09965_));
 sg13g2_xnor2_1 _16798_ (.Y(_09966_),
    .A(\cpu.intr.r_timer_count[15] ),
    .B(_09918_));
 sg13g2_nor2_1 _16799_ (.A(\cpu.intr.r_timer_reload[15] ),
    .B(net63),
    .Y(_09967_));
 sg13g2_a21oi_1 _16800_ (.A1(_09933_),
    .A2(_09966_),
    .Y(_00061_),
    .B1(_09967_));
 sg13g2_buf_1 _16801_ (.A(\cpu.dcache.wdata[0] ),
    .X(_09968_));
 sg13g2_inv_1 _16802_ (.Y(_09969_),
    .A(_09968_));
 sg13g2_buf_1 _16803_ (.A(_09969_),
    .X(_09970_));
 sg13g2_buf_1 _16804_ (.A(net922),
    .X(_09971_));
 sg13g2_buf_1 _16805_ (.A(_09900_),
    .X(_09972_));
 sg13g2_buf_1 _16806_ (.A(_09900_),
    .X(_09973_));
 sg13g2_nor4_1 _16807_ (.A(_09903_),
    .B(_09901_),
    .C(_09902_),
    .D(\cpu.intr.r_timer_reload[16] ),
    .Y(_09974_));
 sg13g2_a21oi_1 _16808_ (.A1(_09928_),
    .A2(_09974_),
    .Y(_09975_),
    .B1(_09904_));
 sg13g2_mux2_1 _16809_ (.A0(_09975_),
    .A1(_09904_),
    .S(_09919_),
    .X(_09976_));
 sg13g2_nor2_1 _16810_ (.A(net184),
    .B(_09976_),
    .Y(_09977_));
 sg13g2_a21oi_1 _16811_ (.A1(net797),
    .A2(net185),
    .Y(_00062_),
    .B1(_09977_));
 sg13g2_buf_2 _16812_ (.A(\cpu.dcache.wdata[1] ),
    .X(_09978_));
 sg13g2_buf_1 _16813_ (.A(_09978_),
    .X(_09979_));
 sg13g2_nor2_1 _16814_ (.A(\cpu.intr.r_timer_reload[17] ),
    .B(_09930_),
    .Y(_09980_));
 sg13g2_o21ai_1 _16815_ (.B1(_09903_),
    .Y(_09981_),
    .A1(_09904_),
    .A2(_09919_));
 sg13g2_nor2b_1 _16816_ (.A(_09920_),
    .B_N(_09981_),
    .Y(_09982_));
 sg13g2_nor3_1 _16817_ (.A(_09900_),
    .B(_09980_),
    .C(_09982_),
    .Y(_09983_));
 sg13g2_a21o_1 _16818_ (.A2(_09972_),
    .A1(net1060),
    .B1(_09983_),
    .X(_00063_));
 sg13g2_buf_1 _16819_ (.A(\cpu.dcache.wdata[2] ),
    .X(_09984_));
 sg13g2_buf_1 _16820_ (.A(_09984_),
    .X(_09985_));
 sg13g2_buf_1 _16821_ (.A(net1059),
    .X(_09986_));
 sg13g2_nor2_1 _16822_ (.A(\cpu.intr.r_timer_reload[18] ),
    .B(_09930_),
    .Y(_09987_));
 sg13g2_xnor2_1 _16823_ (.Y(_09988_),
    .A(_09902_),
    .B(_09920_));
 sg13g2_nor3_1 _16824_ (.A(_09900_),
    .B(_09987_),
    .C(_09988_),
    .Y(_09989_));
 sg13g2_a21o_1 _16825_ (.A2(net184),
    .A1(net921),
    .B1(_09989_),
    .X(_00064_));
 sg13g2_xnor2_1 _16826_ (.Y(_09990_),
    .A(_09901_),
    .B(_09921_));
 sg13g2_o21ai_1 _16827_ (.B1(_09990_),
    .Y(_09991_),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .A2(_09930_));
 sg13g2_buf_1 _16828_ (.A(\cpu.dcache.wdata[3] ),
    .X(_09992_));
 sg13g2_buf_1 _16829_ (.A(net1144),
    .X(_09993_));
 sg13g2_nand2_1 _16830_ (.Y(_09994_),
    .A(net1058),
    .B(net184));
 sg13g2_o21ai_1 _16831_ (.B1(_09994_),
    .Y(_00065_),
    .A1(net185),
    .A2(_09991_));
 sg13g2_inv_1 _16832_ (.Y(_09995_),
    .A(\cpu.intr.r_timer_reload[20] ));
 sg13g2_and2_1 _16833_ (.A(_09995_),
    .B(_09928_),
    .X(_09996_));
 sg13g2_nor3_1 _16834_ (.A(_09925_),
    .B(_09923_),
    .C(_09996_),
    .Y(_09997_));
 sg13g2_a21oi_1 _16835_ (.A1(_09925_),
    .A2(_09923_),
    .Y(_09998_),
    .B1(_09997_));
 sg13g2_buf_2 _16836_ (.A(\cpu.dcache.wdata[4] ),
    .X(_09999_));
 sg13g2_buf_1 _16837_ (.A(_09999_),
    .X(_10000_));
 sg13g2_nand2_1 _16838_ (.Y(_10001_),
    .A(net1057),
    .B(net184));
 sg13g2_o21ai_1 _16839_ (.B1(_10001_),
    .Y(_00067_),
    .A1(net185),
    .A2(_09998_));
 sg13g2_nor2_1 _16840_ (.A(_09925_),
    .B(_09923_),
    .Y(_10002_));
 sg13g2_xor2_1 _16841_ (.B(_10002_),
    .A(_09924_),
    .X(_10003_));
 sg13g2_o21ai_1 _16842_ (.B1(_10003_),
    .Y(_10004_),
    .A1(\cpu.intr.r_timer_reload[21] ),
    .A2(_09930_));
 sg13g2_buf_1 _16843_ (.A(\cpu.dcache.wdata[5] ),
    .X(_10005_));
 sg13g2_nand2_1 _16844_ (.Y(_10006_),
    .A(_10005_),
    .B(net184));
 sg13g2_o21ai_1 _16845_ (.B1(_10006_),
    .Y(_00068_),
    .A1(net185),
    .A2(_10004_));
 sg13g2_nor3_1 _16846_ (.A(_09924_),
    .B(_09925_),
    .C(_09923_),
    .Y(_10007_));
 sg13g2_xor2_1 _16847_ (.B(_10007_),
    .A(_09927_),
    .X(_10008_));
 sg13g2_o21ai_1 _16848_ (.B1(_10008_),
    .Y(_10009_),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .A2(_09930_));
 sg13g2_buf_1 _16849_ (.A(\cpu.dcache.wdata[6] ),
    .X(_10010_));
 sg13g2_nand2_1 _16850_ (.Y(_10011_),
    .A(_10010_),
    .B(_09900_));
 sg13g2_o21ai_1 _16851_ (.B1(_10011_),
    .Y(_00069_),
    .A1(net185),
    .A2(_10009_));
 sg13g2_nor2b_1 _16852_ (.A(_09926_),
    .B_N(\cpu.intr.r_timer_reload[23] ),
    .Y(_10012_));
 sg13g2_nor2b_1 _16853_ (.A(_09927_),
    .B_N(_10007_),
    .Y(_10013_));
 sg13g2_mux2_1 _16854_ (.A0(_09926_),
    .A1(_10012_),
    .S(_10013_),
    .X(_10014_));
 sg13g2_buf_2 _16855_ (.A(\cpu.dcache.wdata[7] ),
    .X(_10015_));
 sg13g2_buf_1 _16856_ (.A(_10015_),
    .X(_10016_));
 sg13g2_mux2_1 _16857_ (.A0(_10014_),
    .A1(net1056),
    .S(_09973_),
    .X(_00070_));
 sg13g2_buf_1 _16858_ (.A(net640),
    .X(_10017_));
 sg13g2_buf_1 _16859_ (.A(_10017_),
    .X(_10018_));
 sg13g2_buf_1 _16860_ (.A(net491),
    .X(_10019_));
 sg13g2_and2_1 _16861_ (.A(_09195_),
    .B(_09897_),
    .X(_10020_));
 sg13g2_buf_1 _16862_ (.A(_10020_),
    .X(_10021_));
 sg13g2_nand2_1 _16863_ (.Y(_10022_),
    .A(net441),
    .B(net234));
 sg13g2_buf_1 _16864_ (.A(_10022_),
    .X(_10023_));
 sg13g2_buf_1 _16865_ (.A(_10023_),
    .X(_10024_));
 sg13g2_buf_1 _16866_ (.A(_09179_),
    .X(_10025_));
 sg13g2_buf_1 _16867_ (.A(_10025_),
    .X(_10026_));
 sg13g2_buf_1 _16868_ (.A(_10026_),
    .X(_10027_));
 sg13g2_buf_1 _16869_ (.A(net636),
    .X(_10028_));
 sg13g2_nor3_1 _16870_ (.A(net566),
    .B(net922),
    .C(net153),
    .Y(_10029_));
 sg13g2_a21o_1 _16871_ (.A2(net153),
    .A1(_00279_),
    .B1(_10029_),
    .X(_00036_));
 sg13g2_nand2b_1 _16872_ (.Y(_10030_),
    .B(_09346_),
    .A_N(net715));
 sg13g2_buf_1 _16873_ (.A(_10030_),
    .X(_10031_));
 sg13g2_nor2_1 _16874_ (.A(_10031_),
    .B(_09898_),
    .Y(_10032_));
 sg13g2_buf_2 _16875_ (.A(_10032_),
    .X(_10033_));
 sg13g2_buf_1 _16876_ (.A(_10033_),
    .X(_10034_));
 sg13g2_buf_1 _16877_ (.A(net183),
    .X(_10035_));
 sg13g2_buf_2 _16878_ (.A(\cpu.intr.r_clock_count[0] ),
    .X(_10036_));
 sg13g2_buf_2 _16879_ (.A(\cpu.intr.r_clock_count[1] ),
    .X(_10037_));
 sg13g2_xnor2_1 _16880_ (.Y(_10038_),
    .A(_10036_),
    .B(_10037_));
 sg13g2_buf_1 _16881_ (.A(net798),
    .X(_10039_));
 sg13g2_buf_1 _16882_ (.A(net694),
    .X(_10040_));
 sg13g2_buf_1 _16883_ (.A(_10040_),
    .X(_10041_));
 sg13g2_buf_1 _16884_ (.A(_09978_),
    .X(_10042_));
 sg13g2_buf_1 _16885_ (.A(_10033_),
    .X(_10043_));
 sg13g2_nand3_1 _16886_ (.B(_10042_),
    .C(net182),
    .A(net565),
    .Y(_10044_));
 sg13g2_o21ai_1 _16887_ (.B1(_10044_),
    .Y(_00043_),
    .A1(net152),
    .A2(_10038_));
 sg13g2_buf_2 _16888_ (.A(\cpu.intr.r_clock_count[2] ),
    .X(_10045_));
 sg13g2_nand2_1 _16889_ (.Y(_10046_),
    .A(_10036_),
    .B(_10037_));
 sg13g2_xor2_1 _16890_ (.B(_10046_),
    .A(_10045_),
    .X(_10047_));
 sg13g2_nand3_1 _16891_ (.B(net1059),
    .C(net182),
    .A(net565),
    .Y(_10048_));
 sg13g2_o21ai_1 _16892_ (.B1(_10048_),
    .Y(_00044_),
    .A1(net152),
    .A2(_10047_));
 sg13g2_buf_1 _16893_ (.A(\cpu.intr.r_clock_count[3] ),
    .X(_10049_));
 sg13g2_nand3b_1 _16894_ (.B(_10045_),
    .C(_10037_),
    .Y(_10050_),
    .A_N(_00279_));
 sg13g2_xor2_1 _16895_ (.B(_10050_),
    .A(_10049_),
    .X(_10051_));
 sg13g2_nand3_1 _16896_ (.B(_09993_),
    .C(net182),
    .A(net565),
    .Y(_10052_));
 sg13g2_o21ai_1 _16897_ (.B1(_10052_),
    .Y(_00045_),
    .A1(net152),
    .A2(_10051_));
 sg13g2_buf_2 _16898_ (.A(\cpu.intr.r_clock_count[4] ),
    .X(_10053_));
 sg13g2_inv_1 _16899_ (.Y(_10054_),
    .A(_10036_));
 sg13g2_nand3_1 _16900_ (.B(_10045_),
    .C(_10049_),
    .A(_10037_),
    .Y(_10055_));
 sg13g2_nor2_1 _16901_ (.A(_10054_),
    .B(_10055_),
    .Y(_10056_));
 sg13g2_xnor2_1 _16902_ (.Y(_10057_),
    .A(_10053_),
    .B(_10056_));
 sg13g2_nand3_1 _16903_ (.B(net1057),
    .C(net182),
    .A(net565),
    .Y(_10058_));
 sg13g2_o21ai_1 _16904_ (.B1(_10058_),
    .Y(_00046_),
    .A1(net152),
    .A2(_10057_));
 sg13g2_buf_2 _16905_ (.A(\cpu.intr.r_clock_count[5] ),
    .X(_10059_));
 sg13g2_inv_1 _16906_ (.Y(_10060_),
    .A(_10053_));
 sg13g2_nor3_2 _16907_ (.A(_10060_),
    .B(_00279_),
    .C(_10055_),
    .Y(_10061_));
 sg13g2_xnor2_1 _16908_ (.Y(_10062_),
    .A(_10059_),
    .B(_10061_));
 sg13g2_buf_1 _16909_ (.A(_10005_),
    .X(_10063_));
 sg13g2_nand3_1 _16910_ (.B(net1054),
    .C(net182),
    .A(net565),
    .Y(_10064_));
 sg13g2_o21ai_1 _16911_ (.B1(_10064_),
    .Y(_00047_),
    .A1(net152),
    .A2(_10062_));
 sg13g2_buf_1 _16912_ (.A(\cpu.intr.r_clock_count[6] ),
    .X(_10065_));
 sg13g2_and2_1 _16913_ (.A(_10053_),
    .B(_10056_),
    .X(_10066_));
 sg13g2_nand2_1 _16914_ (.Y(_10067_),
    .A(_10059_),
    .B(_10066_));
 sg13g2_xor2_1 _16915_ (.B(_10067_),
    .A(_10065_),
    .X(_10068_));
 sg13g2_buf_1 _16916_ (.A(_10010_),
    .X(_10069_));
 sg13g2_buf_1 _16917_ (.A(net183),
    .X(_10070_));
 sg13g2_nand3_1 _16918_ (.B(net1053),
    .C(net151),
    .A(net565),
    .Y(_10071_));
 sg13g2_o21ai_1 _16919_ (.B1(_10071_),
    .Y(_00048_),
    .A1(net152),
    .A2(_10068_));
 sg13g2_buf_1 _16920_ (.A(\cpu.intr.r_clock_count[7] ),
    .X(_10072_));
 sg13g2_nand3_1 _16921_ (.B(_10065_),
    .C(_10061_),
    .A(_10059_),
    .Y(_10073_));
 sg13g2_xor2_1 _16922_ (.B(_10073_),
    .A(_10072_),
    .X(_10074_));
 sg13g2_nand3_1 _16923_ (.B(_10015_),
    .C(net151),
    .A(net565),
    .Y(_10075_));
 sg13g2_o21ai_1 _16924_ (.B1(_10075_),
    .Y(_00049_),
    .A1(net152),
    .A2(_10074_));
 sg13g2_buf_2 _16925_ (.A(\cpu.intr.r_clock_count[8] ),
    .X(_10076_));
 sg13g2_nand2_1 _16926_ (.Y(_10077_),
    .A(_10053_),
    .B(_10056_));
 sg13g2_nand3_1 _16927_ (.B(_10065_),
    .C(_10072_),
    .A(_10059_),
    .Y(_10078_));
 sg13g2_nor2_1 _16928_ (.A(_10077_),
    .B(_10078_),
    .Y(_10079_));
 sg13g2_xnor2_1 _16929_ (.Y(_10080_),
    .A(_10076_),
    .B(_10079_));
 sg13g2_buf_2 _16930_ (.A(\cpu.dcache.wdata[8] ),
    .X(_10081_));
 sg13g2_nand3_1 _16931_ (.B(_10081_),
    .C(net151),
    .A(net565),
    .Y(_10082_));
 sg13g2_o21ai_1 _16932_ (.B1(_10082_),
    .Y(_00050_),
    .A1(_10035_),
    .A2(_10080_));
 sg13g2_buf_2 _16933_ (.A(\cpu.intr.r_clock_count[9] ),
    .X(_10083_));
 sg13g2_nand2_1 _16934_ (.Y(_10084_),
    .A(_10076_),
    .B(_10079_));
 sg13g2_xor2_1 _16935_ (.B(_10084_),
    .A(_10083_),
    .X(_10085_));
 sg13g2_buf_2 _16936_ (.A(\cpu.dcache.wdata[9] ),
    .X(_10086_));
 sg13g2_nand3_1 _16937_ (.B(_10086_),
    .C(net151),
    .A(net635),
    .Y(_10087_));
 sg13g2_o21ai_1 _16938_ (.B1(_10087_),
    .Y(_00051_),
    .A1(net152),
    .A2(_10085_));
 sg13g2_buf_1 _16939_ (.A(\cpu.intr.r_clock_count[10] ),
    .X(_10088_));
 sg13g2_nand3_1 _16940_ (.B(_10083_),
    .C(_10079_),
    .A(_10076_),
    .Y(_10089_));
 sg13g2_xor2_1 _16941_ (.B(_10089_),
    .A(_10088_),
    .X(_10090_));
 sg13g2_buf_2 _16942_ (.A(\cpu.dcache.wdata[10] ),
    .X(_10091_));
 sg13g2_nand3_1 _16943_ (.B(_10091_),
    .C(net151),
    .A(net635),
    .Y(_10092_));
 sg13g2_o21ai_1 _16944_ (.B1(_10092_),
    .Y(_00037_),
    .A1(_10035_),
    .A2(_10090_));
 sg13g2_buf_2 _16945_ (.A(\cpu.intr.r_clock_count[11] ),
    .X(_10093_));
 sg13g2_nand3_1 _16946_ (.B(_10083_),
    .C(_10088_),
    .A(_10076_),
    .Y(_10094_));
 sg13g2_nor2_1 _16947_ (.A(_10078_),
    .B(_10094_),
    .Y(_10095_));
 sg13g2_and2_1 _16948_ (.A(_10061_),
    .B(_10095_),
    .X(_10096_));
 sg13g2_xnor2_1 _16949_ (.Y(_10097_),
    .A(_10093_),
    .B(_10096_));
 sg13g2_buf_2 _16950_ (.A(\cpu.dcache.wdata[11] ),
    .X(_10098_));
 sg13g2_nand3_1 _16951_ (.B(_10098_),
    .C(net151),
    .A(net635),
    .Y(_10099_));
 sg13g2_o21ai_1 _16952_ (.B1(_10099_),
    .Y(_00038_),
    .A1(net182),
    .A2(_10097_));
 sg13g2_buf_2 _16953_ (.A(\cpu.intr.r_clock_count[12] ),
    .X(_10100_));
 sg13g2_nand3_1 _16954_ (.B(_10066_),
    .C(_10095_),
    .A(_10093_),
    .Y(_10101_));
 sg13g2_xor2_1 _16955_ (.B(_10101_),
    .A(_10100_),
    .X(_10102_));
 sg13g2_buf_1 _16956_ (.A(\cpu.dcache.wdata[12] ),
    .X(_10103_));
 sg13g2_nand3_1 _16957_ (.B(_10103_),
    .C(net151),
    .A(net635),
    .Y(_10104_));
 sg13g2_o21ai_1 _16958_ (.B1(_10104_),
    .Y(_00039_),
    .A1(net182),
    .A2(_10102_));
 sg13g2_buf_1 _16959_ (.A(\cpu.intr.r_clock_count[13] ),
    .X(_10105_));
 sg13g2_nand4_1 _16960_ (.B(_10100_),
    .C(_10061_),
    .A(_10093_),
    .Y(_10106_),
    .D(_10095_));
 sg13g2_xor2_1 _16961_ (.B(_10106_),
    .A(_10105_),
    .X(_10107_));
 sg13g2_buf_1 _16962_ (.A(\cpu.dcache.wdata[13] ),
    .X(_10108_));
 sg13g2_nand3_1 _16963_ (.B(_10108_),
    .C(_10070_),
    .A(net635),
    .Y(_10109_));
 sg13g2_o21ai_1 _16964_ (.B1(_10109_),
    .Y(_00040_),
    .A1(_10043_),
    .A2(_10107_));
 sg13g2_buf_1 _16965_ (.A(\cpu.intr.r_clock_count[14] ),
    .X(_10110_));
 sg13g2_nand4_1 _16966_ (.B(_10100_),
    .C(_10105_),
    .A(_10093_),
    .Y(_10111_),
    .D(_10095_));
 sg13g2_nor2_1 _16967_ (.A(_10077_),
    .B(_10111_),
    .Y(_10112_));
 sg13g2_xnor2_1 _16968_ (.Y(_10113_),
    .A(_10110_),
    .B(_10112_));
 sg13g2_buf_2 _16969_ (.A(\cpu.dcache.wdata[14] ),
    .X(_10114_));
 sg13g2_nand3_1 _16970_ (.B(_10114_),
    .C(net151),
    .A(net635),
    .Y(_10115_));
 sg13g2_o21ai_1 _16971_ (.B1(_10115_),
    .Y(_00041_),
    .A1(_10043_),
    .A2(_10113_));
 sg13g2_buf_1 _16972_ (.A(\cpu.intr.r_clock_count[15] ),
    .X(_10116_));
 sg13g2_inv_1 _16973_ (.Y(_10117_),
    .A(_10116_));
 sg13g2_inv_1 _16974_ (.Y(_10118_),
    .A(_10110_));
 sg13g2_nor2_1 _16975_ (.A(_10118_),
    .B(_10111_),
    .Y(_10119_));
 sg13g2_nand2_1 _16976_ (.Y(_10120_),
    .A(_10061_),
    .B(_10119_));
 sg13g2_xnor2_1 _16977_ (.Y(_10121_),
    .A(_10117_),
    .B(_10120_));
 sg13g2_buf_2 _16978_ (.A(\cpu.dcache.wdata[15] ),
    .X(_10122_));
 sg13g2_nand3_1 _16979_ (.B(_10122_),
    .C(_10070_),
    .A(net635),
    .Y(_10123_));
 sg13g2_o21ai_1 _16980_ (.B1(_10123_),
    .Y(_00042_),
    .A1(net182),
    .A2(_10121_));
 sg13g2_inv_1 _16981_ (.Y(_10124_),
    .A(_09272_));
 sg13g2_nand2_1 _16982_ (.Y(_10125_),
    .A(_09277_),
    .B(net814));
 sg13g2_buf_2 _16983_ (.A(_10125_),
    .X(_10126_));
 sg13g2_buf_1 _16984_ (.A(_10126_),
    .X(_10127_));
 sg13g2_a21oi_1 _16985_ (.A1(_10124_),
    .A2(net564),
    .Y(_10128_),
    .B1(net492));
 sg13g2_buf_1 _16986_ (.A(_10128_),
    .X(_10129_));
 sg13g2_buf_1 _16987_ (.A(net386),
    .X(_10130_));
 sg13g2_buf_1 _16988_ (.A(\cpu.ex.r_mult[25] ),
    .X(_10131_));
 sg13g2_buf_1 _16989_ (.A(_10131_),
    .X(_10132_));
 sg13g2_buf_1 _16990_ (.A(\cpu.dec.r_rs2_pc ),
    .X(_10133_));
 sg13g2_inv_2 _16991_ (.Y(_10134_),
    .A(_10133_));
 sg13g2_buf_1 _16992_ (.A(_10134_),
    .X(_10135_));
 sg13g2_buf_1 _16993_ (.A(_00286_),
    .X(_10136_));
 sg13g2_nor2_1 _16994_ (.A(net920),
    .B(_10136_),
    .Y(_10137_));
 sg13g2_buf_1 _16995_ (.A(_10133_),
    .X(_10138_));
 sg13g2_buf_1 _16996_ (.A(_10138_),
    .X(_10139_));
 sg13g2_buf_1 _16997_ (.A(\cpu.dec.needs_rs2 ),
    .X(_10140_));
 sg13g2_buf_1 _16998_ (.A(_10140_),
    .X(_10141_));
 sg13g2_nor2_1 _16999_ (.A(net1050),
    .B(\cpu.dec.imm[10] ),
    .Y(_10142_));
 sg13g2_buf_1 _17000_ (.A(\cpu.addr[10] ),
    .X(_10143_));
 sg13g2_buf_8 _17001_ (.A(\cpu.ex.r_wb_addr[1] ),
    .X(_10144_));
 sg13g2_buf_8 _17002_ (.A(\cpu.ex.r_wb_addr[0] ),
    .X(_10145_));
 sg13g2_nor2_1 _17003_ (.A(net1142),
    .B(_10145_),
    .Y(_10146_));
 sg13g2_buf_1 _17004_ (.A(\cpu.ex.r_wb_addr[3] ),
    .X(_10147_));
 sg13g2_buf_8 _17005_ (.A(\cpu.ex.r_wb_addr[2] ),
    .X(_10148_));
 sg13g2_nor2_1 _17006_ (.A(net1141),
    .B(_10148_),
    .Y(_10149_));
 sg13g2_buf_8 _17007_ (.A(\cpu.ex.r_wb_valid ),
    .X(_10150_));
 sg13g2_inv_1 _17008_ (.Y(_10151_),
    .A(_10150_));
 sg13g2_a21o_1 _17009_ (.A2(_10149_),
    .A1(_10146_),
    .B1(_10151_),
    .X(_10152_));
 sg13g2_buf_1 _17010_ (.A(_10152_),
    .X(_10153_));
 sg13g2_buf_8 _17011_ (.A(\cpu.dec.r_rs2[2] ),
    .X(_10154_));
 sg13g2_xor2_1 _17012_ (.B(net1140),
    .A(_10148_),
    .X(_10155_));
 sg13g2_buf_8 _17013_ (.A(\cpu.dec.r_rs2[1] ),
    .X(_10156_));
 sg13g2_xor2_1 _17014_ (.B(net1139),
    .A(net1142),
    .X(_10157_));
 sg13g2_buf_8 _17015_ (.A(\cpu.dec.r_rs2[3] ),
    .X(_10158_));
 sg13g2_xnor2_1 _17016_ (.Y(_10159_),
    .A(net1141),
    .B(net1138));
 sg13g2_buf_8 _17017_ (.A(\cpu.dec.r_rs2[0] ),
    .X(_10160_));
 sg13g2_xnor2_1 _17018_ (.Y(_10161_),
    .A(_10145_),
    .B(_10160_));
 sg13g2_nand2_1 _17019_ (.Y(_10162_),
    .A(_10159_),
    .B(_10161_));
 sg13g2_nor4_2 _17020_ (.A(_10153_),
    .B(_10155_),
    .C(_10157_),
    .Y(_10163_),
    .D(_10162_));
 sg13g2_buf_8 _17021_ (.A(_10163_),
    .X(_10164_));
 sg13g2_buf_1 _17022_ (.A(_10164_),
    .X(_10165_));
 sg13g2_nor2_1 _17023_ (.A(_10160_),
    .B(net1139),
    .Y(_10166_));
 sg13g2_buf_1 _17024_ (.A(_10166_),
    .X(_10167_));
 sg13g2_nor2_2 _17025_ (.A(_10158_),
    .B(_10154_),
    .Y(_10168_));
 sg13g2_buf_1 _17026_ (.A(_10168_),
    .X(_10169_));
 sg13g2_a21oi_1 _17027_ (.A1(net918),
    .A2(net917),
    .Y(_10170_),
    .B1(_10164_));
 sg13g2_buf_1 _17028_ (.A(_10170_),
    .X(_10171_));
 sg13g2_and2_1 _17029_ (.A(_10160_),
    .B(_10156_),
    .X(_10172_));
 sg13g2_buf_2 _17030_ (.A(_10172_),
    .X(_10173_));
 sg13g2_a22oi_1 _17031_ (.Y(_10174_),
    .B1(_10173_),
    .B2(\cpu.ex.r_11[10] ),
    .A2(net918),
    .A1(\cpu.ex.r_8[10] ));
 sg13g2_nor2b_1 _17032_ (.A(net1140),
    .B_N(net1138),
    .Y(_10175_));
 sg13g2_buf_1 _17033_ (.A(_10175_),
    .X(_10176_));
 sg13g2_nand2b_1 _17034_ (.Y(_10177_),
    .B(net916),
    .A_N(_10174_));
 sg13g2_nor2b_1 _17035_ (.A(net1138),
    .B_N(net1139),
    .Y(_10178_));
 sg13g2_buf_2 _17036_ (.A(_10178_),
    .X(_10179_));
 sg13g2_buf_1 _17037_ (.A(_10179_),
    .X(_10180_));
 sg13g2_inv_1 _17038_ (.Y(_10181_),
    .A(\cpu.ex.r_epc[10] ));
 sg13g2_buf_8 _17039_ (.A(net1140),
    .X(_10182_));
 sg13g2_buf_8 _17040_ (.A(_10160_),
    .X(_10183_));
 sg13g2_buf_8 _17041_ (.A(net1048),
    .X(_10184_));
 sg13g2_nand2b_1 _17042_ (.Y(_10185_),
    .B(net915),
    .A_N(net1049));
 sg13g2_buf_8 _17043_ (.A(_10185_),
    .X(_10186_));
 sg13g2_buf_8 _17044_ (.A(net915),
    .X(_10187_));
 sg13g2_buf_1 _17045_ (.A(net794),
    .X(_10188_));
 sg13g2_buf_8 _17046_ (.A(net1049),
    .X(_10189_));
 sg13g2_buf_1 _17047_ (.A(net914),
    .X(_10190_));
 sg13g2_buf_1 _17048_ (.A(_10190_),
    .X(_10191_));
 sg13g2_nand3b_1 _17049_ (.B(net692),
    .C(\cpu.ex.r_stmp[10] ),
    .Y(_10192_),
    .A_N(net693));
 sg13g2_o21ai_1 _17050_ (.B1(_10192_),
    .Y(_10193_),
    .A1(_10181_),
    .A2(_10186_));
 sg13g2_buf_8 _17051_ (.A(_10156_),
    .X(_10194_));
 sg13g2_buf_8 _17052_ (.A(_10194_),
    .X(_10195_));
 sg13g2_buf_8 _17053_ (.A(net913),
    .X(_10196_));
 sg13g2_buf_8 _17054_ (.A(_10196_),
    .X(_10197_));
 sg13g2_buf_8 _17055_ (.A(net1138),
    .X(_10198_));
 sg13g2_buf_8 _17056_ (.A(net1046),
    .X(_10199_));
 sg13g2_buf_1 _17057_ (.A(net912),
    .X(_10200_));
 sg13g2_buf_8 _17058_ (.A(net692),
    .X(_10201_));
 sg13g2_and3_1 _17059_ (.X(_10202_),
    .A(net691),
    .B(net791),
    .C(net634));
 sg13g2_inv_1 _17060_ (.Y(_10203_),
    .A(_00260_));
 sg13g2_inv_1 _17061_ (.Y(_10204_),
    .A(net794));
 sg13g2_buf_1 _17062_ (.A(_10204_),
    .X(_10205_));
 sg13g2_mux2_1 _17063_ (.A0(_10203_),
    .A1(\cpu.ex.r_14[10] ),
    .S(_10205_),
    .X(_10206_));
 sg13g2_inv_1 _17064_ (.Y(_10207_),
    .A(net1049));
 sg13g2_buf_1 _17065_ (.A(_10207_),
    .X(_10208_));
 sg13g2_nor2b_1 _17066_ (.A(net1048),
    .B_N(net1139),
    .Y(_10209_));
 sg13g2_buf_1 _17067_ (.A(_10209_),
    .X(_10210_));
 sg13g2_buf_1 _17068_ (.A(\cpu.ex.r_sp[10] ),
    .X(_10211_));
 sg13g2_mux2_1 _17069_ (.A0(_10211_),
    .A1(\cpu.ex.r_10[10] ),
    .S(net791),
    .X(_10212_));
 sg13g2_and3_1 _17070_ (.X(_10213_),
    .A(net790),
    .B(net789),
    .C(_10212_));
 sg13g2_a221oi_1 _17071_ (.B2(_10206_),
    .C1(_10213_),
    .B1(_10202_),
    .A1(net795),
    .Y(_10214_),
    .A2(_10193_));
 sg13g2_buf_1 _17072_ (.A(\cpu.ex.r_mult[26] ),
    .X(_10215_));
 sg13g2_buf_1 _17073_ (.A(net693),
    .X(_10216_));
 sg13g2_nand3_1 _17074_ (.B(net632),
    .C(net795),
    .A(_10215_),
    .Y(_10217_));
 sg13g2_buf_1 _17075_ (.A(net791),
    .X(_10218_));
 sg13g2_nand3_1 _17076_ (.B(_10218_),
    .C(net918),
    .A(\cpu.ex.r_12[10] ),
    .Y(_10219_));
 sg13g2_a21o_1 _17077_ (.A2(_10219_),
    .A1(_10217_),
    .B1(net790),
    .X(_10220_));
 sg13g2_mux2_1 _17078_ (.A0(\cpu.ex.r_9[10] ),
    .A1(\cpu.ex.r_13[10] ),
    .S(net692),
    .X(_10221_));
 sg13g2_a22oi_1 _17079_ (.Y(_10222_),
    .B1(_10221_),
    .B2(_10218_),
    .A2(net917),
    .A1(\cpu.ex.r_lr[10] ));
 sg13g2_nor2b_1 _17080_ (.A(net1139),
    .B_N(_10160_),
    .Y(_10223_));
 sg13g2_buf_2 _17081_ (.A(_10223_),
    .X(_10224_));
 sg13g2_nand2b_1 _17082_ (.Y(_10225_),
    .B(_10224_),
    .A_N(_10222_));
 sg13g2_nand4_1 _17083_ (.B(_10214_),
    .C(_10220_),
    .A(_10177_),
    .Y(_10226_),
    .D(_10225_));
 sg13g2_inv_1 _17084_ (.Y(_10227_),
    .A(_10140_));
 sg13g2_buf_1 _17085_ (.A(_10227_),
    .X(_10228_));
 sg13g2_a221oi_1 _17086_ (.B2(_10226_),
    .C1(net911),
    .B1(_10171_),
    .A1(net1143),
    .Y(_10229_),
    .A2(net563));
 sg13g2_nor3_1 _17087_ (.A(net919),
    .B(_10142_),
    .C(_10229_),
    .Y(_10230_));
 sg13g2_or2_1 _17088_ (.X(_10231_),
    .B(_10230_),
    .A(_10137_));
 sg13g2_buf_2 _17089_ (.A(_10231_),
    .X(_10232_));
 sg13g2_buf_1 _17090_ (.A(\cpu.ex.r_mult[24] ),
    .X(_10233_));
 sg13g2_buf_2 _17091_ (.A(\cpu.addr[9] ),
    .X(_10234_));
 sg13g2_buf_1 _17092_ (.A(_10165_),
    .X(_10235_));
 sg13g2_nand2_1 _17093_ (.Y(_10236_),
    .A(_10234_),
    .B(_10235_));
 sg13g2_nor3_1 _17094_ (.A(net1139),
    .B(net1138),
    .C(net1140),
    .Y(_10237_));
 sg13g2_nand2_1 _17095_ (.Y(_10238_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_10237_));
 sg13g2_nor2b_1 _17096_ (.A(_00259_),
    .B_N(net791),
    .Y(_10239_));
 sg13g2_nor2b_1 _17097_ (.A(net690),
    .B_N(_10131_),
    .Y(_10240_));
 sg13g2_and2_1 _17098_ (.A(_10194_),
    .B(_10182_),
    .X(_10241_));
 sg13g2_buf_2 _17099_ (.A(_10241_),
    .X(_10242_));
 sg13g2_o21ai_1 _17100_ (.B1(_10242_),
    .Y(_10243_),
    .A1(_10239_),
    .A2(_10240_));
 sg13g2_inv_1 _17101_ (.Y(_10244_),
    .A(net1047));
 sg13g2_buf_1 _17102_ (.A(_10244_),
    .X(_10245_));
 sg13g2_and2_1 _17103_ (.A(net1138),
    .B(\cpu.dec.r_rs2[2] ),
    .X(_10246_));
 sg13g2_buf_1 _17104_ (.A(_10246_),
    .X(_10247_));
 sg13g2_buf_1 _17105_ (.A(_10247_),
    .X(_10248_));
 sg13g2_nand3_1 _17106_ (.B(_10245_),
    .C(net787),
    .A(\cpu.ex.r_13[9] ),
    .Y(_10249_));
 sg13g2_buf_1 _17107_ (.A(net691),
    .X(_10250_));
 sg13g2_nand3_1 _17108_ (.B(net631),
    .C(_10169_),
    .A(\cpu.ex.r_epc[9] ),
    .Y(_10251_));
 sg13g2_nand4_1 _17109_ (.B(_10243_),
    .C(_10249_),
    .A(_10238_),
    .Y(_10252_),
    .D(_10251_));
 sg13g2_mux2_1 _17110_ (.A0(\cpu.ex.r_stmp[9] ),
    .A1(\cpu.ex.r_14[9] ),
    .S(net791),
    .X(_10253_));
 sg13g2_a22oi_1 _17111_ (.Y(_10254_),
    .B1(_10253_),
    .B2(_10201_),
    .A2(net916),
    .A1(\cpu.ex.r_10[9] ));
 sg13g2_nand3_1 _17112_ (.B(net788),
    .C(net916),
    .A(\cpu.ex.r_8[9] ),
    .Y(_10255_));
 sg13g2_o21ai_1 _17113_ (.B1(_10255_),
    .Y(_10256_),
    .A1(net788),
    .A2(_10254_));
 sg13g2_buf_1 _17114_ (.A(net633),
    .X(_10257_));
 sg13g2_mux2_1 _17115_ (.A0(_10252_),
    .A1(_10256_),
    .S(net562),
    .X(_10258_));
 sg13g2_nor2b_1 _17116_ (.A(net913),
    .B_N(_10182_),
    .Y(_10259_));
 sg13g2_buf_2 _17117_ (.A(_10259_),
    .X(_10260_));
 sg13g2_nand3_1 _17118_ (.B(_10257_),
    .C(_10260_),
    .A(\cpu.ex.r_12[9] ),
    .Y(_10261_));
 sg13g2_nand3_1 _17119_ (.B(net790),
    .C(_10173_),
    .A(\cpu.ex.r_11[9] ),
    .Y(_10262_));
 sg13g2_inv_2 _17120_ (.Y(_10263_),
    .A(net1046));
 sg13g2_a21oi_1 _17121_ (.A1(_10261_),
    .A2(_10262_),
    .Y(_10264_),
    .B1(_10263_));
 sg13g2_buf_1 _17122_ (.A(\cpu.ex.r_sp[9] ),
    .X(_10265_));
 sg13g2_nand3_1 _17123_ (.B(net562),
    .C(net795),
    .A(_10265_),
    .Y(_10266_));
 sg13g2_nor2b_1 _17124_ (.A(net913),
    .B_N(net1046),
    .Y(_10267_));
 sg13g2_buf_1 _17125_ (.A(_10267_),
    .X(_10268_));
 sg13g2_nand3_1 _17126_ (.B(_10216_),
    .C(_10268_),
    .A(\cpu.ex.r_9[9] ),
    .Y(_10269_));
 sg13g2_buf_1 _17127_ (.A(net634),
    .X(_10270_));
 sg13g2_a21oi_1 _17128_ (.A1(_10266_),
    .A2(_10269_),
    .Y(_10271_),
    .B1(net561));
 sg13g2_or2_1 _17129_ (.X(_10272_),
    .B(_10271_),
    .A(_10264_));
 sg13g2_buf_1 _17130_ (.A(_10171_),
    .X(_10273_));
 sg13g2_o21ai_1 _17131_ (.B1(net440),
    .Y(_10274_),
    .A1(_10258_),
    .A2(_10272_));
 sg13g2_nand2_2 _17132_ (.Y(_10275_),
    .A(_10134_),
    .B(_10140_));
 sg13g2_a21oi_1 _17133_ (.A1(_10236_),
    .A2(_10274_),
    .Y(_10276_),
    .B1(_10275_));
 sg13g2_inv_1 _17134_ (.Y(_10277_),
    .A(_00287_));
 sg13g2_nor2_1 _17135_ (.A(net1051),
    .B(_10140_),
    .Y(_10278_));
 sg13g2_buf_2 _17136_ (.A(_10278_),
    .X(_10279_));
 sg13g2_a22oi_1 _17137_ (.Y(_10280_),
    .B1(\cpu.dec.imm[9] ),
    .B2(_10279_),
    .A2(_10277_),
    .A1(net919));
 sg13g2_nor2b_1 _17138_ (.A(_10276_),
    .B_N(_10280_),
    .Y(_10281_));
 sg13g2_buf_2 _17139_ (.A(_10281_),
    .X(_10282_));
 sg13g2_nor2_1 _17140_ (.A(net1137),
    .B(_10282_),
    .Y(_10283_));
 sg13g2_and2_1 _17141_ (.A(net1048),
    .B(net1140),
    .X(_10284_));
 sg13g2_buf_2 _17142_ (.A(_10284_),
    .X(_10285_));
 sg13g2_inv_1 _17143_ (.Y(_10286_),
    .A(_00258_));
 sg13g2_mux2_1 _17144_ (.A0(_10286_),
    .A1(\cpu.ex.r_13[8] ),
    .S(net788),
    .X(_10287_));
 sg13g2_nor2b_1 _17145_ (.A(net632),
    .B_N(\cpu.ex.r_8[8] ),
    .Y(_10288_));
 sg13g2_nor2_2 _17146_ (.A(net913),
    .B(_10189_),
    .Y(_10289_));
 sg13g2_a22oi_1 _17147_ (.Y(_10290_),
    .B1(_10288_),
    .B2(_10289_),
    .A2(_10287_),
    .A1(_10285_));
 sg13g2_buf_1 _17148_ (.A(net690),
    .X(_10291_));
 sg13g2_nand2b_1 _17149_ (.Y(_10292_),
    .B(_10291_),
    .A_N(_10290_));
 sg13g2_mux2_1 _17150_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net1137),
    .S(net692),
    .X(_10293_));
 sg13g2_nand3_1 _17151_ (.B(_10180_),
    .C(_10293_),
    .A(net632),
    .Y(_10294_));
 sg13g2_nand4_1 _17152_ (.B(net562),
    .C(net788),
    .A(\cpu.ex.r_12[8] ),
    .Y(_10295_),
    .D(net787));
 sg13g2_and2_1 _17153_ (.A(_10294_),
    .B(_10295_),
    .X(_10296_));
 sg13g2_a22oi_1 _17154_ (.Y(_10297_),
    .B1(_10224_),
    .B2(\cpu.ex.r_9[8] ),
    .A2(_10173_),
    .A1(\cpu.ex.r_11[8] ));
 sg13g2_inv_1 _17155_ (.Y(_10298_),
    .A(_10297_));
 sg13g2_and2_1 _17156_ (.A(net917),
    .B(_10224_),
    .X(_10299_));
 sg13g2_a22oi_1 _17157_ (.Y(_10300_),
    .B1(_10299_),
    .B2(\cpu.ex.r_lr[8] ),
    .A2(_10298_),
    .A1(net916));
 sg13g2_buf_1 _17158_ (.A(\cpu.ex.r_sp[8] ),
    .X(_10301_));
 sg13g2_mux4_1 _17159_ (.S0(net634),
    .A0(_10301_),
    .A1(\cpu.ex.r_stmp[8] ),
    .A2(\cpu.ex.r_10[8] ),
    .A3(\cpu.ex.r_14[8] ),
    .S1(net690),
    .X(_10302_));
 sg13g2_nand2_1 _17160_ (.Y(_10303_),
    .A(net789),
    .B(_10302_));
 sg13g2_nand4_1 _17161_ (.B(_10296_),
    .C(_10300_),
    .A(_10292_),
    .Y(_10304_),
    .D(_10303_));
 sg13g2_and2_1 _17162_ (.A(_09165_),
    .B(net563),
    .X(_10305_));
 sg13g2_a21o_1 _17163_ (.A2(_10304_),
    .A1(_10273_),
    .B1(_10305_),
    .X(_10306_));
 sg13g2_nor2_1 _17164_ (.A(_10133_),
    .B(_10227_),
    .Y(_10307_));
 sg13g2_buf_2 _17165_ (.A(_10307_),
    .X(_10308_));
 sg13g2_nor2_1 _17166_ (.A(net920),
    .B(_00282_),
    .Y(_10309_));
 sg13g2_a221oi_1 _17167_ (.B2(_10308_),
    .C1(_10309_),
    .B1(_10306_),
    .A1(\cpu.dec.imm[8] ),
    .Y(_10310_),
    .A2(_10279_));
 sg13g2_buf_1 _17168_ (.A(_10310_),
    .X(_10311_));
 sg13g2_buf_1 _17169_ (.A(\cpu.ex.r_mult[23] ),
    .X(_10312_));
 sg13g2_a22oi_1 _17170_ (.Y(_10313_),
    .B1(_10311_),
    .B2(net1136),
    .A2(_10282_),
    .A1(net1137));
 sg13g2_nor3_1 _17171_ (.A(_10232_),
    .B(_10283_),
    .C(_10313_),
    .Y(_10314_));
 sg13g2_nor2_1 _17172_ (.A(_10132_),
    .B(_10314_),
    .Y(_10315_));
 sg13g2_buf_1 _17173_ (.A(_10215_),
    .X(_10316_));
 sg13g2_o21ai_1 _17174_ (.B1(_10232_),
    .Y(_10317_),
    .A1(_10283_),
    .A2(_10313_));
 sg13g2_nand2_1 _17175_ (.Y(_10318_),
    .A(net1045),
    .B(_10317_));
 sg13g2_buf_1 _17176_ (.A(_00285_),
    .X(_10319_));
 sg13g2_nor2_1 _17177_ (.A(net920),
    .B(_10319_),
    .Y(_10320_));
 sg13g2_nor2_1 _17178_ (.A(_10141_),
    .B(\cpu.dec.imm[11] ),
    .Y(_10321_));
 sg13g2_buf_1 _17179_ (.A(\cpu.addr[11] ),
    .X(_10322_));
 sg13g2_nor2b_1 _17180_ (.A(net915),
    .B_N(net1046),
    .Y(_10323_));
 sg13g2_buf_2 _17181_ (.A(_10323_),
    .X(_10324_));
 sg13g2_inv_1 _17182_ (.Y(_10325_),
    .A(_10324_));
 sg13g2_a22oi_1 _17183_ (.Y(_10326_),
    .B1(_10242_),
    .B2(\cpu.ex.r_14[11] ),
    .A2(_10289_),
    .A1(\cpu.ex.r_8[11] ));
 sg13g2_nor2b_1 _17184_ (.A(_00261_),
    .B_N(net691),
    .Y(_10327_));
 sg13g2_nor2b_1 _17185_ (.A(net691),
    .B_N(\cpu.ex.r_13[11] ),
    .Y(_10328_));
 sg13g2_and3_1 _17186_ (.X(_10329_),
    .A(_10188_),
    .B(net791),
    .C(net692));
 sg13g2_o21ai_1 _17187_ (.B1(_10329_),
    .Y(_10330_),
    .A1(_10327_),
    .A2(_10328_));
 sg13g2_o21ai_1 _17188_ (.B1(_10330_),
    .Y(_10331_),
    .A1(_10325_),
    .A2(_10326_));
 sg13g2_nand3_1 _17189_ (.B(net632),
    .C(_10169_),
    .A(\cpu.ex.r_lr[11] ),
    .Y(_10332_));
 sg13g2_nand3_1 _17190_ (.B(net633),
    .C(_10248_),
    .A(\cpu.ex.r_12[11] ),
    .Y(_10333_));
 sg13g2_a21oi_1 _17191_ (.A1(_10332_),
    .A2(_10333_),
    .Y(_10334_),
    .B1(net631));
 sg13g2_nand2b_1 _17192_ (.Y(_10335_),
    .B(net1138),
    .A_N(_10154_));
 sg13g2_buf_2 _17193_ (.A(_10335_),
    .X(_10336_));
 sg13g2_a22oi_1 _17194_ (.Y(_10337_),
    .B1(net789),
    .B2(\cpu.ex.r_10[11] ),
    .A2(_10224_),
    .A1(\cpu.ex.r_9[11] ));
 sg13g2_buf_1 _17195_ (.A(\cpu.ex.r_mult[27] ),
    .X(_10338_));
 sg13g2_nand3b_1 _17196_ (.B(_10191_),
    .C(net1134),
    .Y(_10339_),
    .A_N(net791));
 sg13g2_nand3b_1 _17197_ (.B(net791),
    .C(\cpu.ex.r_11[11] ),
    .Y(_10340_),
    .A_N(net692));
 sg13g2_nand2_1 _17198_ (.Y(_10341_),
    .A(net794),
    .B(net792));
 sg13g2_a21o_1 _17199_ (.A2(_10340_),
    .A1(_10339_),
    .B1(_10341_),
    .X(_10342_));
 sg13g2_o21ai_1 _17200_ (.B1(_10342_),
    .Y(_10343_),
    .A1(_10336_),
    .A2(_10337_));
 sg13g2_nand2b_1 _17201_ (.Y(_10344_),
    .B(net913),
    .A_N(net912));
 sg13g2_buf_2 _17202_ (.A(_10344_),
    .X(_10345_));
 sg13g2_nor2b_1 _17203_ (.A(net793),
    .B_N(_10187_),
    .Y(_10346_));
 sg13g2_buf_1 _17204_ (.A(\cpu.ex.r_sp[11] ),
    .X(_10347_));
 sg13g2_mux2_1 _17205_ (.A0(_10347_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net692),
    .X(_10348_));
 sg13g2_a22oi_1 _17206_ (.Y(_10349_),
    .B1(_10348_),
    .B2(net562),
    .A2(_10346_),
    .A1(\cpu.ex.r_epc[11] ));
 sg13g2_nor2_1 _17207_ (.A(_10345_),
    .B(_10349_),
    .Y(_10350_));
 sg13g2_or4_1 _17208_ (.A(_10331_),
    .B(_10334_),
    .C(_10343_),
    .D(_10350_),
    .X(_10351_));
 sg13g2_a221oi_1 _17209_ (.B2(_10351_),
    .C1(net911),
    .B1(_10171_),
    .A1(net1135),
    .Y(_10352_),
    .A2(net563));
 sg13g2_nor3_2 _17210_ (.A(net1051),
    .B(_10321_),
    .C(_10352_),
    .Y(_10353_));
 sg13g2_or2_1 _17211_ (.X(_10354_),
    .B(_10353_),
    .A(_10320_));
 sg13g2_buf_2 _17212_ (.A(_10354_),
    .X(_10355_));
 sg13g2_o21ai_1 _17213_ (.B1(_10355_),
    .Y(_10356_),
    .A1(_10315_),
    .A2(_10318_));
 sg13g2_a21oi_1 _17214_ (.A1(_10132_),
    .A2(_10317_),
    .Y(_10357_),
    .B1(net1045));
 sg13g2_nor2_1 _17215_ (.A(net568),
    .B(_10357_),
    .Y(_10358_));
 sg13g2_nand2b_1 _17216_ (.Y(_10359_),
    .B(_10280_),
    .A_N(_10276_));
 sg13g2_buf_2 _17217_ (.A(_10359_),
    .X(_10360_));
 sg13g2_a22oi_1 _17218_ (.Y(_10361_),
    .B1(net440),
    .B2(_10304_),
    .A2(net490),
    .A1(_09165_));
 sg13g2_a21oi_1 _17219_ (.A1(\cpu.dec.imm[8] ),
    .A2(_10279_),
    .Y(_10362_),
    .B1(_10309_));
 sg13g2_o21ai_1 _17220_ (.B1(_10362_),
    .Y(_10363_),
    .A1(_10275_),
    .A2(_10361_));
 sg13g2_buf_1 _17221_ (.A(_10363_),
    .X(_10364_));
 sg13g2_buf_1 _17222_ (.A(_10364_),
    .X(_10365_));
 sg13g2_nor2_2 _17223_ (.A(_10360_),
    .B(net233),
    .Y(_10366_));
 sg13g2_nor2_1 _17224_ (.A(_10355_),
    .B(_10232_),
    .Y(_10367_));
 sg13g2_nor2_1 _17225_ (.A(net1136),
    .B(_10311_),
    .Y(_10368_));
 sg13g2_inv_2 _17226_ (.Y(_10369_),
    .A(_10355_));
 sg13g2_o21ai_1 _17227_ (.B1(net564),
    .Y(_10370_),
    .A1(_10316_),
    .A2(_10369_));
 sg13g2_nor2_1 _17228_ (.A(_10137_),
    .B(_10230_),
    .Y(_10371_));
 sg13g2_a21oi_1 _17229_ (.A1(net1045),
    .A2(_10371_),
    .Y(_10372_),
    .B1(_10131_));
 sg13g2_nor4_1 _17230_ (.A(_10283_),
    .B(_10368_),
    .C(_10370_),
    .D(_10372_),
    .Y(_10373_));
 sg13g2_a21o_1 _17231_ (.A2(_10367_),
    .A1(_10366_),
    .B1(_10373_),
    .X(_10374_));
 sg13g2_buf_1 _17232_ (.A(\cpu.ex.r_mult[21] ),
    .X(_10375_));
 sg13g2_buf_1 _17233_ (.A(\cpu.ex.r_mult[22] ),
    .X(_10376_));
 sg13g2_inv_2 _17234_ (.Y(_10377_),
    .A(net1132));
 sg13g2_nand2_1 _17235_ (.Y(_10378_),
    .A(_09166_),
    .B(net563));
 sg13g2_mux4_1 _17236_ (.S0(net691),
    .A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_10[7] ),
    .A2(\cpu.ex.r_12[7] ),
    .A3(\cpu.ex.r_14[7] ),
    .S1(net634),
    .X(_10379_));
 sg13g2_nor2_1 _17237_ (.A(net1047),
    .B(_10336_),
    .Y(_10380_));
 sg13g2_and3_1 _17238_ (.X(_10381_),
    .A(_10312_),
    .B(_10191_),
    .C(_10180_));
 sg13g2_a21o_1 _17239_ (.A2(_10380_),
    .A1(\cpu.ex.r_9[7] ),
    .B1(_10381_),
    .X(_10382_));
 sg13g2_buf_1 _17240_ (.A(net632),
    .X(_10383_));
 sg13g2_a22oi_1 _17241_ (.Y(_10384_),
    .B1(_10382_),
    .B2(net560),
    .A2(_10379_),
    .A1(_10324_));
 sg13g2_nor2b_1 _17242_ (.A(net1048),
    .B_N(net1140),
    .Y(_10385_));
 sg13g2_a22oi_1 _17243_ (.Y(_10386_),
    .B1(_10385_),
    .B2(\cpu.ex.r_stmp[7] ),
    .A2(_10346_),
    .A1(\cpu.ex.r_epc[7] ));
 sg13g2_nor2_1 _17244_ (.A(_10345_),
    .B(_10386_),
    .Y(_10387_));
 sg13g2_buf_1 _17245_ (.A(net912),
    .X(_10388_));
 sg13g2_and2_1 _17246_ (.A(net693),
    .B(net786),
    .X(_10389_));
 sg13g2_nor2_2 _17247_ (.A(net1048),
    .B(net1046),
    .Y(_10390_));
 sg13g2_buf_1 _17248_ (.A(\cpu.ex.r_sp[7] ),
    .X(_10391_));
 sg13g2_a22oi_1 _17249_ (.Y(_10392_),
    .B1(_10390_),
    .B2(_10391_),
    .A2(_10389_),
    .A1(\cpu.ex.r_11[7] ));
 sg13g2_nor2b_1 _17250_ (.A(net793),
    .B_N(net691),
    .Y(_10393_));
 sg13g2_nor2b_1 _17251_ (.A(_10392_),
    .B_N(_10393_),
    .Y(_10394_));
 sg13g2_nand2b_1 _17252_ (.Y(_10395_),
    .B(net693),
    .A_N(net792));
 sg13g2_a22oi_1 _17253_ (.Y(_10396_),
    .B1(net787),
    .B2(\cpu.ex.r_13[7] ),
    .A2(net917),
    .A1(\cpu.ex.r_lr[7] ));
 sg13g2_nor2_1 _17254_ (.A(_10395_),
    .B(_10396_),
    .Y(_10397_));
 sg13g2_inv_1 _17255_ (.Y(_10398_),
    .A(_00257_));
 sg13g2_and2_1 _17256_ (.A(net1139),
    .B(_10158_),
    .X(_10399_));
 sg13g2_buf_1 _17257_ (.A(_10399_),
    .X(_10400_));
 sg13g2_nand3_1 _17258_ (.B(net693),
    .C(_10400_),
    .A(_10398_),
    .Y(_10401_));
 sg13g2_buf_1 _17259_ (.A(\cpu.dec.user_io ),
    .X(_10402_));
 sg13g2_nor2_2 _17260_ (.A(net792),
    .B(_10388_),
    .Y(_10403_));
 sg13g2_nand3_1 _17261_ (.B(net633),
    .C(_10403_),
    .A(_10402_),
    .Y(_10404_));
 sg13g2_a21oi_1 _17262_ (.A1(_10401_),
    .A2(_10404_),
    .Y(_10405_),
    .B1(net790));
 sg13g2_nor4_1 _17263_ (.A(_10387_),
    .B(_10394_),
    .C(_10397_),
    .D(_10405_),
    .Y(_10406_));
 sg13g2_a21o_1 _17264_ (.A2(_10168_),
    .A1(net918),
    .B1(_10164_),
    .X(_10407_));
 sg13g2_buf_8 _17265_ (.A(_10407_),
    .X(_10408_));
 sg13g2_a21o_1 _17266_ (.A2(_10406_),
    .A1(_10384_),
    .B1(_10408_),
    .X(_10409_));
 sg13g2_a21oi_2 _17267_ (.B1(_10275_),
    .Y(_10410_),
    .A2(_10409_),
    .A1(_10378_));
 sg13g2_buf_2 _17268_ (.A(_00288_),
    .X(_10411_));
 sg13g2_nand2_1 _17269_ (.Y(_10412_),
    .A(\cpu.dec.imm[7] ),
    .B(_10279_));
 sg13g2_o21ai_1 _17270_ (.B1(_10412_),
    .Y(_10413_),
    .A1(net920),
    .A2(_10411_));
 sg13g2_buf_1 _17271_ (.A(_10413_),
    .X(_10414_));
 sg13g2_nor2_1 _17272_ (.A(_10410_),
    .B(_10414_),
    .Y(_10415_));
 sg13g2_mux2_1 _17273_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_10[6] ),
    .S(_10196_),
    .X(_10416_));
 sg13g2_a221oi_1 _17274_ (.B2(net633),
    .C1(_10263_),
    .B1(_10416_),
    .A1(\cpu.ex.r_9[6] ),
    .Y(_10417_),
    .A2(_10224_));
 sg13g2_a221oi_1 _17275_ (.B2(\cpu.ex.r_sp[6] ),
    .C1(_10200_),
    .B1(net789),
    .A1(\cpu.ex.r_lr[6] ),
    .Y(_10418_),
    .A2(_10224_));
 sg13g2_nor3_1 _17276_ (.A(_10201_),
    .B(_10417_),
    .C(_10418_),
    .Y(_10419_));
 sg13g2_inv_1 _17277_ (.Y(_10420_),
    .A(_00256_));
 sg13g2_mux2_1 _17278_ (.A0(\cpu.ex.r_epc[6] ),
    .A1(net1132),
    .S(net793),
    .X(_10421_));
 sg13g2_a22oi_1 _17279_ (.Y(_10422_),
    .B1(_10421_),
    .B2(_10263_),
    .A2(net787),
    .A1(_10420_));
 sg13g2_nor2_1 _17280_ (.A(_10341_),
    .B(_10422_),
    .Y(_10423_));
 sg13g2_nand3_1 _17281_ (.B(net633),
    .C(net795),
    .A(\cpu.ex.r_stmp[6] ),
    .Y(_10424_));
 sg13g2_nand3_1 _17282_ (.B(_10216_),
    .C(_10268_),
    .A(\cpu.ex.r_13[6] ),
    .Y(_10425_));
 sg13g2_a21oi_1 _17283_ (.A1(_10424_),
    .A2(_10425_),
    .Y(_10426_),
    .B1(_10208_));
 sg13g2_nand3_1 _17284_ (.B(net790),
    .C(_10173_),
    .A(\cpu.ex.r_11[6] ),
    .Y(_10427_));
 sg13g2_mux2_1 _17285_ (.A0(\cpu.ex.r_12[6] ),
    .A1(\cpu.ex.r_14[6] ),
    .S(_10197_),
    .X(_10428_));
 sg13g2_nand2_1 _17286_ (.Y(_10429_),
    .A(_10385_),
    .B(_10428_));
 sg13g2_a21oi_1 _17287_ (.A1(_10427_),
    .A2(_10429_),
    .Y(_10430_),
    .B1(_10263_));
 sg13g2_or4_1 _17288_ (.A(_10419_),
    .B(_10423_),
    .C(_10426_),
    .D(_10430_),
    .X(_10431_));
 sg13g2_a221oi_1 _17289_ (.B2(_10431_),
    .C1(net911),
    .B1(_10171_),
    .A1(_09164_),
    .Y(_10432_),
    .A2(net563));
 sg13g2_o21ai_1 _17290_ (.B1(_10135_),
    .Y(_10433_),
    .A1(net1050),
    .A2(\cpu.dec.imm[6] ));
 sg13g2_inv_2 _17291_ (.Y(_10434_),
    .A(_00289_));
 sg13g2_nand2_1 _17292_ (.Y(_10435_),
    .A(net1051),
    .B(_10434_));
 sg13g2_o21ai_1 _17293_ (.B1(_10435_),
    .Y(_10436_),
    .A1(_10432_),
    .A2(_10433_));
 sg13g2_buf_2 _17294_ (.A(_10436_),
    .X(_10437_));
 sg13g2_nor4_1 _17295_ (.A(net1133),
    .B(_10377_),
    .C(_10415_),
    .D(_10437_),
    .Y(_10438_));
 sg13g2_o21ai_1 _17296_ (.B1(_10376_),
    .Y(_10439_),
    .A1(_10410_),
    .A2(_10414_));
 sg13g2_or3_1 _17297_ (.A(_10376_),
    .B(_10410_),
    .C(_10414_),
    .X(_10440_));
 sg13g2_nand2_1 _17298_ (.Y(_10441_),
    .A(_10375_),
    .B(_10437_));
 sg13g2_a21oi_1 _17299_ (.A1(_10439_),
    .A2(_10440_),
    .Y(_10442_),
    .B1(_10441_));
 sg13g2_o21ai_1 _17300_ (.B1(_10126_),
    .Y(_10443_),
    .A1(_10438_),
    .A2(_10442_));
 sg13g2_buf_1 _17301_ (.A(_10415_),
    .X(_10444_));
 sg13g2_nor2_1 _17302_ (.A(_10432_),
    .B(_10433_),
    .Y(_10445_));
 sg13g2_a21oi_1 _17303_ (.A1(_10139_),
    .A2(_10434_),
    .Y(_10446_),
    .B1(_10445_));
 sg13g2_buf_1 _17304_ (.A(_10446_),
    .X(_10447_));
 sg13g2_o21ai_1 _17305_ (.B1(_10126_),
    .Y(_10448_),
    .A1(net1133),
    .A2(net1132));
 sg13g2_nand3_1 _17306_ (.B(net260),
    .C(_10448_),
    .A(net261),
    .Y(_10449_));
 sg13g2_buf_1 _17307_ (.A(\cpu.ex.r_mult[19] ),
    .X(_10450_));
 sg13g2_nand3_1 _17308_ (.B(_10268_),
    .C(_10285_),
    .A(\cpu.ex.r_13[4] ),
    .Y(_10451_));
 sg13g2_mux2_1 _17309_ (.A0(\cpu.ex.r_10[4] ),
    .A1(\cpu.ex.r_14[4] ),
    .S(net914),
    .X(_10452_));
 sg13g2_nand3_1 _17310_ (.B(net789),
    .C(_10452_),
    .A(net786),
    .Y(_10453_));
 sg13g2_nand2_1 _17311_ (.Y(_10454_),
    .A(_10451_),
    .B(_10453_));
 sg13g2_buf_1 _17312_ (.A(\cpu.ex.r_mult[20] ),
    .X(_10455_));
 sg13g2_nor2_1 _17313_ (.A(net794),
    .B(net914),
    .Y(_10456_));
 sg13g2_buf_1 _17314_ (.A(\cpu.ex.r_sp[4] ),
    .X(_10457_));
 sg13g2_a22oi_1 _17315_ (.Y(_10458_),
    .B1(_10456_),
    .B2(_10457_),
    .A2(_10285_),
    .A1(net1130));
 sg13g2_nor2_1 _17316_ (.A(_10345_),
    .B(_10458_),
    .Y(_10459_));
 sg13g2_and2_1 _17317_ (.A(\cpu.ex.r_lr[4] ),
    .B(net915),
    .X(_10460_));
 sg13g2_nor2b_1 _17318_ (.A(net794),
    .B_N(\cpu.ex.r_stmp[4] ),
    .Y(_10461_));
 sg13g2_a22oi_1 _17319_ (.Y(_10462_),
    .B1(_10461_),
    .B2(_10242_),
    .A2(_10460_),
    .A1(_10289_));
 sg13g2_nand3b_1 _17320_ (.B(net912),
    .C(\cpu.ex.r_9[4] ),
    .Y(_10463_),
    .A_N(net913));
 sg13g2_nand3b_1 _17321_ (.B(_10195_),
    .C(\cpu.ex.r_epc[4] ),
    .Y(_10464_),
    .A_N(net912));
 sg13g2_a21o_1 _17322_ (.A2(_10464_),
    .A1(_10463_),
    .B1(_10186_),
    .X(_10465_));
 sg13g2_o21ai_1 _17323_ (.B1(_10465_),
    .Y(_10466_),
    .A1(net786),
    .A2(_10462_));
 sg13g2_or2_1 _17324_ (.X(_10467_),
    .B(net1139),
    .A(_10183_));
 sg13g2_nor2b_1 _17325_ (.A(_10198_),
    .B_N(net1049),
    .Y(_10468_));
 sg13g2_mux2_1 _17326_ (.A0(\cpu.ex.r_8[4] ),
    .A1(\cpu.ex.r_12[4] ),
    .S(_10189_),
    .X(_10469_));
 sg13g2_a22oi_1 _17327_ (.Y(_10470_),
    .B1(_10469_),
    .B2(net786),
    .A2(_10468_),
    .A1(_08274_));
 sg13g2_nor2b_1 _17328_ (.A(_00254_),
    .B_N(net914),
    .Y(_10471_));
 sg13g2_nor2b_1 _17329_ (.A(net914),
    .B_N(\cpu.ex.r_11[4] ),
    .Y(_10472_));
 sg13g2_and3_1 _17330_ (.X(_10473_),
    .A(net794),
    .B(_10195_),
    .C(net912));
 sg13g2_o21ai_1 _17331_ (.B1(_10473_),
    .Y(_10474_),
    .A1(_10471_),
    .A2(_10472_));
 sg13g2_o21ai_1 _17332_ (.B1(_10474_),
    .Y(_10475_),
    .A1(_10467_),
    .A2(_10470_));
 sg13g2_or4_1 _17333_ (.A(_10454_),
    .B(_10459_),
    .C(_10466_),
    .D(_10475_),
    .X(_10476_));
 sg13g2_a221oi_1 _17334_ (.B2(_10476_),
    .C1(net911),
    .B1(_10171_),
    .A1(_09500_),
    .Y(_10477_),
    .A2(net563));
 sg13g2_o21ai_1 _17335_ (.B1(_10134_),
    .Y(_10478_),
    .A1(_10140_),
    .A2(\cpu.dec.imm[4] ));
 sg13g2_nand2_1 _17336_ (.Y(_10479_),
    .A(net1076),
    .B(net1051));
 sg13g2_o21ai_1 _17337_ (.B1(_10479_),
    .Y(_10480_),
    .A1(_10477_),
    .A2(_10478_));
 sg13g2_buf_2 _17338_ (.A(_10480_),
    .X(_10481_));
 sg13g2_nand2_1 _17339_ (.Y(_10482_),
    .A(net1131),
    .B(_10481_));
 sg13g2_nor2b_1 _17340_ (.A(_00255_),
    .B_N(net794),
    .Y(_10483_));
 sg13g2_buf_1 _17341_ (.A(\cpu.ex.r_sp[5] ),
    .X(_10484_));
 sg13g2_nor2b_1 _17342_ (.A(net693),
    .B_N(_10484_),
    .Y(_10485_));
 sg13g2_a22oi_1 _17343_ (.Y(_10486_),
    .B1(_10485_),
    .B2(_10168_),
    .A2(_10483_),
    .A1(_10248_));
 sg13g2_nand3b_1 _17344_ (.B(net914),
    .C(\cpu.ex.r_13[5] ),
    .Y(_10487_),
    .A_N(net792));
 sg13g2_nand3b_1 _17345_ (.B(net792),
    .C(\cpu.ex.r_11[5] ),
    .Y(_10488_),
    .A_N(net914));
 sg13g2_nand2_1 _17346_ (.Y(_10489_),
    .A(net794),
    .B(_10199_));
 sg13g2_a21o_1 _17347_ (.A2(_10488_),
    .A1(_10487_),
    .B1(_10489_),
    .X(_10490_));
 sg13g2_o21ai_1 _17348_ (.B1(_10490_),
    .Y(_10491_),
    .A1(_10245_),
    .A2(_10486_));
 sg13g2_mux2_1 _17349_ (.A0(\cpu.ex.r_stmp[5] ),
    .A1(\cpu.ex.r_14[5] ),
    .S(net912),
    .X(_10492_));
 sg13g2_a22oi_1 _17350_ (.Y(_10493_),
    .B1(_10492_),
    .B2(_10197_),
    .A2(_10268_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_nor2b_1 _17351_ (.A(_10493_),
    .B_N(_10385_),
    .Y(_10494_));
 sg13g2_nand3_1 _17352_ (.B(net793),
    .C(_10179_),
    .A(_10375_),
    .Y(_10495_));
 sg13g2_nand3_1 _17353_ (.B(net788),
    .C(_10176_),
    .A(\cpu.ex.r_9[5] ),
    .Y(_10496_));
 sg13g2_a21oi_1 _17354_ (.A1(_10495_),
    .A2(_10496_),
    .Y(_10497_),
    .B1(net633));
 sg13g2_nor2b_1 _17355_ (.A(_10199_),
    .B_N(_10184_),
    .Y(_10498_));
 sg13g2_mux2_1 _17356_ (.A0(\cpu.ex.r_lr[5] ),
    .A1(\cpu.ex.r_epc[5] ),
    .S(net792),
    .X(_10499_));
 sg13g2_mux2_1 _17357_ (.A0(\cpu.ex.r_8[5] ),
    .A1(\cpu.ex.r_10[5] ),
    .S(net792),
    .X(_10500_));
 sg13g2_a22oi_1 _17358_ (.Y(_10501_),
    .B1(_10500_),
    .B2(_10324_),
    .A2(_10499_),
    .A1(_10498_));
 sg13g2_nor2_1 _17359_ (.A(net692),
    .B(_10501_),
    .Y(_10502_));
 sg13g2_nor4_1 _17360_ (.A(_10491_),
    .B(_10494_),
    .C(_10497_),
    .D(_10502_),
    .Y(_10503_));
 sg13g2_nand2_1 _17361_ (.Y(_10504_),
    .A(_09893_),
    .B(_10165_));
 sg13g2_o21ai_1 _17362_ (.B1(_10504_),
    .Y(_10505_),
    .A1(_10408_),
    .A2(_10503_));
 sg13g2_buf_2 _17363_ (.A(_10505_),
    .X(_10506_));
 sg13g2_buf_2 _17364_ (.A(_00290_),
    .X(_10507_));
 sg13g2_nand2_1 _17365_ (.Y(_10508_),
    .A(\cpu.dec.imm[5] ),
    .B(_10279_));
 sg13g2_o21ai_1 _17366_ (.B1(_10508_),
    .Y(_10509_),
    .A1(net920),
    .A2(_10507_));
 sg13g2_a21oi_1 _17367_ (.A1(_10308_),
    .A2(_10506_),
    .Y(_10510_),
    .B1(_10509_));
 sg13g2_buf_1 _17368_ (.A(_10510_),
    .X(_10511_));
 sg13g2_xnor2_1 _17369_ (.Y(_10512_),
    .A(net1130),
    .B(_10511_));
 sg13g2_inv_2 _17370_ (.Y(_10513_),
    .A(net1130));
 sg13g2_or4_1 _17371_ (.A(net1131),
    .B(_10513_),
    .C(_10481_),
    .D(_10511_),
    .X(_10514_));
 sg13g2_o21ai_1 _17372_ (.B1(_10514_),
    .Y(_10515_),
    .A1(_10482_),
    .A2(_10512_));
 sg13g2_o21ai_1 _17373_ (.B1(_10126_),
    .Y(_10516_),
    .A1(_10450_),
    .A2(net1130));
 sg13g2_buf_1 _17374_ (.A(_10481_),
    .X(_10517_));
 sg13g2_a21o_1 _17375_ (.A2(_10506_),
    .A1(_10308_),
    .B1(_10509_),
    .X(_10518_));
 sg13g2_buf_2 _17376_ (.A(_10518_),
    .X(_10519_));
 sg13g2_buf_1 _17377_ (.A(_10519_),
    .X(_10520_));
 sg13g2_nor2_1 _17378_ (.A(net303),
    .B(net232),
    .Y(_10521_));
 sg13g2_a22oi_1 _17379_ (.Y(_10522_),
    .B1(_10516_),
    .B2(_10521_),
    .A2(_10515_),
    .A1(_10126_));
 sg13g2_buf_1 _17380_ (.A(_10522_),
    .X(_10523_));
 sg13g2_a21o_1 _17381_ (.A2(_10449_),
    .A1(_10443_),
    .B1(_10523_),
    .X(_10524_));
 sg13g2_and2_1 _17382_ (.A(\cpu.ex.r_lr[2] ),
    .B(_10237_),
    .X(_10525_));
 sg13g2_nand2_1 _17383_ (.Y(_10526_),
    .A(net1046),
    .B(net1049));
 sg13g2_nor3_1 _17384_ (.A(_00252_),
    .B(_10244_),
    .C(_10526_),
    .Y(_10527_));
 sg13g2_o21ai_1 _17385_ (.B1(_10187_),
    .Y(_10528_),
    .A1(_10525_),
    .A2(_10527_));
 sg13g2_buf_1 _17386_ (.A(\cpu.ex.r_sp[2] ),
    .X(_10529_));
 sg13g2_nand3_1 _17387_ (.B(net1047),
    .C(_10168_),
    .A(_10529_),
    .Y(_10530_));
 sg13g2_nand3_1 _17388_ (.B(_10244_),
    .C(_10247_),
    .A(\cpu.ex.r_12[2] ),
    .Y(_10531_));
 sg13g2_a21o_1 _17389_ (.A2(_10531_),
    .A1(_10530_),
    .B1(net915),
    .X(_10532_));
 sg13g2_buf_1 _17390_ (.A(\cpu.ex.mmu_read[2] ),
    .X(_10533_));
 sg13g2_mux2_1 _17391_ (.A0(_10533_),
    .A1(\cpu.ex.r_13[2] ),
    .S(net1046),
    .X(_10534_));
 sg13g2_nand3_1 _17392_ (.B(_10224_),
    .C(_10534_),
    .A(net1049),
    .Y(_10535_));
 sg13g2_mux2_1 _17393_ (.A0(\cpu.ex.r_epc[2] ),
    .A1(\cpu.ex.r_11[2] ),
    .S(net1138),
    .X(_10536_));
 sg13g2_nand3_1 _17394_ (.B(_10173_),
    .C(_10536_),
    .A(_10207_),
    .Y(_10537_));
 sg13g2_nand3_1 _17395_ (.B(_10179_),
    .C(_10385_),
    .A(\cpu.ex.r_stmp[2] ),
    .Y(_10538_));
 sg13g2_and3_1 _17396_ (.X(_10539_),
    .A(_10535_),
    .B(_10537_),
    .C(_10538_));
 sg13g2_buf_1 _17397_ (.A(\cpu.ex.r_mult[18] ),
    .X(_10540_));
 sg13g2_nand3_1 _17398_ (.B(_10183_),
    .C(net1047),
    .A(_10540_),
    .Y(_10541_));
 sg13g2_o21ai_1 _17399_ (.B1(_10541_),
    .Y(_10542_),
    .A1(_08437_),
    .A2(_10467_));
 sg13g2_mux2_1 _17400_ (.A0(\cpu.ex.r_8[2] ),
    .A1(\cpu.ex.r_9[2] ),
    .S(_10184_),
    .X(_10543_));
 sg13g2_mux2_1 _17401_ (.A0(\cpu.ex.r_10[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net1140),
    .X(_10544_));
 sg13g2_and3_1 _17402_ (.X(_10545_),
    .A(_10198_),
    .B(_10209_),
    .C(_10544_));
 sg13g2_a221oi_1 _17403_ (.B2(_10380_),
    .C1(_10545_),
    .B1(_10543_),
    .A1(_10468_),
    .Y(_10546_),
    .A2(_10542_));
 sg13g2_and4_1 _17404_ (.A(_10528_),
    .B(_10532_),
    .C(_10539_),
    .D(_10546_),
    .X(_10547_));
 sg13g2_nand2_1 _17405_ (.Y(_10548_),
    .A(_09173_),
    .B(_10164_));
 sg13g2_o21ai_1 _17406_ (.B1(_10548_),
    .Y(_10549_),
    .A1(_10408_),
    .A2(_10547_));
 sg13g2_buf_2 _17407_ (.A(_10549_),
    .X(_10550_));
 sg13g2_buf_1 _17408_ (.A(\cpu.dec.imm[2] ),
    .X(_10551_));
 sg13g2_nand3_1 _17409_ (.B(_10134_),
    .C(net911),
    .A(_10551_),
    .Y(_10552_));
 sg13g2_o21ai_1 _17410_ (.B1(_10552_),
    .Y(_10553_),
    .A1(_10134_),
    .A2(_00283_));
 sg13g2_a21o_1 _17411_ (.A2(_10550_),
    .A1(_10308_),
    .B1(_10553_),
    .X(_10554_));
 sg13g2_buf_2 _17412_ (.A(_10554_),
    .X(_10555_));
 sg13g2_buf_1 _17413_ (.A(\cpu.ex.r_mult[17] ),
    .X(_10556_));
 sg13g2_buf_1 _17414_ (.A(_10556_),
    .X(_10557_));
 sg13g2_nand2_1 _17415_ (.Y(_10558_),
    .A(net1044),
    .B(_10126_));
 sg13g2_or2_1 _17416_ (.X(_10559_),
    .B(_10558_),
    .A(_10555_));
 sg13g2_buf_1 _17417_ (.A(_10559_),
    .X(_10560_));
 sg13g2_buf_2 _17418_ (.A(\cpu.ex.r_mult[16] ),
    .X(_10561_));
 sg13g2_inv_1 _17419_ (.Y(_10562_),
    .A(_10561_));
 sg13g2_buf_1 _17420_ (.A(_00198_),
    .X(_10563_));
 sg13g2_nand2b_1 _17421_ (.Y(_10564_),
    .B(net1051),
    .A_N(_10563_));
 sg13g2_buf_1 _17422_ (.A(_10564_),
    .X(_10565_));
 sg13g2_mux2_1 _17423_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(net1140),
    .X(_10566_));
 sg13g2_a22oi_1 _17424_ (.Y(_10567_),
    .B1(_10566_),
    .B2(_10263_),
    .A2(net916),
    .A1(\cpu.ex.r_9[1] ));
 sg13g2_nand3b_1 _17425_ (.B(net1047),
    .C(net787),
    .Y(_10568_),
    .A_N(_00251_));
 sg13g2_o21ai_1 _17426_ (.B1(_10568_),
    .Y(_10569_),
    .A1(net913),
    .A2(_10567_));
 sg13g2_buf_1 _17427_ (.A(\cpu.ex.r_sp[1] ),
    .X(_10570_));
 sg13g2_mux2_1 _17428_ (.A0(_10570_),
    .A1(\cpu.ex.r_epc[1] ),
    .S(net1048),
    .X(_10571_));
 sg13g2_mux2_1 _17429_ (.A0(\cpu.ex.r_10[1] ),
    .A1(\cpu.ex.r_11[1] ),
    .S(net1048),
    .X(_10572_));
 sg13g2_a22oi_1 _17430_ (.Y(_10573_),
    .B1(_10400_),
    .B2(_10572_),
    .A2(_10571_),
    .A1(_10179_));
 sg13g2_inv_1 _17431_ (.Y(_10574_),
    .A(_10573_));
 sg13g2_nand3b_1 _17432_ (.B(net1047),
    .C(\cpu.ex.r_14[1] ),
    .Y(_10575_),
    .A_N(net1048));
 sg13g2_nand3b_1 _17433_ (.B(net915),
    .C(\cpu.ex.r_13[1] ),
    .Y(_10576_),
    .A_N(net1047));
 sg13g2_a21o_1 _17434_ (.A2(_10576_),
    .A1(_10575_),
    .B1(_10526_),
    .X(_10577_));
 sg13g2_mux2_1 _17435_ (.A0(\cpu.ex.r_8[1] ),
    .A1(\cpu.ex.r_12[1] ),
    .S(net1049),
    .X(_10578_));
 sg13g2_nand3_1 _17436_ (.B(net918),
    .C(_10578_),
    .A(net1046),
    .Y(_10579_));
 sg13g2_buf_1 _17437_ (.A(\cpu.ex.r_prev_ie ),
    .X(_10580_));
 sg13g2_mux2_1 _17438_ (.A0(_10580_),
    .A1(\cpu.ex.r_stmp[1] ),
    .S(net1047),
    .X(_10581_));
 sg13g2_nand3_1 _17439_ (.B(_10390_),
    .C(_10581_),
    .A(net1049),
    .Y(_10582_));
 sg13g2_nand3_1 _17440_ (.B(_10179_),
    .C(_10285_),
    .A(_10556_),
    .Y(_10583_));
 sg13g2_nand4_1 _17441_ (.B(_10579_),
    .C(_10582_),
    .A(_10577_),
    .Y(_10584_),
    .D(_10583_));
 sg13g2_a221oi_1 _17442_ (.B2(_10207_),
    .C1(_10584_),
    .B1(_10574_),
    .A1(_10188_),
    .Y(_10585_),
    .A2(_10569_));
 sg13g2_nand2_1 _17443_ (.Y(_10586_),
    .A(_09177_),
    .B(_10164_));
 sg13g2_o21ai_1 _17444_ (.B1(_10586_),
    .Y(_10587_),
    .A1(_10408_),
    .A2(_10585_));
 sg13g2_buf_1 _17445_ (.A(_10587_),
    .X(_10588_));
 sg13g2_buf_1 _17446_ (.A(\cpu.dec.imm[1] ),
    .X(_10589_));
 sg13g2_inv_1 _17447_ (.Y(_10590_),
    .A(_10589_));
 sg13g2_a21oi_1 _17448_ (.A1(_10590_),
    .A2(net911),
    .Y(_10591_),
    .B1(net1051));
 sg13g2_o21ai_1 _17449_ (.B1(_10591_),
    .Y(_10592_),
    .A1(net911),
    .A2(_10588_));
 sg13g2_nand2_1 _17450_ (.Y(_10593_),
    .A(_10565_),
    .B(_10592_));
 sg13g2_buf_2 _17451_ (.A(_10593_),
    .X(_10594_));
 sg13g2_a21oi_1 _17452_ (.A1(_10308_),
    .A2(_10550_),
    .Y(_10595_),
    .B1(_10553_));
 sg13g2_buf_8 _17453_ (.A(_10595_),
    .X(_10596_));
 sg13g2_nand3_1 _17454_ (.B(_10565_),
    .C(_10592_),
    .A(_10596_),
    .Y(_10597_));
 sg13g2_buf_2 _17455_ (.A(_10597_),
    .X(_10598_));
 sg13g2_nor2_1 _17456_ (.A(net1044),
    .B(_10596_),
    .Y(_10599_));
 sg13g2_a221oi_1 _17457_ (.B2(_09290_),
    .C1(_10599_),
    .B1(_10598_),
    .A1(_10562_),
    .Y(_10600_),
    .A2(_10594_));
 sg13g2_buf_1 _17458_ (.A(_10600_),
    .X(_10601_));
 sg13g2_inv_1 _17459_ (.Y(_10602_),
    .A(_10601_));
 sg13g2_nand2_1 _17460_ (.Y(_10603_),
    .A(_10540_),
    .B(_10126_));
 sg13g2_a21oi_1 _17461_ (.A1(_10560_),
    .A2(_10602_),
    .Y(_10604_),
    .B1(_10603_));
 sg13g2_nand2b_1 _17462_ (.Y(_10605_),
    .B(_08357_),
    .A_N(_08351_));
 sg13g2_buf_8 _17463_ (.A(_10605_),
    .X(_10606_));
 sg13g2_nand4_1 _17464_ (.B(_08386_),
    .C(_08401_),
    .A(_08373_),
    .Y(_10607_),
    .D(_08413_));
 sg13g2_buf_8 _17465_ (.A(_10607_),
    .X(_10608_));
 sg13g2_buf_1 _17466_ (.A(_00266_),
    .X(_10609_));
 sg13g2_buf_8 _17467_ (.A(\cpu.dec.r_rs1[0] ),
    .X(_10610_));
 sg13g2_buf_2 _17468_ (.A(\cpu.dec.r_rs1[1] ),
    .X(_10611_));
 sg13g2_buf_8 _17469_ (.A(\cpu.dec.r_rs1[3] ),
    .X(_10612_));
 sg13g2_buf_8 _17470_ (.A(\cpu.dec.r_rs1[2] ),
    .X(_10613_));
 sg13g2_nor4_2 _17471_ (.A(_10610_),
    .B(_10611_),
    .C(net1129),
    .Y(_10614_),
    .D(net1128));
 sg13g2_nor3_1 _17472_ (.A(_09110_),
    .B(_10609_),
    .C(_10614_),
    .Y(_10615_));
 sg13g2_nand4_1 _17473_ (.B(_09135_),
    .C(_09154_),
    .A(_09123_),
    .Y(_10616_),
    .D(_10615_));
 sg13g2_nor4_1 _17474_ (.A(_09110_),
    .B(_09155_),
    .C(_10609_),
    .D(_10614_),
    .Y(_10617_));
 sg13g2_nor4_1 _17475_ (.A(_09110_),
    .B(_09158_),
    .C(_10609_),
    .D(_10614_),
    .Y(_10618_));
 sg13g2_a21oi_1 _17476_ (.A1(_09123_),
    .A2(_10617_),
    .Y(_10619_),
    .B1(_10618_));
 sg13g2_nand2_1 _17477_ (.Y(_10620_),
    .A(_10616_),
    .B(_10619_));
 sg13g2_buf_8 _17478_ (.A(_10620_),
    .X(_10621_));
 sg13g2_and2_1 _17479_ (.A(_08299_),
    .B(_10621_),
    .X(_10622_));
 sg13g2_buf_8 _17480_ (.A(_10622_),
    .X(_10623_));
 sg13g2_nand3_1 _17481_ (.B(net438),
    .C(_10623_),
    .A(net439),
    .Y(_10624_));
 sg13g2_buf_8 _17482_ (.A(_10624_),
    .X(_10625_));
 sg13g2_buf_1 _17483_ (.A(\cpu.br ),
    .X(_10626_));
 sg13g2_inv_1 _17484_ (.Y(_10627_),
    .A(net1127));
 sg13g2_buf_1 _17485_ (.A(_10627_),
    .X(_10628_));
 sg13g2_nor2_1 _17486_ (.A(net910),
    .B(_00193_),
    .Y(_10629_));
 sg13g2_inv_1 _17487_ (.Y(_10630_),
    .A(_10621_));
 sg13g2_buf_1 _17488_ (.A(_10630_),
    .X(_10631_));
 sg13g2_xnor2_1 _17489_ (.Y(_10632_),
    .A(net1141),
    .B(_10612_));
 sg13g2_buf_8 _17490_ (.A(_10145_),
    .X(_10633_));
 sg13g2_xnor2_1 _17491_ (.Y(_10634_),
    .A(net1043),
    .B(_10610_));
 sg13g2_xnor2_1 _17492_ (.Y(_10635_),
    .A(_10148_),
    .B(net1128));
 sg13g2_xnor2_1 _17493_ (.Y(_10636_),
    .A(net1142),
    .B(_10611_));
 sg13g2_nand4_1 _17494_ (.B(_10634_),
    .C(_10635_),
    .A(_10632_),
    .Y(_10637_),
    .D(_10636_));
 sg13g2_nor2_1 _17495_ (.A(_10153_),
    .B(_10637_),
    .Y(_10638_));
 sg13g2_buf_1 _17496_ (.A(_10638_),
    .X(_10639_));
 sg13g2_buf_8 _17497_ (.A(_10612_),
    .X(_10640_));
 sg13g2_inv_1 _17498_ (.Y(_10641_),
    .A(net1042));
 sg13g2_buf_1 _17499_ (.A(_10641_),
    .X(_10642_));
 sg13g2_nor2b_1 _17500_ (.A(_10611_),
    .B_N(_10610_),
    .Y(_10643_));
 sg13g2_buf_1 _17501_ (.A(_10643_),
    .X(_10644_));
 sg13g2_nand3_1 _17502_ (.B(\cpu.ex.mmu_read[14] ),
    .C(net909),
    .A(_10642_),
    .Y(_10645_));
 sg13g2_buf_8 _17503_ (.A(net1042),
    .X(_10646_));
 sg13g2_buf_1 _17504_ (.A(net908),
    .X(_10647_));
 sg13g2_nor2b_1 _17505_ (.A(_10610_),
    .B_N(_10611_),
    .Y(_10648_));
 sg13g2_buf_1 _17506_ (.A(_10648_),
    .X(_10649_));
 sg13g2_buf_1 _17507_ (.A(_10649_),
    .X(_10650_));
 sg13g2_nand3_1 _17508_ (.B(\cpu.ex.r_14[14] ),
    .C(net783),
    .A(net784),
    .Y(_10651_));
 sg13g2_inv_2 _17509_ (.Y(_10652_),
    .A(net1128));
 sg13g2_buf_1 _17510_ (.A(_10652_),
    .X(_10653_));
 sg13g2_buf_8 _17511_ (.A(net907),
    .X(_10654_));
 sg13g2_buf_1 _17512_ (.A(net782),
    .X(_10655_));
 sg13g2_a21oi_1 _17513_ (.A1(_10645_),
    .A2(_10651_),
    .Y(_10656_),
    .B1(_10655_));
 sg13g2_nor2b_1 _17514_ (.A(_10610_),
    .B_N(net1129),
    .Y(_10657_));
 sg13g2_buf_2 _17515_ (.A(_10657_),
    .X(_10658_));
 sg13g2_and3_1 _17516_ (.X(_10659_),
    .A(_10653_),
    .B(\cpu.ex.r_10[14] ),
    .C(_10658_));
 sg13g2_buf_8 _17517_ (.A(_10610_),
    .X(_10660_));
 sg13g2_buf_8 _17518_ (.A(net1041),
    .X(_10661_));
 sg13g2_buf_1 _17519_ (.A(\cpu.ex.r_mult[30] ),
    .X(_10662_));
 sg13g2_nor2b_1 _17520_ (.A(net1129),
    .B_N(net1128),
    .Y(_10663_));
 sg13g2_buf_2 _17521_ (.A(_10663_),
    .X(_10664_));
 sg13g2_and3_1 _17522_ (.X(_10665_),
    .A(net906),
    .B(net1126),
    .C(_10664_));
 sg13g2_buf_8 _17523_ (.A(_10611_),
    .X(_10666_));
 sg13g2_buf_8 _17524_ (.A(net1040),
    .X(_10667_));
 sg13g2_buf_8 _17525_ (.A(net905),
    .X(_10668_));
 sg13g2_o21ai_1 _17526_ (.B1(net781),
    .Y(_10669_),
    .A1(_10659_),
    .A2(_10665_));
 sg13g2_inv_1 _17527_ (.Y(_10670_),
    .A(\cpu.ex.r_11[14] ));
 sg13g2_buf_8 _17528_ (.A(_10613_),
    .X(_10671_));
 sg13g2_buf_8 _17529_ (.A(net1041),
    .X(_10672_));
 sg13g2_nand3b_1 _17530_ (.B(net1040),
    .C(net904),
    .Y(_10673_),
    .A_N(_10671_));
 sg13g2_nor2_1 _17531_ (.A(_10670_),
    .B(_10673_),
    .Y(_10674_));
 sg13g2_buf_8 _17532_ (.A(net1039),
    .X(_10675_));
 sg13g2_buf_8 _17533_ (.A(_10675_),
    .X(_10676_));
 sg13g2_nor2_1 _17534_ (.A(_10660_),
    .B(_10666_),
    .Y(_10677_));
 sg13g2_buf_2 _17535_ (.A(_10677_),
    .X(_10678_));
 sg13g2_and3_1 _17536_ (.X(_10679_),
    .A(net780),
    .B(\cpu.ex.r_12[14] ),
    .C(_10678_));
 sg13g2_buf_1 _17537_ (.A(net908),
    .X(_10680_));
 sg13g2_o21ai_1 _17538_ (.B1(net779),
    .Y(_10681_),
    .A1(_10674_),
    .A2(_10679_));
 sg13g2_nor2_1 _17539_ (.A(net904),
    .B(net1042),
    .Y(_10682_));
 sg13g2_and2_1 _17540_ (.A(net1041),
    .B(net1042),
    .X(_10683_));
 sg13g2_buf_2 _17541_ (.A(_10683_),
    .X(_10684_));
 sg13g2_inv_1 _17542_ (.Y(_10685_),
    .A(_00264_));
 sg13g2_a22oi_1 _17543_ (.Y(_10686_),
    .B1(_10684_),
    .B2(_10685_),
    .A2(_10682_),
    .A1(\cpu.ex.r_stmp[14] ));
 sg13g2_and2_1 _17544_ (.A(net1040),
    .B(net1039),
    .X(_10687_));
 sg13g2_buf_2 _17545_ (.A(_10687_),
    .X(_10688_));
 sg13g2_nand2b_1 _17546_ (.Y(_10689_),
    .B(_10688_),
    .A_N(_10686_));
 sg13g2_nor2b_1 _17547_ (.A(net1040),
    .B_N(net1129),
    .Y(_10690_));
 sg13g2_buf_2 _17548_ (.A(_10690_),
    .X(_10691_));
 sg13g2_nor2_1 _17549_ (.A(_10660_),
    .B(net1039),
    .Y(_10692_));
 sg13g2_buf_2 _17550_ (.A(_10692_),
    .X(_10693_));
 sg13g2_and3_1 _17551_ (.X(_10694_),
    .A(_10672_),
    .B(net1039),
    .C(\cpu.ex.r_13[14] ));
 sg13g2_a21o_1 _17552_ (.A2(_10693_),
    .A1(\cpu.ex.r_8[14] ),
    .B1(_10694_),
    .X(_10695_));
 sg13g2_buf_8 _17553_ (.A(net1040),
    .X(_10696_));
 sg13g2_buf_1 _17554_ (.A(\cpu.ex.r_sp[14] ),
    .X(_10697_));
 sg13g2_nand3b_1 _17555_ (.B(net902),
    .C(_10697_),
    .Y(_10698_),
    .A_N(net904));
 sg13g2_nand3b_1 _17556_ (.B(\cpu.ex.r_lr[14] ),
    .C(_10661_),
    .Y(_10699_),
    .A_N(net902));
 sg13g2_or2_1 _17557_ (.X(_10700_),
    .B(_10671_),
    .A(_10640_));
 sg13g2_buf_1 _17558_ (.A(_10700_),
    .X(_10701_));
 sg13g2_a21oi_1 _17559_ (.A1(_10698_),
    .A2(_10699_),
    .Y(_10702_),
    .B1(_10701_));
 sg13g2_a21oi_1 _17560_ (.A1(_10691_),
    .A2(_10695_),
    .Y(_10703_),
    .B1(_10702_));
 sg13g2_nand4_1 _17561_ (.B(_10681_),
    .C(_10689_),
    .A(_10669_),
    .Y(_10704_),
    .D(_10703_));
 sg13g2_buf_1 _17562_ (.A(_10691_),
    .X(_10705_));
 sg13g2_nor2b_1 _17563_ (.A(net1129),
    .B_N(_10611_),
    .Y(_10706_));
 sg13g2_buf_2 _17564_ (.A(_10706_),
    .X(_10707_));
 sg13g2_a22oi_1 _17565_ (.Y(_10708_),
    .B1(_10707_),
    .B2(\cpu.ex.r_epc[14] ),
    .A2(net688),
    .A1(\cpu.ex.r_9[14] ));
 sg13g2_nor2b_1 _17566_ (.A(net1039),
    .B_N(net1041),
    .Y(_10709_));
 sg13g2_nor2b_1 _17567_ (.A(_10708_),
    .B_N(_10709_),
    .Y(_10710_));
 sg13g2_nor4_2 _17568_ (.A(net629),
    .B(_10656_),
    .C(_10704_),
    .Y(_10711_),
    .D(_10710_));
 sg13g2_or2_1 _17569_ (.X(_10712_),
    .B(_10637_),
    .A(_10153_));
 sg13g2_buf_2 _17570_ (.A(_10712_),
    .X(_10713_));
 sg13g2_nor2_1 _17571_ (.A(net809),
    .B(_10713_),
    .Y(_10714_));
 sg13g2_nor4_1 _17572_ (.A(_09108_),
    .B(net437),
    .C(_10711_),
    .D(_10714_),
    .Y(_10715_));
 sg13g2_nor3_1 _17573_ (.A(net1127),
    .B(_10711_),
    .C(_10714_),
    .Y(_10716_));
 sg13g2_a221oi_1 _17574_ (.B2(net358),
    .C1(_10716_),
    .B1(_10715_),
    .A1(_10625_),
    .Y(_10717_),
    .A2(_10629_));
 sg13g2_buf_1 _17575_ (.A(_10717_),
    .X(_10718_));
 sg13g2_and2_1 _17576_ (.A(_09276_),
    .B(_09273_),
    .X(_10719_));
 sg13g2_nor2_1 _17577_ (.A(_09276_),
    .B(_09273_),
    .Y(_10720_));
 sg13g2_inv_1 _17578_ (.Y(_10721_),
    .A(_10720_));
 sg13g2_nand4_1 _17579_ (.B(_09275_),
    .C(net646),
    .A(_09274_),
    .Y(_10722_),
    .D(_10721_));
 sg13g2_a21o_1 _17580_ (.A2(_10719_),
    .A1(_10718_),
    .B1(_10722_),
    .X(_10723_));
 sg13g2_buf_1 _17581_ (.A(net910),
    .X(_10724_));
 sg13g2_nor4_1 _17582_ (.A(_09108_),
    .B(_08359_),
    .C(_08415_),
    .D(net437),
    .Y(_10725_));
 sg13g2_buf_2 _17583_ (.A(_10725_),
    .X(_10726_));
 sg13g2_nor3_1 _17584_ (.A(net778),
    .B(_00192_),
    .C(_10726_),
    .Y(_10727_));
 sg13g2_buf_1 _17585_ (.A(_10626_),
    .X(_10728_));
 sg13g2_buf_8 _17586_ (.A(_10625_),
    .X(_10729_));
 sg13g2_buf_1 _17587_ (.A(net808),
    .X(_10730_));
 sg13g2_buf_1 _17588_ (.A(_10713_),
    .X(_10731_));
 sg13g2_buf_1 _17589_ (.A(_10661_),
    .X(_10732_));
 sg13g2_buf_8 _17590_ (.A(net777),
    .X(_10733_));
 sg13g2_buf_1 _17591_ (.A(\cpu.ex.r_sp[15] ),
    .X(_10734_));
 sg13g2_and2_1 _17592_ (.A(net779),
    .B(\cpu.ex.r_10[15] ),
    .X(_10735_));
 sg13g2_a21oi_1 _17593_ (.A1(net785),
    .A2(_10734_),
    .Y(_10736_),
    .B1(_10735_));
 sg13g2_buf_2 _17594_ (.A(net785),
    .X(_10737_));
 sg13g2_nand3_1 _17595_ (.B(net685),
    .C(\cpu.ex.r_epc[15] ),
    .A(net686),
    .Y(_10738_));
 sg13g2_o21ai_1 _17596_ (.B1(_10738_),
    .Y(_10739_),
    .A1(net686),
    .A2(_10736_));
 sg13g2_nor2b_2 _17597_ (.A(_10676_),
    .B_N(net905),
    .Y(_10740_));
 sg13g2_nand2b_1 _17598_ (.Y(_10741_),
    .B(net904),
    .A_N(net902));
 sg13g2_buf_1 _17599_ (.A(_10741_),
    .X(_10742_));
 sg13g2_buf_1 _17600_ (.A(\cpu.ex.mmu_read[15] ),
    .X(_10743_));
 sg13g2_buf_1 _17601_ (.A(net780),
    .X(_10744_));
 sg13g2_mux2_1 _17602_ (.A0(\cpu.ex.r_lr[15] ),
    .A1(net1125),
    .S(net684),
    .X(_10745_));
 sg13g2_and2_1 _17603_ (.A(net1129),
    .B(net1128),
    .X(_10746_));
 sg13g2_buf_2 _17604_ (.A(_10746_),
    .X(_10747_));
 sg13g2_a22oi_1 _17605_ (.Y(_10748_),
    .B1(_10747_),
    .B2(\cpu.ex.r_13[15] ),
    .A2(_10745_),
    .A1(net685));
 sg13g2_nor2_1 _17606_ (.A(_10742_),
    .B(_10748_),
    .Y(_10749_));
 sg13g2_a21oi_1 _17607_ (.A1(_10739_),
    .A2(_10740_),
    .Y(_10750_),
    .B1(_10749_));
 sg13g2_and2_1 _17608_ (.A(net1041),
    .B(net1040),
    .X(_10751_));
 sg13g2_buf_2 _17609_ (.A(_10751_),
    .X(_10752_));
 sg13g2_buf_8 _17610_ (.A(_10752_),
    .X(_10753_));
 sg13g2_a22oi_1 _17611_ (.Y(_10754_),
    .B1(net683),
    .B2(\cpu.ex.r_11[15] ),
    .A2(_10678_),
    .A1(\cpu.ex.r_8[15] ));
 sg13g2_nor2_1 _17612_ (.A(net684),
    .B(_10754_),
    .Y(_10755_));
 sg13g2_buf_1 _17613_ (.A(net905),
    .X(_10756_));
 sg13g2_buf_8 _17614_ (.A(_10675_),
    .X(_10757_));
 sg13g2_nor2b_1 _17615_ (.A(net777),
    .B_N(net775),
    .Y(_10758_));
 sg13g2_a22oi_1 _17616_ (.Y(_10759_),
    .B1(_10758_),
    .B2(\cpu.ex.r_12[15] ),
    .A2(_10709_),
    .A1(\cpu.ex.r_9[15] ));
 sg13g2_nor2_1 _17617_ (.A(net776),
    .B(_10759_),
    .Y(_10760_));
 sg13g2_buf_1 _17618_ (.A(_10680_),
    .X(_10761_));
 sg13g2_o21ai_1 _17619_ (.B1(net682),
    .Y(_10762_),
    .A1(_10755_),
    .A2(_10760_));
 sg13g2_inv_1 _17620_ (.Y(_10763_),
    .A(_00265_));
 sg13g2_inv_2 _17621_ (.Y(_10764_),
    .A(net904));
 sg13g2_buf_8 _17622_ (.A(_10764_),
    .X(_10765_));
 sg13g2_mux4_1 _17623_ (.S0(net681),
    .A0(_10763_),
    .A1(\cpu.ex.r_14[15] ),
    .A2(\cpu.ex.r_mult[31] ),
    .A3(\cpu.ex.r_stmp[15] ),
    .S1(net685),
    .X(_10766_));
 sg13g2_nand2_1 _17624_ (.Y(_10767_),
    .A(_10688_),
    .B(_10766_));
 sg13g2_nand4_1 _17625_ (.B(_10750_),
    .C(_10762_),
    .A(net559),
    .Y(_10768_),
    .D(_10767_));
 sg13g2_o21ai_1 _17626_ (.B1(_10768_),
    .Y(_10769_),
    .A1(net687),
    .A2(net559));
 sg13g2_a21oi_1 _17627_ (.A1(_10728_),
    .A2(net301),
    .Y(_10770_),
    .B1(_10769_));
 sg13g2_nand2b_1 _17628_ (.Y(_10771_),
    .B(_10720_),
    .A_N(_09274_));
 sg13g2_o21ai_1 _17629_ (.B1(_09284_),
    .Y(_10772_),
    .A1(_09275_),
    .A2(_10771_));
 sg13g2_o21ai_1 _17630_ (.B1(_10772_),
    .Y(_10773_),
    .A1(_10727_),
    .A2(_10770_));
 sg13g2_xor2_1 _17631_ (.B(_09273_),
    .A(_09276_),
    .X(_10774_));
 sg13g2_and2_1 _17632_ (.A(_09283_),
    .B(_10774_),
    .X(_10775_));
 sg13g2_buf_2 _17633_ (.A(_10775_),
    .X(_10776_));
 sg13g2_buf_1 _17634_ (.A(_00194_),
    .X(_10777_));
 sg13g2_buf_1 _17635_ (.A(_00284_),
    .X(_10778_));
 sg13g2_buf_8 _17636_ (.A(net629),
    .X(_10779_));
 sg13g2_and2_1 _17637_ (.A(net689),
    .B(net683),
    .X(_10780_));
 sg13g2_or2_1 _17638_ (.X(_10781_),
    .B(net902),
    .A(net904));
 sg13g2_buf_1 _17639_ (.A(_10781_),
    .X(_10782_));
 sg13g2_nor2_1 _17640_ (.A(net689),
    .B(_10782_),
    .Y(_10783_));
 sg13g2_a22oi_1 _17641_ (.Y(_10784_),
    .B1(_10783_),
    .B2(\cpu.ex.r_12[13] ),
    .A2(_10780_),
    .A1(\cpu.ex.r_11[13] ));
 sg13g2_buf_1 _17642_ (.A(_10664_),
    .X(_10785_));
 sg13g2_mux2_1 _17643_ (.A0(\cpu.ex.r_10[13] ),
    .A1(\cpu.ex.r_14[13] ),
    .S(net684),
    .X(_10786_));
 sg13g2_a22oi_1 _17644_ (.Y(_10787_),
    .B1(_10786_),
    .B2(_10761_),
    .A2(net774),
    .A1(\cpu.ex.r_stmp[13] ));
 sg13g2_nand2b_1 _17645_ (.Y(_10788_),
    .B(net783),
    .A_N(_10787_));
 sg13g2_o21ai_1 _17646_ (.B1(_10788_),
    .Y(_10789_),
    .A1(_10737_),
    .A2(_10784_));
 sg13g2_a221oi_1 _17647_ (.B2(\cpu.ex.r_epc[13] ),
    .C1(net681),
    .B1(_10707_),
    .A1(\cpu.ex.r_9[13] ),
    .Y(_10790_),
    .A2(net688));
 sg13g2_buf_1 _17648_ (.A(\cpu.ex.r_sp[13] ),
    .X(_10791_));
 sg13g2_a221oi_1 _17649_ (.B2(_10791_),
    .C1(net686),
    .B1(_10707_),
    .A1(\cpu.ex.r_8[13] ),
    .Y(_10792_),
    .A2(net688));
 sg13g2_nor3_1 _17650_ (.A(net684),
    .B(_10790_),
    .C(_10792_),
    .Y(_10793_));
 sg13g2_nor2_2 _17651_ (.A(_10666_),
    .B(net1039),
    .Y(_10794_));
 sg13g2_buf_1 _17652_ (.A(\cpu.ex.r_mult[29] ),
    .X(_10795_));
 sg13g2_a22oi_1 _17653_ (.Y(_10796_),
    .B1(_10688_),
    .B2(_10795_),
    .A2(_10794_),
    .A1(\cpu.ex.r_lr[13] ));
 sg13g2_or2_1 _17654_ (.X(_10797_),
    .B(_10796_),
    .A(net682));
 sg13g2_buf_1 _17655_ (.A(\cpu.ex.mmu_read[13] ),
    .X(_10798_));
 sg13g2_inv_2 _17656_ (.Y(_10799_),
    .A(net1124));
 sg13g2_nand2_1 _17657_ (.Y(_10800_),
    .A(net682),
    .B(\cpu.ex.r_13[13] ));
 sg13g2_o21ai_1 _17658_ (.B1(_10800_),
    .Y(_10801_),
    .A1(net682),
    .A2(_10799_));
 sg13g2_nand2b_1 _17659_ (.Y(_10802_),
    .B(net779),
    .A_N(_00263_));
 sg13g2_a21oi_1 _17660_ (.A1(net776),
    .A2(_10802_),
    .Y(_10803_),
    .B1(net689));
 sg13g2_o21ai_1 _17661_ (.B1(_10803_),
    .Y(_10804_),
    .A1(net776),
    .A2(_10801_));
 sg13g2_a21oi_1 _17662_ (.A1(_10797_),
    .A2(_10804_),
    .Y(_10805_),
    .B1(net681));
 sg13g2_or4_1 _17663_ (.A(net558),
    .B(_10789_),
    .C(_10793_),
    .D(_10805_),
    .X(_10806_));
 sg13g2_buf_1 _17664_ (.A(net701),
    .X(_10807_));
 sg13g2_nand2b_1 _17665_ (.Y(_10808_),
    .B(net558),
    .A_N(net628));
 sg13g2_nand2_1 _17666_ (.Y(_10809_),
    .A(_10806_),
    .B(_10808_));
 sg13g2_buf_1 _17667_ (.A(net702),
    .X(_10810_));
 sg13g2_inv_1 _17668_ (.Y(_10811_),
    .A(net902));
 sg13g2_buf_1 _17669_ (.A(\cpu.ex.r_mult[28] ),
    .X(_10812_));
 sg13g2_and2_1 _17670_ (.A(net1041),
    .B(net1128),
    .X(_10813_));
 sg13g2_buf_2 _17671_ (.A(_10813_),
    .X(_10814_));
 sg13g2_a221oi_1 _17672_ (.B2(\cpu.ex.r_sp[12] ),
    .C1(net682),
    .B1(_10693_),
    .A1(_10812_),
    .Y(_10815_),
    .A2(_10814_));
 sg13g2_inv_1 _17673_ (.Y(_10816_),
    .A(_00262_));
 sg13g2_a221oi_1 _17674_ (.B2(\cpu.ex.r_10[12] ),
    .C1(net685),
    .B1(_10693_),
    .A1(_10816_),
    .Y(_10817_),
    .A2(_10814_));
 sg13g2_or3_1 _17675_ (.A(_10811_),
    .B(_10815_),
    .C(_10817_),
    .X(_10818_));
 sg13g2_mux2_1 _17676_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_9[12] ),
    .S(net686),
    .X(_10819_));
 sg13g2_nor2b_1 _17677_ (.A(net686),
    .B_N(\cpu.ex.r_14[12] ),
    .Y(_10820_));
 sg13g2_a22oi_1 _17678_ (.Y(_10821_),
    .B1(_10820_),
    .B2(_10688_),
    .A2(_10819_),
    .A1(_10794_));
 sg13g2_nand2_1 _17679_ (.Y(_10822_),
    .A(\cpu.ex.r_12[12] ),
    .B(_10783_));
 sg13g2_a21o_1 _17680_ (.A2(_10822_),
    .A1(_10821_),
    .B1(net685),
    .X(_10823_));
 sg13g2_inv_1 _17681_ (.Y(_10824_),
    .A(\cpu.ex.r_epc[12] ));
 sg13g2_nand2_1 _17682_ (.Y(_10825_),
    .A(net682),
    .B(\cpu.ex.r_11[12] ));
 sg13g2_o21ai_1 _17683_ (.B1(_10825_),
    .Y(_10826_),
    .A1(net682),
    .A2(_10824_));
 sg13g2_and2_1 _17684_ (.A(_10649_),
    .B(_10664_),
    .X(_10827_));
 sg13g2_nor2_1 _17685_ (.A(_10640_),
    .B(net1039),
    .Y(_10828_));
 sg13g2_buf_1 _17686_ (.A(_10828_),
    .X(_10829_));
 sg13g2_a22oi_1 _17687_ (.Y(_10830_),
    .B1(_10747_),
    .B2(\cpu.ex.r_13[12] ),
    .A2(net773),
    .A1(\cpu.ex.r_lr[12] ));
 sg13g2_buf_1 _17688_ (.A(\cpu.ex.mmu_read[12] ),
    .X(_10831_));
 sg13g2_nand2_1 _17689_ (.Y(_10832_),
    .A(_10831_),
    .B(net774));
 sg13g2_a21oi_1 _17690_ (.A1(_10830_),
    .A2(_10832_),
    .Y(_10833_),
    .B1(_10742_));
 sg13g2_a221oi_1 _17691_ (.B2(\cpu.ex.r_stmp[12] ),
    .C1(_10833_),
    .B1(_10827_),
    .A1(_10780_),
    .Y(_10834_),
    .A2(_10826_));
 sg13g2_nand4_1 _17692_ (.B(_10818_),
    .C(_10823_),
    .A(net559),
    .Y(_10835_),
    .D(_10834_));
 sg13g2_o21ai_1 _17693_ (.B1(_10835_),
    .Y(_10836_),
    .A1(net627),
    .A2(net559));
 sg13g2_nand2_1 _17694_ (.Y(_10837_),
    .A(net1127),
    .B(_10625_));
 sg13g2_buf_2 _17695_ (.A(_10837_),
    .X(_10838_));
 sg13g2_mux4_1 _17696_ (.S0(_09286_),
    .A0(_10777_),
    .A1(_10778_),
    .A2(_10809_),
    .A3(_10836_),
    .S1(_10838_),
    .X(_10839_));
 sg13g2_a22oi_1 _17697_ (.Y(_10840_),
    .B1(_10776_),
    .B2(_10839_),
    .A2(_10773_),
    .A1(_10723_));
 sg13g2_buf_1 _17698_ (.A(_10840_),
    .X(_10841_));
 sg13g2_nand2b_1 _17699_ (.Y(_10842_),
    .B(_10639_),
    .A_N(net1135));
 sg13g2_a22oi_1 _17700_ (.Y(_10843_),
    .B1(_10752_),
    .B2(\cpu.ex.r_11[11] ),
    .A2(_10678_),
    .A1(\cpu.ex.r_8[11] ));
 sg13g2_nor2b_1 _17701_ (.A(net1128),
    .B_N(net1129),
    .Y(_10844_));
 sg13g2_buf_2 _17702_ (.A(_10844_),
    .X(_10845_));
 sg13g2_nor2b_1 _17703_ (.A(_10843_),
    .B_N(_10845_),
    .Y(_10846_));
 sg13g2_mux2_1 _17704_ (.A0(\cpu.ex.r_12[11] ),
    .A1(\cpu.ex.r_13[11] ),
    .S(net1041),
    .X(_10847_));
 sg13g2_nand3_1 _17705_ (.B(_10691_),
    .C(_10847_),
    .A(net903),
    .Y(_10848_));
 sg13g2_mux2_1 _17706_ (.A0(\cpu.ex.r_lr[11] ),
    .A1(\cpu.ex.r_9[11] ),
    .S(net1042),
    .X(_10849_));
 sg13g2_nand3_1 _17707_ (.B(net909),
    .C(_10849_),
    .A(_10653_),
    .Y(_10850_));
 sg13g2_nor2b_1 _17708_ (.A(_00261_),
    .B_N(net1041),
    .Y(_10851_));
 sg13g2_nor2b_1 _17709_ (.A(_10672_),
    .B_N(\cpu.ex.r_14[11] ),
    .Y(_10852_));
 sg13g2_and3_1 _17710_ (.X(_10853_),
    .A(net1040),
    .B(net1129),
    .C(net1128));
 sg13g2_buf_1 _17711_ (.A(_10853_),
    .X(_10854_));
 sg13g2_o21ai_1 _17712_ (.B1(_10854_),
    .Y(_10855_),
    .A1(_10851_),
    .A2(_10852_));
 sg13g2_nand3_1 _17713_ (.B(net783),
    .C(_10664_),
    .A(\cpu.ex.r_stmp[11] ),
    .Y(_10856_));
 sg13g2_nand4_1 _17714_ (.B(_10850_),
    .C(_10855_),
    .A(_10848_),
    .Y(_10857_),
    .D(_10856_));
 sg13g2_nor2b_1 _17715_ (.A(net1039),
    .B_N(\cpu.ex.r_10[11] ),
    .Y(_10858_));
 sg13g2_nand2_1 _17716_ (.Y(_10859_),
    .A(_10658_),
    .B(_10858_));
 sg13g2_a22oi_1 _17717_ (.Y(_10860_),
    .B1(_10693_),
    .B2(_10347_),
    .A2(_10814_),
    .A1(net1134));
 sg13g2_a22oi_1 _17718_ (.Y(_10861_),
    .B1(_10858_),
    .B2(_10658_),
    .A2(_10709_),
    .A1(\cpu.ex.r_epc[11] ));
 sg13g2_a221oi_1 _17719_ (.B2(_10861_),
    .C1(_10811_),
    .B1(_10860_),
    .A1(net784),
    .Y(_10862_),
    .A2(_10859_));
 sg13g2_or4_1 _17720_ (.A(net629),
    .B(_10846_),
    .C(_10857_),
    .D(_10862_),
    .X(_10863_));
 sg13g2_and4_1 _17721_ (.A(_08299_),
    .B(_10621_),
    .C(_10842_),
    .D(_10863_),
    .X(_10864_));
 sg13g2_nand3_1 _17722_ (.B(net438),
    .C(_10864_),
    .A(net439),
    .Y(_10865_));
 sg13g2_nor2_1 _17723_ (.A(_10627_),
    .B(_10319_),
    .Y(_10866_));
 sg13g2_o21ai_1 _17724_ (.B1(_10866_),
    .Y(_10867_),
    .A1(_08359_),
    .A2(_08415_));
 sg13g2_and2_1 _17725_ (.A(_10842_),
    .B(_10863_),
    .X(_10868_));
 sg13g2_nor2b_1 _17726_ (.A(net498),
    .B_N(_10866_),
    .Y(_10869_));
 sg13g2_a221oi_1 _17727_ (.B2(_10631_),
    .C1(_10869_),
    .B1(_10866_),
    .A1(_10627_),
    .Y(_10870_),
    .A2(_10868_));
 sg13g2_nand3_1 _17728_ (.B(_10867_),
    .C(_10870_),
    .A(_10865_),
    .Y(_10871_));
 sg13g2_buf_2 _17729_ (.A(_10871_),
    .X(_10872_));
 sg13g2_and2_1 _17730_ (.A(_09274_),
    .B(_10720_),
    .X(_10873_));
 sg13g2_nor2_1 _17731_ (.A(_09274_),
    .B(_10720_),
    .Y(_10874_));
 sg13g2_a21o_1 _17732_ (.A2(_10873_),
    .A1(_10872_),
    .B1(_10874_),
    .X(_10875_));
 sg13g2_inv_1 _17733_ (.Y(_10876_),
    .A(_10234_));
 sg13g2_and2_1 _17734_ (.A(net903),
    .B(\cpu.ex.r_stmp[9] ),
    .X(_10877_));
 sg13g2_nor2b_1 _17735_ (.A(net903),
    .B_N(\cpu.ex.r_8[9] ),
    .Y(_10878_));
 sg13g2_a22oi_1 _17736_ (.Y(_10879_),
    .B1(_10878_),
    .B2(_10691_),
    .A2(_10877_),
    .A1(_10707_));
 sg13g2_nand2b_1 _17737_ (.Y(_10880_),
    .B(_10854_),
    .A_N(_00259_));
 sg13g2_nor3_1 _17738_ (.A(_10696_),
    .B(net1042),
    .C(net903),
    .Y(_10881_));
 sg13g2_a21oi_1 _17739_ (.A1(\cpu.ex.r_lr[9] ),
    .A2(_10881_),
    .Y(_10882_),
    .B1(_10764_));
 sg13g2_a22oi_1 _17740_ (.Y(_10883_),
    .B1(_10880_),
    .B2(_10882_),
    .A2(_10879_),
    .A1(_10765_));
 sg13g2_mux4_1 _17741_ (.S0(net906),
    .A0(_10265_),
    .A1(\cpu.ex.r_epc[9] ),
    .A2(\cpu.ex.r_10[9] ),
    .A3(\cpu.ex.r_11[9] ),
    .S1(net908),
    .X(_10884_));
 sg13g2_and2_1 _17742_ (.A(_10740_),
    .B(_10884_),
    .X(_10885_));
 sg13g2_nand3_1 _17743_ (.B(_10650_),
    .C(_10747_),
    .A(\cpu.ex.r_14[9] ),
    .Y(_10886_));
 sg13g2_mux2_1 _17744_ (.A0(\cpu.ex.r_12[9] ),
    .A1(\cpu.ex.r_13[9] ),
    .S(net904),
    .X(_10887_));
 sg13g2_nand3_1 _17745_ (.B(_10691_),
    .C(_10887_),
    .A(_10757_),
    .Y(_10888_));
 sg13g2_nand3_1 _17746_ (.B(net774),
    .C(_10752_),
    .A(_10131_),
    .Y(_10889_));
 sg13g2_nand3_1 _17747_ (.B(net909),
    .C(_10845_),
    .A(\cpu.ex.r_9[9] ),
    .Y(_10890_));
 sg13g2_nand4_1 _17748_ (.B(_10888_),
    .C(_10889_),
    .A(_10886_),
    .Y(_10891_),
    .D(_10890_));
 sg13g2_nor4_1 _17749_ (.A(net629),
    .B(_10883_),
    .C(_10885_),
    .D(_10891_),
    .Y(_10892_));
 sg13g2_a21oi_1 _17750_ (.A1(_10876_),
    .A2(net558),
    .Y(_10893_),
    .B1(_10892_));
 sg13g2_nor2_1 _17751_ (.A(_10627_),
    .B(_00287_),
    .Y(_10894_));
 sg13g2_nor2b_1 _17752_ (.A(net498),
    .B_N(_10894_),
    .Y(_10895_));
 sg13g2_a221oi_1 _17753_ (.B2(net437),
    .C1(_10895_),
    .B1(_10894_),
    .A1(_10627_),
    .Y(_10896_),
    .A2(_10893_));
 sg13g2_o21ai_1 _17754_ (.B1(_10894_),
    .Y(_10897_),
    .A1(_08359_),
    .A2(_08415_));
 sg13g2_nand4_1 _17755_ (.B(_10608_),
    .C(_10623_),
    .A(_10606_),
    .Y(_10898_),
    .D(_10893_));
 sg13g2_and3_1 _17756_ (.X(_10899_),
    .A(_10896_),
    .B(_10897_),
    .C(_10898_));
 sg13g2_buf_2 _17757_ (.A(_10899_),
    .X(_10900_));
 sg13g2_inv_2 _17758_ (.Y(\cpu.ex.c_mult_off[1] ),
    .A(_10776_));
 sg13g2_nor2_1 _17759_ (.A(_09286_),
    .B(\cpu.ex.c_mult_off[1] ),
    .Y(_10901_));
 sg13g2_nor2_1 _17760_ (.A(\cpu.ex.c_mult_off[0] ),
    .B(\cpu.ex.c_mult_off[1] ),
    .Y(_10902_));
 sg13g2_nor2_1 _17761_ (.A(net910),
    .B(_00282_),
    .Y(_10903_));
 sg13g2_a22oi_1 _17762_ (.Y(_10904_),
    .B1(_10693_),
    .B2(\cpu.ex.r_8[8] ),
    .A2(_10814_),
    .A1(\cpu.ex.r_13[8] ));
 sg13g2_nand2b_1 _17763_ (.Y(_10905_),
    .B(_10705_),
    .A_N(_10904_));
 sg13g2_nand3_1 _17764_ (.B(net783),
    .C(_10845_),
    .A(\cpu.ex.r_10[8] ),
    .Y(_10906_));
 sg13g2_nand4_1 _17765_ (.B(_10654_),
    .C(\cpu.ex.r_lr[8] ),
    .A(net785),
    .Y(_10907_),
    .D(_10644_));
 sg13g2_and2_1 _17766_ (.A(_10649_),
    .B(_10747_),
    .X(_10908_));
 sg13g2_and4_1 _17767_ (.A(net908),
    .B(net907),
    .C(\cpu.ex.r_9[8] ),
    .D(net909),
    .X(_10909_));
 sg13g2_a221oi_1 _17768_ (.B2(\cpu.ex.r_14[8] ),
    .C1(_10909_),
    .B1(_10908_),
    .A1(\cpu.ex.r_stmp[8] ),
    .Y(_10910_),
    .A2(_10827_));
 sg13g2_nand4_1 _17769_ (.B(_10906_),
    .C(_10907_),
    .A(_10905_),
    .Y(_10911_),
    .D(_10910_));
 sg13g2_mux2_1 _17770_ (.A0(\cpu.ex.r_epc[8] ),
    .A1(net1137),
    .S(net903),
    .X(_10912_));
 sg13g2_nand3_1 _17771_ (.B(_10753_),
    .C(_10912_),
    .A(net785),
    .Y(_10913_));
 sg13g2_mux2_1 _17772_ (.A0(_10286_),
    .A1(\cpu.ex.r_11[8] ),
    .S(net907),
    .X(_10914_));
 sg13g2_nand3_1 _17773_ (.B(_10753_),
    .C(_10914_),
    .A(net779),
    .Y(_10915_));
 sg13g2_and4_1 _17774_ (.A(_10764_),
    .B(net907),
    .C(_10301_),
    .D(_10707_),
    .X(_10916_));
 sg13g2_nand4_1 _17775_ (.B(net780),
    .C(\cpu.ex.r_12[8] ),
    .A(_10764_),
    .Y(_10917_),
    .D(_10691_));
 sg13g2_nor2b_1 _17776_ (.A(_10916_),
    .B_N(_10917_),
    .Y(_10918_));
 sg13g2_nand4_1 _17777_ (.B(_10913_),
    .C(_10915_),
    .A(_10713_),
    .Y(_10919_),
    .D(_10918_));
 sg13g2_inv_2 _17778_ (.Y(_10920_),
    .A(_09165_));
 sg13g2_nand2_1 _17779_ (.Y(_10921_),
    .A(_10920_),
    .B(net629));
 sg13g2_o21ai_1 _17780_ (.B1(_10921_),
    .Y(_10922_),
    .A1(_10911_),
    .A2(_10919_));
 sg13g2_buf_1 _17781_ (.A(_10922_),
    .X(_10923_));
 sg13g2_nor3_1 _17782_ (.A(_09108_),
    .B(net437),
    .C(_10923_),
    .Y(_10924_));
 sg13g2_nor2_1 _17783_ (.A(net1127),
    .B(_10923_),
    .Y(_10925_));
 sg13g2_a221oi_1 _17784_ (.B2(net358),
    .C1(_10925_),
    .B1(_10924_),
    .A1(_10625_),
    .Y(_10926_),
    .A2(_10903_));
 sg13g2_buf_2 _17785_ (.A(_10926_),
    .X(_10927_));
 sg13g2_a22oi_1 _17786_ (.Y(_10928_),
    .B1(_10902_),
    .B2(_10927_),
    .A2(_10901_),
    .A1(_10900_));
 sg13g2_nand3b_1 _17787_ (.B(net301),
    .C(net1038),
    .Y(_10929_),
    .A_N(_10136_));
 sg13g2_a22oi_1 _17788_ (.Y(_10930_),
    .B1(_10684_),
    .B2(\cpu.ex.r_11[10] ),
    .A2(_10682_),
    .A1(_10211_));
 sg13g2_nand2b_1 _17789_ (.Y(_10931_),
    .B(_10740_),
    .A_N(_10930_));
 sg13g2_nand3_1 _17790_ (.B(\cpu.ex.r_10[10] ),
    .C(net783),
    .A(_10761_),
    .Y(_10932_));
 sg13g2_nand3_1 _17791_ (.B(\cpu.ex.r_lr[10] ),
    .C(net909),
    .A(net685),
    .Y(_10933_));
 sg13g2_a21oi_1 _17792_ (.A1(_10932_),
    .A2(_10933_),
    .Y(_10934_),
    .B1(_10744_));
 sg13g2_nand2b_1 _17793_ (.Y(_10935_),
    .B(net775),
    .A_N(net906));
 sg13g2_mux2_1 _17794_ (.A0(\cpu.ex.r_stmp[10] ),
    .A1(\cpu.ex.r_14[10] ),
    .S(net779),
    .X(_10936_));
 sg13g2_a22oi_1 _17795_ (.Y(_10937_),
    .B1(_10936_),
    .B2(net776),
    .A2(net688),
    .A1(\cpu.ex.r_12[10] ));
 sg13g2_nor2_1 _17796_ (.A(_10935_),
    .B(_10937_),
    .Y(_10938_));
 sg13g2_nor2_1 _17797_ (.A(_10934_),
    .B(_10938_),
    .Y(_10939_));
 sg13g2_nand2_1 _17798_ (.Y(_10940_),
    .A(_10811_),
    .B(_10680_));
 sg13g2_a22oi_1 _17799_ (.Y(_10941_),
    .B1(_10693_),
    .B2(\cpu.ex.r_8[10] ),
    .A2(_10814_),
    .A1(\cpu.ex.r_13[10] ));
 sg13g2_nor2_1 _17800_ (.A(_10940_),
    .B(_10941_),
    .Y(_10942_));
 sg13g2_a22oi_1 _17801_ (.Y(_10943_),
    .B1(_10747_),
    .B2(_10203_),
    .A2(net773),
    .A1(\cpu.ex.r_epc[10] ));
 sg13g2_nor2b_1 _17802_ (.A(_10943_),
    .B_N(net683),
    .Y(_10944_));
 sg13g2_nand3_1 _17803_ (.B(_10215_),
    .C(_10785_),
    .A(_10756_),
    .Y(_10945_));
 sg13g2_nand3_1 _17804_ (.B(\cpu.ex.r_9[10] ),
    .C(net688),
    .A(_10655_),
    .Y(_10946_));
 sg13g2_a21oi_1 _17805_ (.A1(_10945_),
    .A2(_10946_),
    .Y(_10947_),
    .B1(net681));
 sg13g2_nor3_1 _17806_ (.A(_10942_),
    .B(_10944_),
    .C(_10947_),
    .Y(_10948_));
 sg13g2_nand4_1 _17807_ (.B(_10931_),
    .C(_10939_),
    .A(_10731_),
    .Y(_10949_),
    .D(_10948_));
 sg13g2_o21ai_1 _17808_ (.B1(_10949_),
    .Y(_10950_),
    .A1(net1143),
    .A2(net559));
 sg13g2_a21o_1 _17809_ (.A2(net301),
    .A1(_10728_),
    .B1(_10950_),
    .X(_10951_));
 sg13g2_nand3_1 _17810_ (.B(_10929_),
    .C(_10951_),
    .A(_10719_),
    .Y(_10952_));
 sg13g2_and2_1 _17811_ (.A(_09278_),
    .B(net814),
    .X(_10953_));
 sg13g2_buf_1 _17812_ (.A(_10953_),
    .X(_10954_));
 sg13g2_xor2_1 _17813_ (.B(_10771_),
    .A(_09275_),
    .X(_10955_));
 sg13g2_nor3_1 _17814_ (.A(_09290_),
    .B(net626),
    .C(_10955_),
    .Y(_10956_));
 sg13g2_and4_1 _17815_ (.A(_10875_),
    .B(_10928_),
    .C(_10952_),
    .D(_10956_),
    .X(_10957_));
 sg13g2_buf_1 _17816_ (.A(_10957_),
    .X(_10958_));
 sg13g2_nor2_1 _17817_ (.A(net782),
    .B(_10742_),
    .Y(_10959_));
 sg13g2_nand2b_1 _17818_ (.Y(_10960_),
    .B(_10696_),
    .A_N(net904));
 sg13g2_nor2_1 _17819_ (.A(net780),
    .B(_10960_),
    .Y(_10961_));
 sg13g2_a221oi_1 _17820_ (.B2(_10529_),
    .C1(net682),
    .B1(_10961_),
    .A1(_10533_),
    .Y(_10962_),
    .A2(_10959_));
 sg13g2_a221oi_1 _17821_ (.B2(\cpu.ex.r_10[2] ),
    .C1(net685),
    .B1(_10961_),
    .A1(\cpu.ex.r_13[2] ),
    .Y(_10963_),
    .A2(_10959_));
 sg13g2_nor2_1 _17822_ (.A(net681),
    .B(_10701_),
    .Y(_10964_));
 sg13g2_mux2_1 _17823_ (.A0(\cpu.ex.r_lr[2] ),
    .A1(\cpu.ex.r_epc[2] ),
    .S(net776),
    .X(_10965_));
 sg13g2_nand3_1 _17824_ (.B(net781),
    .C(_10540_),
    .A(_10732_),
    .Y(_10966_));
 sg13g2_o21ai_1 _17825_ (.B1(_10966_),
    .Y(_10967_),
    .A1(_08437_),
    .A2(_10782_));
 sg13g2_a22oi_1 _17826_ (.Y(_10968_),
    .B1(_10967_),
    .B2(net774),
    .A2(_10965_),
    .A1(_10964_));
 sg13g2_o21ai_1 _17827_ (.B1(_10968_),
    .Y(_10969_),
    .A1(_10962_),
    .A2(_10963_));
 sg13g2_nand3_1 _17828_ (.B(\cpu.ex.r_8[2] ),
    .C(net688),
    .A(net689),
    .Y(_10970_));
 sg13g2_nand3_1 _17829_ (.B(\cpu.ex.r_stmp[2] ),
    .C(net774),
    .A(net776),
    .Y(_10971_));
 sg13g2_a21oi_1 _17830_ (.A1(_10970_),
    .A2(_10971_),
    .Y(_10972_),
    .B1(net686));
 sg13g2_nand2_1 _17831_ (.Y(_10973_),
    .A(net777),
    .B(net779));
 sg13g2_inv_1 _17832_ (.Y(_10974_),
    .A(_00252_));
 sg13g2_a22oi_1 _17833_ (.Y(_10975_),
    .B1(_10688_),
    .B2(_10974_),
    .A2(_10794_),
    .A1(\cpu.ex.r_9[2] ));
 sg13g2_nor2_1 _17834_ (.A(_10973_),
    .B(_10975_),
    .Y(_10976_));
 sg13g2_nand3_1 _17835_ (.B(\cpu.ex.r_11[2] ),
    .C(net683),
    .A(net689),
    .Y(_10977_));
 sg13g2_mux2_1 _17836_ (.A0(\cpu.ex.r_12[2] ),
    .A1(\cpu.ex.r_14[2] ),
    .S(net905),
    .X(_10978_));
 sg13g2_nand2_1 _17837_ (.Y(_10979_),
    .A(_10758_),
    .B(_10978_));
 sg13g2_a21oi_1 _17838_ (.A1(_10977_),
    .A2(_10979_),
    .Y(_10980_),
    .B1(net685));
 sg13g2_or4_1 _17839_ (.A(net558),
    .B(_10972_),
    .C(_10976_),
    .D(_10980_),
    .X(_10981_));
 sg13g2_nand2_1 _17840_ (.Y(_10982_),
    .A(_09455_),
    .B(_10779_));
 sg13g2_o21ai_1 _17841_ (.B1(_10982_),
    .Y(_10983_),
    .A1(_10969_),
    .A2(_10981_));
 sg13g2_inv_2 _17842_ (.Y(_10984_),
    .A(net1162));
 sg13g2_nand2_1 _17843_ (.Y(_10985_),
    .A(_10984_),
    .B(net558));
 sg13g2_a22oi_1 _17844_ (.Y(_10986_),
    .B1(_10688_),
    .B2(\cpu.ex.r_15[0] ),
    .A2(_10794_),
    .A1(\cpu.ex.r_9[0] ));
 sg13g2_and2_1 _17845_ (.A(net905),
    .B(net1042),
    .X(_10987_));
 sg13g2_buf_1 _17846_ (.A(_10987_),
    .X(_10988_));
 sg13g2_mux2_1 _17847_ (.A0(\cpu.ex.r_10[0] ),
    .A1(\cpu.ex.r_11[0] ),
    .S(net906),
    .X(_10989_));
 sg13g2_nand3_1 _17848_ (.B(_10988_),
    .C(_10989_),
    .A(net689),
    .Y(_10990_));
 sg13g2_o21ai_1 _17849_ (.B1(_10990_),
    .Y(_10991_),
    .A1(_10973_),
    .A2(_10986_));
 sg13g2_a22oi_1 _17850_ (.Y(_10992_),
    .B1(_10845_),
    .B2(\cpu.ex.r_8[0] ),
    .A2(net774),
    .A1(_09158_));
 sg13g2_nand3b_1 _17851_ (.B(net775),
    .C(\cpu.ex.r_stmp[0] ),
    .Y(_10993_),
    .A_N(net906));
 sg13g2_buf_1 _17852_ (.A(\cpu.ex.genblk3.r_prev_supmode ),
    .X(_10994_));
 sg13g2_nand3b_1 _17853_ (.B(net777),
    .C(_10994_),
    .Y(_10995_),
    .A_N(net780));
 sg13g2_nand2b_1 _17854_ (.Y(_10996_),
    .B(net781),
    .A_N(net908));
 sg13g2_a21o_1 _17855_ (.A2(_10995_),
    .A1(_10993_),
    .B1(_10996_),
    .X(_10997_));
 sg13g2_o21ai_1 _17856_ (.B1(_10997_),
    .Y(_10998_),
    .A1(_10782_),
    .A2(_10992_));
 sg13g2_mux2_1 _17857_ (.A0(\cpu.ex.r_12[0] ),
    .A1(\cpu.ex.r_14[0] ),
    .S(net905),
    .X(_10999_));
 sg13g2_nand2_1 _17858_ (.Y(_11000_),
    .A(_10658_),
    .B(_10999_));
 sg13g2_and2_1 _17859_ (.A(net784),
    .B(\cpu.ex.r_13[0] ),
    .X(_11001_));
 sg13g2_nor2b_1 _17860_ (.A(net784),
    .B_N(_10561_),
    .Y(_11002_));
 sg13g2_a22oi_1 _17861_ (.Y(_11003_),
    .B1(_11002_),
    .B2(net683),
    .A2(_11001_),
    .A1(net909));
 sg13g2_a21oi_1 _17862_ (.A1(_11000_),
    .A2(_11003_),
    .Y(_11004_),
    .B1(net689));
 sg13g2_or4_1 _17863_ (.A(net558),
    .B(_10991_),
    .C(_10998_),
    .D(_11004_),
    .X(_11005_));
 sg13g2_buf_1 _17864_ (.A(_11005_),
    .X(_11006_));
 sg13g2_nand3_1 _17865_ (.B(_10985_),
    .C(_11006_),
    .A(_10776_),
    .Y(_11007_));
 sg13g2_o21ai_1 _17866_ (.B1(_11007_),
    .Y(_11008_),
    .A1(_10776_),
    .A2(_10983_));
 sg13g2_o21ai_1 _17867_ (.B1(_11008_),
    .Y(_11009_),
    .A1(net778),
    .A2(_10726_));
 sg13g2_or4_1 _17868_ (.A(net910),
    .B(_00283_),
    .C(_10726_),
    .D(_10776_),
    .X(_11010_));
 sg13g2_inv_1 _17869_ (.Y(_11011_),
    .A(_09110_));
 sg13g2_and3_1 _17870_ (.X(_11012_),
    .A(_11011_),
    .B(net498),
    .C(_09160_));
 sg13g2_nand3_1 _17871_ (.B(_10608_),
    .C(_11012_),
    .A(_10606_),
    .Y(_11013_));
 sg13g2_buf_1 _17872_ (.A(_11013_),
    .X(_11014_));
 sg13g2_nor2_1 _17873_ (.A(_08265_),
    .B(net910),
    .Y(_11015_));
 sg13g2_nand3_1 _17874_ (.B(_11014_),
    .C(_11015_),
    .A(_10776_),
    .Y(_11016_));
 sg13g2_nand4_1 _17875_ (.B(_11009_),
    .C(_11010_),
    .A(_09286_),
    .Y(_11017_),
    .D(_11016_));
 sg13g2_nand2_1 _17876_ (.Y(\cpu.ex.c_mult_off[3] ),
    .A(net646),
    .B(_10955_));
 sg13g2_or2_1 _17877_ (.X(_11018_),
    .B(_10873_),
    .A(_10874_));
 sg13g2_nand2_1 _17878_ (.Y(\cpu.ex.c_mult_off[2] ),
    .A(_09284_),
    .B(_11018_));
 sg13g2_nand3b_1 _17879_ (.B(_10752_),
    .C(net784),
    .Y(_11019_),
    .A_N(_00251_));
 sg13g2_nand3_1 _17880_ (.B(_10580_),
    .C(_10678_),
    .A(net785),
    .Y(_11020_));
 sg13g2_a21oi_1 _17881_ (.A1(_11019_),
    .A2(_11020_),
    .Y(_11021_),
    .B1(net689));
 sg13g2_a22oi_1 _17882_ (.Y(_11022_),
    .B1(net683),
    .B2(\cpu.ex.r_11[1] ),
    .A2(_10678_),
    .A1(\cpu.ex.r_8[1] ));
 sg13g2_nor2b_1 _17883_ (.A(_11022_),
    .B_N(_10845_),
    .Y(_11023_));
 sg13g2_a22oi_1 _17884_ (.Y(_11024_),
    .B1(_10845_),
    .B2(\cpu.ex.r_10[1] ),
    .A2(_10785_),
    .A1(\cpu.ex.r_stmp[1] ));
 sg13g2_nand3b_1 _17885_ (.B(net908),
    .C(\cpu.ex.r_14[1] ),
    .Y(_11025_),
    .A_N(net906));
 sg13g2_nand3b_1 _17886_ (.B(_10556_),
    .C(net906),
    .Y(_11026_),
    .A_N(net908));
 sg13g2_nand2_1 _17887_ (.Y(_11027_),
    .A(net905),
    .B(net780));
 sg13g2_a21o_1 _17888_ (.A2(_11026_),
    .A1(_11025_),
    .B1(_11027_),
    .X(_11028_));
 sg13g2_o21ai_1 _17889_ (.B1(_11028_),
    .Y(_11029_),
    .A1(_10960_),
    .A2(_11024_));
 sg13g2_mux2_1 _17890_ (.A0(\cpu.ex.r_9[1] ),
    .A1(\cpu.ex.r_13[1] ),
    .S(net903),
    .X(_11030_));
 sg13g2_nand3_1 _17891_ (.B(net909),
    .C(_11030_),
    .A(net784),
    .Y(_11031_));
 sg13g2_mux2_1 _17892_ (.A0(_10570_),
    .A1(\cpu.ex.r_epc[1] ),
    .S(net906),
    .X(_11032_));
 sg13g2_nand3_1 _17893_ (.B(_10707_),
    .C(_11032_),
    .A(net782),
    .Y(_11033_));
 sg13g2_mux2_1 _17894_ (.A0(\cpu.ex.r_lr[1] ),
    .A1(\cpu.ex.mmu_read[1] ),
    .S(net903),
    .X(_11034_));
 sg13g2_nand3_1 _17895_ (.B(net909),
    .C(_11034_),
    .A(_10642_),
    .Y(_11035_));
 sg13g2_nand3_1 _17896_ (.B(_10678_),
    .C(_10747_),
    .A(\cpu.ex.r_12[1] ),
    .Y(_11036_));
 sg13g2_nand4_1 _17897_ (.B(_11033_),
    .C(_11035_),
    .A(_11031_),
    .Y(_11037_),
    .D(_11036_));
 sg13g2_nor4_1 _17898_ (.A(_11021_),
    .B(_11023_),
    .C(_11029_),
    .D(_11037_),
    .Y(_11038_));
 sg13g2_nor2_1 _17899_ (.A(_09177_),
    .B(_10713_),
    .Y(_11039_));
 sg13g2_a21oi_2 _17900_ (.B1(_11039_),
    .Y(_11040_),
    .A2(_11038_),
    .A1(_10713_));
 sg13g2_and2_1 _17901_ (.A(net777),
    .B(\cpu.ex.r_epc[3] ),
    .X(_11041_));
 sg13g2_a21oi_1 _17902_ (.A1(net681),
    .A2(\cpu.ex.r_sp[3] ),
    .Y(_11042_),
    .B1(_11041_));
 sg13g2_nor3_1 _17903_ (.A(net684),
    .B(_10996_),
    .C(_11042_),
    .Y(_11043_));
 sg13g2_nor2b_1 _17904_ (.A(net775),
    .B_N(\cpu.ex.r_8[3] ),
    .Y(_11044_));
 sg13g2_nor2b_1 _17905_ (.A(net781),
    .B_N(net1165),
    .Y(_11045_));
 sg13g2_a22oi_1 _17906_ (.Y(_11046_),
    .B1(_11045_),
    .B2(net774),
    .A2(_11044_),
    .A1(_10705_));
 sg13g2_nor2b_1 _17907_ (.A(net775),
    .B_N(\cpu.ex.r_10[3] ),
    .Y(_11047_));
 sg13g2_and2_1 _17908_ (.A(net775),
    .B(\cpu.ex.r_stmp[3] ),
    .X(_11048_));
 sg13g2_a22oi_1 _17909_ (.Y(_11049_),
    .B1(_11048_),
    .B2(_10707_),
    .A2(_11047_),
    .A1(_10988_));
 sg13g2_a21oi_1 _17910_ (.A1(_11046_),
    .A2(_11049_),
    .Y(_11050_),
    .B1(net686));
 sg13g2_nor2b_1 _17911_ (.A(net781),
    .B_N(\cpu.ex.r_13[3] ),
    .Y(_11051_));
 sg13g2_nor2b_1 _17912_ (.A(_00253_),
    .B_N(net781),
    .Y(_11052_));
 sg13g2_o21ai_1 _17913_ (.B1(net684),
    .Y(_11053_),
    .A1(_11051_),
    .A2(_11052_));
 sg13g2_nand2_1 _17914_ (.Y(_11054_),
    .A(\cpu.ex.r_11[3] ),
    .B(_10740_));
 sg13g2_a21oi_1 _17915_ (.A1(_11053_),
    .A2(_11054_),
    .Y(_11055_),
    .B1(_10973_));
 sg13g2_nor3_1 _17916_ (.A(_11043_),
    .B(_11050_),
    .C(_11055_),
    .Y(_11056_));
 sg13g2_and3_1 _17917_ (.X(_11057_),
    .A(net779),
    .B(\cpu.ex.r_14[3] ),
    .C(net783));
 sg13g2_inv_2 _17918_ (.Y(_11058_),
    .A(\cpu.ex.mmu_read[3] ));
 sg13g2_nor3_1 _17919_ (.A(net779),
    .B(_11058_),
    .C(_10742_),
    .Y(_11059_));
 sg13g2_o21ai_1 _17920_ (.B1(net684),
    .Y(_11060_),
    .A1(_11057_),
    .A2(_11059_));
 sg13g2_nand3_1 _17921_ (.B(\cpu.ex.r_12[3] ),
    .C(_10658_),
    .A(net684),
    .Y(_11061_));
 sg13g2_nand3_1 _17922_ (.B(\cpu.ex.r_lr[3] ),
    .C(net773),
    .A(net777),
    .Y(_11062_));
 sg13g2_a21o_1 _17923_ (.A2(_11062_),
    .A1(_11061_),
    .B1(net776),
    .X(_11063_));
 sg13g2_and3_1 _17924_ (.X(_11064_),
    .A(net782),
    .B(\cpu.ex.r_9[3] ),
    .C(net688));
 sg13g2_inv_2 _17925_ (.Y(_11065_),
    .A(net1131));
 sg13g2_nor3_1 _17926_ (.A(net782),
    .B(_11065_),
    .C(_10996_),
    .Y(_11066_));
 sg13g2_o21ai_1 _17927_ (.B1(net686),
    .Y(_11067_),
    .A1(_11064_),
    .A2(_11066_));
 sg13g2_and4_1 _17928_ (.A(_10713_),
    .B(_11060_),
    .C(_11063_),
    .D(_11067_),
    .X(_11068_));
 sg13g2_nor2_1 _17929_ (.A(_09190_),
    .B(_10731_),
    .Y(_11069_));
 sg13g2_a21oi_1 _17930_ (.A1(_11056_),
    .A2(_11068_),
    .Y(_11070_),
    .B1(_11069_));
 sg13g2_mux2_1 _17931_ (.A0(_11040_),
    .A1(_11070_),
    .S(\cpu.ex.c_mult_off[1] ),
    .X(_11071_));
 sg13g2_a221oi_1 _17932_ (.B2(net1038),
    .C1(_11071_),
    .B1(net301),
    .A1(_09276_),
    .Y(_11072_),
    .A2(net646));
 sg13g2_buf_1 _17933_ (.A(_00189_),
    .X(_11073_));
 sg13g2_and2_1 _17934_ (.A(_10563_),
    .B(_10776_),
    .X(_11074_));
 sg13g2_a21oi_1 _17935_ (.A1(_11073_),
    .A2(\cpu.ex.c_mult_off[1] ),
    .Y(_11075_),
    .B1(_11074_));
 sg13g2_nor4_1 _17936_ (.A(net778),
    .B(_09286_),
    .C(_10726_),
    .D(_11075_),
    .Y(_11076_));
 sg13g2_nor4_1 _17937_ (.A(\cpu.ex.c_mult_off[3] ),
    .B(\cpu.ex.c_mult_off[2] ),
    .C(_11072_),
    .D(_11076_),
    .Y(_11077_));
 sg13g2_mux4_1 _17938_ (.S0(_09286_),
    .A0(_10411_),
    .A1(_00289_),
    .A2(_10507_),
    .A3(_08448_),
    .S1(_10776_),
    .X(_11078_));
 sg13g2_nand3b_1 _17939_ (.B(net1038),
    .C(net301),
    .Y(_11079_),
    .A_N(_11078_));
 sg13g2_inv_2 _17940_ (.Y(_11080_),
    .A(_09893_));
 sg13g2_a22oi_1 _17941_ (.Y(_11081_),
    .B1(_10747_),
    .B2(\cpu.ex.r_14[5] ),
    .A2(net773),
    .A1(_10484_));
 sg13g2_nor2_1 _17942_ (.A(_10960_),
    .B(_11081_),
    .Y(_11082_));
 sg13g2_a22oi_1 _17943_ (.Y(_11083_),
    .B1(_10693_),
    .B2(\cpu.ex.r_8[5] ),
    .A2(_10814_),
    .A1(\cpu.ex.r_13[5] ));
 sg13g2_nor2_1 _17944_ (.A(_10940_),
    .B(_11083_),
    .Y(_11084_));
 sg13g2_a22oi_1 _17945_ (.Y(_11085_),
    .B1(_10707_),
    .B2(\cpu.ex.r_stmp[5] ),
    .A2(_10691_),
    .A1(\cpu.ex.r_12[5] ));
 sg13g2_mux2_1 _17946_ (.A0(\cpu.ex.r_lr[5] ),
    .A1(\cpu.ex.r_epc[5] ),
    .S(net905),
    .X(_11086_));
 sg13g2_nand3_1 _17947_ (.B(_10829_),
    .C(_11086_),
    .A(net777),
    .Y(_11087_));
 sg13g2_o21ai_1 _17948_ (.B1(_11087_),
    .Y(_11088_),
    .A1(_10935_),
    .A2(_11085_));
 sg13g2_nor3_1 _17949_ (.A(_11082_),
    .B(_11084_),
    .C(_11088_),
    .Y(_11089_));
 sg13g2_nor2b_1 _17950_ (.A(_00255_),
    .B_N(_10676_),
    .Y(_11090_));
 sg13g2_a21oi_1 _17951_ (.A1(net782),
    .A2(\cpu.ex.r_11[5] ),
    .Y(_11091_),
    .B1(_11090_));
 sg13g2_nor2b_1 _17952_ (.A(_10757_),
    .B_N(\cpu.ex.r_10[5] ),
    .Y(_11092_));
 sg13g2_o21ai_1 _17953_ (.B1(_10988_),
    .Y(_11093_),
    .A1(net777),
    .A2(_11092_));
 sg13g2_a21oi_1 _17954_ (.A1(_10733_),
    .A2(_11091_),
    .Y(_11094_),
    .B1(_11093_));
 sg13g2_nand3_1 _17955_ (.B(net774),
    .C(net683),
    .A(\cpu.ex.r_mult[21] ),
    .Y(_11095_));
 sg13g2_nand4_1 _17956_ (.B(net782),
    .C(\cpu.ex.r_9[5] ),
    .A(_10732_),
    .Y(_11096_),
    .D(net688));
 sg13g2_nand2_1 _17957_ (.Y(_11097_),
    .A(_11095_),
    .B(_11096_));
 sg13g2_nor3_1 _17958_ (.A(net629),
    .B(_11094_),
    .C(_11097_),
    .Y(_11098_));
 sg13g2_a22oi_1 _17959_ (.Y(_11099_),
    .B1(_11089_),
    .B2(_11098_),
    .A2(_10779_),
    .A1(_11080_));
 sg13g2_buf_1 _17960_ (.A(_11099_),
    .X(_11100_));
 sg13g2_nand2_1 _17961_ (.Y(_11101_),
    .A(_09167_),
    .B(net629));
 sg13g2_nand3_1 _17962_ (.B(net783),
    .C(_10664_),
    .A(\cpu.ex.r_stmp[7] ),
    .Y(_11102_));
 sg13g2_nand3_1 _17963_ (.B(net773),
    .C(_10650_),
    .A(_10391_),
    .Y(_11103_));
 sg13g2_mux2_1 _17964_ (.A0(\cpu.ex.r_8[7] ),
    .A1(\cpu.ex.r_10[7] ),
    .S(net1040),
    .X(_11104_));
 sg13g2_nand3_1 _17965_ (.B(_10658_),
    .C(_11104_),
    .A(net907),
    .Y(_11105_));
 sg13g2_nand4_1 _17966_ (.B(net780),
    .C(_10402_),
    .A(net785),
    .Y(_11106_),
    .D(_10678_));
 sg13g2_nand4_1 _17967_ (.B(_11103_),
    .C(_11105_),
    .A(_11102_),
    .Y(_11107_),
    .D(_11106_));
 sg13g2_mux2_1 _17968_ (.A0(\cpu.ex.r_9[7] ),
    .A1(\cpu.ex.r_11[7] ),
    .S(net902),
    .X(_11108_));
 sg13g2_nand3_1 _17969_ (.B(_10684_),
    .C(_11108_),
    .A(_10654_),
    .Y(_11109_));
 sg13g2_nand3_1 _17970_ (.B(net773),
    .C(_10752_),
    .A(\cpu.ex.r_epc[7] ),
    .Y(_11110_));
 sg13g2_mux2_1 _17971_ (.A0(\cpu.ex.r_12[7] ),
    .A1(\cpu.ex.r_14[7] ),
    .S(net902),
    .X(_11111_));
 sg13g2_nand3_1 _17972_ (.B(_10658_),
    .C(_11111_),
    .A(net775),
    .Y(_11112_));
 sg13g2_nand3_1 _17973_ (.B(_11110_),
    .C(_11112_),
    .A(_11109_),
    .Y(_11113_));
 sg13g2_a22oi_1 _17974_ (.Y(_11114_),
    .B1(_10881_),
    .B2(\cpu.ex.r_lr[7] ),
    .A2(_10854_),
    .A1(_10398_));
 sg13g2_nand3b_1 _17975_ (.B(_10646_),
    .C(\cpu.ex.r_13[7] ),
    .Y(_11115_),
    .A_N(net902));
 sg13g2_nand3b_1 _17976_ (.B(_10312_),
    .C(_10667_),
    .Y(_11116_),
    .A_N(net1042));
 sg13g2_a21o_1 _17977_ (.A2(_11116_),
    .A1(_11115_),
    .B1(net907),
    .X(_11117_));
 sg13g2_a21oi_1 _17978_ (.A1(_11114_),
    .A2(_11117_),
    .Y(_11118_),
    .B1(net681));
 sg13g2_or4_1 _17979_ (.A(net629),
    .B(_11107_),
    .C(_11113_),
    .D(_11118_),
    .X(_11119_));
 sg13g2_and2_1 _17980_ (.A(_11101_),
    .B(_11119_),
    .X(_11120_));
 sg13g2_buf_1 _17981_ (.A(_11120_),
    .X(_11121_));
 sg13g2_a22oi_1 _17982_ (.Y(_11122_),
    .B1(_10845_),
    .B2(\cpu.ex.r_8[4] ),
    .A2(_10664_),
    .A1(_08274_));
 sg13g2_nor2_1 _17983_ (.A(_10782_),
    .B(_11122_),
    .Y(_11123_));
 sg13g2_a22oi_1 _17984_ (.Y(_11124_),
    .B1(_10688_),
    .B2(net1130),
    .A2(_10794_),
    .A1(\cpu.ex.r_lr[4] ));
 sg13g2_nor3_1 _17985_ (.A(net681),
    .B(_10647_),
    .C(_11124_),
    .Y(_11125_));
 sg13g2_nand3_1 _17986_ (.B(\cpu.ex.r_11[4] ),
    .C(_10684_),
    .A(net907),
    .Y(_11126_));
 sg13g2_nand3_1 _17987_ (.B(\cpu.ex.r_stmp[4] ),
    .C(_10664_),
    .A(_10764_),
    .Y(_11127_));
 sg13g2_a21oi_1 _17988_ (.A1(_11126_),
    .A2(_11127_),
    .Y(_11128_),
    .B1(_10811_));
 sg13g2_nand2_1 _17989_ (.Y(_11129_),
    .A(net785),
    .B(\cpu.ex.r_epc[4] ));
 sg13g2_nand3_1 _17990_ (.B(_10678_),
    .C(_10747_),
    .A(\cpu.ex.r_12[4] ),
    .Y(_11130_));
 sg13g2_o21ai_1 _17991_ (.B1(_11130_),
    .Y(_11131_),
    .A1(_10673_),
    .A2(_11129_));
 sg13g2_nor4_1 _17992_ (.A(_11123_),
    .B(_11125_),
    .C(_11128_),
    .D(_11131_),
    .Y(_11132_));
 sg13g2_nand2b_1 _17993_ (.Y(_11133_),
    .B(\cpu.ex.r_13[4] ),
    .A_N(_10667_));
 sg13g2_o21ai_1 _17994_ (.B1(_11133_),
    .Y(_11134_),
    .A1(_10811_),
    .A2(_00254_));
 sg13g2_nand3_1 _17995_ (.B(_10684_),
    .C(_11134_),
    .A(net775),
    .Y(_11135_));
 sg13g2_nand2_1 _17996_ (.Y(_11136_),
    .A(\cpu.ex.r_14[4] ),
    .B(_10908_));
 sg13g2_and2_1 _17997_ (.A(_10644_),
    .B(_10845_),
    .X(_11137_));
 sg13g2_mux2_1 _17998_ (.A0(_10457_),
    .A1(\cpu.ex.r_10[4] ),
    .S(_10646_),
    .X(_11138_));
 sg13g2_a22oi_1 _17999_ (.Y(_11139_),
    .B1(_10961_),
    .B2(_11138_),
    .A2(_11137_),
    .A1(\cpu.ex.r_9[4] ));
 sg13g2_and4_1 _18000_ (.A(_10713_),
    .B(_11135_),
    .C(_11136_),
    .D(_11139_),
    .X(_11140_));
 sg13g2_a22oi_1 _18001_ (.Y(_11141_),
    .B1(_11132_),
    .B2(_11140_),
    .A2(net558),
    .A1(_09454_));
 sg13g2_buf_1 _18002_ (.A(_11141_),
    .X(_11142_));
 sg13g2_inv_1 _18003_ (.Y(_11143_),
    .A(\cpu.ex.r_11[6] ));
 sg13g2_inv_1 _18004_ (.Y(_11144_),
    .A(\cpu.ex.r_epc[6] ));
 sg13g2_mux4_1 _18005_ (.S0(net907),
    .A0(_00256_),
    .A1(_11143_),
    .A2(_10377_),
    .A3(_11144_),
    .S1(net785),
    .X(_11145_));
 sg13g2_mux2_1 _18006_ (.A0(\cpu.ex.r_9[6] ),
    .A1(\cpu.ex.r_13[6] ),
    .S(net903),
    .X(_11146_));
 sg13g2_a221oi_1 _18007_ (.B2(net784),
    .C1(_10668_),
    .B1(_11146_),
    .A1(\cpu.ex.r_lr[6] ),
    .Y(_11147_),
    .A2(net773));
 sg13g2_a21o_1 _18008_ (.A2(_11145_),
    .A1(net776),
    .B1(_11147_),
    .X(_11148_));
 sg13g2_inv_1 _18009_ (.Y(_11149_),
    .A(\cpu.ex.r_sp[6] ));
 sg13g2_nand3_1 _18010_ (.B(net780),
    .C(\cpu.ex.r_14[6] ),
    .A(net784),
    .Y(_11150_));
 sg13g2_o21ai_1 _18011_ (.B1(_11150_),
    .Y(_11151_),
    .A1(_11149_),
    .A2(_10701_));
 sg13g2_mux2_1 _18012_ (.A0(\cpu.ex.r_8[6] ),
    .A1(\cpu.ex.r_10[6] ),
    .S(net781),
    .X(_11152_));
 sg13g2_and2_1 _18013_ (.A(net782),
    .B(_10658_),
    .X(_11153_));
 sg13g2_nand3b_1 _18014_ (.B(_10647_),
    .C(\cpu.ex.r_12[6] ),
    .Y(_11154_),
    .A_N(_10668_));
 sg13g2_nand3b_1 _18015_ (.B(\cpu.ex.r_stmp[6] ),
    .C(net781),
    .Y(_11155_),
    .A_N(net908));
 sg13g2_a21oi_1 _18016_ (.A1(_11154_),
    .A2(_11155_),
    .Y(_11156_),
    .B1(_10935_));
 sg13g2_a221oi_1 _18017_ (.B2(_11153_),
    .C1(_11156_),
    .B1(_11152_),
    .A1(net783),
    .Y(_11157_),
    .A2(_11151_));
 sg13g2_o21ai_1 _18018_ (.B1(_11157_),
    .Y(_11158_),
    .A1(_10765_),
    .A2(_11148_));
 sg13g2_mux2_1 _18019_ (.A0(_09164_),
    .A1(_11158_),
    .S(net559),
    .X(_11159_));
 sg13g2_mux4_1 _18020_ (.S0(\cpu.ex.c_mult_off[1] ),
    .A0(_11100_),
    .A1(_11121_),
    .A2(_11142_),
    .A3(_11159_),
    .S1(_09286_),
    .X(_11160_));
 sg13g2_o21ai_1 _18021_ (.B1(_11160_),
    .Y(_11161_),
    .A1(net778),
    .A2(_10726_));
 sg13g2_a221oi_1 _18022_ (.B2(_11161_),
    .C1(\cpu.ex.c_mult_off[3] ),
    .B1(_11079_),
    .A1(net646),
    .Y(_11162_),
    .A2(_11018_));
 sg13g2_a21o_1 _18023_ (.A2(_11077_),
    .A1(_11017_),
    .B1(_11162_),
    .X(_11163_));
 sg13g2_buf_1 _18024_ (.A(_11163_),
    .X(_11164_));
 sg13g2_and2_1 _18025_ (.A(_10565_),
    .B(_10592_),
    .X(_11165_));
 sg13g2_buf_1 _18026_ (.A(_11165_),
    .X(_11166_));
 sg13g2_nor2_1 _18027_ (.A(_10562_),
    .B(_09290_),
    .Y(_11167_));
 sg13g2_buf_1 _18028_ (.A(\cpu.dec.imm[0] ),
    .X(_11168_));
 sg13g2_nor2_1 _18029_ (.A(_11168_),
    .B(_10141_),
    .Y(_11169_));
 sg13g2_a22oi_1 _18030_ (.Y(_11170_),
    .B1(_10242_),
    .B2(\cpu.ex.r_15[0] ),
    .A2(_10289_),
    .A1(\cpu.ex.r_9[0] ));
 sg13g2_nor2_1 _18031_ (.A(_10489_),
    .B(_11170_),
    .Y(_11171_));
 sg13g2_a22oi_1 _18032_ (.Y(_11172_),
    .B1(_10173_),
    .B2(\cpu.ex.r_11[0] ),
    .A2(net918),
    .A1(\cpu.ex.r_8[0] ));
 sg13g2_nor2_1 _18033_ (.A(_10336_),
    .B(_11172_),
    .Y(_11173_));
 sg13g2_mux2_1 _18034_ (.A0(\cpu.ex.r_12[0] ),
    .A1(\cpu.ex.r_13[0] ),
    .S(net915),
    .X(_11174_));
 sg13g2_nand3_1 _18035_ (.B(net787),
    .C(_11174_),
    .A(_10244_),
    .Y(_11175_));
 sg13g2_mux2_1 _18036_ (.A0(_09158_),
    .A1(\cpu.ex.r_stmp[0] ),
    .S(net913),
    .X(_11176_));
 sg13g2_nand3_1 _18037_ (.B(_10390_),
    .C(_11176_),
    .A(net793),
    .Y(_11177_));
 sg13g2_nand2_1 _18038_ (.Y(_11178_),
    .A(_11175_),
    .B(_11177_));
 sg13g2_a221oi_1 _18039_ (.B2(_10994_),
    .C1(_10190_),
    .B1(_10498_),
    .A1(\cpu.ex.r_10[0] ),
    .Y(_11179_),
    .A2(_10324_));
 sg13g2_a221oi_1 _18040_ (.B2(_10561_),
    .C1(_10208_),
    .B1(_10498_),
    .A1(\cpu.ex.r_14[0] ),
    .Y(_11180_),
    .A2(_10324_));
 sg13g2_nor3_1 _18041_ (.A(net788),
    .B(_11179_),
    .C(_11180_),
    .Y(_11181_));
 sg13g2_nor4_1 _18042_ (.A(_11171_),
    .B(_11173_),
    .C(_11178_),
    .D(_11181_),
    .Y(_11182_));
 sg13g2_nand2_1 _18043_ (.Y(_11183_),
    .A(net1162),
    .B(net563));
 sg13g2_o21ai_1 _18044_ (.B1(_11183_),
    .Y(_11184_),
    .A1(_10408_),
    .A2(_11182_));
 sg13g2_nor2_1 _18045_ (.A(net911),
    .B(_11184_),
    .Y(_11185_));
 sg13g2_or3_1 _18046_ (.A(_10138_),
    .B(_11169_),
    .C(_11185_),
    .X(_11186_));
 sg13g2_buf_2 _18047_ (.A(_11186_),
    .X(_11187_));
 sg13g2_a21o_1 _18048_ (.A2(_11167_),
    .A1(_11166_),
    .B1(_11187_),
    .X(_11188_));
 sg13g2_nand2b_1 _18049_ (.Y(_11189_),
    .B(_10560_),
    .A_N(_11188_));
 sg13g2_or4_1 _18050_ (.A(_10841_),
    .B(_10958_),
    .C(_11164_),
    .D(_11189_),
    .X(_11190_));
 sg13g2_nand2_1 _18051_ (.Y(_11191_),
    .A(_10603_),
    .B(_10560_));
 sg13g2_or2_1 _18052_ (.X(_11192_),
    .B(_11191_),
    .A(_11188_));
 sg13g2_or4_1 _18053_ (.A(_10841_),
    .B(_10958_),
    .C(_11164_),
    .D(_11192_),
    .X(_11193_));
 sg13g2_nor2_1 _18054_ (.A(net790),
    .B(_10341_),
    .Y(_11194_));
 sg13g2_nand2b_1 _18055_ (.Y(_11195_),
    .B(net786),
    .A_N(_00253_));
 sg13g2_o21ai_1 _18056_ (.B1(_11195_),
    .Y(_11196_),
    .A1(_11065_),
    .A2(net786));
 sg13g2_inv_1 _18057_ (.Y(_11197_),
    .A(\cpu.ex.r_sp[3] ));
 sg13g2_or2_1 _18058_ (.X(_11198_),
    .B(net912),
    .A(net915));
 sg13g2_buf_1 _18059_ (.A(_11198_),
    .X(_11199_));
 sg13g2_nand3_1 _18060_ (.B(net693),
    .C(net786),
    .A(\cpu.ex.r_11[3] ),
    .Y(_11200_));
 sg13g2_o21ai_1 _18061_ (.B1(_11200_),
    .Y(_11201_),
    .A1(_11197_),
    .A2(_11199_));
 sg13g2_nand3b_1 _18062_ (.B(net793),
    .C(\cpu.ex.mmu_read[3] ),
    .Y(_11202_),
    .A_N(_10388_));
 sg13g2_nand3b_1 _18063_ (.B(net786),
    .C(\cpu.ex.r_9[3] ),
    .Y(_11203_),
    .A_N(net793));
 sg13g2_a21oi_1 _18064_ (.A1(_11202_),
    .A2(_11203_),
    .Y(_11204_),
    .B1(_10395_));
 sg13g2_a221oi_1 _18065_ (.B2(_11201_),
    .C1(_11204_),
    .B1(_10393_),
    .A1(_11194_),
    .Y(_11205_),
    .A2(_11196_));
 sg13g2_nand3_1 _18066_ (.B(net793),
    .C(net795),
    .A(\cpu.ex.r_stmp[3] ),
    .Y(_11206_));
 sg13g2_nand3_1 _18067_ (.B(net788),
    .C(net916),
    .A(\cpu.ex.r_8[3] ),
    .Y(_11207_));
 sg13g2_a21o_1 _18068_ (.A2(_11207_),
    .A1(_11206_),
    .B1(net632),
    .X(_11208_));
 sg13g2_mux2_1 _18069_ (.A0(\cpu.ex.r_10[3] ),
    .A1(\cpu.ex.r_14[3] ),
    .S(net914),
    .X(_11209_));
 sg13g2_a221oi_1 _18070_ (.B2(net691),
    .C1(net693),
    .B1(_11209_),
    .A1(\cpu.ex.r_12[3] ),
    .Y(_11210_),
    .A2(_10260_));
 sg13g2_a21oi_1 _18071_ (.A1(\cpu.ex.r_13[3] ),
    .A2(_10260_),
    .Y(_11211_),
    .B1(net633));
 sg13g2_or3_1 _18072_ (.A(_10263_),
    .B(_11210_),
    .C(_11211_),
    .X(_11212_));
 sg13g2_nand3_1 _18073_ (.B(net633),
    .C(_10260_),
    .A(net1165),
    .Y(_11213_));
 sg13g2_mux2_1 _18074_ (.A0(\cpu.ex.r_lr[3] ),
    .A1(\cpu.ex.r_epc[3] ),
    .S(net792),
    .X(_11214_));
 sg13g2_nand2_1 _18075_ (.Y(_11215_),
    .A(_10346_),
    .B(_11214_));
 sg13g2_a21o_1 _18076_ (.A2(_11215_),
    .A1(_11213_),
    .B1(_10200_),
    .X(_11216_));
 sg13g2_and4_1 _18077_ (.A(_11205_),
    .B(_11208_),
    .C(_11212_),
    .D(_11216_),
    .X(_11217_));
 sg13g2_nand2_1 _18078_ (.Y(_11218_),
    .A(_09190_),
    .B(net563));
 sg13g2_o21ai_1 _18079_ (.B1(_11218_),
    .Y(_11219_),
    .A1(_10408_),
    .A2(_11217_));
 sg13g2_buf_2 _18080_ (.A(_11219_),
    .X(_11220_));
 sg13g2_buf_1 _18081_ (.A(\cpu.dec.imm[3] ),
    .X(_11221_));
 sg13g2_nand3_1 _18082_ (.B(_10134_),
    .C(_10228_),
    .A(_11221_),
    .Y(_11222_));
 sg13g2_o21ai_1 _18083_ (.B1(_11222_),
    .Y(_11223_),
    .A1(_10135_),
    .A2(_11073_));
 sg13g2_a21o_1 _18084_ (.A2(_10308_),
    .A1(_11220_),
    .B1(_11223_),
    .X(_11224_));
 sg13g2_buf_2 _18085_ (.A(_11224_),
    .X(_11225_));
 sg13g2_buf_8 _18086_ (.A(_11225_),
    .X(_11226_));
 sg13g2_nor2_1 _18087_ (.A(_10601_),
    .B(_11191_),
    .Y(_11227_));
 sg13g2_nor2_1 _18088_ (.A(net231),
    .B(_11227_),
    .Y(_11228_));
 sg13g2_a22oi_1 _18089_ (.Y(_11229_),
    .B1(_11193_),
    .B2(_11228_),
    .A2(_11190_),
    .A1(_10604_));
 sg13g2_buf_1 _18090_ (.A(_11229_),
    .X(_11230_));
 sg13g2_nand2_1 _18091_ (.Y(_11231_),
    .A(_10513_),
    .B(_10519_));
 sg13g2_nor2_1 _18092_ (.A(_11065_),
    .B(net303),
    .Y(_11232_));
 sg13g2_nor2_1 _18093_ (.A(_10513_),
    .B(_10519_),
    .Y(_11233_));
 sg13g2_a221oi_1 _18094_ (.B2(_11232_),
    .C1(_11233_),
    .B1(_11231_),
    .A1(net1133),
    .Y(_11234_),
    .A2(net260));
 sg13g2_inv_1 _18095_ (.Y(_11235_),
    .A(net1133));
 sg13g2_nand2_1 _18096_ (.Y(_11236_),
    .A(_11235_),
    .B(_10437_));
 sg13g2_o21ai_1 _18097_ (.B1(_11236_),
    .Y(_11237_),
    .A1(net1132),
    .A2(net261));
 sg13g2_nand2_1 _18098_ (.Y(_11238_),
    .A(net1132),
    .B(net261));
 sg13g2_o21ai_1 _18099_ (.B1(_11238_),
    .Y(_11239_),
    .A1(_11234_),
    .A2(_11237_));
 sg13g2_and2_1 _18100_ (.A(net564),
    .B(_11239_),
    .X(_11240_));
 sg13g2_inv_1 _18101_ (.Y(_11241_),
    .A(_11240_));
 sg13g2_o21ai_1 _18102_ (.B1(_11241_),
    .Y(_11242_),
    .A1(_10524_),
    .A2(_11230_));
 sg13g2_buf_2 _18103_ (.A(_11242_),
    .X(_11243_));
 sg13g2_a22oi_1 _18104_ (.Y(_11244_),
    .B1(_10374_),
    .B2(_11243_),
    .A2(_10358_),
    .A1(_10356_));
 sg13g2_buf_1 _18105_ (.A(_10232_),
    .X(_11245_));
 sg13g2_nor3_1 _18106_ (.A(net568),
    .B(_10355_),
    .C(net230),
    .Y(_11246_));
 sg13g2_buf_1 _18107_ (.A(_10311_),
    .X(_11247_));
 sg13g2_nor3_1 _18108_ (.A(net1137),
    .B(net229),
    .C(_11240_),
    .Y(_11248_));
 sg13g2_o21ai_1 _18109_ (.B1(_11248_),
    .Y(_11249_),
    .A1(_10524_),
    .A2(_11230_));
 sg13g2_or2_1 _18110_ (.X(_11250_),
    .B(net1137),
    .A(net1136));
 sg13g2_nand2_1 _18111_ (.Y(_11251_),
    .A(net1137),
    .B(net564));
 sg13g2_nor2_1 _18112_ (.A(net233),
    .B(_11251_),
    .Y(_11252_));
 sg13g2_and2_1 _18113_ (.A(net1136),
    .B(net1137),
    .X(_11253_));
 sg13g2_and2_1 _18114_ (.A(net564),
    .B(_11253_),
    .X(_11254_));
 sg13g2_o21ai_1 _18115_ (.B1(_11239_),
    .Y(_11255_),
    .A1(_11252_),
    .A2(_11254_));
 sg13g2_buf_1 _18116_ (.A(_10282_),
    .X(_11256_));
 sg13g2_a21oi_1 _18117_ (.A1(_10311_),
    .A2(_11253_),
    .Y(_11257_),
    .B1(net208));
 sg13g2_a21oi_1 _18118_ (.A1(_10443_),
    .A2(_10449_),
    .Y(_11258_),
    .B1(_10523_));
 sg13g2_inv_1 _18119_ (.Y(_11259_),
    .A(_10233_));
 sg13g2_nor2_1 _18120_ (.A(_11259_),
    .B(_10368_),
    .Y(_11260_));
 sg13g2_nand4_1 _18121_ (.B(_10604_),
    .C(_11190_),
    .A(_11258_),
    .Y(_11261_),
    .D(_11260_));
 sg13g2_inv_1 _18122_ (.Y(_11262_),
    .A(_11227_));
 sg13g2_nor3_1 _18123_ (.A(_11259_),
    .B(net231),
    .C(_10368_),
    .Y(_11263_));
 sg13g2_nand4_1 _18124_ (.B(_11193_),
    .C(_11262_),
    .A(_11258_),
    .Y(_11264_),
    .D(_11263_));
 sg13g2_nand4_1 _18125_ (.B(_11257_),
    .C(_11261_),
    .A(_11255_),
    .Y(_11265_),
    .D(_11264_));
 sg13g2_nand4_1 _18126_ (.B(_11249_),
    .C(_11250_),
    .A(_11246_),
    .Y(_11266_),
    .D(_11265_));
 sg13g2_inv_1 _18127_ (.Y(_11267_),
    .A(net1134));
 sg13g2_inv_1 _18128_ (.Y(_11268_),
    .A(_10831_));
 sg13g2_nor2_1 _18129_ (.A(_11268_),
    .B(net562),
    .Y(_11269_));
 sg13g2_nor2b_1 _18130_ (.A(net560),
    .B_N(\cpu.ex.r_14[12] ),
    .Y(_11270_));
 sg13g2_a22oi_1 _18131_ (.Y(_11271_),
    .B1(_11270_),
    .B2(_10400_),
    .A2(_11269_),
    .A1(_10403_));
 sg13g2_inv_1 _18132_ (.Y(_11272_),
    .A(\cpu.ex.r_sp[12] ));
 sg13g2_nand3_1 _18133_ (.B(net632),
    .C(net690),
    .A(\cpu.ex.r_11[12] ),
    .Y(_11273_));
 sg13g2_o21ai_1 _18134_ (.B1(_11273_),
    .Y(_11274_),
    .A1(_11272_),
    .A2(_11199_));
 sg13g2_nand3b_1 _18135_ (.B(net690),
    .C(\cpu.ex.r_9[12] ),
    .Y(_11275_),
    .A_N(net631));
 sg13g2_o21ai_1 _18136_ (.B1(_11275_),
    .Y(_11276_),
    .A1(_10824_),
    .A2(_10345_));
 sg13g2_a221oi_1 _18137_ (.B2(net560),
    .C1(net561),
    .B1(_11276_),
    .A1(net631),
    .Y(_11277_),
    .A2(_11274_));
 sg13g2_a21oi_1 _18138_ (.A1(net561),
    .A2(_11271_),
    .Y(_11278_),
    .B1(_11277_));
 sg13g2_a22oi_1 _18139_ (.Y(_11279_),
    .B1(net787),
    .B2(\cpu.ex.r_13[12] ),
    .A2(net917),
    .A1(\cpu.ex.r_lr[12] ));
 sg13g2_mux2_1 _18140_ (.A0(_10816_),
    .A1(_10812_),
    .S(_10263_),
    .X(_11280_));
 sg13g2_inv_1 _18141_ (.Y(_11281_),
    .A(\cpu.ex.r_10[12] ));
 sg13g2_nand3b_1 _18142_ (.B(net634),
    .C(\cpu.ex.r_stmp[12] ),
    .Y(_11282_),
    .A_N(net690));
 sg13g2_o21ai_1 _18143_ (.B1(_11282_),
    .Y(_11283_),
    .A1(_11281_),
    .A2(_10336_));
 sg13g2_mux2_1 _18144_ (.A0(\cpu.ex.r_8[12] ),
    .A1(\cpu.ex.r_12[12] ),
    .S(net634),
    .X(_11284_));
 sg13g2_and3_1 _18145_ (.X(_11285_),
    .A(net630),
    .B(net918),
    .C(_11284_));
 sg13g2_a221oi_1 _18146_ (.B2(net789),
    .C1(_11285_),
    .B1(_11283_),
    .A1(_11194_),
    .Y(_11286_),
    .A2(_11280_));
 sg13g2_o21ai_1 _18147_ (.B1(_11286_),
    .Y(_11287_),
    .A1(_10395_),
    .A2(_11279_));
 sg13g2_nor2_1 _18148_ (.A(_11278_),
    .B(_11287_),
    .Y(_11288_));
 sg13g2_nand2_1 _18149_ (.Y(_11289_),
    .A(net627),
    .B(net490));
 sg13g2_o21ai_1 _18150_ (.B1(_11289_),
    .Y(_11290_),
    .A1(_10408_),
    .A2(_11288_));
 sg13g2_inv_1 _18151_ (.Y(_11291_),
    .A(\cpu.dec.imm[12] ));
 sg13g2_nor2_1 _18152_ (.A(net1050),
    .B(_11291_),
    .Y(_11292_));
 sg13g2_a21oi_1 _18153_ (.A1(net1050),
    .A2(_11290_),
    .Y(_11293_),
    .B1(_11292_));
 sg13g2_mux2_1 _18154_ (.A0(_10778_),
    .A1(_11293_),
    .S(net920),
    .X(_11294_));
 sg13g2_buf_1 _18155_ (.A(_11294_),
    .X(_11295_));
 sg13g2_buf_1 _18156_ (.A(_11295_),
    .X(_11296_));
 sg13g2_buf_1 _18157_ (.A(_10812_),
    .X(_11297_));
 sg13g2_inv_1 _18158_ (.Y(_11298_),
    .A(\cpu.dec.imm[13] ));
 sg13g2_nand3_1 _18159_ (.B(net560),
    .C(net917),
    .A(\cpu.ex.r_lr[13] ),
    .Y(_11299_));
 sg13g2_nand3_1 _18160_ (.B(net562),
    .C(net787),
    .A(\cpu.ex.r_12[13] ),
    .Y(_11300_));
 sg13g2_a21o_1 _18161_ (.A2(_11300_),
    .A1(_11299_),
    .B1(net631),
    .X(_11301_));
 sg13g2_and3_1 _18162_ (.X(_11302_),
    .A(\cpu.ex.r_14[13] ),
    .B(net690),
    .C(net634));
 sg13g2_a21o_1 _18163_ (.A2(net917),
    .A1(_10791_),
    .B1(_11302_),
    .X(_11303_));
 sg13g2_inv_1 _18164_ (.Y(_11304_),
    .A(\cpu.ex.r_stmp[13] ));
 sg13g2_nand3b_1 _18165_ (.B(net632),
    .C(net690),
    .Y(_11305_),
    .A_N(_00263_));
 sg13g2_o21ai_1 _18166_ (.B1(_11305_),
    .Y(_11306_),
    .A1(_11304_),
    .A2(_11199_));
 sg13g2_mux2_1 _18167_ (.A0(\cpu.ex.r_8[13] ),
    .A1(\cpu.ex.r_10[13] ),
    .S(net691),
    .X(_11307_));
 sg13g2_and3_1 _18168_ (.X(_11308_),
    .A(net790),
    .B(_10324_),
    .C(_11307_));
 sg13g2_a221oi_1 _18169_ (.B2(_10242_),
    .C1(_11308_),
    .B1(_11306_),
    .A1(net789),
    .Y(_11309_),
    .A2(_11303_));
 sg13g2_a221oi_1 _18170_ (.B2(\cpu.ex.r_epc[13] ),
    .C1(net630),
    .B1(_10393_),
    .A1(_10798_),
    .Y(_11310_),
    .A2(_10260_));
 sg13g2_a221oi_1 _18171_ (.B2(\cpu.ex.r_11[13] ),
    .C1(_10263_),
    .B1(_10393_),
    .A1(\cpu.ex.r_13[13] ),
    .Y(_11311_),
    .A2(_10260_));
 sg13g2_or3_1 _18172_ (.A(net562),
    .B(_11310_),
    .C(_11311_),
    .X(_11312_));
 sg13g2_and3_1 _18173_ (.X(_11313_),
    .A(\cpu.ex.r_9[13] ),
    .B(net788),
    .C(net916));
 sg13g2_and3_1 _18174_ (.X(_11314_),
    .A(_10795_),
    .B(net561),
    .C(net795));
 sg13g2_o21ai_1 _18175_ (.B1(net560),
    .Y(_11315_),
    .A1(_11313_),
    .A2(_11314_));
 sg13g2_nand4_1 _18176_ (.B(_11309_),
    .C(_11312_),
    .A(_11301_),
    .Y(_11316_),
    .D(_11315_));
 sg13g2_a22oi_1 _18177_ (.Y(_11317_),
    .B1(_10273_),
    .B2(_11316_),
    .A2(_10235_),
    .A1(net628));
 sg13g2_mux2_1 _18178_ (.A0(_11298_),
    .A1(_11317_),
    .S(net1050),
    .X(_11318_));
 sg13g2_mux2_1 _18179_ (.A0(_10777_),
    .A1(_11318_),
    .S(net920),
    .X(_11319_));
 sg13g2_buf_1 _18180_ (.A(_11319_),
    .X(_11320_));
 sg13g2_buf_1 _18181_ (.A(_11320_),
    .X(_11321_));
 sg13g2_xnor2_1 _18182_ (.Y(_11322_),
    .A(net1037),
    .B(net207));
 sg13g2_nor3_1 _18183_ (.A(_11267_),
    .B(net181),
    .C(_11322_),
    .Y(_11323_));
 sg13g2_inv_1 _18184_ (.Y(_11324_),
    .A(_10777_));
 sg13g2_nand2_1 _18185_ (.Y(_11325_),
    .A(net919),
    .B(_11324_));
 sg13g2_o21ai_1 _18186_ (.B1(_11325_),
    .Y(_11326_),
    .A1(net919),
    .A2(_11318_));
 sg13g2_buf_1 _18187_ (.A(_11326_),
    .X(_11327_));
 sg13g2_buf_1 _18188_ (.A(_11327_),
    .X(_11328_));
 sg13g2_and4_1 _18189_ (.A(_11267_),
    .B(net1037),
    .C(net206),
    .D(net181),
    .X(_11329_));
 sg13g2_o21ai_1 _18190_ (.B1(_10127_),
    .Y(_11330_),
    .A1(_11323_),
    .A2(_11329_));
 sg13g2_buf_1 _18191_ (.A(_11296_),
    .X(_11331_));
 sg13g2_o21ai_1 _18192_ (.B1(net564),
    .Y(_11332_),
    .A1(net1134),
    .A2(net1037));
 sg13g2_nand3_1 _18193_ (.B(net150),
    .C(_11332_),
    .A(net207),
    .Y(_11333_));
 sg13g2_buf_1 _18194_ (.A(_10795_),
    .X(_11334_));
 sg13g2_inv_1 _18195_ (.Y(_11335_),
    .A(\cpu.dec.imm[15] ));
 sg13g2_inv_1 _18196_ (.Y(_11336_),
    .A(net1125));
 sg13g2_nand2_1 _18197_ (.Y(_11337_),
    .A(\cpu.ex.r_13[15] ),
    .B(net630));
 sg13g2_o21ai_1 _18198_ (.B1(_11337_),
    .Y(_11338_),
    .A1(net1035),
    .A2(net630));
 sg13g2_nor2b_1 _18199_ (.A(net560),
    .B_N(\cpu.ex.r_8[15] ),
    .Y(_11339_));
 sg13g2_a22oi_1 _18200_ (.Y(_11340_),
    .B1(_11339_),
    .B2(net916),
    .A2(_11338_),
    .A1(_10285_));
 sg13g2_mux2_1 _18201_ (.A0(\cpu.ex.r_10[15] ),
    .A1(\cpu.ex.r_14[15] ),
    .S(net634),
    .X(_11341_));
 sg13g2_a22oi_1 _18202_ (.Y(_11342_),
    .B1(_11341_),
    .B2(net630),
    .A2(net917),
    .A1(_10734_));
 sg13g2_nand2b_1 _18203_ (.Y(_11343_),
    .B(net789),
    .A_N(_11342_));
 sg13g2_o21ai_1 _18204_ (.B1(_11343_),
    .Y(_11344_),
    .A1(net631),
    .A2(_11340_));
 sg13g2_a22oi_1 _18205_ (.Y(_11345_),
    .B1(_10403_),
    .B2(\cpu.ex.r_lr[15] ),
    .A2(_10400_),
    .A1(\cpu.ex.r_11[15] ));
 sg13g2_nor2_1 _18206_ (.A(_10186_),
    .B(_11345_),
    .Y(_11346_));
 sg13g2_a22oi_1 _18207_ (.Y(_11347_),
    .B1(_10390_),
    .B2(\cpu.ex.r_stmp[15] ),
    .A2(_10389_),
    .A1(_10763_));
 sg13g2_nor2b_1 _18208_ (.A(_11347_),
    .B_N(_10242_),
    .Y(_11348_));
 sg13g2_a22oi_1 _18209_ (.Y(_11349_),
    .B1(net795),
    .B2(\cpu.ex.r_epc[15] ),
    .A2(_10268_),
    .A1(\cpu.ex.r_9[15] ));
 sg13g2_nor2_1 _18210_ (.A(_10186_),
    .B(_11349_),
    .Y(_11350_));
 sg13g2_nand3_1 _18211_ (.B(net630),
    .C(net918),
    .A(\cpu.ex.r_12[15] ),
    .Y(_11351_));
 sg13g2_nand3_1 _18212_ (.B(net560),
    .C(net795),
    .A(\cpu.ex.r_mult[31] ),
    .Y(_11352_));
 sg13g2_a21oi_1 _18213_ (.A1(_11351_),
    .A2(_11352_),
    .Y(_11353_),
    .B1(net790));
 sg13g2_nor4_1 _18214_ (.A(_11346_),
    .B(_11348_),
    .C(_11350_),
    .D(_11353_),
    .Y(_11354_));
 sg13g2_nand2b_1 _18215_ (.Y(_11355_),
    .B(_11354_),
    .A_N(_11344_));
 sg13g2_a22oi_1 _18216_ (.Y(_11356_),
    .B1(net440),
    .B2(_11355_),
    .A2(net490),
    .A1(net687));
 sg13g2_mux2_1 _18217_ (.A0(_11335_),
    .A1(_11356_),
    .S(net1050),
    .X(_11357_));
 sg13g2_nand2b_1 _18218_ (.Y(_11358_),
    .B(net919),
    .A_N(_00192_));
 sg13g2_o21ai_1 _18219_ (.B1(_11358_),
    .Y(_11359_),
    .A1(net919),
    .A2(_11357_));
 sg13g2_buf_2 _18220_ (.A(_11359_),
    .X(_11360_));
 sg13g2_buf_1 _18221_ (.A(_11360_),
    .X(_11361_));
 sg13g2_inv_1 _18222_ (.Y(_11362_),
    .A(_00193_));
 sg13g2_mux2_1 _18223_ (.A0(\cpu.ex.r_9[14] ),
    .A1(\cpu.ex.r_11[14] ),
    .S(net631),
    .X(_11363_));
 sg13g2_a22oi_1 _18224_ (.Y(_11364_),
    .B1(_11363_),
    .B2(net560),
    .A2(_10210_),
    .A1(\cpu.ex.r_10[14] ));
 sg13g2_nor2_1 _18225_ (.A(_10336_),
    .B(_11364_),
    .Y(_11365_));
 sg13g2_mux2_1 _18226_ (.A0(_10697_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(net561),
    .X(_11366_));
 sg13g2_a22oi_1 _18227_ (.Y(_11367_),
    .B1(_11366_),
    .B2(_10257_),
    .A2(_10285_),
    .A1(net1126));
 sg13g2_nor2_1 _18228_ (.A(_10345_),
    .B(_11367_),
    .Y(_11368_));
 sg13g2_nor2b_1 _18229_ (.A(net561),
    .B_N(\cpu.ex.r_lr[14] ),
    .Y(_11369_));
 sg13g2_a22oi_1 _18230_ (.Y(_11370_),
    .B1(_10403_),
    .B2(_11369_),
    .A2(_10202_),
    .A1(_10685_));
 sg13g2_mux2_1 _18231_ (.A0(\cpu.ex.r_8[14] ),
    .A1(\cpu.ex.r_12[14] ),
    .S(net561),
    .X(_11371_));
 sg13g2_nand3_1 _18232_ (.B(_10167_),
    .C(_11371_),
    .A(net630),
    .Y(_11372_));
 sg13g2_o21ai_1 _18233_ (.B1(_11372_),
    .Y(_11373_),
    .A1(net562),
    .A2(_11370_));
 sg13g2_a22oi_1 _18234_ (.Y(_11374_),
    .B1(_10210_),
    .B2(\cpu.ex.r_14[14] ),
    .A2(_10224_),
    .A1(\cpu.ex.r_13[14] ));
 sg13g2_buf_1 _18235_ (.A(\cpu.ex.mmu_read[14] ),
    .X(_11375_));
 sg13g2_nand3b_1 _18236_ (.B(_10270_),
    .C(net1123),
    .Y(_11376_),
    .A_N(_10250_));
 sg13g2_nand3b_1 _18237_ (.B(net631),
    .C(\cpu.ex.r_epc[14] ),
    .Y(_11377_),
    .A_N(net561));
 sg13g2_nand2b_1 _18238_ (.Y(_11378_),
    .B(_10383_),
    .A_N(net630));
 sg13g2_a21o_1 _18239_ (.A2(_11377_),
    .A1(_11376_),
    .B1(_11378_),
    .X(_11379_));
 sg13g2_o21ai_1 _18240_ (.B1(_11379_),
    .Y(_11380_),
    .A1(_10526_),
    .A2(_11374_));
 sg13g2_or4_1 _18241_ (.A(_11365_),
    .B(_11368_),
    .C(_11373_),
    .D(_11380_),
    .X(_11381_));
 sg13g2_a22oi_1 _18242_ (.Y(_11382_),
    .B1(net440),
    .B2(_11381_),
    .A2(net490),
    .A1(net698));
 sg13g2_nor2_1 _18243_ (.A(net1050),
    .B(\cpu.dec.imm[14] ),
    .Y(_11383_));
 sg13g2_a21oi_1 _18244_ (.A1(net1050),
    .A2(_11382_),
    .Y(_11384_),
    .B1(_11383_));
 sg13g2_mux2_1 _18245_ (.A0(_11362_),
    .A1(_11384_),
    .S(net920),
    .X(_11385_));
 sg13g2_buf_2 _18246_ (.A(_11385_),
    .X(_11386_));
 sg13g2_inv_1 _18247_ (.Y(_11387_),
    .A(_11386_));
 sg13g2_nand3_1 _18248_ (.B(net180),
    .C(_11387_),
    .A(net1126),
    .Y(_11388_));
 sg13g2_buf_1 _18249_ (.A(_11386_),
    .X(_11389_));
 sg13g2_xnor2_1 _18250_ (.Y(_11390_),
    .A(net1126),
    .B(net180));
 sg13g2_nand3_1 _18251_ (.B(net179),
    .C(_11390_),
    .A(net1036),
    .Y(_11391_));
 sg13g2_o21ai_1 _18252_ (.B1(_11391_),
    .Y(_11392_),
    .A1(net1036),
    .A2(_11388_));
 sg13g2_o21ai_1 _18253_ (.B1(net564),
    .Y(_11393_),
    .A1(net1036),
    .A2(net1126));
 sg13g2_nor2_1 _18254_ (.A(net180),
    .B(_11386_),
    .Y(_11394_));
 sg13g2_a22oi_1 _18255_ (.Y(_11395_),
    .B1(_11393_),
    .B2(_11394_),
    .A2(_11392_),
    .A1(net564));
 sg13g2_a221oi_1 _18256_ (.B2(_11333_),
    .C1(_11395_),
    .B1(_11330_),
    .A1(_11244_),
    .Y(_11396_),
    .A2(_11266_));
 sg13g2_buf_1 _18257_ (.A(_11396_),
    .X(_11397_));
 sg13g2_nand2b_1 _18258_ (.Y(_11398_),
    .B(_11386_),
    .A_N(_11334_));
 sg13g2_inv_1 _18259_ (.Y(_11399_),
    .A(_10778_));
 sg13g2_nand2_1 _18260_ (.Y(_11400_),
    .A(net919),
    .B(_11399_));
 sg13g2_o21ai_1 _18261_ (.B1(_11400_),
    .Y(_11401_),
    .A1(net919),
    .A2(_11293_));
 sg13g2_buf_2 _18262_ (.A(_11401_),
    .X(_11402_));
 sg13g2_o21ai_1 _18263_ (.B1(net1134),
    .Y(_11403_),
    .A1(_11297_),
    .A2(_11320_));
 sg13g2_nand2_1 _18264_ (.Y(_11404_),
    .A(_11297_),
    .B(_11320_));
 sg13g2_o21ai_1 _18265_ (.B1(_11404_),
    .Y(_11405_),
    .A1(_11402_),
    .A2(_11403_));
 sg13g2_and2_1 _18266_ (.A(_11334_),
    .B(_11387_),
    .X(_11406_));
 sg13g2_a21oi_1 _18267_ (.A1(_11398_),
    .A2(_11405_),
    .Y(_11407_),
    .B1(_11406_));
 sg13g2_nand2_1 _18268_ (.Y(_11408_),
    .A(net180),
    .B(_11407_));
 sg13g2_nor2_1 _18269_ (.A(net180),
    .B(_11407_),
    .Y(_11409_));
 sg13g2_a21oi_1 _18270_ (.A1(net1126),
    .A2(_11408_),
    .Y(_11410_),
    .B1(_11409_));
 sg13g2_nor2_1 _18271_ (.A(net568),
    .B(_11410_),
    .Y(_11411_));
 sg13g2_nor3_1 _18272_ (.A(net1051),
    .B(_11169_),
    .C(_11185_),
    .Y(_11412_));
 sg13g2_buf_2 _18273_ (.A(_11412_),
    .X(_11413_));
 sg13g2_a21oi_1 _18274_ (.A1(_11220_),
    .A2(_10308_),
    .Y(_11414_),
    .B1(_11223_));
 sg13g2_buf_2 _18275_ (.A(_11414_),
    .X(_11415_));
 sg13g2_buf_1 _18276_ (.A(net302),
    .X(_11416_));
 sg13g2_nand2_1 _18277_ (.Y(_11417_),
    .A(_11415_),
    .B(net259));
 sg13g2_buf_1 _18278_ (.A(_11417_),
    .X(_11418_));
 sg13g2_buf_1 _18279_ (.A(_10594_),
    .X(_11419_));
 sg13g2_nor3_2 _18280_ (.A(_11413_),
    .B(net205),
    .C(net228),
    .Y(_11420_));
 sg13g2_nand4_1 _18281_ (.B(_10366_),
    .C(_10367_),
    .A(_11420_),
    .Y(_11421_),
    .D(_10521_));
 sg13g2_nand2_1 _18282_ (.Y(_11422_),
    .A(_11320_),
    .B(net181));
 sg13g2_nand3_1 _18283_ (.B(net261),
    .C(net260),
    .A(_11394_),
    .Y(_11423_));
 sg13g2_nor3_1 _18284_ (.A(_11421_),
    .B(_11422_),
    .C(_11423_),
    .Y(_11424_));
 sg13g2_buf_2 _18285_ (.A(_11424_),
    .X(_11425_));
 sg13g2_buf_1 _18286_ (.A(_11425_),
    .X(_11426_));
 sg13g2_inv_1 _18287_ (.Y(_11427_),
    .A(net74));
 sg13g2_o21ai_1 _18288_ (.B1(_11427_),
    .Y(_11428_),
    .A1(_11397_),
    .A2(_11411_));
 sg13g2_nand2_1 _18289_ (.Y(_11429_),
    .A(_10150_),
    .B(\cpu.dec.r_set_cc ));
 sg13g2_inv_1 _18290_ (.Y(_11430_),
    .A(_10148_));
 sg13g2_nor2_1 _18291_ (.A(net1141),
    .B(_11430_),
    .Y(_11431_));
 sg13g2_nand4_1 _18292_ (.B(net1043),
    .C(_10150_),
    .A(net1142),
    .Y(_11432_),
    .D(_11431_));
 sg13g2_buf_2 _18293_ (.A(_11432_),
    .X(_11433_));
 sg13g2_and2_1 _18294_ (.A(_11429_),
    .B(_11433_),
    .X(_11434_));
 sg13g2_buf_2 _18295_ (.A(_11434_),
    .X(_11435_));
 sg13g2_buf_1 _18296_ (.A(_11187_),
    .X(_11436_));
 sg13g2_nor3_1 _18297_ (.A(_10841_),
    .B(_10958_),
    .C(_11164_),
    .Y(_11437_));
 sg13g2_buf_1 _18298_ (.A(_11437_),
    .X(_11438_));
 sg13g2_buf_1 _18299_ (.A(net110),
    .X(_11439_));
 sg13g2_o21ai_1 _18300_ (.B1(net492),
    .Y(_11440_),
    .A1(net258),
    .A2(net91));
 sg13g2_inv_1 _18301_ (.Y(_11441_),
    .A(\cpu.ex.r_mult[0] ));
 sg13g2_buf_1 _18302_ (.A(_10127_),
    .X(_11442_));
 sg13g2_buf_1 _18303_ (.A(net626),
    .X(_11443_));
 sg13g2_buf_1 _18304_ (.A(net557),
    .X(_11444_));
 sg13g2_nor2_2 _18305_ (.A(_09293_),
    .B(net488),
    .Y(_11445_));
 sg13g2_nand4_1 _18306_ (.B(_11441_),
    .C(net489),
    .A(_10124_),
    .Y(_11446_),
    .D(_11445_));
 sg13g2_nand3_1 _18307_ (.B(_11440_),
    .C(_11446_),
    .A(_11435_),
    .Y(_11447_));
 sg13g2_a21o_1 _18308_ (.A2(_11428_),
    .A1(net348),
    .B1(_11447_),
    .X(_11448_));
 sg13g2_nand2_1 _18309_ (.Y(_11449_),
    .A(net1142),
    .B(net1043));
 sg13g2_inv_1 _18310_ (.Y(_11450_),
    .A(_11431_));
 sg13g2_nor3_1 _18311_ (.A(_10151_),
    .B(_11449_),
    .C(_11450_),
    .Y(_11451_));
 sg13g2_buf_1 _18312_ (.A(_11451_),
    .X(_11452_));
 sg13g2_buf_1 _18313_ (.A(_11452_),
    .X(_11453_));
 sg13g2_or2_1 _18314_ (.X(_11454_),
    .B(_10770_),
    .A(_10727_));
 sg13g2_buf_2 _18315_ (.A(_11454_),
    .X(_11455_));
 sg13g2_and2_1 _18316_ (.A(_11455_),
    .B(net180),
    .X(_11456_));
 sg13g2_buf_1 _18317_ (.A(_11456_),
    .X(_11457_));
 sg13g2_nor2_1 _18318_ (.A(_11429_),
    .B(_11453_),
    .Y(_11458_));
 sg13g2_a22oi_1 _18319_ (.Y(_11459_),
    .B1(_11457_),
    .B2(_11458_),
    .A2(net556),
    .A1(\cpu.ex.r_mult[0] ));
 sg13g2_buf_1 _18320_ (.A(_11455_),
    .X(_11460_));
 sg13g2_or2_1 _18321_ (.X(_11461_),
    .B(net180),
    .A(_11460_));
 sg13g2_buf_1 _18322_ (.A(_11461_),
    .X(_11462_));
 sg13g2_a21oi_1 _18323_ (.A1(_11441_),
    .A2(_11452_),
    .Y(_11463_),
    .B1(_11429_));
 sg13g2_nor2_1 _18324_ (.A(_10724_),
    .B(_10726_),
    .Y(_11464_));
 sg13g2_nand2_1 _18325_ (.Y(_11465_),
    .A(_11399_),
    .B(_11464_));
 sg13g2_o21ai_1 _18326_ (.B1(_11465_),
    .Y(_11466_),
    .A1(_11464_),
    .A2(_10836_));
 sg13g2_buf_1 _18327_ (.A(_11466_),
    .X(_11467_));
 sg13g2_buf_1 _18328_ (.A(_11402_),
    .X(_11468_));
 sg13g2_nor2_1 _18329_ (.A(net204),
    .B(net177),
    .Y(_11469_));
 sg13g2_nand2_1 _18330_ (.Y(_11470_),
    .A(net301),
    .B(_10903_));
 sg13g2_o21ai_1 _18331_ (.B1(_11470_),
    .Y(_11471_),
    .A1(_11464_),
    .A2(_10923_));
 sg13g2_buf_1 _18332_ (.A(_11471_),
    .X(_11472_));
 sg13g2_nor2_1 _18333_ (.A(_10900_),
    .B(_10282_),
    .Y(_11473_));
 sg13g2_a21oi_1 _18334_ (.A1(_11472_),
    .A2(net233),
    .Y(_11474_),
    .B1(_11473_));
 sg13g2_buf_8 _18335_ (.A(_11166_),
    .X(_11475_));
 sg13g2_nor2_1 _18336_ (.A(_10627_),
    .B(_10563_),
    .Y(_11476_));
 sg13g2_o21ai_1 _18337_ (.B1(_11476_),
    .Y(_11477_),
    .A1(_08359_),
    .A2(_08415_));
 sg13g2_nand4_1 _18338_ (.B(net438),
    .C(_10623_),
    .A(net439),
    .Y(_11478_),
    .D(_11040_));
 sg13g2_nor2b_1 _18339_ (.A(net498),
    .B_N(_11476_),
    .Y(_11479_));
 sg13g2_a221oi_1 _18340_ (.B2(_10631_),
    .C1(_11479_),
    .B1(_11476_),
    .A1(_10628_),
    .Y(_11480_),
    .A2(_11040_));
 sg13g2_and3_1 _18341_ (.X(_11481_),
    .A(_11477_),
    .B(_11478_),
    .C(_11480_));
 sg13g2_buf_8 _18342_ (.A(_11481_),
    .X(_11482_));
 sg13g2_nor2_1 _18343_ (.A(net227),
    .B(_11482_),
    .Y(_11483_));
 sg13g2_buf_2 _18344_ (.A(_11483_),
    .X(_11484_));
 sg13g2_nand2_1 _18345_ (.Y(_11485_),
    .A(_10985_),
    .B(_11006_));
 sg13g2_inv_1 _18346_ (.Y(_11486_),
    .A(_11485_));
 sg13g2_o21ai_1 _18347_ (.B1(_11486_),
    .Y(_11487_),
    .A1(net778),
    .A2(_10726_));
 sg13g2_nand2_1 _18348_ (.Y(_11488_),
    .A(net347),
    .B(_11015_));
 sg13g2_a221oi_1 _18349_ (.B2(_11488_),
    .C1(_11187_),
    .B1(_11487_),
    .A1(net227),
    .Y(_11489_),
    .A2(_11482_));
 sg13g2_buf_1 _18350_ (.A(_11489_),
    .X(_11490_));
 sg13g2_nor2_1 _18351_ (.A(_10477_),
    .B(_10478_),
    .Y(_11491_));
 sg13g2_a21oi_1 _18352_ (.A1(net1076),
    .A2(net1051),
    .Y(_11492_),
    .B1(_11491_));
 sg13g2_buf_2 _18353_ (.A(_11492_),
    .X(_11493_));
 sg13g2_nand2_1 _18354_ (.Y(_11494_),
    .A(net1076),
    .B(net1127));
 sg13g2_a21oi_1 _18355_ (.A1(net439),
    .A2(net438),
    .Y(_11495_),
    .B1(_11494_));
 sg13g2_and4_1 _18356_ (.A(net439),
    .B(net438),
    .C(_10623_),
    .D(_11142_),
    .X(_11496_));
 sg13g2_buf_1 _18357_ (.A(_11496_),
    .X(_11497_));
 sg13g2_a21oi_1 _18358_ (.A1(net498),
    .A2(_10621_),
    .Y(_11498_),
    .B1(_08448_));
 sg13g2_mux2_1 _18359_ (.A0(_11142_),
    .A1(_11498_),
    .S(_10626_),
    .X(_11499_));
 sg13g2_buf_1 _18360_ (.A(_11499_),
    .X(_11500_));
 sg13g2_nor3_1 _18361_ (.A(_11495_),
    .B(_11497_),
    .C(_11500_),
    .Y(_11501_));
 sg13g2_buf_1 _18362_ (.A(_11501_),
    .X(_11502_));
 sg13g2_nor2_1 _18363_ (.A(net910),
    .B(_00283_),
    .Y(_11503_));
 sg13g2_nor2_1 _18364_ (.A(_09174_),
    .B(net559),
    .Y(_11504_));
 sg13g2_nor2_1 _18365_ (.A(_10969_),
    .B(_10981_),
    .Y(_11505_));
 sg13g2_nor4_1 _18366_ (.A(_09108_),
    .B(net437),
    .C(_11504_),
    .D(_11505_),
    .Y(_11506_));
 sg13g2_nor3_1 _18367_ (.A(net1038),
    .B(_11504_),
    .C(_11505_),
    .Y(_11507_));
 sg13g2_a221oi_1 _18368_ (.B2(net358),
    .C1(_11507_),
    .B1(_11506_),
    .A1(_10729_),
    .Y(_11508_),
    .A2(_11503_));
 sg13g2_buf_2 _18369_ (.A(_11508_),
    .X(_11509_));
 sg13g2_buf_8 _18370_ (.A(_11509_),
    .X(_11510_));
 sg13g2_nor2_1 _18371_ (.A(_10628_),
    .B(_11073_),
    .Y(_11511_));
 sg13g2_and2_1 _18372_ (.A(_11056_),
    .B(_11068_),
    .X(_11512_));
 sg13g2_nor4_1 _18373_ (.A(_09108_),
    .B(net437),
    .C(_11069_),
    .D(_11512_),
    .Y(_11513_));
 sg13g2_nor3_1 _18374_ (.A(net1127),
    .B(_11069_),
    .C(_11512_),
    .Y(_11514_));
 sg13g2_a221oi_1 _18375_ (.B2(net358),
    .C1(_11514_),
    .B1(_11513_),
    .A1(net301),
    .Y(_11515_),
    .A2(_11511_));
 sg13g2_buf_1 _18376_ (.A(_11515_),
    .X(_11516_));
 sg13g2_buf_8 _18377_ (.A(_11516_),
    .X(_11517_));
 sg13g2_a221oi_1 _18378_ (.B2(net302),
    .C1(net202),
    .B1(net203),
    .A1(_11493_),
    .Y(_11518_),
    .A2(net257));
 sg13g2_o21ai_1 _18379_ (.B1(_11518_),
    .Y(_11519_),
    .A1(_11484_),
    .A2(_11490_));
 sg13g2_a221oi_1 _18380_ (.B2(net302),
    .C1(_11415_),
    .B1(_11509_),
    .A1(_11493_),
    .Y(_11520_),
    .A2(net257));
 sg13g2_o21ai_1 _18381_ (.B1(_11520_),
    .Y(_11521_),
    .A1(_11484_),
    .A2(_11490_));
 sg13g2_nor4_2 _18382_ (.A(_10481_),
    .B(_11495_),
    .C(_11497_),
    .Y(_11522_),
    .D(_11500_));
 sg13g2_nor4_1 _18383_ (.A(net302),
    .B(_11522_),
    .C(net202),
    .D(_11509_),
    .Y(_11523_));
 sg13g2_nor4_1 _18384_ (.A(_11415_),
    .B(net302),
    .C(_11522_),
    .D(_11509_),
    .Y(_11524_));
 sg13g2_nor3_1 _18385_ (.A(_11415_),
    .B(_11522_),
    .C(net202),
    .Y(_11525_));
 sg13g2_nor3_1 _18386_ (.A(_11523_),
    .B(_11524_),
    .C(_11525_),
    .Y(_11526_));
 sg13g2_nand3_1 _18387_ (.B(_11521_),
    .C(_11526_),
    .A(_11519_),
    .Y(_11527_));
 sg13g2_or2_1 _18388_ (.X(_11528_),
    .B(_10414_),
    .A(_10410_));
 sg13g2_buf_2 _18389_ (.A(_11528_),
    .X(_11529_));
 sg13g2_and4_1 _18390_ (.A(net498),
    .B(_10621_),
    .C(_11101_),
    .D(_11119_),
    .X(_11530_));
 sg13g2_nand3_1 _18391_ (.B(net438),
    .C(_11530_),
    .A(net439),
    .Y(_11531_));
 sg13g2_nor2_1 _18392_ (.A(net910),
    .B(_10411_),
    .Y(_11532_));
 sg13g2_o21ai_1 _18393_ (.B1(_11532_),
    .Y(_11533_),
    .A1(_08359_),
    .A2(_08415_));
 sg13g2_nand2_1 _18394_ (.Y(_11534_),
    .A(_09108_),
    .B(_11532_));
 sg13g2_a22oi_1 _18395_ (.Y(_11535_),
    .B1(_11532_),
    .B2(net437),
    .A2(_11121_),
    .A1(net910));
 sg13g2_nand4_1 _18396_ (.B(_11533_),
    .C(_11534_),
    .A(_11531_),
    .Y(_11536_),
    .D(_11535_));
 sg13g2_buf_1 _18397_ (.A(_11536_),
    .X(_11537_));
 sg13g2_and2_1 _18398_ (.A(_11529_),
    .B(net300),
    .X(_11538_));
 sg13g2_buf_1 _18399_ (.A(_11538_),
    .X(_11539_));
 sg13g2_mux2_1 _18400_ (.A0(_10434_),
    .A1(_11159_),
    .S(_10838_),
    .X(_11540_));
 sg13g2_buf_2 _18401_ (.A(_11540_),
    .X(_11541_));
 sg13g2_nand2_1 _18402_ (.Y(_11542_),
    .A(_10437_),
    .B(_11541_));
 sg13g2_nor2_1 _18403_ (.A(_11493_),
    .B(net257),
    .Y(_11543_));
 sg13g2_nand2b_1 _18404_ (.Y(_11544_),
    .B(net1127),
    .A_N(_10507_));
 sg13g2_a21oi_1 _18405_ (.A1(net439),
    .A2(net438),
    .Y(_11545_),
    .B1(_11544_));
 sg13g2_and4_1 _18406_ (.A(net439),
    .B(net438),
    .C(_10623_),
    .D(_11100_),
    .X(_11546_));
 sg13g2_a21oi_1 _18407_ (.A1(_08300_),
    .A2(_10621_),
    .Y(_11547_),
    .B1(_10507_));
 sg13g2_mux2_1 _18408_ (.A0(_11100_),
    .A1(_11547_),
    .S(net1127),
    .X(_11548_));
 sg13g2_nor3_2 _18409_ (.A(_11545_),
    .B(_11546_),
    .C(_11548_),
    .Y(_11549_));
 sg13g2_nor2_1 _18410_ (.A(_10511_),
    .B(_11549_),
    .Y(_11550_));
 sg13g2_buf_8 _18411_ (.A(_11549_),
    .X(_11551_));
 sg13g2_nand2_1 _18412_ (.Y(_11552_),
    .A(_10511_),
    .B(net256));
 sg13g2_o21ai_1 _18413_ (.B1(_11552_),
    .Y(_11553_),
    .A1(_11543_),
    .A2(_11550_));
 sg13g2_nand3b_1 _18414_ (.B(_11542_),
    .C(_11553_),
    .Y(_11554_),
    .A_N(_11539_));
 sg13g2_nor2_1 _18415_ (.A(net778),
    .B(_00289_),
    .Y(_11555_));
 sg13g2_nor2_1 _18416_ (.A(_09164_),
    .B(net559),
    .Y(_11556_));
 sg13g2_nor2_1 _18417_ (.A(net558),
    .B(_11158_),
    .Y(_11557_));
 sg13g2_nor4_1 _18418_ (.A(_09108_),
    .B(net437),
    .C(_11556_),
    .D(_11557_),
    .Y(_11558_));
 sg13g2_nor3_1 _18419_ (.A(net1038),
    .B(_11556_),
    .C(_11557_),
    .Y(_11559_));
 sg13g2_a221oi_1 _18420_ (.B2(net358),
    .C1(_11559_),
    .B1(_11558_),
    .A1(_10729_),
    .Y(_11560_),
    .A2(_11555_));
 sg13g2_buf_1 _18421_ (.A(_11560_),
    .X(_11561_));
 sg13g2_nand2_1 _18422_ (.Y(_11562_),
    .A(_10447_),
    .B(_11561_));
 sg13g2_nor4_1 _18423_ (.A(net232),
    .B(_11545_),
    .C(_11546_),
    .D(_11548_),
    .Y(_11563_));
 sg13g2_o21ai_1 _18424_ (.B1(_11563_),
    .Y(_11564_),
    .A1(net260),
    .A2(_11561_));
 sg13g2_a21oi_1 _18425_ (.A1(_11562_),
    .A2(_11564_),
    .Y(_11565_),
    .B1(_11539_));
 sg13g2_inv_1 _18426_ (.Y(_11566_),
    .A(_11565_));
 sg13g2_o21ai_1 _18427_ (.B1(_11566_),
    .Y(_11567_),
    .A1(_11527_),
    .A2(_11554_));
 sg13g2_buf_1 _18428_ (.A(_11567_),
    .X(_11568_));
 sg13g2_nor2_2 _18429_ (.A(_11529_),
    .B(net300),
    .Y(_11569_));
 sg13g2_nor2_1 _18430_ (.A(_10364_),
    .B(_11529_),
    .Y(_11570_));
 sg13g2_inv_1 _18431_ (.Y(_11571_),
    .A(net300));
 sg13g2_and2_1 _18432_ (.A(_10927_),
    .B(_10311_),
    .X(_11572_));
 sg13g2_a221oi_1 _18433_ (.B2(_11571_),
    .C1(_11572_),
    .B1(_11570_),
    .A1(_10927_),
    .Y(_11573_),
    .A2(_11569_));
 sg13g2_nand2_1 _18434_ (.Y(_11574_),
    .A(_10900_),
    .B(_10282_));
 sg13g2_o21ai_1 _18435_ (.B1(_11574_),
    .Y(_11575_),
    .A1(_11473_),
    .A2(_11573_));
 sg13g2_a21oi_2 _18436_ (.B1(_11575_),
    .Y(_11576_),
    .A2(_11568_),
    .A1(_11474_));
 sg13g2_nor2_1 _18437_ (.A(_10355_),
    .B(_11402_),
    .Y(_11577_));
 sg13g2_inv_1 _18438_ (.Y(_11578_),
    .A(_11577_));
 sg13g2_nand2b_1 _18439_ (.Y(_11579_),
    .B(_10369_),
    .A_N(net204));
 sg13g2_buf_1 _18440_ (.A(_10371_),
    .X(_11580_));
 sg13g2_and2_1 _18441_ (.A(_11580_),
    .B(_11474_),
    .X(_11581_));
 sg13g2_nor2_1 _18442_ (.A(_11527_),
    .B(_11554_),
    .Y(_11582_));
 sg13g2_a21o_1 _18443_ (.A2(_11565_),
    .A1(_11474_),
    .B1(_11575_),
    .X(_11583_));
 sg13g2_and2_1 _18444_ (.A(_10929_),
    .B(_10951_),
    .X(_11584_));
 sg13g2_buf_2 _18445_ (.A(_11584_),
    .X(_11585_));
 sg13g2_a221oi_1 _18446_ (.B2(net255),
    .C1(_11585_),
    .B1(_11583_),
    .A1(_11581_),
    .Y(_11586_),
    .A2(_11582_));
 sg13g2_buf_1 _18447_ (.A(_11586_),
    .X(_11587_));
 sg13g2_a221oi_1 _18448_ (.B2(_11579_),
    .C1(_11587_),
    .B1(_11578_),
    .A1(net230),
    .Y(_11588_),
    .A2(_11576_));
 sg13g2_and3_1 _18449_ (.X(_11589_),
    .A(_10865_),
    .B(_10867_),
    .C(_10870_));
 sg13g2_buf_1 _18450_ (.A(_11589_),
    .X(_11590_));
 sg13g2_nand2_1 _18451_ (.Y(_11591_),
    .A(net299),
    .B(net181));
 sg13g2_nand2b_1 _18452_ (.Y(_11592_),
    .B(net299),
    .A_N(net204));
 sg13g2_a221oi_1 _18453_ (.B2(_11592_),
    .C1(_11587_),
    .B1(_11591_),
    .A1(_11245_),
    .Y(_11593_),
    .A2(_11576_));
 sg13g2_buf_1 _18454_ (.A(_10355_),
    .X(_11594_));
 sg13g2_a21oi_1 _18455_ (.A1(_11591_),
    .A2(_11592_),
    .Y(_11595_),
    .B1(net201));
 sg13g2_or4_1 _18456_ (.A(_11469_),
    .B(_11588_),
    .C(_11593_),
    .D(_11595_),
    .X(_11596_));
 sg13g2_buf_8 _18457_ (.A(_11596_),
    .X(_11597_));
 sg13g2_and2_1 _18458_ (.A(_10806_),
    .B(_10808_),
    .X(_11598_));
 sg13g2_nand2_1 _18459_ (.Y(_11599_),
    .A(_10838_),
    .B(_11598_));
 sg13g2_o21ai_1 _18460_ (.B1(_11599_),
    .Y(_11600_),
    .A1(_10777_),
    .A2(_10838_));
 sg13g2_buf_1 _18461_ (.A(_11600_),
    .X(_11601_));
 sg13g2_buf_1 _18462_ (.A(_11601_),
    .X(_11602_));
 sg13g2_nand2_2 _18463_ (.Y(_11603_),
    .A(net149),
    .B(_11328_));
 sg13g2_buf_1 _18464_ (.A(net149),
    .X(_11604_));
 sg13g2_nor2_2 _18465_ (.A(net109),
    .B(_11328_),
    .Y(_11605_));
 sg13g2_a21oi_2 _18466_ (.B1(_11605_),
    .Y(_11606_),
    .A2(_11603_),
    .A1(_11597_));
 sg13g2_nand4_1 _18467_ (.B(_11462_),
    .C(_11463_),
    .A(net179),
    .Y(_11607_),
    .D(_11606_));
 sg13g2_a21oi_1 _18468_ (.A1(_08417_),
    .A2(_10715_),
    .Y(_11608_),
    .B1(_10716_));
 sg13g2_o21ai_1 _18469_ (.B1(_11608_),
    .Y(_11609_),
    .A1(_00193_),
    .A2(_10838_));
 sg13g2_buf_1 _18470_ (.A(_11609_),
    .X(_11610_));
 sg13g2_buf_1 _18471_ (.A(_11610_),
    .X(_11611_));
 sg13g2_buf_1 _18472_ (.A(net176),
    .X(_11612_));
 sg13g2_and3_1 _18473_ (.X(_11613_),
    .A(net148),
    .B(_11462_),
    .C(_11463_));
 sg13g2_o21ai_1 _18474_ (.B1(_11613_),
    .Y(_11614_),
    .A1(net179),
    .A2(_11606_));
 sg13g2_nand4_1 _18475_ (.B(_11459_),
    .C(_11607_),
    .A(_11448_),
    .Y(_11615_),
    .D(_11614_));
 sg13g2_buf_1 _18476_ (.A(_11615_),
    .X(\cpu.ex.c_mult[0] ));
 sg13g2_buf_1 _18477_ (.A(\cpu.dec.load ),
    .X(_11616_));
 sg13g2_nand2_2 _18478_ (.Y(_11617_),
    .A(net1164),
    .B(_08419_));
 sg13g2_nor2_1 _18479_ (.A(\cpu.ex.c_div_running ),
    .B(\cpu.ex.c_mult_running ),
    .Y(_11618_));
 sg13g2_buf_1 _18480_ (.A(_00250_),
    .X(_11619_));
 sg13g2_nand2_1 _18481_ (.Y(_11620_),
    .A(net1038),
    .B(\cpu.cond[2] ));
 sg13g2_a21o_1 _18482_ (.A2(_11620_),
    .A1(_11619_),
    .B1(_08375_),
    .X(_11621_));
 sg13g2_buf_1 _18483_ (.A(_11621_),
    .X(_11622_));
 sg13g2_or2_1 _18484_ (.X(_11623_),
    .B(\cpu.dec.jmp ),
    .A(net1038));
 sg13g2_nand2_1 _18485_ (.Y(_11624_),
    .A(net1161),
    .B(net814));
 sg13g2_a221oi_1 _18486_ (.B2(_11623_),
    .C1(_11624_),
    .B1(_11622_),
    .A1(_10994_),
    .Y(_11625_),
    .A2(\cpu.dec.r_swapsp ));
 sg13g2_nor2_2 _18487_ (.A(_09272_),
    .B(_09293_),
    .Y(_11626_));
 sg13g2_nand2b_1 _18488_ (.Y(_11627_),
    .B(net1071),
    .A_N(_09287_));
 sg13g2_nor2b_1 _18489_ (.A(_11626_),
    .B_N(_11627_),
    .Y(_11628_));
 sg13g2_buf_1 _18490_ (.A(_11628_),
    .X(_11629_));
 sg13g2_a21oi_1 _18491_ (.A1(_11618_),
    .A2(_11625_),
    .Y(_11630_),
    .B1(_11629_));
 sg13g2_a21oi_1 _18492_ (.A1(_11617_),
    .A2(_11630_),
    .Y(_11631_),
    .B1(_09257_));
 sg13g2_buf_1 _18493_ (.A(_11631_),
    .X(_11632_));
 sg13g2_nand2_1 _18494_ (.Y(_11633_),
    .A(_00291_),
    .B(net175));
 sg13g2_and2_1 _18495_ (.A(_09740_),
    .B(_09742_),
    .X(_11634_));
 sg13g2_nor2_1 _18496_ (.A(_09747_),
    .B(_11634_),
    .Y(_11635_));
 sg13g2_nor2_2 _18497_ (.A(_08383_),
    .B(_11635_),
    .Y(_11636_));
 sg13g2_inv_1 _18498_ (.Y(_11637_),
    .A(_11636_));
 sg13g2_o21ai_1 _18499_ (.B1(_11633_),
    .Y(_11638_),
    .A1(net175),
    .A2(_11637_));
 sg13g2_nand2_1 _18500_ (.Y(_11639_),
    .A(net1081),
    .B(_11638_));
 sg13g2_o21ai_1 _18501_ (.B1(_11639_),
    .Y(_00054_),
    .A1(_11616_),
    .A2(_11633_));
 sg13g2_buf_1 _18502_ (.A(\cpu.ex.r_mult[1] ),
    .X(_11640_));
 sg13g2_inv_1 _18503_ (.Y(_11641_),
    .A(_11640_));
 sg13g2_or3_1 _18504_ (.A(_10841_),
    .B(_10958_),
    .C(_11164_),
    .X(_11642_));
 sg13g2_buf_2 _18505_ (.A(_11642_),
    .X(_11643_));
 sg13g2_buf_1 _18506_ (.A(_11643_),
    .X(_11644_));
 sg13g2_buf_1 _18507_ (.A(_11419_),
    .X(_11645_));
 sg13g2_nand2_1 _18508_ (.Y(_11646_),
    .A(net90),
    .B(net200));
 sg13g2_buf_1 _18509_ (.A(_00091_),
    .X(_11647_));
 sg13g2_nor2_1 _18510_ (.A(_11647_),
    .B(net488),
    .Y(_11648_));
 sg13g2_xnor2_1 _18511_ (.Y(_11649_),
    .A(_11646_),
    .B(_11648_));
 sg13g2_or2_1 _18512_ (.X(_11650_),
    .B(_11425_),
    .A(_11647_));
 sg13g2_and2_1 _18513_ (.A(net646),
    .B(_11626_),
    .X(_11651_));
 sg13g2_buf_1 _18514_ (.A(_11651_),
    .X(_11652_));
 sg13g2_buf_1 _18515_ (.A(_11652_),
    .X(_11653_));
 sg13g2_nand2_1 _18516_ (.Y(_11654_),
    .A(_11429_),
    .B(_11433_));
 sg13g2_buf_1 _18517_ (.A(_11654_),
    .X(_11655_));
 sg13g2_a221oi_1 _18518_ (.B2(_00092_),
    .C1(_11655_),
    .B1(net436),
    .A1(_10129_),
    .Y(_11656_),
    .A2(_11650_));
 sg13g2_o21ai_1 _18519_ (.B1(_11656_),
    .Y(_11657_),
    .A1(_11445_),
    .A2(_11649_));
 sg13g2_o21ai_1 _18520_ (.B1(_11657_),
    .Y(\cpu.ex.c_mult[1] ),
    .A1(_11641_),
    .A2(_11433_));
 sg13g2_buf_1 _18521_ (.A(net645),
    .X(_11658_));
 sg13g2_buf_1 _18522_ (.A(_11658_),
    .X(_11659_));
 sg13g2_buf_1 _18523_ (.A(net487),
    .X(_11660_));
 sg13g2_buf_1 _18524_ (.A(_09293_),
    .X(_11661_));
 sg13g2_buf_8 _18525_ (.A(_10555_),
    .X(_11662_));
 sg13g2_buf_1 _18526_ (.A(net254),
    .X(_11663_));
 sg13g2_nor2_1 _18527_ (.A(_11647_),
    .B(_10275_),
    .Y(_11664_));
 sg13g2_nand2_1 _18528_ (.Y(_11665_),
    .A(_10589_),
    .B(_10279_));
 sg13g2_a21oi_1 _18529_ (.A1(_10565_),
    .A2(_11665_),
    .Y(_11666_),
    .B1(_11647_));
 sg13g2_a21o_1 _18530_ (.A2(_11664_),
    .A1(_10588_),
    .B1(_11666_),
    .X(_11667_));
 sg13g2_buf_1 _18531_ (.A(_11667_),
    .X(_11668_));
 sg13g2_xnor2_1 _18532_ (.Y(_11669_),
    .A(net226),
    .B(_11668_));
 sg13g2_o21ai_1 _18533_ (.B1(_11640_),
    .Y(_11670_),
    .A1(net110),
    .A2(_11669_));
 sg13g2_nand2_1 _18534_ (.Y(_11671_),
    .A(net1034),
    .B(_11670_));
 sg13g2_or2_1 _18535_ (.X(_11672_),
    .B(_11668_),
    .A(net259));
 sg13g2_nand3_1 _18536_ (.B(net259),
    .C(_11668_),
    .A(net487),
    .Y(_11673_));
 sg13g2_a21oi_1 _18537_ (.A1(_11672_),
    .A2(_11673_),
    .Y(_11674_),
    .B1(_11640_));
 sg13g2_a21o_1 _18538_ (.A2(net226),
    .A1(net488),
    .B1(_11674_),
    .X(_11675_));
 sg13g2_buf_1 _18539_ (.A(net90),
    .X(_11676_));
 sg13g2_a22oi_1 _18540_ (.Y(_11677_),
    .B1(_11675_),
    .B2(net82),
    .A2(_11671_),
    .A1(net435));
 sg13g2_o21ai_1 _18541_ (.B1(net386),
    .Y(_11678_),
    .A1(_00092_),
    .A2(net74));
 sg13g2_a21oi_1 _18542_ (.A1(_00103_),
    .A2(_11652_),
    .Y(_11679_),
    .B1(net555));
 sg13g2_nand2_1 _18543_ (.Y(_11680_),
    .A(_11678_),
    .B(_11679_));
 sg13g2_buf_1 _18544_ (.A(\cpu.ex.r_mult[2] ),
    .X(_11681_));
 sg13g2_nand2_1 _18545_ (.Y(_11682_),
    .A(_11681_),
    .B(net556));
 sg13g2_o21ai_1 _18546_ (.B1(_11682_),
    .Y(\cpu.ex.c_mult[2] ),
    .A1(_11677_),
    .A2(_11680_));
 sg13g2_buf_1 _18547_ (.A(\cpu.ex.r_mult[3] ),
    .X(_11683_));
 sg13g2_buf_1 _18548_ (.A(net231),
    .X(_11684_));
 sg13g2_nand2_1 _18549_ (.Y(_11685_),
    .A(_11640_),
    .B(net254));
 sg13g2_buf_2 _18550_ (.A(_11685_),
    .X(_11686_));
 sg13g2_o21ai_1 _18551_ (.B1(_11668_),
    .Y(_11687_),
    .A1(_11640_),
    .A2(net254));
 sg13g2_buf_1 _18552_ (.A(_11687_),
    .X(_11688_));
 sg13g2_a21o_1 _18553_ (.A2(_11688_),
    .A1(_11686_),
    .B1(_11443_),
    .X(_11689_));
 sg13g2_nand3_1 _18554_ (.B(_11686_),
    .C(_11688_),
    .A(_11684_),
    .Y(_11690_));
 sg13g2_o21ai_1 _18555_ (.B1(_11690_),
    .Y(_11691_),
    .A1(net199),
    .A2(_11689_));
 sg13g2_inv_1 _18556_ (.Y(_11692_),
    .A(_11681_));
 sg13g2_a22oi_1 _18557_ (.Y(_11693_),
    .B1(_11691_),
    .B2(_11692_),
    .A2(net199),
    .A1(net488));
 sg13g2_buf_1 _18558_ (.A(_11415_),
    .X(_11694_));
 sg13g2_a21oi_1 _18559_ (.A1(_11686_),
    .A2(_11688_),
    .Y(_11695_),
    .B1(net225));
 sg13g2_nand3_1 _18560_ (.B(_11686_),
    .C(_11688_),
    .A(net225),
    .Y(_11696_));
 sg13g2_nand2b_1 _18561_ (.Y(_11697_),
    .B(_11696_),
    .A_N(_11695_));
 sg13g2_o21ai_1 _18562_ (.B1(_11681_),
    .Y(_11698_),
    .A1(net110),
    .A2(_11697_));
 sg13g2_a21o_1 _18563_ (.A2(_11698_),
    .A1(net1034),
    .B1(net488),
    .X(_11699_));
 sg13g2_o21ai_1 _18564_ (.B1(_11699_),
    .Y(_11700_),
    .A1(net91),
    .A2(_11693_));
 sg13g2_or2_1 _18565_ (.X(_11701_),
    .B(_11425_),
    .A(_00103_));
 sg13g2_a221oi_1 _18566_ (.B2(net386),
    .C1(net555),
    .B1(_11701_),
    .A1(_00113_),
    .Y(_11702_),
    .A2(net436));
 sg13g2_a22oi_1 _18567_ (.Y(_11703_),
    .B1(_11700_),
    .B2(_11702_),
    .A2(net556),
    .A1(_11683_));
 sg13g2_inv_1 _18568_ (.Y(\cpu.ex.c_mult[3] ),
    .A(_11703_));
 sg13g2_buf_1 _18569_ (.A(net303),
    .X(_11704_));
 sg13g2_a21oi_1 _18570_ (.A1(_11681_),
    .A2(_11696_),
    .Y(_11705_),
    .B1(_11695_));
 sg13g2_xnor2_1 _18571_ (.Y(_11706_),
    .A(net253),
    .B(_11705_));
 sg13g2_nand2_1 _18572_ (.Y(_11707_),
    .A(net82),
    .B(_11706_));
 sg13g2_inv_1 _18573_ (.Y(_11708_),
    .A(_11683_));
 sg13g2_nor2_1 _18574_ (.A(_11708_),
    .B(net488),
    .Y(_11709_));
 sg13g2_nor3_1 _18575_ (.A(_11443_),
    .B(net303),
    .C(_11705_),
    .Y(_11710_));
 sg13g2_a21oi_1 _18576_ (.A1(net253),
    .A2(_11705_),
    .Y(_11711_),
    .B1(_11710_));
 sg13g2_nand2_1 _18577_ (.Y(_11712_),
    .A(net488),
    .B(net253));
 sg13g2_o21ai_1 _18578_ (.B1(_11712_),
    .Y(_11713_),
    .A1(_11683_),
    .A2(_11711_));
 sg13g2_a221oi_1 _18579_ (.B2(net82),
    .C1(_11445_),
    .B1(_11713_),
    .A1(_11707_),
    .Y(_11714_),
    .A2(_11709_));
 sg13g2_o21ai_1 _18580_ (.B1(net386),
    .Y(_11715_),
    .A1(_00113_),
    .A2(_11425_));
 sg13g2_a21oi_1 _18581_ (.A1(_00120_),
    .A2(_11652_),
    .Y(_11716_),
    .B1(_11654_));
 sg13g2_nand2_1 _18582_ (.Y(_11717_),
    .A(_11715_),
    .B(_11716_));
 sg13g2_buf_1 _18583_ (.A(\cpu.ex.r_mult[4] ),
    .X(_11718_));
 sg13g2_nand2_1 _18584_ (.Y(_11719_),
    .A(_11718_),
    .B(_11452_));
 sg13g2_o21ai_1 _18585_ (.B1(_11719_),
    .Y(\cpu.ex.c_mult[4] ),
    .A1(_11714_),
    .A2(_11717_));
 sg13g2_buf_1 _18586_ (.A(\cpu.ex.r_mult[5] ),
    .X(_11720_));
 sg13g2_buf_1 _18587_ (.A(net488),
    .X(_11721_));
 sg13g2_buf_1 _18588_ (.A(_10511_),
    .X(_11722_));
 sg13g2_nand2_1 _18589_ (.Y(_11723_),
    .A(net645),
    .B(_11225_));
 sg13g2_a221oi_1 _18590_ (.B2(_11688_),
    .C1(_11723_),
    .B1(_11686_),
    .A1(_11708_),
    .Y(_11724_),
    .A2(_11493_));
 sg13g2_nand2_1 _18591_ (.Y(_11725_),
    .A(_11681_),
    .B(_09295_));
 sg13g2_a221oi_1 _18592_ (.B2(_11688_),
    .C1(_11725_),
    .B1(_11686_),
    .A1(_11708_),
    .Y(_11726_),
    .A2(_11493_));
 sg13g2_nor2_1 _18593_ (.A(_11683_),
    .B(_10481_),
    .Y(_11727_));
 sg13g2_nand2_1 _18594_ (.Y(_11728_),
    .A(_11681_),
    .B(_11225_));
 sg13g2_nand2_1 _18595_ (.Y(_11729_),
    .A(_11683_),
    .B(net303));
 sg13g2_o21ai_1 _18596_ (.B1(_11729_),
    .Y(_11730_),
    .A1(_11727_),
    .A2(_11728_));
 sg13g2_or3_1 _18597_ (.A(_11724_),
    .B(_11726_),
    .C(_11730_),
    .X(_11731_));
 sg13g2_buf_1 _18598_ (.A(_11731_),
    .X(_11732_));
 sg13g2_nand3_1 _18599_ (.B(net224),
    .C(_11732_),
    .A(net487),
    .Y(_11733_));
 sg13g2_o21ai_1 _18600_ (.B1(_11733_),
    .Y(_11734_),
    .A1(net224),
    .A2(_11732_));
 sg13g2_inv_1 _18601_ (.Y(_11735_),
    .A(_11718_));
 sg13g2_a22oi_1 _18602_ (.Y(_11736_),
    .B1(_11734_),
    .B2(_11735_),
    .A2(net232),
    .A1(net434));
 sg13g2_xnor2_1 _18603_ (.Y(_11737_),
    .A(net224),
    .B(_11732_));
 sg13g2_a21oi_1 _18604_ (.A1(net82),
    .A2(_11737_),
    .Y(_11738_),
    .B1(_11735_));
 sg13g2_o21ai_1 _18605_ (.B1(net487),
    .Y(_11739_),
    .A1(_09294_),
    .A2(_11738_));
 sg13g2_o21ai_1 _18606_ (.B1(_11739_),
    .Y(_11740_),
    .A1(net91),
    .A2(_11736_));
 sg13g2_or2_1 _18607_ (.X(_11741_),
    .B(_11425_),
    .A(_00120_));
 sg13g2_a221oi_1 _18608_ (.B2(net348),
    .C1(net555),
    .B1(_11741_),
    .A1(_00132_),
    .Y(_11742_),
    .A2(net436));
 sg13g2_a22oi_1 _18609_ (.Y(_11743_),
    .B1(_11740_),
    .B2(_11742_),
    .A2(net556),
    .A1(net1122));
 sg13g2_inv_1 _18610_ (.Y(\cpu.ex.c_mult[5] ),
    .A(_11743_));
 sg13g2_buf_1 _18611_ (.A(\cpu.ex.r_mult[6] ),
    .X(_11744_));
 sg13g2_buf_1 _18612_ (.A(_11453_),
    .X(_11745_));
 sg13g2_or2_1 _18613_ (.X(_11746_),
    .B(net74),
    .A(_00132_));
 sg13g2_buf_1 _18614_ (.A(net555),
    .X(_11747_));
 sg13g2_a221oi_1 _18615_ (.B2(net348),
    .C1(net485),
    .B1(_11746_),
    .A1(_00144_),
    .Y(_11748_),
    .A2(_11653_));
 sg13g2_buf_1 _18616_ (.A(_10437_),
    .X(_11749_));
 sg13g2_nor3_2 _18617_ (.A(_11724_),
    .B(_11726_),
    .C(_11730_),
    .Y(_11750_));
 sg13g2_nand2_1 _18618_ (.Y(_11751_),
    .A(net224),
    .B(_11750_));
 sg13g2_o21ai_1 _18619_ (.B1(_11735_),
    .Y(_11752_),
    .A1(net224),
    .A2(_11750_));
 sg13g2_nand2_1 _18620_ (.Y(_11753_),
    .A(_11751_),
    .B(_11752_));
 sg13g2_xnor2_1 _18621_ (.Y(_11754_),
    .A(net252),
    .B(_11753_));
 sg13g2_inv_1 _18622_ (.Y(_11755_),
    .A(net1122));
 sg13g2_a21oi_1 _18623_ (.A1(net82),
    .A2(_11754_),
    .Y(_11756_),
    .B1(_11755_));
 sg13g2_o21ai_1 _18624_ (.B1(net435),
    .Y(_11757_),
    .A1(_09294_),
    .A2(_11756_));
 sg13g2_nand2_1 _18625_ (.Y(_11758_),
    .A(net487),
    .B(net260));
 sg13g2_mux2_1 _18626_ (.A0(_11758_),
    .A1(_10447_),
    .S(_11753_),
    .X(_11759_));
 sg13g2_nand2_1 _18627_ (.Y(_11760_),
    .A(net434),
    .B(_11749_));
 sg13g2_o21ai_1 _18628_ (.B1(_11760_),
    .Y(_11761_),
    .A1(net1122),
    .A2(_11759_));
 sg13g2_nand2_1 _18629_ (.Y(_11762_),
    .A(net82),
    .B(_11761_));
 sg13g2_nand2_1 _18630_ (.Y(_11763_),
    .A(_11757_),
    .B(_11762_));
 sg13g2_a22oi_1 _18631_ (.Y(_11764_),
    .B1(_11748_),
    .B2(_11763_),
    .A2(net486),
    .A1(_11744_));
 sg13g2_inv_1 _18632_ (.Y(\cpu.ex.c_mult[6] ),
    .A(_11764_));
 sg13g2_buf_2 _18633_ (.A(\cpu.ex.r_mult[7] ),
    .X(_11765_));
 sg13g2_or2_1 _18634_ (.X(_11766_),
    .B(_11425_),
    .A(_00144_));
 sg13g2_a221oi_1 _18635_ (.B2(net348),
    .C1(net485),
    .B1(_11766_),
    .A1(_00156_),
    .Y(_11767_),
    .A2(net436));
 sg13g2_and2_1 _18636_ (.A(_11744_),
    .B(net645),
    .X(_11768_));
 sg13g2_buf_1 _18637_ (.A(_11768_),
    .X(_11769_));
 sg13g2_nor2_1 _18638_ (.A(net1122),
    .B(_10437_),
    .Y(_11770_));
 sg13g2_a21oi_1 _18639_ (.A1(_11735_),
    .A2(net224),
    .Y(_11771_),
    .B1(_11770_));
 sg13g2_nand2_1 _18640_ (.Y(_11772_),
    .A(_11718_),
    .B(net232));
 sg13g2_nand2_1 _18641_ (.Y(_11773_),
    .A(net1122),
    .B(net252));
 sg13g2_o21ai_1 _18642_ (.B1(_11773_),
    .Y(_11774_),
    .A1(_11770_),
    .A2(_11772_));
 sg13g2_a21o_1 _18643_ (.A2(_11771_),
    .A1(_11732_),
    .B1(_11774_),
    .X(_11775_));
 sg13g2_buf_2 _18644_ (.A(_11529_),
    .X(_11776_));
 sg13g2_a21oi_1 _18645_ (.A1(net487),
    .A2(_11775_),
    .Y(_11777_),
    .B1(net223));
 sg13g2_a21oi_1 _18646_ (.A1(_11732_),
    .A2(_11771_),
    .Y(_11778_),
    .B1(_11774_));
 sg13g2_nor3_1 _18647_ (.A(_11444_),
    .B(_10444_),
    .C(_11778_),
    .Y(_11779_));
 sg13g2_nor3_1 _18648_ (.A(_11439_),
    .B(_11777_),
    .C(_11779_),
    .Y(_11780_));
 sg13g2_xnor2_1 _18649_ (.Y(_11781_),
    .A(_11769_),
    .B(_11780_));
 sg13g2_nand2_1 _18650_ (.Y(_11782_),
    .A(net492),
    .B(_11781_));
 sg13g2_a22oi_1 _18651_ (.Y(_11783_),
    .B1(_11767_),
    .B2(_11782_),
    .A2(net556),
    .A1(_11765_));
 sg13g2_inv_1 _18652_ (.Y(\cpu.ex.c_mult[7] ),
    .A(_11783_));
 sg13g2_buf_1 _18653_ (.A(\cpu.ex.r_mult[8] ),
    .X(_11784_));
 sg13g2_buf_1 _18654_ (.A(net436),
    .X(_11785_));
 sg13g2_or2_1 _18655_ (.X(_11786_),
    .B(net74),
    .A(_00156_));
 sg13g2_a221oi_1 _18656_ (.B2(net348),
    .C1(_11747_),
    .B1(_11786_),
    .A1(_00157_),
    .Y(_11787_),
    .A2(_11785_));
 sg13g2_nand2_1 _18657_ (.Y(_11788_),
    .A(net223),
    .B(_11769_));
 sg13g2_nor2_1 _18658_ (.A(net223),
    .B(_11769_),
    .Y(_11789_));
 sg13g2_nor3_1 _18659_ (.A(net626),
    .B(net260),
    .C(_11789_),
    .Y(_11790_));
 sg13g2_nand3_1 _18660_ (.B(_11752_),
    .C(_11790_),
    .A(_11751_),
    .Y(_11791_));
 sg13g2_nand4_1 _18661_ (.B(_09296_),
    .C(_10520_),
    .A(_11720_),
    .Y(_11792_),
    .D(net223));
 sg13g2_nand4_1 _18662_ (.B(\cpu.ex.r_mult[5] ),
    .C(net645),
    .A(_11718_),
    .Y(_11793_),
    .D(_11529_));
 sg13g2_a21oi_1 _18663_ (.A1(_11792_),
    .A2(_11793_),
    .Y(_11794_),
    .B1(_11750_));
 sg13g2_nand4_1 _18664_ (.B(net645),
    .C(net223),
    .A(net1122),
    .Y(_11795_),
    .D(_10437_));
 sg13g2_o21ai_1 _18665_ (.B1(_11795_),
    .Y(_11796_),
    .A1(net224),
    .A2(_11793_));
 sg13g2_nand3_1 _18666_ (.B(_10520_),
    .C(_11769_),
    .A(_11720_),
    .Y(_11797_));
 sg13g2_nand4_1 _18667_ (.B(net1122),
    .C(_11744_),
    .A(_11718_),
    .Y(_11798_),
    .D(net645));
 sg13g2_a21oi_1 _18668_ (.A1(_11797_),
    .A2(_11798_),
    .Y(_11799_),
    .B1(_11750_));
 sg13g2_nand3_1 _18669_ (.B(_10437_),
    .C(_11769_),
    .A(net1122),
    .Y(_11800_));
 sg13g2_o21ai_1 _18670_ (.B1(_11800_),
    .Y(_11801_),
    .A1(net224),
    .A2(_11798_));
 sg13g2_nor4_1 _18671_ (.A(_11794_),
    .B(_11796_),
    .C(_11799_),
    .D(_11801_),
    .Y(_11802_));
 sg13g2_nand3_1 _18672_ (.B(_11791_),
    .C(_11802_),
    .A(_11788_),
    .Y(_11803_));
 sg13g2_xnor2_1 _18673_ (.Y(_11804_),
    .A(net233),
    .B(_11803_));
 sg13g2_nor2_1 _18674_ (.A(net91),
    .B(_11804_),
    .Y(_11805_));
 sg13g2_inv_1 _18675_ (.Y(_11806_),
    .A(_11765_));
 sg13g2_nor2_1 _18676_ (.A(_11806_),
    .B(net434),
    .Y(_11807_));
 sg13g2_xnor2_1 _18677_ (.Y(_11808_),
    .A(_11805_),
    .B(_11807_));
 sg13g2_nand2_1 _18678_ (.Y(_11809_),
    .A(_09298_),
    .B(_11808_));
 sg13g2_a22oi_1 _18679_ (.Y(_11810_),
    .B1(_11787_),
    .B2(_11809_),
    .A2(_11745_),
    .A1(_11784_));
 sg13g2_inv_1 _18680_ (.Y(\cpu.ex.c_mult[8] ),
    .A(_11810_));
 sg13g2_and4_1 _18681_ (.A(_11744_),
    .B(_11765_),
    .C(_11658_),
    .D(_11775_),
    .X(_11811_));
 sg13g2_nor4_1 _18682_ (.A(net557),
    .B(net110),
    .C(net261),
    .D(_11778_),
    .Y(_11812_));
 sg13g2_o21ai_1 _18683_ (.B1(_11788_),
    .Y(_11813_),
    .A1(net557),
    .A2(_11247_));
 sg13g2_o21ai_1 _18684_ (.B1(_11765_),
    .Y(_11814_),
    .A1(_11812_),
    .A2(_11813_));
 sg13g2_or4_1 _18685_ (.A(net557),
    .B(_11437_),
    .C(_11778_),
    .D(_11789_),
    .X(_11815_));
 sg13g2_a21o_1 _18686_ (.A2(_11815_),
    .A1(_11788_),
    .B1(_11247_),
    .X(_11816_));
 sg13g2_nand3b_1 _18687_ (.B(_11814_),
    .C(_11816_),
    .Y(_11817_),
    .A_N(_11811_));
 sg13g2_xnor2_1 _18688_ (.Y(_11818_),
    .A(_11256_),
    .B(_11817_));
 sg13g2_inv_1 _18689_ (.Y(_11819_),
    .A(_11784_));
 sg13g2_nand2_1 _18690_ (.Y(_11820_),
    .A(net1034),
    .B(_11819_));
 sg13g2_buf_1 _18691_ (.A(\cpu.ex.r_mult[9] ),
    .X(_11821_));
 sg13g2_inv_1 _18692_ (.Y(_11822_),
    .A(_11821_));
 sg13g2_nor2_1 _18693_ (.A(_11822_),
    .B(_11433_),
    .Y(_11823_));
 sg13g2_a221oi_1 _18694_ (.B2(net435),
    .C1(_11823_),
    .B1(_11820_),
    .A1(net82),
    .Y(_11824_),
    .A2(_11818_));
 sg13g2_o21ai_1 _18695_ (.B1(net348),
    .Y(_11825_),
    .A1(_00157_),
    .A2(net74));
 sg13g2_a21oi_1 _18696_ (.A1(_00158_),
    .A2(net436),
    .Y(_11826_),
    .B1(net555));
 sg13g2_a21oi_1 _18697_ (.A1(_11825_),
    .A2(_11826_),
    .Y(_11827_),
    .B1(_11823_));
 sg13g2_nor2_1 _18698_ (.A(_09294_),
    .B(_11819_),
    .Y(_11828_));
 sg13g2_nor2_1 _18699_ (.A(net434),
    .B(_11823_),
    .Y(_11829_));
 sg13g2_and4_1 _18700_ (.A(net82),
    .B(_11818_),
    .C(_11828_),
    .D(_11829_),
    .X(_11830_));
 sg13g2_nor3_1 _18701_ (.A(_11824_),
    .B(_11827_),
    .C(_11830_),
    .Y(\cpu.ex.c_mult[9] ));
 sg13g2_buf_1 _18702_ (.A(\cpu.ex.r_mult[10] ),
    .X(_11831_));
 sg13g2_nand2_1 _18703_ (.Y(_11832_),
    .A(net1034),
    .B(_11822_));
 sg13g2_nor2_1 _18704_ (.A(net110),
    .B(net230),
    .Y(_11833_));
 sg13g2_nor2_1 _18705_ (.A(net110),
    .B(_11580_),
    .Y(_11834_));
 sg13g2_xnor2_1 _18706_ (.Y(_11835_),
    .A(_11784_),
    .B(_10282_));
 sg13g2_nor2_1 _18707_ (.A(_11806_),
    .B(_10364_),
    .Y(_11836_));
 sg13g2_nor4_1 _18708_ (.A(_11765_),
    .B(_11819_),
    .C(_10360_),
    .D(_10311_),
    .Y(_11837_));
 sg13g2_a21oi_1 _18709_ (.A1(_11835_),
    .A2(_11836_),
    .Y(_11838_),
    .B1(_11837_));
 sg13g2_o21ai_1 _18710_ (.B1(net645),
    .Y(_11839_),
    .A1(_11765_),
    .A2(_11784_));
 sg13g2_nand3_1 _18711_ (.B(net233),
    .C(_11839_),
    .A(_10360_),
    .Y(_11840_));
 sg13g2_o21ai_1 _18712_ (.B1(_11840_),
    .Y(_11841_),
    .A1(net626),
    .A2(_11838_));
 sg13g2_nand2_1 _18713_ (.Y(_11842_),
    .A(_11784_),
    .B(_10360_));
 sg13g2_nand2_1 _18714_ (.Y(_11843_),
    .A(_11819_),
    .B(_10282_));
 sg13g2_nand3_1 _18715_ (.B(net233),
    .C(_11843_),
    .A(_11765_),
    .Y(_11844_));
 sg13g2_a21oi_1 _18716_ (.A1(_11842_),
    .A2(_11844_),
    .Y(_11845_),
    .B1(net626));
 sg13g2_a21oi_1 _18717_ (.A1(_11803_),
    .A2(_11841_),
    .Y(_11846_),
    .B1(_11845_));
 sg13g2_mux2_1 _18718_ (.A0(_11833_),
    .A1(_11834_),
    .S(_11846_),
    .X(_11847_));
 sg13g2_a221oi_1 _18719_ (.B2(net435),
    .C1(_11847_),
    .B1(_11832_),
    .A1(_11831_),
    .Y(_11848_),
    .A2(_11452_));
 sg13g2_o21ai_1 _18720_ (.B1(net386),
    .Y(_11849_),
    .A1(_00158_),
    .A2(net74));
 sg13g2_a21oi_1 _18721_ (.A1(_00159_),
    .A2(_11653_),
    .Y(_11850_),
    .B1(net555));
 sg13g2_a22oi_1 _18722_ (.Y(_11851_),
    .B1(_11849_),
    .B2(_11850_),
    .A2(net556),
    .A1(_11831_));
 sg13g2_a21oi_1 _18723_ (.A1(net1121),
    .A2(_11452_),
    .Y(_11852_),
    .B1(_11721_));
 sg13g2_and4_1 _18724_ (.A(net1034),
    .B(_11821_),
    .C(_11847_),
    .D(_11852_),
    .X(_11853_));
 sg13g2_nor3_1 _18725_ (.A(_11848_),
    .B(_11851_),
    .C(_11853_),
    .Y(\cpu.ex.c_mult[10] ));
 sg13g2_or2_1 _18726_ (.X(_11854_),
    .B(_11425_),
    .A(_00159_));
 sg13g2_a221oi_1 _18727_ (.B2(net386),
    .C1(net555),
    .B1(_11854_),
    .A1(_00160_),
    .Y(_11855_),
    .A2(net436));
 sg13g2_inv_1 _18728_ (.Y(_11856_),
    .A(_11855_));
 sg13g2_nor2_1 _18729_ (.A(_11821_),
    .B(net230),
    .Y(_11857_));
 sg13g2_o21ai_1 _18730_ (.B1(_11821_),
    .Y(_11858_),
    .A1(_10137_),
    .A2(_10230_));
 sg13g2_buf_1 _18731_ (.A(_11858_),
    .X(_11859_));
 sg13g2_o21ai_1 _18732_ (.B1(_11859_),
    .Y(_11860_),
    .A1(_11842_),
    .A2(_11857_));
 sg13g2_a22oi_1 _18733_ (.Y(_11861_),
    .B1(_11860_),
    .B2(_11659_),
    .A2(_11811_),
    .A1(net90));
 sg13g2_nand3_1 _18734_ (.B(_11816_),
    .C(_11861_),
    .A(_11814_),
    .Y(_11862_));
 sg13g2_buf_1 _18735_ (.A(_11862_),
    .X(_11863_));
 sg13g2_nor2_1 _18736_ (.A(_11822_),
    .B(net557),
    .Y(_11864_));
 sg13g2_and2_1 _18737_ (.A(_11819_),
    .B(_11859_),
    .X(_11865_));
 sg13g2_o21ai_1 _18738_ (.B1(_11256_),
    .Y(_11866_),
    .A1(net557),
    .A2(_11865_));
 sg13g2_o21ai_1 _18739_ (.B1(_11866_),
    .Y(_11867_),
    .A1(net230),
    .A2(_11864_));
 sg13g2_nor2_1 _18740_ (.A(net110),
    .B(_11867_),
    .Y(_11868_));
 sg13g2_nand2_1 _18741_ (.Y(_11869_),
    .A(_11863_),
    .B(_11868_));
 sg13g2_nand2_1 _18742_ (.Y(_11870_),
    .A(net1121),
    .B(net487));
 sg13g2_nand2_1 _18743_ (.Y(_11871_),
    .A(_11676_),
    .B(net201));
 sg13g2_xnor2_1 _18744_ (.Y(_11872_),
    .A(_11870_),
    .B(_11871_));
 sg13g2_xnor2_1 _18745_ (.Y(_11873_),
    .A(_11869_),
    .B(_11872_));
 sg13g2_buf_1 _18746_ (.A(\cpu.ex.r_mult[11] ),
    .X(_11874_));
 sg13g2_a22oi_1 _18747_ (.Y(_11875_),
    .B1(_11855_),
    .B2(_11445_),
    .A2(net556),
    .A1(_11874_));
 sg13g2_o21ai_1 _18748_ (.B1(_11875_),
    .Y(\cpu.ex.c_mult[11] ),
    .A1(_11856_),
    .A2(_11873_));
 sg13g2_or2_1 _18749_ (.X(_11876_),
    .B(_11426_),
    .A(_00160_));
 sg13g2_a221oi_1 _18750_ (.B2(_10130_),
    .C1(_11747_),
    .B1(_11876_),
    .A1(_00161_),
    .Y(_11877_),
    .A2(_11785_));
 sg13g2_nand2_1 _18751_ (.Y(_11878_),
    .A(net554),
    .B(_11643_));
 sg13g2_buf_1 _18752_ (.A(_11878_),
    .X(_11879_));
 sg13g2_nor3_1 _18753_ (.A(net1121),
    .B(_10320_),
    .C(_10353_),
    .Y(_11880_));
 sg13g2_o21ai_1 _18754_ (.B1(net1121),
    .Y(_11881_),
    .A1(_10320_),
    .A2(_10353_));
 sg13g2_buf_1 _18755_ (.A(_11881_),
    .X(_11882_));
 sg13g2_o21ai_1 _18756_ (.B1(_11882_),
    .Y(_11883_),
    .A1(_11859_),
    .A2(_11880_));
 sg13g2_buf_1 _18757_ (.A(_11883_),
    .X(_11884_));
 sg13g2_nor2_1 _18758_ (.A(net1120),
    .B(net177),
    .Y(_11885_));
 sg13g2_or2_1 _18759_ (.X(_11886_),
    .B(_10355_),
    .A(net1121));
 sg13g2_nand4_1 _18760_ (.B(_10371_),
    .C(_11886_),
    .A(_11821_),
    .Y(_11887_),
    .D(_11882_));
 sg13g2_nand4_1 _18761_ (.B(net1121),
    .C(_10369_),
    .A(_11822_),
    .Y(_11888_),
    .D(_10232_));
 sg13g2_a21oi_1 _18762_ (.A1(_11887_),
    .A2(_11888_),
    .Y(_11889_),
    .B1(net626));
 sg13g2_o21ai_1 _18763_ (.B1(net554),
    .Y(_11890_),
    .A1(_11821_),
    .A2(net1121));
 sg13g2_and3_1 _18764_ (.X(_11891_),
    .A(_10355_),
    .B(_10232_),
    .C(_11890_));
 sg13g2_o21ai_1 _18765_ (.B1(_11643_),
    .Y(_11892_),
    .A1(_11889_),
    .A2(_11891_));
 sg13g2_nor2_1 _18766_ (.A(_11841_),
    .B(_11845_),
    .Y(_11893_));
 sg13g2_nor2_1 _18767_ (.A(_11892_),
    .B(_11893_),
    .Y(_11894_));
 sg13g2_inv_1 _18768_ (.Y(_11895_),
    .A(_11845_));
 sg13g2_nand4_1 _18769_ (.B(_11791_),
    .C(_11802_),
    .A(_11788_),
    .Y(_11896_),
    .D(_11895_));
 sg13g2_and2_1 _18770_ (.A(_11894_),
    .B(_11896_),
    .X(_11897_));
 sg13g2_buf_1 _18771_ (.A(_11897_),
    .X(_11898_));
 sg13g2_or2_1 _18772_ (.X(_11899_),
    .B(_11898_),
    .A(_11884_));
 sg13g2_inv_1 _18773_ (.Y(_11900_),
    .A(net1120));
 sg13g2_nor2_1 _18774_ (.A(_11900_),
    .B(net181),
    .Y(_11901_));
 sg13g2_a22oi_1 _18775_ (.Y(_11902_),
    .B1(_11899_),
    .B2(_11901_),
    .A2(_11885_),
    .A1(_11884_));
 sg13g2_nor2_1 _18776_ (.A(net91),
    .B(net150),
    .Y(_11903_));
 sg13g2_nand2_1 _18777_ (.Y(_11904_),
    .A(net1120),
    .B(net554));
 sg13g2_nor2b_1 _18778_ (.A(_11903_),
    .B_N(_11904_),
    .Y(_11905_));
 sg13g2_o21ai_1 _18779_ (.B1(net487),
    .Y(_11906_),
    .A1(net1120),
    .A2(_11884_));
 sg13g2_nand2_1 _18780_ (.Y(_11907_),
    .A(_11859_),
    .B(_11882_));
 sg13g2_nand2_1 _18781_ (.Y(_11908_),
    .A(_11886_),
    .B(_11907_));
 sg13g2_nand2_1 _18782_ (.Y(_11909_),
    .A(net150),
    .B(_11908_));
 sg13g2_a21oi_1 _18783_ (.A1(net90),
    .A2(_11909_),
    .Y(_11910_),
    .B1(_11904_));
 sg13g2_a21oi_1 _18784_ (.A1(_11906_),
    .A2(_11903_),
    .Y(_11911_),
    .B1(_11910_));
 sg13g2_nor2_1 _18785_ (.A(_11911_),
    .B(_11898_),
    .Y(_11912_));
 sg13g2_a221oi_1 _18786_ (.B2(_11905_),
    .C1(_11912_),
    .B1(_11898_),
    .A1(_09294_),
    .Y(_11913_),
    .A2(net435));
 sg13g2_o21ai_1 _18787_ (.B1(_11913_),
    .Y(_11914_),
    .A1(_11879_),
    .A2(_11902_));
 sg13g2_buf_2 _18788_ (.A(\cpu.ex.r_mult[12] ),
    .X(_11915_));
 sg13g2_inv_1 _18789_ (.Y(_11916_),
    .A(_11915_));
 sg13g2_nor2_1 _18790_ (.A(_11916_),
    .B(_11433_),
    .Y(_11917_));
 sg13g2_a21o_1 _18791_ (.A2(_11914_),
    .A1(_11877_),
    .B1(_11917_),
    .X(\cpu.ex.c_mult[12] ));
 sg13g2_a21oi_1 _18792_ (.A1(_11900_),
    .A2(net181),
    .Y(_11918_),
    .B1(_11882_));
 sg13g2_nor2_1 _18793_ (.A(_11901_),
    .B(_11918_),
    .Y(_11919_));
 sg13g2_o21ai_1 _18794_ (.B1(net207),
    .Y(_11920_),
    .A1(_11879_),
    .A2(_11919_));
 sg13g2_o21ai_1 _18795_ (.B1(net1120),
    .Y(_11921_),
    .A1(net110),
    .A2(_11577_));
 sg13g2_nand3_1 _18796_ (.B(_10369_),
    .C(_11402_),
    .A(_11900_),
    .Y(_11922_));
 sg13g2_a21oi_1 _18797_ (.A1(_11921_),
    .A2(_11922_),
    .Y(_11923_),
    .B1(_11870_));
 sg13g2_mux2_1 _18798_ (.A0(net1120),
    .A1(_11904_),
    .S(net181),
    .X(_11924_));
 sg13g2_nand2_1 _18799_ (.Y(_11925_),
    .A(net557),
    .B(_11402_));
 sg13g2_o21ai_1 _18800_ (.B1(_11925_),
    .Y(_11926_),
    .A1(net1121),
    .A2(_11924_));
 sg13g2_nand2_1 _18801_ (.Y(_11927_),
    .A(net201),
    .B(_11926_));
 sg13g2_inv_1 _18802_ (.Y(_11928_),
    .A(_11927_));
 sg13g2_nor3_1 _18803_ (.A(_11438_),
    .B(net207),
    .C(_11867_),
    .Y(_11929_));
 sg13g2_o21ai_1 _18804_ (.B1(_11929_),
    .Y(_11930_),
    .A1(_11923_),
    .A2(_11928_));
 sg13g2_mux2_1 _18805_ (.A0(_11920_),
    .A1(_11930_),
    .S(_11863_),
    .X(_11931_));
 sg13g2_nor3_1 _18806_ (.A(_11923_),
    .B(_11928_),
    .C(_11920_),
    .Y(_11932_));
 sg13g2_nor2_1 _18807_ (.A(_11879_),
    .B(_11919_),
    .Y(_11933_));
 sg13g2_nand2_1 _18808_ (.Y(_11934_),
    .A(net207),
    .B(_11867_));
 sg13g2_o21ai_1 _18809_ (.B1(_11676_),
    .Y(_11935_),
    .A1(_11933_),
    .A2(_11934_));
 sg13g2_nor4_1 _18810_ (.A(_11444_),
    .B(_11439_),
    .C(net207),
    .D(_11919_),
    .Y(_11936_));
 sg13g2_nor3_1 _18811_ (.A(_11932_),
    .B(_11935_),
    .C(_11936_),
    .Y(_11937_));
 sg13g2_buf_2 _18812_ (.A(\cpu.ex.r_mult[13] ),
    .X(_11938_));
 sg13g2_nand2_1 _18813_ (.Y(_11939_),
    .A(_11938_),
    .B(_11452_));
 sg13g2_nand2_1 _18814_ (.Y(_11940_),
    .A(_11721_),
    .B(_11939_));
 sg13g2_nand3_1 _18815_ (.B(_11916_),
    .C(_11939_),
    .A(_11661_),
    .Y(_11941_));
 sg13g2_a22oi_1 _18816_ (.Y(_11942_),
    .B1(_11940_),
    .B2(_11941_),
    .A2(_11937_),
    .A1(_11931_));
 sg13g2_nand2_1 _18817_ (.Y(_11943_),
    .A(_11931_),
    .B(_11937_));
 sg13g2_nand4_1 _18818_ (.B(_11915_),
    .C(_11660_),
    .A(_11661_),
    .Y(_11944_),
    .D(_11939_));
 sg13g2_o21ai_1 _18819_ (.B1(_10130_),
    .Y(_11945_),
    .A1(_00161_),
    .A2(_11426_));
 sg13g2_a21oi_1 _18820_ (.A1(_00162_),
    .A2(net436),
    .Y(_11946_),
    .B1(_11655_));
 sg13g2_nand2_1 _18821_ (.Y(_11947_),
    .A(_11945_),
    .B(_11946_));
 sg13g2_nand2_1 _18822_ (.Y(_11948_),
    .A(_11939_),
    .B(_11947_));
 sg13g2_o21ai_1 _18823_ (.B1(_11948_),
    .Y(_11949_),
    .A1(_11943_),
    .A2(_11944_));
 sg13g2_nor2_1 _18824_ (.A(_11942_),
    .B(_11949_),
    .Y(\cpu.ex.c_mult[13] ));
 sg13g2_o21ai_1 _18825_ (.B1(net386),
    .Y(_11950_),
    .A1(_00162_),
    .A2(_11425_));
 sg13g2_buf_1 _18826_ (.A(_00163_),
    .X(_11951_));
 sg13g2_a21oi_1 _18827_ (.A1(_11951_),
    .A2(_11652_),
    .Y(_11952_),
    .B1(_11654_));
 sg13g2_nand2_1 _18828_ (.Y(_11953_),
    .A(_11950_),
    .B(_11952_));
 sg13g2_nand2_1 _18829_ (.Y(_11954_),
    .A(_11938_),
    .B(net554));
 sg13g2_buf_1 _18830_ (.A(_11387_),
    .X(_11955_));
 sg13g2_nor2_1 _18831_ (.A(net91),
    .B(net147),
    .Y(_11956_));
 sg13g2_xnor2_1 _18832_ (.Y(_11957_),
    .A(_11954_),
    .B(_11956_));
 sg13g2_nor2b_1 _18833_ (.A(_11953_),
    .B_N(_11957_),
    .Y(_11958_));
 sg13g2_nor2_1 _18834_ (.A(_11953_),
    .B(_11957_),
    .Y(_11959_));
 sg13g2_nand2_1 _18835_ (.Y(_11960_),
    .A(net645),
    .B(_11320_));
 sg13g2_nand2_1 _18836_ (.Y(_11961_),
    .A(_11916_),
    .B(_11327_));
 sg13g2_o21ai_1 _18837_ (.B1(_11961_),
    .Y(_11962_),
    .A1(_11916_),
    .A2(_11960_));
 sg13g2_a22oi_1 _18838_ (.Y(_11963_),
    .B1(_11962_),
    .B2(_11900_),
    .A2(_11327_),
    .A1(_10954_));
 sg13g2_or4_1 _18839_ (.A(_11915_),
    .B(_11320_),
    .C(_11402_),
    .D(_11904_),
    .X(_11964_));
 sg13g2_o21ai_1 _18840_ (.B1(_11964_),
    .Y(_11965_),
    .A1(net181),
    .A2(_11963_));
 sg13g2_nand3_1 _18841_ (.B(_11915_),
    .C(net554),
    .A(net1120),
    .Y(_11966_));
 sg13g2_a21oi_1 _18842_ (.A1(_11643_),
    .A2(_11422_),
    .Y(_11967_),
    .B1(_11966_));
 sg13g2_a21o_1 _18843_ (.A2(_11965_),
    .A1(net90),
    .B1(_11967_),
    .X(_11968_));
 sg13g2_nand3_1 _18844_ (.B(_11896_),
    .C(_11968_),
    .A(_11894_),
    .Y(_11969_));
 sg13g2_o21ai_1 _18845_ (.B1(net1120),
    .Y(_11970_),
    .A1(_11402_),
    .A2(_11884_));
 sg13g2_o21ai_1 _18846_ (.B1(_11970_),
    .Y(_11971_),
    .A1(_11295_),
    .A2(_11908_));
 sg13g2_o21ai_1 _18847_ (.B1(_11971_),
    .Y(_11972_),
    .A1(_11915_),
    .A2(_11327_));
 sg13g2_nand2_1 _18848_ (.Y(_11973_),
    .A(_11915_),
    .B(net206));
 sg13g2_a21o_1 _18849_ (.A2(_11973_),
    .A1(_11972_),
    .B1(_11879_),
    .X(_11974_));
 sg13g2_nand2_1 _18850_ (.Y(_11975_),
    .A(_11969_),
    .B(_11974_));
 sg13g2_mux2_1 _18851_ (.A0(_11958_),
    .A1(_11959_),
    .S(_11975_),
    .X(_11976_));
 sg13g2_nand2_1 _18852_ (.Y(_11977_),
    .A(\cpu.ex.r_mult[14] ),
    .B(net556));
 sg13g2_o21ai_1 _18853_ (.B1(_11977_),
    .Y(_11978_),
    .A1(net492),
    .A2(_11953_));
 sg13g2_or2_1 _18854_ (.X(\cpu.ex.c_mult[14] ),
    .B(_11978_),
    .A(_11976_));
 sg13g2_nand2_1 _18855_ (.Y(_11979_),
    .A(net90),
    .B(net180));
 sg13g2_nor2_1 _18856_ (.A(_11951_),
    .B(net626),
    .Y(_11980_));
 sg13g2_xnor2_1 _18857_ (.Y(_11981_),
    .A(_11979_),
    .B(_11980_));
 sg13g2_nand2_1 _18858_ (.Y(_11982_),
    .A(net492),
    .B(_11981_));
 sg13g2_nand2b_1 _18859_ (.Y(_11983_),
    .B(net492),
    .A_N(_11981_));
 sg13g2_a21o_1 _18860_ (.A2(_11922_),
    .A1(_11921_),
    .B1(_11870_),
    .X(_11984_));
 sg13g2_nand2_1 _18861_ (.Y(_11985_),
    .A(net147),
    .B(net207));
 sg13g2_nand3_1 _18862_ (.B(_11938_),
    .C(_11659_),
    .A(_11915_),
    .Y(_11986_));
 sg13g2_a21oi_1 _18863_ (.A1(_11644_),
    .A2(_11985_),
    .Y(_11987_),
    .B1(_11986_));
 sg13g2_mux2_1 _18864_ (.A0(_11954_),
    .A1(_11938_),
    .S(_11386_),
    .X(_11988_));
 sg13g2_nand2_1 _18865_ (.Y(_11989_),
    .A(net557),
    .B(net179));
 sg13g2_o21ai_1 _18866_ (.B1(_11989_),
    .Y(_11990_),
    .A1(_11915_),
    .A2(_11988_));
 sg13g2_nor4_1 _18867_ (.A(_11916_),
    .B(_11938_),
    .C(net147),
    .D(_11960_),
    .Y(_11991_));
 sg13g2_a21oi_1 _18868_ (.A1(net206),
    .A2(_11990_),
    .Y(_11992_),
    .B1(_11991_));
 sg13g2_nor2_1 _18869_ (.A(_11438_),
    .B(_11992_),
    .Y(_11993_));
 sg13g2_o21ai_1 _18870_ (.B1(_11868_),
    .Y(_11994_),
    .A1(_11987_),
    .A2(_11993_));
 sg13g2_a21oi_1 _18871_ (.A1(_11984_),
    .A2(_11927_),
    .Y(_11995_),
    .B1(_11994_));
 sg13g2_inv_1 _18872_ (.Y(_11996_),
    .A(_11938_));
 sg13g2_nor3_1 _18873_ (.A(net179),
    .B(_11901_),
    .C(_11918_),
    .Y(_11997_));
 sg13g2_o21ai_1 _18874_ (.B1(_11916_),
    .Y(_11998_),
    .A1(_11996_),
    .A2(_11997_));
 sg13g2_nor3_1 _18875_ (.A(net206),
    .B(_11901_),
    .C(_11918_),
    .Y(_11999_));
 sg13g2_o21ai_1 _18876_ (.B1(_11996_),
    .Y(_12000_),
    .A1(net147),
    .A2(_11999_));
 sg13g2_nand3_1 _18877_ (.B(_11998_),
    .C(_12000_),
    .A(_11985_),
    .Y(_12001_));
 sg13g2_nand3_1 _18878_ (.B(net179),
    .C(net206),
    .A(_11644_),
    .Y(_12002_));
 sg13g2_a21o_1 _18879_ (.A2(_12002_),
    .A1(_11986_),
    .B1(_11919_),
    .X(_12003_));
 sg13g2_a21oi_1 _18880_ (.A1(_12001_),
    .A2(_12003_),
    .Y(_12004_),
    .B1(_11879_));
 sg13g2_a21oi_1 _18881_ (.A1(_11863_),
    .A2(_11995_),
    .Y(_12005_),
    .B1(_12004_));
 sg13g2_mux2_1 _18882_ (.A0(_11982_),
    .A1(_11983_),
    .S(_12005_),
    .X(_12006_));
 sg13g2_o21ai_1 _18883_ (.B1(net386),
    .Y(_12007_),
    .A1(_11951_),
    .A2(net74));
 sg13g2_nand2_1 _18884_ (.Y(_12008_),
    .A(_11435_),
    .B(_12007_));
 sg13g2_nor2_1 _18885_ (.A(net385),
    .B(_12008_),
    .Y(_12009_));
 sg13g2_a21oi_1 _18886_ (.A1(_12006_),
    .A2(_12009_),
    .Y(_12010_),
    .B1(\cpu.ex.r_mult[15] ));
 sg13g2_inv_1 _18887_ (.Y(_12011_),
    .A(_12008_));
 sg13g2_a21oi_1 _18888_ (.A1(_12006_),
    .A2(_12011_),
    .Y(_12012_),
    .B1(_11745_));
 sg13g2_nor2_1 _18889_ (.A(_12010_),
    .B(_12012_),
    .Y(\cpu.ex.c_mult[15] ));
 sg13g2_inv_1 _18890_ (.Y(_00000_),
    .A(net2));
 sg13g2_inv_1 _18891_ (.Y(_12013_),
    .A(_09779_));
 sg13g2_nor3_1 _18892_ (.A(_12013_),
    .B(net714),
    .C(_09778_),
    .Y(_00008_));
 sg13g2_buf_1 _18893_ (.A(net818),
    .X(_12014_));
 sg13g2_and3_1 _18894_ (.X(_00005_),
    .A(net1148),
    .B(net680),
    .C(_09768_));
 sg13g2_buf_2 _18895_ (.A(\cpu.qspi.r_state[3] ),
    .X(_12015_));
 sg13g2_and2_1 _18896_ (.A(_12015_),
    .B(net680),
    .X(_00009_));
 sg13g2_buf_1 _18897_ (.A(\cpu.qspi.r_state[11] ),
    .X(_12016_));
 sg13g2_inv_1 _18898_ (.Y(_12017_),
    .A(_12016_));
 sg13g2_nor2_1 _18899_ (.A(_12017_),
    .B(net647),
    .Y(_00004_));
 sg13g2_buf_2 _18900_ (.A(\cpu.qspi.r_state[10] ),
    .X(_12018_));
 sg13g2_and2_1 _18901_ (.A(_12018_),
    .B(net680),
    .X(_00003_));
 sg13g2_buf_1 _18902_ (.A(\cpu.qspi.r_state[15] ),
    .X(_12019_));
 sg13g2_and2_1 _18903_ (.A(_12019_),
    .B(_12014_),
    .X(_00002_));
 sg13g2_inv_1 _18904_ (.Y(_12020_),
    .A(net1149));
 sg13g2_nor3_1 _18905_ (.A(_12020_),
    .B(net714),
    .C(net799),
    .Y(_00001_));
 sg13g2_nand2b_1 _18906_ (.Y(_12021_),
    .B(_09805_),
    .A_N(_09803_));
 sg13g2_nor2_1 _18907_ (.A(net647),
    .B(_12021_),
    .Y(_00007_));
 sg13g2_nand2_1 _18908_ (.Y(_12022_),
    .A(\cpu.dec.iready ),
    .B(_00197_));
 sg13g2_nor2_1 _18909_ (.A(\cpu.ex.r_branch_stall ),
    .B(_12022_),
    .Y(_12023_));
 sg13g2_buf_2 _18910_ (.A(_12023_),
    .X(_12024_));
 sg13g2_nand2_1 _18911_ (.Y(_12025_),
    .A(_09105_),
    .B(_12024_));
 sg13g2_o21ai_1 _18912_ (.B1(_10923_),
    .Y(_12026_),
    .A1(_10711_),
    .A2(_10714_));
 sg13g2_or2_1 _18913_ (.X(_12027_),
    .B(_11142_),
    .A(_10868_));
 sg13g2_nand2_1 _18914_ (.Y(_12028_),
    .A(_10836_),
    .B(_10983_));
 sg13g2_or4_1 _18915_ (.A(_11159_),
    .B(_12026_),
    .C(_12027_),
    .D(_12028_),
    .X(_12029_));
 sg13g2_nor3_1 _18916_ (.A(_10893_),
    .B(_11100_),
    .C(_11121_),
    .Y(_12030_));
 sg13g2_nor2_1 _18917_ (.A(_11486_),
    .B(_11040_),
    .Y(_12031_));
 sg13g2_nand3_1 _18918_ (.B(_12030_),
    .C(_12031_),
    .A(_10950_),
    .Y(_12032_));
 sg13g2_nor4_1 _18919_ (.A(_11598_),
    .B(_11070_),
    .C(_12029_),
    .D(_12032_),
    .Y(_12033_));
 sg13g2_o21ai_1 _18920_ (.B1(_10769_),
    .Y(_12034_),
    .A1(\cpu.cond[1] ),
    .A2(_12033_));
 sg13g2_xnor2_1 _18921_ (.Y(_12035_),
    .A(_08375_),
    .B(_12034_));
 sg13g2_a21o_1 _18922_ (.A2(_12035_),
    .A1(_10609_),
    .B1(_10724_),
    .X(_12036_));
 sg13g2_nor2b_1 _18923_ (.A(\cpu.dec.jmp ),
    .B_N(_12036_),
    .Y(_12037_));
 sg13g2_nor2_1 _18924_ (.A(_12025_),
    .B(_12037_),
    .Y(_00053_));
 sg13g2_buf_2 _18925_ (.A(\cpu.qspi.r_state[6] ),
    .X(_12038_));
 sg13g2_and2_1 _18926_ (.A(_12038_),
    .B(net680),
    .X(_00010_));
 sg13g2_buf_1 _18927_ (.A(\cpu.qspi.r_state[13] ),
    .X(_12039_));
 sg13g2_and2_1 _18928_ (.A(_12039_),
    .B(net680),
    .X(_00006_));
 sg13g2_or3_1 _18929_ (.A(_08245_),
    .B(_08419_),
    .C(_09757_),
    .X(_12040_));
 sg13g2_buf_1 _18930_ (.A(_12040_),
    .X(_12041_));
 sg13g2_buf_1 _18931_ (.A(_12041_),
    .X(_12042_));
 sg13g2_nor2_1 _18932_ (.A(_12042_),
    .B(net647),
    .Y(_00052_));
 sg13g2_or2_1 _18933_ (.X(_12043_),
    .B(_09254_),
    .A(net1151));
 sg13g2_buf_1 _18934_ (.A(_12043_),
    .X(_12044_));
 sg13g2_nor3_1 _18935_ (.A(net1150),
    .B(_09265_),
    .C(_12044_),
    .Y(_12045_));
 sg13g2_a21oi_1 _18936_ (.A1(_09249_),
    .A2(_12044_),
    .Y(_12046_),
    .B1(_12045_));
 sg13g2_nand2_1 _18937_ (.Y(_12047_),
    .A(_09302_),
    .B(_12046_));
 sg13g2_inv_1 _18938_ (.Y(_12048_),
    .A(_00219_));
 sg13g2_or3_1 _18939_ (.A(_09254_),
    .B(net1150),
    .C(_12048_),
    .X(_12049_));
 sg13g2_buf_1 _18940_ (.A(_12049_),
    .X(_12050_));
 sg13g2_buf_2 _18941_ (.A(\cpu.spi.r_sel[0] ),
    .X(_12051_));
 sg13g2_buf_1 _18942_ (.A(_00275_),
    .X(_12052_));
 sg13g2_buf_1 _18943_ (.A(\cpu.spi.r_sel[1] ),
    .X(_12053_));
 sg13g2_buf_1 _18944_ (.A(net1119),
    .X(_12054_));
 sg13g2_mux2_1 _18945_ (.A0(_00276_),
    .A1(_12052_),
    .S(_12054_),
    .X(_12055_));
 sg13g2_buf_1 _18946_ (.A(\cpu.spi.r_src[2] ),
    .X(_12056_));
 sg13g2_nand2_1 _18947_ (.Y(_12057_),
    .A(net1119),
    .B(_12056_));
 sg13g2_o21ai_1 _18948_ (.B1(_12057_),
    .Y(_12058_),
    .A1(net1033),
    .A2(_12052_));
 sg13g2_nor2_1 _18949_ (.A(_12051_),
    .B(_12058_),
    .Y(_12059_));
 sg13g2_a21oi_2 _18950_ (.B1(_12059_),
    .Y(_12060_),
    .A2(_12055_),
    .A1(_12051_));
 sg13g2_and2_1 _18951_ (.A(_12050_),
    .B(_12060_),
    .X(_12061_));
 sg13g2_nor2_1 _18952_ (.A(net1151),
    .B(_09247_),
    .Y(_12062_));
 sg13g2_inv_1 _18953_ (.Y(_12063_),
    .A(_12051_));
 sg13g2_buf_1 _18954_ (.A(_12063_),
    .X(_12064_));
 sg13g2_buf_1 _18955_ (.A(net901),
    .X(_12065_));
 sg13g2_buf_1 _18956_ (.A(\cpu.spi.r_mode[0][1] ),
    .X(_12066_));
 sg13g2_buf_1 _18957_ (.A(\cpu.spi.r_mode[2][1] ),
    .X(_12067_));
 sg13g2_buf_1 _18958_ (.A(net1119),
    .X(_12068_));
 sg13g2_mux2_1 _18959_ (.A0(_12066_),
    .A1(_12067_),
    .S(net1032),
    .X(_12069_));
 sg13g2_nor2_1 _18960_ (.A(net901),
    .B(_12053_),
    .Y(_12070_));
 sg13g2_buf_1 _18961_ (.A(\cpu.spi.r_mode[1][1] ),
    .X(_12071_));
 sg13g2_a22oi_1 _18962_ (.Y(_12072_),
    .B1(_12070_),
    .B2(_12071_),
    .A2(_12069_),
    .A1(_12065_));
 sg13g2_xnor2_1 _18963_ (.Y(_12073_),
    .A(_12062_),
    .B(_12072_));
 sg13g2_buf_1 _18964_ (.A(_11080_),
    .X(_12074_));
 sg13g2_buf_1 _18965_ (.A(_09454_),
    .X(_12075_));
 sg13g2_buf_1 _18966_ (.A(net771),
    .X(_12076_));
 sg13g2_buf_1 _18967_ (.A(net925),
    .X(_12077_));
 sg13g2_and2_1 _18968_ (.A(net770),
    .B(_00276_),
    .X(_12078_));
 sg13g2_a21oi_1 _18969_ (.A1(net679),
    .A2(_12052_),
    .Y(_12079_),
    .B1(_12078_));
 sg13g2_nor2_1 _18970_ (.A(net900),
    .B(net770),
    .Y(_12080_));
 sg13g2_a22oi_1 _18971_ (.Y(_12081_),
    .B1(_12080_),
    .B2(_12056_),
    .A2(_12079_),
    .A1(net900));
 sg13g2_nor2_1 _18972_ (.A(_12050_),
    .B(_12081_),
    .Y(_12082_));
 sg13g2_buf_1 _18973_ (.A(net1061),
    .X(_12083_));
 sg13g2_buf_1 _18974_ (.A(net899),
    .X(_12084_));
 sg13g2_buf_1 _18975_ (.A(net769),
    .X(_12085_));
 sg13g2_buf_1 _18976_ (.A(net770),
    .X(_12086_));
 sg13g2_nand2b_1 _18977_ (.Y(_12087_),
    .B(net677),
    .A_N(_12066_));
 sg13g2_o21ai_1 _18978_ (.B1(_12087_),
    .Y(_12088_),
    .A1(net677),
    .A2(_12067_));
 sg13g2_mux2_1 _18979_ (.A0(_12066_),
    .A1(_12071_),
    .S(net677),
    .X(_12089_));
 sg13g2_nor2_1 _18980_ (.A(net678),
    .B(_12089_),
    .Y(_12090_));
 sg13g2_a21oi_1 _18981_ (.A1(_12085_),
    .A2(_12088_),
    .Y(_12091_),
    .B1(_12090_));
 sg13g2_a22oi_1 _18982_ (.Y(_12092_),
    .B1(_12082_),
    .B2(_12091_),
    .A2(_12073_),
    .A1(_12061_));
 sg13g2_nor2_1 _18983_ (.A(_12061_),
    .B(_12082_),
    .Y(_12093_));
 sg13g2_buf_1 _18984_ (.A(\cpu.gpio.genblk1[3].srcs_o[5] ),
    .X(_12094_));
 sg13g2_o21ai_1 _18985_ (.B1(_12094_),
    .Y(_12095_),
    .A1(_12047_),
    .A2(_12093_));
 sg13g2_o21ai_1 _18986_ (.B1(_12095_),
    .Y(_00309_),
    .A1(_12047_),
    .A2(_12092_));
 sg13g2_nor2b_1 _18987_ (.A(_12047_),
    .B_N(_12093_),
    .Y(_12096_));
 sg13g2_buf_1 _18988_ (.A(_12050_),
    .X(_12097_));
 sg13g2_nor2b_1 _18989_ (.A(_12097_),
    .B_N(_12091_),
    .Y(_12098_));
 sg13g2_a21oi_1 _18990_ (.A1(net768),
    .A2(_12073_),
    .Y(_12099_),
    .B1(_12098_));
 sg13g2_buf_1 _18991_ (.A(\cpu.gpio.genblk1[3].srcs_o[4] ),
    .X(_12100_));
 sg13g2_nor2_1 _18992_ (.A(_12100_),
    .B(_12096_),
    .Y(_12101_));
 sg13g2_a21oi_1 _18993_ (.A1(_12096_),
    .A2(_12099_),
    .Y(_00310_),
    .B1(_12101_));
 sg13g2_buf_1 _18994_ (.A(net1152),
    .X(_12102_));
 sg13g2_mux2_1 _18995_ (.A0(\cpu.spi.r_out[7] ),
    .A1(_10015_),
    .S(_12102_),
    .X(_12103_));
 sg13g2_buf_1 _18996_ (.A(\cpu.gpio.genblk1[3].srcs_o[3] ),
    .X(_12104_));
 sg13g2_inv_1 _18997_ (.Y(_12105_),
    .A(_00217_));
 sg13g2_mux2_1 _18998_ (.A0(_12105_),
    .A1(\cpu.spi.r_mode[2][0] ),
    .S(net1119),
    .X(_12106_));
 sg13g2_a22oi_1 _18999_ (.Y(_12107_),
    .B1(_12106_),
    .B2(_12064_),
    .A2(_12070_),
    .A1(\cpu.spi.r_mode[1][0] ));
 sg13g2_buf_1 _19000_ (.A(_12107_),
    .X(_12108_));
 sg13g2_buf_1 _19001_ (.A(_12108_),
    .X(_12109_));
 sg13g2_a21oi_1 _19002_ (.A1(_09245_),
    .A2(net553),
    .Y(_12110_),
    .B1(_09261_));
 sg13g2_or3_1 _19003_ (.A(net1152),
    .B(net1150),
    .C(_12044_),
    .X(_12111_));
 sg13g2_nand2_1 _19004_ (.Y(_12112_),
    .A(_09239_),
    .B(_12108_));
 sg13g2_a21o_1 _19005_ (.A2(_09206_),
    .A1(_00213_),
    .B1(_09254_),
    .X(_12113_));
 sg13g2_o21ai_1 _19006_ (.B1(_09254_),
    .Y(_12114_),
    .A1(_09249_),
    .A2(_12108_));
 sg13g2_nand2_1 _19007_ (.Y(_12115_),
    .A(_09251_),
    .B(_12114_));
 sg13g2_o21ai_1 _19008_ (.B1(_12115_),
    .Y(_12116_),
    .A1(_12112_),
    .A2(_12113_));
 sg13g2_nand3_1 _19009_ (.B(_12111_),
    .C(_12116_),
    .A(net933),
    .Y(_12117_));
 sg13g2_nor2_1 _19010_ (.A(_12110_),
    .B(_12117_),
    .Y(_12118_));
 sg13g2_nand2_1 _19011_ (.Y(_12119_),
    .A(_12060_),
    .B(_12118_));
 sg13g2_mux2_1 _19012_ (.A0(_12103_),
    .A1(_12104_),
    .S(_12119_),
    .X(_00311_));
 sg13g2_buf_1 _19013_ (.A(\cpu.gpio.genblk1[3].srcs_o[2] ),
    .X(_12120_));
 sg13g2_nor3_1 _19014_ (.A(_12060_),
    .B(_12110_),
    .C(_12117_),
    .Y(_12121_));
 sg13g2_mux2_1 _19015_ (.A0(_12120_),
    .A1(_12103_),
    .S(_12121_),
    .X(_00312_));
 sg13g2_buf_1 _19016_ (.A(net926),
    .X(_12122_));
 sg13g2_nand2_1 _19017_ (.Y(_12123_),
    .A(net767),
    .B(_09351_));
 sg13g2_nor3_1 _19018_ (.A(_09303_),
    .B(_08355_),
    .C(_09747_),
    .Y(_12124_));
 sg13g2_buf_1 _19019_ (.A(\cpu.dcache.r_offset[2] ),
    .X(_12125_));
 sg13g2_buf_1 _19020_ (.A(\cpu.d_wstrobe_d ),
    .X(_12126_));
 sg13g2_buf_2 _19021_ (.A(\cpu.dcache.r_offset[0] ),
    .X(_12127_));
 sg13g2_and2_1 _19022_ (.A(\cpu.dcache.r_offset[1] ),
    .B(_12127_),
    .X(_12128_));
 sg13g2_buf_2 _19023_ (.A(_12128_),
    .X(_12129_));
 sg13g2_nand3_1 _19024_ (.B(_12126_),
    .C(_12129_),
    .A(net1114),
    .Y(_12130_));
 sg13g2_buf_2 _19025_ (.A(_12130_),
    .X(_12131_));
 sg13g2_nand2b_1 _19026_ (.Y(_12132_),
    .B(_12131_),
    .A_N(_09742_));
 sg13g2_and2_1 _19027_ (.A(_12124_),
    .B(_12132_),
    .X(_12133_));
 sg13g2_buf_1 _19028_ (.A(_12133_),
    .X(_12134_));
 sg13g2_nand2b_1 _19029_ (.Y(_12135_),
    .B(_12134_),
    .A_N(_12123_));
 sg13g2_buf_1 _19030_ (.A(_12135_),
    .X(_12136_));
 sg13g2_nand2_1 _19031_ (.Y(_12137_),
    .A(_08267_),
    .B(net1067));
 sg13g2_buf_1 _19032_ (.A(_12137_),
    .X(_12138_));
 sg13g2_buf_2 _19033_ (.A(_00268_),
    .X(_12139_));
 sg13g2_buf_1 _19034_ (.A(_12139_),
    .X(_12140_));
 sg13g2_o21ai_1 _19035_ (.B1(net1030),
    .Y(_12141_),
    .A1(_08268_),
    .A2(_12138_));
 sg13g2_nor2_1 _19036_ (.A(_12136_),
    .B(_12141_),
    .Y(_12142_));
 sg13g2_buf_2 _19037_ (.A(_12142_),
    .X(_12143_));
 sg13g2_buf_1 _19038_ (.A(_12143_),
    .X(_12144_));
 sg13g2_buf_1 _19039_ (.A(uio_in[0]),
    .X(_12145_));
 sg13g2_buf_1 _19040_ (.A(_12145_),
    .X(_12146_));
 sg13g2_buf_1 _19041_ (.A(_12123_),
    .X(_12147_));
 sg13g2_buf_1 _19042_ (.A(_12126_),
    .X(_12148_));
 sg13g2_buf_1 _19043_ (.A(_00269_),
    .X(_12149_));
 sg13g2_buf_1 _19044_ (.A(_12149_),
    .X(_12150_));
 sg13g2_buf_1 _19045_ (.A(\cpu.dcache.r_offset[1] ),
    .X(_12151_));
 sg13g2_nor2b_1 _19046_ (.A(_12151_),
    .B_N(_12127_),
    .Y(_12152_));
 sg13g2_buf_1 _19047_ (.A(_12152_),
    .X(_12153_));
 sg13g2_nand3_1 _19048_ (.B(net1028),
    .C(_12153_),
    .A(net1029),
    .Y(_12154_));
 sg13g2_buf_2 _19049_ (.A(_12154_),
    .X(_12155_));
 sg13g2_nor2_1 _19050_ (.A(net625),
    .B(_12155_),
    .Y(_12156_));
 sg13g2_buf_2 _19051_ (.A(_12156_),
    .X(_12157_));
 sg13g2_mux2_1 _19052_ (.A0(\cpu.dcache.r_data[0][0] ),
    .A1(net1113),
    .S(_12157_),
    .X(_12158_));
 sg13g2_nor2_1 _19053_ (.A(_12143_),
    .B(_12158_),
    .Y(_12159_));
 sg13g2_a21oi_1 _19054_ (.A1(_09971_),
    .A2(net62),
    .Y(_00313_),
    .B1(_12159_));
 sg13g2_inv_1 _19055_ (.Y(_12160_),
    .A(_12139_));
 sg13g2_buf_1 _19056_ (.A(_12160_),
    .X(_12161_));
 sg13g2_mux2_1 _19057_ (.A0(_10026_),
    .A1(net898),
    .S(_08290_),
    .X(_12162_));
 sg13g2_nor3_1 _19058_ (.A(_12136_),
    .B(_12138_),
    .C(_12162_),
    .Y(_12163_));
 sg13g2_buf_2 _19059_ (.A(_12163_),
    .X(_12164_));
 sg13g2_buf_1 _19060_ (.A(_12164_),
    .X(_12165_));
 sg13g2_buf_1 _19061_ (.A(uio_in[2]),
    .X(_12166_));
 sg13g2_buf_1 _19062_ (.A(_12166_),
    .X(_12167_));
 sg13g2_buf_2 _19063_ (.A(net1111),
    .X(_12168_));
 sg13g2_nand3_1 _19064_ (.B(net1028),
    .C(_12129_),
    .A(net1029),
    .Y(_12169_));
 sg13g2_buf_2 _19065_ (.A(_12169_),
    .X(_12170_));
 sg13g2_nor2_1 _19066_ (.A(net625),
    .B(_12170_),
    .Y(_12171_));
 sg13g2_buf_2 _19067_ (.A(_12171_),
    .X(_12172_));
 sg13g2_nor2b_1 _19068_ (.A(_12172_),
    .B_N(\cpu.dcache.r_data[0][10] ),
    .Y(_12173_));
 sg13g2_a21oi_1 _19069_ (.A1(net1027),
    .A2(_12172_),
    .Y(_12174_),
    .B1(_12173_));
 sg13g2_inv_1 _19070_ (.Y(_12175_),
    .A(_09984_));
 sg13g2_nor2_1 _19071_ (.A(_08290_),
    .B(_12138_),
    .Y(_12176_));
 sg13g2_buf_1 _19072_ (.A(_12176_),
    .X(_12177_));
 sg13g2_nand2_1 _19073_ (.Y(_12178_),
    .A(_10091_),
    .B(_12176_));
 sg13g2_o21ai_1 _19074_ (.B1(_12178_),
    .Y(_12179_),
    .A1(_12175_),
    .A2(_12177_));
 sg13g2_buf_2 _19075_ (.A(_12179_),
    .X(_12180_));
 sg13g2_buf_1 _19076_ (.A(_12180_),
    .X(_12181_));
 sg13g2_nand2_1 _19077_ (.Y(_12182_),
    .A(_12181_),
    .B(_12164_));
 sg13g2_o21ai_1 _19078_ (.B1(_12182_),
    .Y(_00314_),
    .A1(net61),
    .A2(_12174_));
 sg13g2_buf_1 _19079_ (.A(uio_in[3]),
    .X(_12183_));
 sg13g2_buf_1 _19080_ (.A(_12183_),
    .X(_12184_));
 sg13g2_buf_2 _19081_ (.A(_12184_),
    .X(_12185_));
 sg13g2_nor2b_1 _19082_ (.A(_12172_),
    .B_N(\cpu.dcache.r_data[0][11] ),
    .Y(_12186_));
 sg13g2_a21oi_1 _19083_ (.A1(net1026),
    .A2(_12172_),
    .Y(_12187_),
    .B1(_12186_));
 sg13g2_mux2_1 _19084_ (.A0(net1144),
    .A1(_10098_),
    .S(net624),
    .X(_12188_));
 sg13g2_buf_2 _19085_ (.A(_12188_),
    .X(_12189_));
 sg13g2_nand2_1 _19086_ (.Y(_12190_),
    .A(net61),
    .B(_12189_));
 sg13g2_o21ai_1 _19087_ (.B1(_12190_),
    .Y(_00315_),
    .A1(_12165_),
    .A2(_12187_));
 sg13g2_inv_1 _19088_ (.Y(_12191_),
    .A(_09999_));
 sg13g2_inv_1 _19089_ (.Y(_12192_),
    .A(_10103_));
 sg13g2_mux2_1 _19090_ (.A0(_12191_),
    .A1(_12192_),
    .S(net624),
    .X(_12193_));
 sg13g2_buf_2 _19091_ (.A(_12193_),
    .X(_12194_));
 sg13g2_buf_1 _19092_ (.A(_12127_),
    .X(_12195_));
 sg13g2_nor2b_1 _19093_ (.A(net1025),
    .B_N(net1112),
    .Y(_12196_));
 sg13g2_nand3_1 _19094_ (.B(_12150_),
    .C(_12196_),
    .A(net1029),
    .Y(_12197_));
 sg13g2_buf_4 _19095_ (.X(_12198_),
    .A(_12197_));
 sg13g2_nor2_2 _19096_ (.A(net625),
    .B(_12198_),
    .Y(_12199_));
 sg13g2_mux2_1 _19097_ (.A0(\cpu.dcache.r_data[0][12] ),
    .A1(_12146_),
    .S(_12199_),
    .X(_12200_));
 sg13g2_nor2_1 _19098_ (.A(_12164_),
    .B(_12200_),
    .Y(_12201_));
 sg13g2_a21oi_1 _19099_ (.A1(net61),
    .A2(_12194_),
    .Y(_00316_),
    .B1(_12201_));
 sg13g2_inv_1 _19100_ (.Y(_12202_),
    .A(_10005_));
 sg13g2_inv_1 _19101_ (.Y(_12203_),
    .A(_10108_));
 sg13g2_mux2_1 _19102_ (.A0(_12202_),
    .A1(_12203_),
    .S(net624),
    .X(_12204_));
 sg13g2_buf_2 _19103_ (.A(_12204_),
    .X(_12205_));
 sg13g2_buf_1 _19104_ (.A(uio_in[1]),
    .X(_12206_));
 sg13g2_buf_2 _19105_ (.A(_12206_),
    .X(_12207_));
 sg13g2_mux2_1 _19106_ (.A0(\cpu.dcache.r_data[0][13] ),
    .A1(net1109),
    .S(_12199_),
    .X(_12208_));
 sg13g2_nor2_1 _19107_ (.A(_12164_),
    .B(_12208_),
    .Y(_12209_));
 sg13g2_a21oi_1 _19108_ (.A1(net61),
    .A2(_12205_),
    .Y(_00317_),
    .B1(_12209_));
 sg13g2_inv_1 _19109_ (.Y(_12210_),
    .A(_10010_));
 sg13g2_nor2_1 _19110_ (.A(_12210_),
    .B(net624),
    .Y(_12211_));
 sg13g2_a21oi_1 _19111_ (.A1(_10114_),
    .A2(net624),
    .Y(_12212_),
    .B1(_12211_));
 sg13g2_buf_2 _19112_ (.A(_12212_),
    .X(_12213_));
 sg13g2_buf_2 _19113_ (.A(_12166_),
    .X(_12214_));
 sg13g2_mux2_1 _19114_ (.A0(\cpu.dcache.r_data[0][14] ),
    .A1(net1108),
    .S(_12199_),
    .X(_12215_));
 sg13g2_nor2_1 _19115_ (.A(_12164_),
    .B(_12215_),
    .Y(_12216_));
 sg13g2_a21oi_1 _19116_ (.A1(net61),
    .A2(_12213_),
    .Y(_00318_),
    .B1(_12216_));
 sg13g2_inv_1 _19117_ (.Y(_12217_),
    .A(_10015_));
 sg13g2_nor2_1 _19118_ (.A(_12217_),
    .B(net624),
    .Y(_12218_));
 sg13g2_a21oi_1 _19119_ (.A1(_10122_),
    .A2(net624),
    .Y(_12219_),
    .B1(_12218_));
 sg13g2_buf_2 _19120_ (.A(_12219_),
    .X(_12220_));
 sg13g2_buf_1 _19121_ (.A(_12183_),
    .X(_12221_));
 sg13g2_mux2_1 _19122_ (.A0(\cpu.dcache.r_data[0][15] ),
    .A1(net1107),
    .S(_12199_),
    .X(_12222_));
 sg13g2_nor2_1 _19123_ (.A(_12164_),
    .B(_12222_),
    .Y(_12223_));
 sg13g2_a21oi_1 _19124_ (.A1(net61),
    .A2(_12220_),
    .Y(_00319_),
    .B1(_12223_));
 sg13g2_buf_1 _19125_ (.A(net796),
    .X(_12224_));
 sg13g2_o21ai_1 _19126_ (.B1(net676),
    .Y(_12225_),
    .A1(_08268_),
    .A2(_12138_));
 sg13g2_nor2_1 _19127_ (.A(_12136_),
    .B(_12225_),
    .Y(_12226_));
 sg13g2_buf_2 _19128_ (.A(_12226_),
    .X(_12227_));
 sg13g2_buf_1 _19129_ (.A(_12227_),
    .X(_12228_));
 sg13g2_nand3_1 _19130_ (.B(net1029),
    .C(_12153_),
    .A(net1114),
    .Y(_12229_));
 sg13g2_buf_2 _19131_ (.A(_12229_),
    .X(_12230_));
 sg13g2_nor2_1 _19132_ (.A(net625),
    .B(_12230_),
    .Y(_12231_));
 sg13g2_buf_2 _19133_ (.A(_12231_),
    .X(_12232_));
 sg13g2_mux2_1 _19134_ (.A0(\cpu.dcache.r_data[0][16] ),
    .A1(net1113),
    .S(_12232_),
    .X(_12233_));
 sg13g2_nor2_1 _19135_ (.A(_12227_),
    .B(_12233_),
    .Y(_12234_));
 sg13g2_a21oi_1 _19136_ (.A1(net797),
    .A2(net60),
    .Y(_00320_),
    .B1(_12234_));
 sg13g2_inv_1 _19137_ (.Y(_12235_),
    .A(_09978_));
 sg13g2_buf_1 _19138_ (.A(_12235_),
    .X(_12236_));
 sg13g2_buf_1 _19139_ (.A(net897),
    .X(_12237_));
 sg13g2_mux2_1 _19140_ (.A0(\cpu.dcache.r_data[0][17] ),
    .A1(net1109),
    .S(_12232_),
    .X(_12238_));
 sg13g2_nor2_1 _19141_ (.A(_12227_),
    .B(_12238_),
    .Y(_12239_));
 sg13g2_a21oi_1 _19142_ (.A1(net766),
    .A2(_12228_),
    .Y(_00321_),
    .B1(_12239_));
 sg13g2_buf_1 _19143_ (.A(_12175_),
    .X(_12240_));
 sg13g2_buf_1 _19144_ (.A(net896),
    .X(_12241_));
 sg13g2_mux2_1 _19145_ (.A0(\cpu.dcache.r_data[0][18] ),
    .A1(net1108),
    .S(_12232_),
    .X(_12242_));
 sg13g2_nor2_1 _19146_ (.A(_12227_),
    .B(_12242_),
    .Y(_12243_));
 sg13g2_a21oi_1 _19147_ (.A1(net765),
    .A2(net60),
    .Y(_00322_),
    .B1(_12243_));
 sg13g2_nor2b_1 _19148_ (.A(_12232_),
    .B_N(\cpu.dcache.r_data[0][19] ),
    .Y(_12244_));
 sg13g2_a21oi_1 _19149_ (.A1(net1026),
    .A2(_12232_),
    .Y(_12245_),
    .B1(_12244_));
 sg13g2_buf_1 _19150_ (.A(net1144),
    .X(_12246_));
 sg13g2_nand2_1 _19151_ (.Y(_12247_),
    .A(net1024),
    .B(net60));
 sg13g2_o21ai_1 _19152_ (.B1(_12247_),
    .Y(_00323_),
    .A1(net60),
    .A2(_12245_));
 sg13g2_mux2_1 _19153_ (.A0(\cpu.dcache.r_data[0][1] ),
    .A1(net1109),
    .S(_12157_),
    .X(_12248_));
 sg13g2_nor2_1 _19154_ (.A(_12143_),
    .B(_12248_),
    .Y(_12249_));
 sg13g2_a21oi_1 _19155_ (.A1(net766),
    .A2(_12144_),
    .Y(_00324_),
    .B1(_12249_));
 sg13g2_buf_1 _19156_ (.A(_12145_),
    .X(_12250_));
 sg13g2_buf_2 _19157_ (.A(net1106),
    .X(_12251_));
 sg13g2_nor2_2 _19158_ (.A(net1112),
    .B(_12127_),
    .Y(_12252_));
 sg13g2_nand3_1 _19159_ (.B(net1029),
    .C(_12252_),
    .A(net1114),
    .Y(_12253_));
 sg13g2_buf_2 _19160_ (.A(_12253_),
    .X(_12254_));
 sg13g2_nor2_1 _19161_ (.A(net625),
    .B(_12254_),
    .Y(_12255_));
 sg13g2_buf_2 _19162_ (.A(_12255_),
    .X(_12256_));
 sg13g2_nor2b_1 _19163_ (.A(_12256_),
    .B_N(\cpu.dcache.r_data[0][20] ),
    .Y(_12257_));
 sg13g2_a21oi_1 _19164_ (.A1(net1023),
    .A2(_12256_),
    .Y(_12258_),
    .B1(_12257_));
 sg13g2_buf_1 _19165_ (.A(_09999_),
    .X(_12259_));
 sg13g2_nand2_1 _19166_ (.Y(_12260_),
    .A(net1022),
    .B(net60));
 sg13g2_o21ai_1 _19167_ (.B1(_12260_),
    .Y(_00325_),
    .A1(net60),
    .A2(_12258_));
 sg13g2_buf_1 _19168_ (.A(_12202_),
    .X(_12261_));
 sg13g2_buf_1 _19169_ (.A(net895),
    .X(_12262_));
 sg13g2_mux2_1 _19170_ (.A0(\cpu.dcache.r_data[0][21] ),
    .A1(net1109),
    .S(_12256_),
    .X(_12263_));
 sg13g2_nor2_1 _19171_ (.A(_12227_),
    .B(_12263_),
    .Y(_12264_));
 sg13g2_a21oi_1 _19172_ (.A1(net764),
    .A2(net60),
    .Y(_00326_),
    .B1(_12264_));
 sg13g2_buf_1 _19173_ (.A(_12210_),
    .X(_12265_));
 sg13g2_buf_1 _19174_ (.A(net894),
    .X(_12266_));
 sg13g2_mux2_1 _19175_ (.A0(\cpu.dcache.r_data[0][22] ),
    .A1(net1108),
    .S(_12256_),
    .X(_12267_));
 sg13g2_nor2_1 _19176_ (.A(_12227_),
    .B(_12267_),
    .Y(_12268_));
 sg13g2_a21oi_1 _19177_ (.A1(net763),
    .A2(_12228_),
    .Y(_00327_),
    .B1(_12268_));
 sg13g2_buf_1 _19178_ (.A(_12217_),
    .X(_12269_));
 sg13g2_buf_1 _19179_ (.A(net893),
    .X(_12270_));
 sg13g2_mux2_1 _19180_ (.A0(\cpu.dcache.r_data[0][23] ),
    .A1(net1107),
    .S(_12256_),
    .X(_12271_));
 sg13g2_nor2_1 _19181_ (.A(_12227_),
    .B(_12271_),
    .Y(_12272_));
 sg13g2_a21oi_1 _19182_ (.A1(_12270_),
    .A2(net60),
    .Y(_00328_),
    .B1(_12272_));
 sg13g2_and3_1 _19183_ (.X(_12273_),
    .A(net1114),
    .B(_12126_),
    .C(_12129_));
 sg13g2_buf_1 _19184_ (.A(_12273_),
    .X(_12274_));
 sg13g2_nand2b_1 _19185_ (.Y(_12275_),
    .B(_12274_),
    .A_N(_12147_));
 sg13g2_buf_1 _19186_ (.A(_12275_),
    .X(_12276_));
 sg13g2_buf_1 _19187_ (.A(_12276_),
    .X(_12277_));
 sg13g2_mux2_1 _19188_ (.A0(net1113),
    .A1(\cpu.dcache.r_data[0][24] ),
    .S(net432),
    .X(_12278_));
 sg13g2_nand2_1 _19189_ (.Y(_12279_),
    .A(_10081_),
    .B(_12176_));
 sg13g2_o21ai_1 _19190_ (.B1(_12279_),
    .Y(_12280_),
    .A1(_09969_),
    .A2(_12177_));
 sg13g2_buf_2 _19191_ (.A(_12280_),
    .X(_12281_));
 sg13g2_buf_1 _19192_ (.A(_12281_),
    .X(_12282_));
 sg13g2_nand2_1 _19193_ (.Y(_12283_),
    .A(_08268_),
    .B(_12139_));
 sg13g2_o21ai_1 _19194_ (.B1(_12283_),
    .Y(_12284_),
    .A1(_08268_),
    .A2(net676));
 sg13g2_nor3_1 _19195_ (.A(_12136_),
    .B(_12138_),
    .C(_12284_),
    .Y(_12285_));
 sg13g2_buf_2 _19196_ (.A(_12285_),
    .X(_12286_));
 sg13g2_mux2_1 _19197_ (.A0(_12278_),
    .A1(net431),
    .S(net73),
    .X(_00329_));
 sg13g2_mux2_1 _19198_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[0][25] ),
    .S(net432),
    .X(_12287_));
 sg13g2_nand2_1 _19199_ (.Y(_12288_),
    .A(_10086_),
    .B(_12176_));
 sg13g2_o21ai_1 _19200_ (.B1(_12288_),
    .Y(_12289_),
    .A1(_12235_),
    .A2(net624));
 sg13g2_buf_2 _19201_ (.A(_12289_),
    .X(_12290_));
 sg13g2_buf_1 _19202_ (.A(_12290_),
    .X(_12291_));
 sg13g2_mux2_1 _19203_ (.A0(_12287_),
    .A1(net430),
    .S(net73),
    .X(_00330_));
 sg13g2_mux2_1 _19204_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[0][26] ),
    .S(net432),
    .X(_12292_));
 sg13g2_mux2_1 _19205_ (.A0(_12292_),
    .A1(net433),
    .S(_12286_),
    .X(_00331_));
 sg13g2_mux2_1 _19206_ (.A0(_12221_),
    .A1(\cpu.dcache.r_data[0][27] ),
    .S(net432),
    .X(_12293_));
 sg13g2_buf_1 _19207_ (.A(_12189_),
    .X(_12294_));
 sg13g2_mux2_1 _19208_ (.A0(_12293_),
    .A1(net429),
    .S(_12286_),
    .X(_00332_));
 sg13g2_buf_1 _19209_ (.A(_12194_),
    .X(_12295_));
 sg13g2_buf_1 _19210_ (.A(_12125_),
    .X(_12296_));
 sg13g2_nand3_1 _19211_ (.B(net1029),
    .C(_12196_),
    .A(net1021),
    .Y(_12297_));
 sg13g2_buf_4 _19212_ (.X(_12298_),
    .A(_12297_));
 sg13g2_nor2_2 _19213_ (.A(net625),
    .B(_12298_),
    .Y(_12299_));
 sg13g2_mux2_1 _19214_ (.A0(\cpu.dcache.r_data[0][28] ),
    .A1(net1113),
    .S(_12299_),
    .X(_12300_));
 sg13g2_nor2_1 _19215_ (.A(net73),
    .B(_12300_),
    .Y(_12301_));
 sg13g2_a21oi_1 _19216_ (.A1(net428),
    .A2(net73),
    .Y(_00333_),
    .B1(_12301_));
 sg13g2_buf_1 _19217_ (.A(_12205_),
    .X(_12302_));
 sg13g2_buf_1 _19218_ (.A(_12206_),
    .X(_12303_));
 sg13g2_buf_1 _19219_ (.A(net1105),
    .X(_12304_));
 sg13g2_mux2_1 _19220_ (.A0(\cpu.dcache.r_data[0][29] ),
    .A1(net1020),
    .S(_12299_),
    .X(_12305_));
 sg13g2_nor2_1 _19221_ (.A(net73),
    .B(_12305_),
    .Y(_12306_));
 sg13g2_a21oi_1 _19222_ (.A1(_12302_),
    .A2(net73),
    .Y(_00334_),
    .B1(_12306_));
 sg13g2_mux2_1 _19223_ (.A0(\cpu.dcache.r_data[0][2] ),
    .A1(net1108),
    .S(_12157_),
    .X(_12307_));
 sg13g2_nor2_1 _19224_ (.A(_12143_),
    .B(_12307_),
    .Y(_12308_));
 sg13g2_a21oi_1 _19225_ (.A1(net765),
    .A2(_12144_),
    .Y(_00335_),
    .B1(_12308_));
 sg13g2_buf_1 _19226_ (.A(_12213_),
    .X(_12309_));
 sg13g2_buf_1 _19227_ (.A(net1111),
    .X(_12310_));
 sg13g2_mux2_1 _19228_ (.A0(\cpu.dcache.r_data[0][30] ),
    .A1(net1019),
    .S(_12299_),
    .X(_12311_));
 sg13g2_nor2_1 _19229_ (.A(_12285_),
    .B(_12311_),
    .Y(_12312_));
 sg13g2_a21oi_1 _19230_ (.A1(net384),
    .A2(net73),
    .Y(_00336_),
    .B1(_12312_));
 sg13g2_buf_1 _19231_ (.A(_12220_),
    .X(_12313_));
 sg13g2_mux2_1 _19232_ (.A0(\cpu.dcache.r_data[0][31] ),
    .A1(net1107),
    .S(_12299_),
    .X(_12314_));
 sg13g2_nor2_1 _19233_ (.A(_12285_),
    .B(_12314_),
    .Y(_12315_));
 sg13g2_a21oi_1 _19234_ (.A1(_12313_),
    .A2(net73),
    .Y(_00337_),
    .B1(_12315_));
 sg13g2_nor2b_1 _19235_ (.A(_12157_),
    .B_N(\cpu.dcache.r_data[0][3] ),
    .Y(_12316_));
 sg13g2_a21oi_1 _19236_ (.A1(net1026),
    .A2(_12157_),
    .Y(_12317_),
    .B1(_12316_));
 sg13g2_nand2_1 _19237_ (.Y(_12318_),
    .A(net1024),
    .B(net62));
 sg13g2_o21ai_1 _19238_ (.B1(_12318_),
    .Y(_00338_),
    .A1(net62),
    .A2(_12317_));
 sg13g2_nand3_1 _19239_ (.B(net1028),
    .C(_12252_),
    .A(net1029),
    .Y(_12319_));
 sg13g2_buf_2 _19240_ (.A(_12319_),
    .X(_12320_));
 sg13g2_nor2_1 _19241_ (.A(net625),
    .B(_12320_),
    .Y(_12321_));
 sg13g2_buf_2 _19242_ (.A(_12321_),
    .X(_12322_));
 sg13g2_nor2b_1 _19243_ (.A(_12322_),
    .B_N(\cpu.dcache.r_data[0][4] ),
    .Y(_12323_));
 sg13g2_a21oi_1 _19244_ (.A1(net1023),
    .A2(_12322_),
    .Y(_12324_),
    .B1(_12323_));
 sg13g2_nand2_1 _19245_ (.Y(_12325_),
    .A(net1022),
    .B(net62));
 sg13g2_o21ai_1 _19246_ (.B1(_12325_),
    .Y(_00339_),
    .A1(net62),
    .A2(_12324_));
 sg13g2_mux2_1 _19247_ (.A0(\cpu.dcache.r_data[0][5] ),
    .A1(net1020),
    .S(_12322_),
    .X(_12326_));
 sg13g2_nor2_1 _19248_ (.A(_12143_),
    .B(_12326_),
    .Y(_12327_));
 sg13g2_a21oi_1 _19249_ (.A1(net764),
    .A2(net62),
    .Y(_00340_),
    .B1(_12327_));
 sg13g2_mux2_1 _19250_ (.A0(\cpu.dcache.r_data[0][6] ),
    .A1(net1019),
    .S(_12322_),
    .X(_12328_));
 sg13g2_nor2_1 _19251_ (.A(_12143_),
    .B(_12328_),
    .Y(_12329_));
 sg13g2_a21oi_1 _19252_ (.A1(net763),
    .A2(net62),
    .Y(_00341_),
    .B1(_12329_));
 sg13g2_mux2_1 _19253_ (.A0(\cpu.dcache.r_data[0][7] ),
    .A1(net1107),
    .S(_12322_),
    .X(_12330_));
 sg13g2_nor2_1 _19254_ (.A(_12143_),
    .B(_12330_),
    .Y(_12331_));
 sg13g2_a21oi_1 _19255_ (.A1(_12270_),
    .A2(net62),
    .Y(_00342_),
    .B1(_12331_));
 sg13g2_nor2b_1 _19256_ (.A(_12172_),
    .B_N(\cpu.dcache.r_data[0][8] ),
    .Y(_12332_));
 sg13g2_a21oi_1 _19257_ (.A1(net1023),
    .A2(_12172_),
    .Y(_12333_),
    .B1(_12332_));
 sg13g2_nand2_1 _19258_ (.Y(_12334_),
    .A(net61),
    .B(_12281_));
 sg13g2_o21ai_1 _19259_ (.B1(_12334_),
    .Y(_00343_),
    .A1(_12165_),
    .A2(_12333_));
 sg13g2_buf_2 _19260_ (.A(net1105),
    .X(_12335_));
 sg13g2_nor2b_1 _19261_ (.A(_12172_),
    .B_N(\cpu.dcache.r_data[0][9] ),
    .Y(_12336_));
 sg13g2_a21oi_1 _19262_ (.A1(net1018),
    .A2(_12172_),
    .Y(_12337_),
    .B1(_12336_));
 sg13g2_nand2_1 _19263_ (.Y(_12338_),
    .A(_12164_),
    .B(_12290_));
 sg13g2_o21ai_1 _19264_ (.B1(_12338_),
    .Y(_00344_),
    .A1(net61),
    .A2(_12337_));
 sg13g2_buf_1 _19265_ (.A(net699),
    .X(_12339_));
 sg13g2_inv_1 _19266_ (.Y(_12340_),
    .A(_12141_));
 sg13g2_nand2_1 _19267_ (.Y(_12341_),
    .A(_12134_),
    .B(_12340_));
 sg13g2_buf_2 _19268_ (.A(_12341_),
    .X(_12342_));
 sg13g2_nor2_1 _19269_ (.A(net623),
    .B(_12342_),
    .Y(_12343_));
 sg13g2_buf_2 _19270_ (.A(_12343_),
    .X(_12344_));
 sg13g2_buf_1 _19271_ (.A(_12344_),
    .X(_12345_));
 sg13g2_nor2_1 _19272_ (.A(net623),
    .B(_12155_),
    .Y(_12346_));
 sg13g2_buf_1 _19273_ (.A(_12346_),
    .X(_12347_));
 sg13g2_mux2_1 _19274_ (.A0(\cpu.dcache.r_data[1][0] ),
    .A1(net1113),
    .S(_12347_),
    .X(_12348_));
 sg13g2_nor2_1 _19275_ (.A(_12344_),
    .B(_12348_),
    .Y(_12349_));
 sg13g2_a21oi_1 _19276_ (.A1(net797),
    .A2(net59),
    .Y(_00345_),
    .B1(_12349_));
 sg13g2_nor2_1 _19277_ (.A(_08289_),
    .B(_08270_),
    .Y(_12350_));
 sg13g2_nand3b_1 _19278_ (.B(_12350_),
    .C(_12134_),
    .Y(_12351_),
    .A_N(_12162_));
 sg13g2_buf_2 _19279_ (.A(_12351_),
    .X(_12352_));
 sg13g2_nor2_1 _19280_ (.A(net623),
    .B(_12352_),
    .Y(_12353_));
 sg13g2_buf_2 _19281_ (.A(_12353_),
    .X(_12354_));
 sg13g2_buf_1 _19282_ (.A(_12354_),
    .X(_12355_));
 sg13g2_nor2_1 _19283_ (.A(net623),
    .B(_12170_),
    .Y(_12356_));
 sg13g2_buf_2 _19284_ (.A(_12356_),
    .X(_12357_));
 sg13g2_nor2b_1 _19285_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[1][10] ),
    .Y(_12358_));
 sg13g2_a21oi_1 _19286_ (.A1(net1027),
    .A2(_12357_),
    .Y(_12359_),
    .B1(_12358_));
 sg13g2_nand2_1 _19287_ (.Y(_12360_),
    .A(net433),
    .B(net58));
 sg13g2_o21ai_1 _19288_ (.B1(_12360_),
    .Y(_00346_),
    .A1(net58),
    .A2(_12359_));
 sg13g2_nor2b_1 _19289_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[1][11] ),
    .Y(_12361_));
 sg13g2_a21oi_1 _19290_ (.A1(net1026),
    .A2(_12357_),
    .Y(_12362_),
    .B1(_12361_));
 sg13g2_nand2_1 _19291_ (.Y(_12363_),
    .A(net429),
    .B(net58));
 sg13g2_o21ai_1 _19292_ (.B1(_12363_),
    .Y(_00347_),
    .A1(_12355_),
    .A2(_12362_));
 sg13g2_nor2_2 _19293_ (.A(net623),
    .B(_12198_),
    .Y(_12364_));
 sg13g2_mux2_1 _19294_ (.A0(\cpu.dcache.r_data[1][12] ),
    .A1(net1113),
    .S(_12364_),
    .X(_12365_));
 sg13g2_nor2_1 _19295_ (.A(_12354_),
    .B(_12365_),
    .Y(_12366_));
 sg13g2_a21oi_1 _19296_ (.A1(net428),
    .A2(net58),
    .Y(_00348_),
    .B1(_12366_));
 sg13g2_mux2_1 _19297_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(net1020),
    .S(_12364_),
    .X(_12367_));
 sg13g2_nor2_1 _19298_ (.A(_12354_),
    .B(_12367_),
    .Y(_12368_));
 sg13g2_a21oi_1 _19299_ (.A1(net427),
    .A2(net58),
    .Y(_00349_),
    .B1(_12368_));
 sg13g2_mux2_1 _19300_ (.A0(\cpu.dcache.r_data[1][14] ),
    .A1(net1019),
    .S(_12364_),
    .X(_12369_));
 sg13g2_nor2_1 _19301_ (.A(_12354_),
    .B(_12369_),
    .Y(_12370_));
 sg13g2_a21oi_1 _19302_ (.A1(net384),
    .A2(net58),
    .Y(_00350_),
    .B1(_12370_));
 sg13g2_mux2_1 _19303_ (.A0(\cpu.dcache.r_data[1][15] ),
    .A1(net1107),
    .S(_12364_),
    .X(_12371_));
 sg13g2_nor2_1 _19304_ (.A(_12354_),
    .B(_12371_),
    .Y(_12372_));
 sg13g2_a21oi_1 _19305_ (.A1(net383),
    .A2(net58),
    .Y(_00351_),
    .B1(_12372_));
 sg13g2_inv_1 _19306_ (.Y(_12373_),
    .A(_12225_));
 sg13g2_nand2_1 _19307_ (.Y(_12374_),
    .A(_12134_),
    .B(_12373_));
 sg13g2_buf_2 _19308_ (.A(_12374_),
    .X(_12375_));
 sg13g2_nor2_1 _19309_ (.A(net623),
    .B(_12375_),
    .Y(_12376_));
 sg13g2_buf_2 _19310_ (.A(_12376_),
    .X(_12377_));
 sg13g2_buf_1 _19311_ (.A(_12377_),
    .X(_12378_));
 sg13g2_nor2_1 _19312_ (.A(net623),
    .B(_12230_),
    .Y(_12379_));
 sg13g2_buf_2 _19313_ (.A(_12379_),
    .X(_12380_));
 sg13g2_mux2_1 _19314_ (.A0(\cpu.dcache.r_data[1][16] ),
    .A1(net1113),
    .S(_12380_),
    .X(_12381_));
 sg13g2_nor2_1 _19315_ (.A(_12377_),
    .B(_12381_),
    .Y(_12382_));
 sg13g2_a21oi_1 _19316_ (.A1(net797),
    .A2(net57),
    .Y(_00352_),
    .B1(_12382_));
 sg13g2_mux2_1 _19317_ (.A0(\cpu.dcache.r_data[1][17] ),
    .A1(net1020),
    .S(_12380_),
    .X(_12383_));
 sg13g2_nor2_1 _19318_ (.A(_12377_),
    .B(_12383_),
    .Y(_12384_));
 sg13g2_a21oi_1 _19319_ (.A1(net766),
    .A2(net57),
    .Y(_00353_),
    .B1(_12384_));
 sg13g2_mux2_1 _19320_ (.A0(\cpu.dcache.r_data[1][18] ),
    .A1(net1019),
    .S(_12380_),
    .X(_12385_));
 sg13g2_nor2_1 _19321_ (.A(_12377_),
    .B(_12385_),
    .Y(_12386_));
 sg13g2_a21oi_1 _19322_ (.A1(net765),
    .A2(net57),
    .Y(_00354_),
    .B1(_12386_));
 sg13g2_nor2b_1 _19323_ (.A(_12380_),
    .B_N(\cpu.dcache.r_data[1][19] ),
    .Y(_12387_));
 sg13g2_a21oi_1 _19324_ (.A1(net1026),
    .A2(_12380_),
    .Y(_12388_),
    .B1(_12387_));
 sg13g2_nand2_1 _19325_ (.Y(_12389_),
    .A(net1024),
    .B(net57));
 sg13g2_o21ai_1 _19326_ (.B1(_12389_),
    .Y(_00355_),
    .A1(net57),
    .A2(_12388_));
 sg13g2_mux2_1 _19327_ (.A0(\cpu.dcache.r_data[1][1] ),
    .A1(net1020),
    .S(_12347_),
    .X(_12390_));
 sg13g2_nor2_1 _19328_ (.A(_12344_),
    .B(_12390_),
    .Y(_12391_));
 sg13g2_a21oi_1 _19329_ (.A1(net766),
    .A2(net59),
    .Y(_00356_),
    .B1(_12391_));
 sg13g2_nor2_1 _19330_ (.A(net699),
    .B(_12254_),
    .Y(_12392_));
 sg13g2_buf_2 _19331_ (.A(_12392_),
    .X(_12393_));
 sg13g2_nor2b_1 _19332_ (.A(_12393_),
    .B_N(\cpu.dcache.r_data[1][20] ),
    .Y(_12394_));
 sg13g2_a21oi_1 _19333_ (.A1(net1023),
    .A2(_12393_),
    .Y(_12395_),
    .B1(_12394_));
 sg13g2_nand2_1 _19334_ (.Y(_12396_),
    .A(net1022),
    .B(net57));
 sg13g2_o21ai_1 _19335_ (.B1(_12396_),
    .Y(_00357_),
    .A1(net57),
    .A2(_12395_));
 sg13g2_mux2_1 _19336_ (.A0(\cpu.dcache.r_data[1][21] ),
    .A1(net1020),
    .S(_12393_),
    .X(_12397_));
 sg13g2_nor2_1 _19337_ (.A(_12377_),
    .B(_12397_),
    .Y(_12398_));
 sg13g2_a21oi_1 _19338_ (.A1(net764),
    .A2(_12378_),
    .Y(_00358_),
    .B1(_12398_));
 sg13g2_mux2_1 _19339_ (.A0(\cpu.dcache.r_data[1][22] ),
    .A1(net1019),
    .S(_12393_),
    .X(_12399_));
 sg13g2_nor2_1 _19340_ (.A(_12377_),
    .B(_12399_),
    .Y(_12400_));
 sg13g2_a21oi_1 _19341_ (.A1(net763),
    .A2(net57),
    .Y(_00359_),
    .B1(_12400_));
 sg13g2_mux2_1 _19342_ (.A0(\cpu.dcache.r_data[1][23] ),
    .A1(net1107),
    .S(_12393_),
    .X(_12401_));
 sg13g2_nor2_1 _19343_ (.A(_12377_),
    .B(_12401_),
    .Y(_12402_));
 sg13g2_a21oi_1 _19344_ (.A1(net762),
    .A2(_12378_),
    .Y(_00360_),
    .B1(_12402_));
 sg13g2_nand3b_1 _19345_ (.B(_12350_),
    .C(_12134_),
    .Y(_12403_),
    .A_N(_12284_));
 sg13g2_buf_2 _19346_ (.A(_12403_),
    .X(_12404_));
 sg13g2_nor2_1 _19347_ (.A(_12339_),
    .B(_12404_),
    .Y(_12405_));
 sg13g2_buf_2 _19348_ (.A(_12405_),
    .X(_12406_));
 sg13g2_buf_1 _19349_ (.A(_12406_),
    .X(_12407_));
 sg13g2_nor2_1 _19350_ (.A(net699),
    .B(_12131_),
    .Y(_12408_));
 sg13g2_buf_1 _19351_ (.A(_12408_),
    .X(_12409_));
 sg13g2_nor2b_1 _19352_ (.A(net552),
    .B_N(\cpu.dcache.r_data[1][24] ),
    .Y(_12410_));
 sg13g2_a21oi_1 _19353_ (.A1(net1023),
    .A2(net552),
    .Y(_12411_),
    .B1(_12410_));
 sg13g2_nand2_1 _19354_ (.Y(_12412_),
    .A(_12282_),
    .B(net56));
 sg13g2_o21ai_1 _19355_ (.B1(_12412_),
    .Y(_00361_),
    .A1(net56),
    .A2(_12411_));
 sg13g2_nor2b_1 _19356_ (.A(net552),
    .B_N(\cpu.dcache.r_data[1][25] ),
    .Y(_12413_));
 sg13g2_a21oi_1 _19357_ (.A1(net1018),
    .A2(net552),
    .Y(_12414_),
    .B1(_12413_));
 sg13g2_nand2_1 _19358_ (.Y(_12415_),
    .A(_12291_),
    .B(net56));
 sg13g2_o21ai_1 _19359_ (.B1(_12415_),
    .Y(_00362_),
    .A1(net56),
    .A2(_12414_));
 sg13g2_nor2b_1 _19360_ (.A(net552),
    .B_N(\cpu.dcache.r_data[1][26] ),
    .Y(_12416_));
 sg13g2_a21oi_1 _19361_ (.A1(net1027),
    .A2(net552),
    .Y(_12417_),
    .B1(_12416_));
 sg13g2_nand2_1 _19362_ (.Y(_12418_),
    .A(net433),
    .B(_12406_));
 sg13g2_o21ai_1 _19363_ (.B1(_12418_),
    .Y(_00363_),
    .A1(_12407_),
    .A2(_12417_));
 sg13g2_nor2b_1 _19364_ (.A(net552),
    .B_N(\cpu.dcache.r_data[1][27] ),
    .Y(_12419_));
 sg13g2_a21oi_1 _19365_ (.A1(net1026),
    .A2(net552),
    .Y(_12420_),
    .B1(_12419_));
 sg13g2_nand2_1 _19366_ (.Y(_12421_),
    .A(_12294_),
    .B(_12406_));
 sg13g2_o21ai_1 _19367_ (.B1(_12421_),
    .Y(_00364_),
    .A1(_12407_),
    .A2(_12420_));
 sg13g2_buf_1 _19368_ (.A(_12250_),
    .X(_12422_));
 sg13g2_nor2_2 _19369_ (.A(net623),
    .B(_12298_),
    .Y(_12423_));
 sg13g2_mux2_1 _19370_ (.A0(\cpu.dcache.r_data[1][28] ),
    .A1(net1017),
    .S(_12423_),
    .X(_12424_));
 sg13g2_nor2_1 _19371_ (.A(_12406_),
    .B(_12424_),
    .Y(_12425_));
 sg13g2_a21oi_1 _19372_ (.A1(_12295_),
    .A2(net56),
    .Y(_00365_),
    .B1(_12425_));
 sg13g2_mux2_1 _19373_ (.A0(\cpu.dcache.r_data[1][29] ),
    .A1(_12304_),
    .S(_12423_),
    .X(_12426_));
 sg13g2_nor2_1 _19374_ (.A(_12406_),
    .B(_12426_),
    .Y(_12427_));
 sg13g2_a21oi_1 _19375_ (.A1(net427),
    .A2(net56),
    .Y(_00366_),
    .B1(_12427_));
 sg13g2_mux2_1 _19376_ (.A0(\cpu.dcache.r_data[1][2] ),
    .A1(net1019),
    .S(_12347_),
    .X(_12428_));
 sg13g2_nor2_1 _19377_ (.A(_12344_),
    .B(_12428_),
    .Y(_12429_));
 sg13g2_a21oi_1 _19378_ (.A1(net765),
    .A2(net59),
    .Y(_00367_),
    .B1(_12429_));
 sg13g2_mux2_1 _19379_ (.A0(\cpu.dcache.r_data[1][30] ),
    .A1(_12310_),
    .S(_12423_),
    .X(_12430_));
 sg13g2_nor2_1 _19380_ (.A(_12406_),
    .B(_12430_),
    .Y(_12431_));
 sg13g2_a21oi_1 _19381_ (.A1(net384),
    .A2(net56),
    .Y(_00368_),
    .B1(_12431_));
 sg13g2_mux2_1 _19382_ (.A0(\cpu.dcache.r_data[1][31] ),
    .A1(net1107),
    .S(_12423_),
    .X(_12432_));
 sg13g2_nor2_1 _19383_ (.A(_12406_),
    .B(_12432_),
    .Y(_12433_));
 sg13g2_a21oi_1 _19384_ (.A1(net383),
    .A2(net56),
    .Y(_00369_),
    .B1(_12433_));
 sg13g2_buf_1 _19385_ (.A(net1110),
    .X(_12434_));
 sg13g2_nor2b_1 _19386_ (.A(_12347_),
    .B_N(\cpu.dcache.r_data[1][3] ),
    .Y(_12435_));
 sg13g2_a21oi_1 _19387_ (.A1(net1016),
    .A2(_12347_),
    .Y(_12436_),
    .B1(_12435_));
 sg13g2_nand2_1 _19388_ (.Y(_12437_),
    .A(net1024),
    .B(net59));
 sg13g2_o21ai_1 _19389_ (.B1(_12437_),
    .Y(_00370_),
    .A1(net59),
    .A2(_12436_));
 sg13g2_nor2_1 _19390_ (.A(net699),
    .B(_12320_),
    .Y(_12438_));
 sg13g2_buf_2 _19391_ (.A(_12438_),
    .X(_12439_));
 sg13g2_nor2b_1 _19392_ (.A(_12439_),
    .B_N(\cpu.dcache.r_data[1][4] ),
    .Y(_12440_));
 sg13g2_a21oi_1 _19393_ (.A1(net1023),
    .A2(_12439_),
    .Y(_12441_),
    .B1(_12440_));
 sg13g2_nand2_1 _19394_ (.Y(_12442_),
    .A(net1022),
    .B(_12345_));
 sg13g2_o21ai_1 _19395_ (.B1(_12442_),
    .Y(_00371_),
    .A1(_12345_),
    .A2(_12441_));
 sg13g2_mux2_1 _19396_ (.A0(\cpu.dcache.r_data[1][5] ),
    .A1(net1020),
    .S(_12439_),
    .X(_12443_));
 sg13g2_nor2_1 _19397_ (.A(_12344_),
    .B(_12443_),
    .Y(_12444_));
 sg13g2_a21oi_1 _19398_ (.A1(_12262_),
    .A2(net59),
    .Y(_00372_),
    .B1(_12444_));
 sg13g2_mux2_1 _19399_ (.A0(\cpu.dcache.r_data[1][6] ),
    .A1(net1019),
    .S(_12439_),
    .X(_12445_));
 sg13g2_nor2_1 _19400_ (.A(_12344_),
    .B(_12445_),
    .Y(_12446_));
 sg13g2_a21oi_1 _19401_ (.A1(net763),
    .A2(net59),
    .Y(_00373_),
    .B1(_12446_));
 sg13g2_buf_1 _19402_ (.A(net1110),
    .X(_12447_));
 sg13g2_mux2_1 _19403_ (.A0(\cpu.dcache.r_data[1][7] ),
    .A1(net1015),
    .S(_12439_),
    .X(_12448_));
 sg13g2_nor2_1 _19404_ (.A(_12344_),
    .B(_12448_),
    .Y(_12449_));
 sg13g2_a21oi_1 _19405_ (.A1(net762),
    .A2(net59),
    .Y(_00374_),
    .B1(_12449_));
 sg13g2_buf_1 _19406_ (.A(net1106),
    .X(_12450_));
 sg13g2_nor2b_1 _19407_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[1][8] ),
    .Y(_12451_));
 sg13g2_a21oi_1 _19408_ (.A1(net1014),
    .A2(_12357_),
    .Y(_12452_),
    .B1(_12451_));
 sg13g2_nand2_1 _19409_ (.Y(_12453_),
    .A(net431),
    .B(_12354_));
 sg13g2_o21ai_1 _19410_ (.B1(_12453_),
    .Y(_00375_),
    .A1(net58),
    .A2(_12452_));
 sg13g2_nor2b_1 _19411_ (.A(_12357_),
    .B_N(\cpu.dcache.r_data[1][9] ),
    .Y(_12454_));
 sg13g2_a21oi_1 _19412_ (.A1(net1018),
    .A2(_12357_),
    .Y(_12455_),
    .B1(_12454_));
 sg13g2_nand2_1 _19413_ (.Y(_12456_),
    .A(net430),
    .B(_12354_));
 sg13g2_o21ai_1 _19414_ (.B1(_12456_),
    .Y(_00376_),
    .A1(_12355_),
    .A2(_12455_));
 sg13g2_buf_1 _19415_ (.A(_09552_),
    .X(_12457_));
 sg13g2_nor2_1 _19416_ (.A(net675),
    .B(_12342_),
    .Y(_12458_));
 sg13g2_buf_1 _19417_ (.A(_12458_),
    .X(_12459_));
 sg13g2_buf_1 _19418_ (.A(_12459_),
    .X(_12460_));
 sg13g2_nor2_1 _19419_ (.A(net675),
    .B(_12155_),
    .Y(_12461_));
 sg13g2_buf_2 _19420_ (.A(_12461_),
    .X(_12462_));
 sg13g2_mux2_1 _19421_ (.A0(\cpu.dcache.r_data[2][0] ),
    .A1(net1017),
    .S(_12462_),
    .X(_12463_));
 sg13g2_nor2_1 _19422_ (.A(_12459_),
    .B(_12463_),
    .Y(_12464_));
 sg13g2_a21oi_1 _19423_ (.A1(net797),
    .A2(net55),
    .Y(_00377_),
    .B1(_12464_));
 sg13g2_nor2_1 _19424_ (.A(net675),
    .B(_12352_),
    .Y(_12465_));
 sg13g2_buf_2 _19425_ (.A(_12465_),
    .X(_12466_));
 sg13g2_buf_1 _19426_ (.A(_12466_),
    .X(_12467_));
 sg13g2_nor2_1 _19427_ (.A(net675),
    .B(_12170_),
    .Y(_12468_));
 sg13g2_buf_2 _19428_ (.A(_12468_),
    .X(_12469_));
 sg13g2_nor2b_1 _19429_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[2][10] ),
    .Y(_12470_));
 sg13g2_a21oi_1 _19430_ (.A1(net1027),
    .A2(_12469_),
    .Y(_12471_),
    .B1(_12470_));
 sg13g2_nand2_1 _19431_ (.Y(_12472_),
    .A(net433),
    .B(net54));
 sg13g2_o21ai_1 _19432_ (.B1(_12472_),
    .Y(_00378_),
    .A1(net54),
    .A2(_12471_));
 sg13g2_nor2b_1 _19433_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[2][11] ),
    .Y(_12473_));
 sg13g2_a21oi_1 _19434_ (.A1(net1016),
    .A2(_12469_),
    .Y(_12474_),
    .B1(_12473_));
 sg13g2_nand2_1 _19435_ (.Y(_12475_),
    .A(net429),
    .B(_12467_));
 sg13g2_o21ai_1 _19436_ (.B1(_12475_),
    .Y(_00379_),
    .A1(net54),
    .A2(_12474_));
 sg13g2_nor2_2 _19437_ (.A(net675),
    .B(_12198_),
    .Y(_12476_));
 sg13g2_mux2_1 _19438_ (.A0(\cpu.dcache.r_data[2][12] ),
    .A1(net1017),
    .S(_12476_),
    .X(_12477_));
 sg13g2_nor2_1 _19439_ (.A(_12466_),
    .B(_12477_),
    .Y(_12478_));
 sg13g2_a21oi_1 _19440_ (.A1(net428),
    .A2(net54),
    .Y(_00380_),
    .B1(_12478_));
 sg13g2_mux2_1 _19441_ (.A0(\cpu.dcache.r_data[2][13] ),
    .A1(_12304_),
    .S(_12476_),
    .X(_12479_));
 sg13g2_nor2_1 _19442_ (.A(_12466_),
    .B(_12479_),
    .Y(_12480_));
 sg13g2_a21oi_1 _19443_ (.A1(net427),
    .A2(net54),
    .Y(_00381_),
    .B1(_12480_));
 sg13g2_mux2_1 _19444_ (.A0(\cpu.dcache.r_data[2][14] ),
    .A1(_12310_),
    .S(_12476_),
    .X(_12481_));
 sg13g2_nor2_1 _19445_ (.A(_12466_),
    .B(_12481_),
    .Y(_12482_));
 sg13g2_a21oi_1 _19446_ (.A1(net384),
    .A2(net54),
    .Y(_00382_),
    .B1(_12482_));
 sg13g2_mux2_1 _19447_ (.A0(\cpu.dcache.r_data[2][15] ),
    .A1(net1015),
    .S(_12476_),
    .X(_12483_));
 sg13g2_nor2_1 _19448_ (.A(_12466_),
    .B(_12483_),
    .Y(_12484_));
 sg13g2_a21oi_1 _19449_ (.A1(net383),
    .A2(net54),
    .Y(_00383_),
    .B1(_12484_));
 sg13g2_nor2_1 _19450_ (.A(net675),
    .B(_12375_),
    .Y(_12485_));
 sg13g2_buf_2 _19451_ (.A(_12485_),
    .X(_12486_));
 sg13g2_buf_1 _19452_ (.A(_12486_),
    .X(_12487_));
 sg13g2_nor2_1 _19453_ (.A(_09552_),
    .B(_12230_),
    .Y(_12488_));
 sg13g2_buf_2 _19454_ (.A(_12488_),
    .X(_12489_));
 sg13g2_mux2_1 _19455_ (.A0(\cpu.dcache.r_data[2][16] ),
    .A1(net1017),
    .S(_12489_),
    .X(_12490_));
 sg13g2_nor2_1 _19456_ (.A(_12486_),
    .B(_12490_),
    .Y(_12491_));
 sg13g2_a21oi_1 _19457_ (.A1(net797),
    .A2(net53),
    .Y(_00384_),
    .B1(_12491_));
 sg13g2_mux2_1 _19458_ (.A0(\cpu.dcache.r_data[2][17] ),
    .A1(net1020),
    .S(_12489_),
    .X(_12492_));
 sg13g2_nor2_1 _19459_ (.A(_12486_),
    .B(_12492_),
    .Y(_12493_));
 sg13g2_a21oi_1 _19460_ (.A1(net766),
    .A2(_12487_),
    .Y(_00385_),
    .B1(_12493_));
 sg13g2_mux2_1 _19461_ (.A0(\cpu.dcache.r_data[2][18] ),
    .A1(net1019),
    .S(_12489_),
    .X(_12494_));
 sg13g2_nor2_1 _19462_ (.A(_12486_),
    .B(_12494_),
    .Y(_12495_));
 sg13g2_a21oi_1 _19463_ (.A1(net765),
    .A2(net53),
    .Y(_00386_),
    .B1(_12495_));
 sg13g2_nor2b_1 _19464_ (.A(_12489_),
    .B_N(\cpu.dcache.r_data[2][19] ),
    .Y(_12496_));
 sg13g2_a21oi_1 _19465_ (.A1(net1016),
    .A2(_12489_),
    .Y(_12497_),
    .B1(_12496_));
 sg13g2_nand2_1 _19466_ (.Y(_12498_),
    .A(net1024),
    .B(_12487_));
 sg13g2_o21ai_1 _19467_ (.B1(_12498_),
    .Y(_00387_),
    .A1(net53),
    .A2(_12497_));
 sg13g2_buf_1 _19468_ (.A(net1105),
    .X(_12499_));
 sg13g2_mux2_1 _19469_ (.A0(\cpu.dcache.r_data[2][1] ),
    .A1(net1013),
    .S(_12462_),
    .X(_12500_));
 sg13g2_nor2_1 _19470_ (.A(_12459_),
    .B(_12500_),
    .Y(_12501_));
 sg13g2_a21oi_1 _19471_ (.A1(_12237_),
    .A2(net55),
    .Y(_00388_),
    .B1(_12501_));
 sg13g2_nor2_1 _19472_ (.A(_09552_),
    .B(_12254_),
    .Y(_12502_));
 sg13g2_buf_2 _19473_ (.A(_12502_),
    .X(_12503_));
 sg13g2_nor2b_1 _19474_ (.A(_12503_),
    .B_N(\cpu.dcache.r_data[2][20] ),
    .Y(_12504_));
 sg13g2_a21oi_1 _19475_ (.A1(net1014),
    .A2(_12503_),
    .Y(_12505_),
    .B1(_12504_));
 sg13g2_nand2_1 _19476_ (.Y(_12506_),
    .A(net1022),
    .B(net53));
 sg13g2_o21ai_1 _19477_ (.B1(_12506_),
    .Y(_00389_),
    .A1(net53),
    .A2(_12505_));
 sg13g2_mux2_1 _19478_ (.A0(\cpu.dcache.r_data[2][21] ),
    .A1(net1013),
    .S(_12503_),
    .X(_12507_));
 sg13g2_nor2_1 _19479_ (.A(_12486_),
    .B(_12507_),
    .Y(_12508_));
 sg13g2_a21oi_1 _19480_ (.A1(net764),
    .A2(net53),
    .Y(_00390_),
    .B1(_12508_));
 sg13g2_buf_1 _19481_ (.A(net1111),
    .X(_12509_));
 sg13g2_mux2_1 _19482_ (.A0(\cpu.dcache.r_data[2][22] ),
    .A1(net1012),
    .S(_12503_),
    .X(_12510_));
 sg13g2_nor2_1 _19483_ (.A(_12486_),
    .B(_12510_),
    .Y(_12511_));
 sg13g2_a21oi_1 _19484_ (.A1(net763),
    .A2(net53),
    .Y(_00391_),
    .B1(_12511_));
 sg13g2_mux2_1 _19485_ (.A0(\cpu.dcache.r_data[2][23] ),
    .A1(net1015),
    .S(_12503_),
    .X(_12512_));
 sg13g2_nor2_1 _19486_ (.A(_12486_),
    .B(_12512_),
    .Y(_12513_));
 sg13g2_a21oi_1 _19487_ (.A1(net762),
    .A2(net53),
    .Y(_00392_),
    .B1(_12513_));
 sg13g2_nor2_1 _19488_ (.A(net675),
    .B(_12404_),
    .Y(_12514_));
 sg13g2_buf_2 _19489_ (.A(_12514_),
    .X(_12515_));
 sg13g2_buf_1 _19490_ (.A(_12515_),
    .X(_12516_));
 sg13g2_nor2_1 _19491_ (.A(_12457_),
    .B(_12131_),
    .Y(_12517_));
 sg13g2_buf_1 _19492_ (.A(_12517_),
    .X(_12518_));
 sg13g2_nor2b_1 _19493_ (.A(net551),
    .B_N(\cpu.dcache.r_data[2][24] ),
    .Y(_12519_));
 sg13g2_a21oi_1 _19494_ (.A1(net1014),
    .A2(net551),
    .Y(_12520_),
    .B1(_12519_));
 sg13g2_nand2_1 _19495_ (.Y(_12521_),
    .A(_12282_),
    .B(net52));
 sg13g2_o21ai_1 _19496_ (.B1(_12521_),
    .Y(_00393_),
    .A1(_12516_),
    .A2(_12520_));
 sg13g2_nor2b_1 _19497_ (.A(net551),
    .B_N(\cpu.dcache.r_data[2][25] ),
    .Y(_12522_));
 sg13g2_a21oi_1 _19498_ (.A1(net1018),
    .A2(net551),
    .Y(_12523_),
    .B1(_12522_));
 sg13g2_nand2_1 _19499_ (.Y(_12524_),
    .A(_12291_),
    .B(net52));
 sg13g2_o21ai_1 _19500_ (.B1(_12524_),
    .Y(_00394_),
    .A1(net52),
    .A2(_12523_));
 sg13g2_nor2b_1 _19501_ (.A(net551),
    .B_N(\cpu.dcache.r_data[2][26] ),
    .Y(_12525_));
 sg13g2_a21oi_1 _19502_ (.A1(net1027),
    .A2(net551),
    .Y(_12526_),
    .B1(_12525_));
 sg13g2_nand2_1 _19503_ (.Y(_12527_),
    .A(net433),
    .B(_12515_));
 sg13g2_o21ai_1 _19504_ (.B1(_12527_),
    .Y(_00395_),
    .A1(_12516_),
    .A2(_12526_));
 sg13g2_nor2b_1 _19505_ (.A(net551),
    .B_N(\cpu.dcache.r_data[2][27] ),
    .Y(_12528_));
 sg13g2_a21oi_1 _19506_ (.A1(net1016),
    .A2(net551),
    .Y(_12529_),
    .B1(_12528_));
 sg13g2_nand2_1 _19507_ (.Y(_12530_),
    .A(_12294_),
    .B(_12515_));
 sg13g2_o21ai_1 _19508_ (.B1(_12530_),
    .Y(_00396_),
    .A1(net52),
    .A2(_12529_));
 sg13g2_nor2_2 _19509_ (.A(net675),
    .B(_12298_),
    .Y(_12531_));
 sg13g2_mux2_1 _19510_ (.A0(\cpu.dcache.r_data[2][28] ),
    .A1(net1017),
    .S(_12531_),
    .X(_12532_));
 sg13g2_nor2_1 _19511_ (.A(_12515_),
    .B(_12532_),
    .Y(_12533_));
 sg13g2_a21oi_1 _19512_ (.A1(net428),
    .A2(net52),
    .Y(_00397_),
    .B1(_12533_));
 sg13g2_mux2_1 _19513_ (.A0(\cpu.dcache.r_data[2][29] ),
    .A1(_12499_),
    .S(_12531_),
    .X(_12534_));
 sg13g2_nor2_1 _19514_ (.A(_12515_),
    .B(_12534_),
    .Y(_12535_));
 sg13g2_a21oi_1 _19515_ (.A1(_12302_),
    .A2(net52),
    .Y(_00398_),
    .B1(_12535_));
 sg13g2_mux2_1 _19516_ (.A0(\cpu.dcache.r_data[2][2] ),
    .A1(_12509_),
    .S(_12462_),
    .X(_12536_));
 sg13g2_nor2_1 _19517_ (.A(_12459_),
    .B(_12536_),
    .Y(_12537_));
 sg13g2_a21oi_1 _19518_ (.A1(_12241_),
    .A2(_12460_),
    .Y(_00399_),
    .B1(_12537_));
 sg13g2_mux2_1 _19519_ (.A0(\cpu.dcache.r_data[2][30] ),
    .A1(net1012),
    .S(_12531_),
    .X(_12538_));
 sg13g2_nor2_1 _19520_ (.A(_12515_),
    .B(_12538_),
    .Y(_12539_));
 sg13g2_a21oi_1 _19521_ (.A1(_12309_),
    .A2(net52),
    .Y(_00400_),
    .B1(_12539_));
 sg13g2_mux2_1 _19522_ (.A0(\cpu.dcache.r_data[2][31] ),
    .A1(net1015),
    .S(_12531_),
    .X(_12540_));
 sg13g2_nor2_1 _19523_ (.A(_12515_),
    .B(_12540_),
    .Y(_12541_));
 sg13g2_a21oi_1 _19524_ (.A1(_12313_),
    .A2(net52),
    .Y(_00401_),
    .B1(_12541_));
 sg13g2_nor2b_1 _19525_ (.A(_12462_),
    .B_N(\cpu.dcache.r_data[2][3] ),
    .Y(_12542_));
 sg13g2_a21oi_1 _19526_ (.A1(net1016),
    .A2(_12462_),
    .Y(_12543_),
    .B1(_12542_));
 sg13g2_nand2_1 _19527_ (.Y(_12544_),
    .A(_12246_),
    .B(net55));
 sg13g2_o21ai_1 _19528_ (.B1(_12544_),
    .Y(_00402_),
    .A1(net55),
    .A2(_12543_));
 sg13g2_nor2_1 _19529_ (.A(_09552_),
    .B(_12320_),
    .Y(_12545_));
 sg13g2_buf_2 _19530_ (.A(_12545_),
    .X(_12546_));
 sg13g2_nor2b_1 _19531_ (.A(_12546_),
    .B_N(\cpu.dcache.r_data[2][4] ),
    .Y(_12547_));
 sg13g2_a21oi_1 _19532_ (.A1(net1014),
    .A2(_12546_),
    .Y(_12548_),
    .B1(_12547_));
 sg13g2_buf_1 _19533_ (.A(_09999_),
    .X(_12549_));
 sg13g2_nand2_1 _19534_ (.Y(_12550_),
    .A(net1011),
    .B(net55));
 sg13g2_o21ai_1 _19535_ (.B1(_12550_),
    .Y(_00403_),
    .A1(net55),
    .A2(_12548_));
 sg13g2_mux2_1 _19536_ (.A0(\cpu.dcache.r_data[2][5] ),
    .A1(net1013),
    .S(_12546_),
    .X(_12551_));
 sg13g2_nor2_1 _19537_ (.A(_12459_),
    .B(_12551_),
    .Y(_12552_));
 sg13g2_a21oi_1 _19538_ (.A1(_12262_),
    .A2(net55),
    .Y(_00404_),
    .B1(_12552_));
 sg13g2_mux2_1 _19539_ (.A0(\cpu.dcache.r_data[2][6] ),
    .A1(net1012),
    .S(_12546_),
    .X(_12553_));
 sg13g2_nor2_1 _19540_ (.A(_12459_),
    .B(_12553_),
    .Y(_12554_));
 sg13g2_a21oi_1 _19541_ (.A1(_12266_),
    .A2(_12460_),
    .Y(_00405_),
    .B1(_12554_));
 sg13g2_mux2_1 _19542_ (.A0(\cpu.dcache.r_data[2][7] ),
    .A1(net1015),
    .S(_12546_),
    .X(_12555_));
 sg13g2_nor2_1 _19543_ (.A(_12459_),
    .B(_12555_),
    .Y(_12556_));
 sg13g2_a21oi_1 _19544_ (.A1(net762),
    .A2(net55),
    .Y(_00406_),
    .B1(_12556_));
 sg13g2_nor2b_1 _19545_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[2][8] ),
    .Y(_12557_));
 sg13g2_a21oi_1 _19546_ (.A1(net1014),
    .A2(_12469_),
    .Y(_12558_),
    .B1(_12557_));
 sg13g2_nand2_1 _19547_ (.Y(_12559_),
    .A(net431),
    .B(_12466_));
 sg13g2_o21ai_1 _19548_ (.B1(_12559_),
    .Y(_00407_),
    .A1(net54),
    .A2(_12558_));
 sg13g2_nor2b_1 _19549_ (.A(_12469_),
    .B_N(\cpu.dcache.r_data[2][9] ),
    .Y(_12560_));
 sg13g2_a21oi_1 _19550_ (.A1(net1018),
    .A2(_12469_),
    .Y(_12561_),
    .B1(_12560_));
 sg13g2_nand2_1 _19551_ (.Y(_12562_),
    .A(net430),
    .B(_12466_));
 sg13g2_o21ai_1 _19552_ (.B1(_12562_),
    .Y(_00408_),
    .A1(_12467_),
    .A2(_12561_));
 sg13g2_buf_1 _19553_ (.A(net716),
    .X(_12563_));
 sg13g2_nand2_1 _19554_ (.Y(_12564_),
    .A(net622),
    .B(_09357_));
 sg13g2_buf_1 _19555_ (.A(_12564_),
    .X(_12565_));
 sg13g2_buf_1 _19556_ (.A(_12565_),
    .X(_12566_));
 sg13g2_nor2_1 _19557_ (.A(net426),
    .B(_12342_),
    .Y(_12567_));
 sg13g2_buf_1 _19558_ (.A(_12567_),
    .X(_12568_));
 sg13g2_buf_1 _19559_ (.A(_12568_),
    .X(_12569_));
 sg13g2_nor2_1 _19560_ (.A(net426),
    .B(_12155_),
    .Y(_12570_));
 sg13g2_buf_2 _19561_ (.A(_12570_),
    .X(_12571_));
 sg13g2_mux2_1 _19562_ (.A0(\cpu.dcache.r_data[3][0] ),
    .A1(net1017),
    .S(_12571_),
    .X(_12572_));
 sg13g2_nor2_1 _19563_ (.A(_12568_),
    .B(_12572_),
    .Y(_12573_));
 sg13g2_a21oi_1 _19564_ (.A1(net797),
    .A2(net51),
    .Y(_00409_),
    .B1(_12573_));
 sg13g2_nor2_1 _19565_ (.A(net426),
    .B(_12352_),
    .Y(_12574_));
 sg13g2_buf_2 _19566_ (.A(_12574_),
    .X(_12575_));
 sg13g2_buf_1 _19567_ (.A(_12575_),
    .X(_12576_));
 sg13g2_nor2_1 _19568_ (.A(_12566_),
    .B(_12170_),
    .Y(_12577_));
 sg13g2_buf_2 _19569_ (.A(_12577_),
    .X(_12578_));
 sg13g2_nor2b_1 _19570_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[3][10] ),
    .Y(_12579_));
 sg13g2_a21oi_1 _19571_ (.A1(net1027),
    .A2(_12578_),
    .Y(_12580_),
    .B1(_12579_));
 sg13g2_nand2_1 _19572_ (.Y(_12581_),
    .A(net433),
    .B(net50));
 sg13g2_o21ai_1 _19573_ (.B1(_12581_),
    .Y(_00410_),
    .A1(_12576_),
    .A2(_12580_));
 sg13g2_nor2b_1 _19574_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[3][11] ),
    .Y(_12582_));
 sg13g2_a21oi_1 _19575_ (.A1(net1016),
    .A2(_12578_),
    .Y(_12583_),
    .B1(_12582_));
 sg13g2_nand2_1 _19576_ (.Y(_12584_),
    .A(net429),
    .B(net50));
 sg13g2_o21ai_1 _19577_ (.B1(_12584_),
    .Y(_00411_),
    .A1(net50),
    .A2(_12583_));
 sg13g2_nor2_2 _19578_ (.A(net426),
    .B(_12198_),
    .Y(_12585_));
 sg13g2_mux2_1 _19579_ (.A0(\cpu.dcache.r_data[3][12] ),
    .A1(_12422_),
    .S(_12585_),
    .X(_12586_));
 sg13g2_nor2_1 _19580_ (.A(_12575_),
    .B(_12586_),
    .Y(_12587_));
 sg13g2_a21oi_1 _19581_ (.A1(net428),
    .A2(net50),
    .Y(_00412_),
    .B1(_12587_));
 sg13g2_mux2_1 _19582_ (.A0(\cpu.dcache.r_data[3][13] ),
    .A1(_12499_),
    .S(_12585_),
    .X(_12588_));
 sg13g2_nor2_1 _19583_ (.A(_12575_),
    .B(_12588_),
    .Y(_12589_));
 sg13g2_a21oi_1 _19584_ (.A1(net427),
    .A2(net50),
    .Y(_00413_),
    .B1(_12589_));
 sg13g2_mux2_1 _19585_ (.A0(\cpu.dcache.r_data[3][14] ),
    .A1(net1012),
    .S(_12585_),
    .X(_12590_));
 sg13g2_nor2_1 _19586_ (.A(_12575_),
    .B(_12590_),
    .Y(_12591_));
 sg13g2_a21oi_1 _19587_ (.A1(net384),
    .A2(net50),
    .Y(_00414_),
    .B1(_12591_));
 sg13g2_mux2_1 _19588_ (.A0(\cpu.dcache.r_data[3][15] ),
    .A1(net1015),
    .S(_12585_),
    .X(_12592_));
 sg13g2_nor2_1 _19589_ (.A(_12575_),
    .B(_12592_),
    .Y(_12593_));
 sg13g2_a21oi_1 _19590_ (.A1(net383),
    .A2(net50),
    .Y(_00415_),
    .B1(_12593_));
 sg13g2_nor2_1 _19591_ (.A(net426),
    .B(_12375_),
    .Y(_12594_));
 sg13g2_buf_1 _19592_ (.A(_12594_),
    .X(_12595_));
 sg13g2_buf_1 _19593_ (.A(_12595_),
    .X(_12596_));
 sg13g2_nor2_1 _19594_ (.A(net426),
    .B(_12230_),
    .Y(_12597_));
 sg13g2_buf_2 _19595_ (.A(_12597_),
    .X(_12598_));
 sg13g2_mux2_1 _19596_ (.A0(\cpu.dcache.r_data[3][16] ),
    .A1(net1017),
    .S(_12598_),
    .X(_12599_));
 sg13g2_nor2_1 _19597_ (.A(_12595_),
    .B(_12599_),
    .Y(_12600_));
 sg13g2_a21oi_1 _19598_ (.A1(net797),
    .A2(_12596_),
    .Y(_00416_),
    .B1(_12600_));
 sg13g2_mux2_1 _19599_ (.A0(\cpu.dcache.r_data[3][17] ),
    .A1(net1013),
    .S(_12598_),
    .X(_12601_));
 sg13g2_nor2_1 _19600_ (.A(_12595_),
    .B(_12601_),
    .Y(_12602_));
 sg13g2_a21oi_1 _19601_ (.A1(net766),
    .A2(_12596_),
    .Y(_00417_),
    .B1(_12602_));
 sg13g2_mux2_1 _19602_ (.A0(\cpu.dcache.r_data[3][18] ),
    .A1(net1012),
    .S(_12598_),
    .X(_12603_));
 sg13g2_nor2_1 _19603_ (.A(_12595_),
    .B(_12603_),
    .Y(_12604_));
 sg13g2_a21oi_1 _19604_ (.A1(net765),
    .A2(net49),
    .Y(_00418_),
    .B1(_12604_));
 sg13g2_nor2b_1 _19605_ (.A(_12598_),
    .B_N(\cpu.dcache.r_data[3][19] ),
    .Y(_12605_));
 sg13g2_a21oi_1 _19606_ (.A1(net1016),
    .A2(_12598_),
    .Y(_12606_),
    .B1(_12605_));
 sg13g2_nand2_1 _19607_ (.Y(_12607_),
    .A(_12246_),
    .B(net49));
 sg13g2_o21ai_1 _19608_ (.B1(_12607_),
    .Y(_00419_),
    .A1(net49),
    .A2(_12606_));
 sg13g2_mux2_1 _19609_ (.A0(\cpu.dcache.r_data[3][1] ),
    .A1(net1013),
    .S(_12571_),
    .X(_12608_));
 sg13g2_nor2_1 _19610_ (.A(_12568_),
    .B(_12608_),
    .Y(_12609_));
 sg13g2_a21oi_1 _19611_ (.A1(net766),
    .A2(net51),
    .Y(_00420_),
    .B1(_12609_));
 sg13g2_nor2_1 _19612_ (.A(_12565_),
    .B(_12254_),
    .Y(_12610_));
 sg13g2_buf_2 _19613_ (.A(_12610_),
    .X(_12611_));
 sg13g2_nor2b_1 _19614_ (.A(_12611_),
    .B_N(\cpu.dcache.r_data[3][20] ),
    .Y(_12612_));
 sg13g2_a21oi_1 _19615_ (.A1(net1014),
    .A2(_12611_),
    .Y(_12613_),
    .B1(_12612_));
 sg13g2_nand2_1 _19616_ (.Y(_12614_),
    .A(net1011),
    .B(net49));
 sg13g2_o21ai_1 _19617_ (.B1(_12614_),
    .Y(_00421_),
    .A1(net49),
    .A2(_12613_));
 sg13g2_mux2_1 _19618_ (.A0(\cpu.dcache.r_data[3][21] ),
    .A1(net1013),
    .S(_12611_),
    .X(_12615_));
 sg13g2_nor2_1 _19619_ (.A(_12595_),
    .B(_12615_),
    .Y(_12616_));
 sg13g2_a21oi_1 _19620_ (.A1(net764),
    .A2(net49),
    .Y(_00422_),
    .B1(_12616_));
 sg13g2_mux2_1 _19621_ (.A0(\cpu.dcache.r_data[3][22] ),
    .A1(net1012),
    .S(_12611_),
    .X(_12617_));
 sg13g2_nor2_1 _19622_ (.A(_12595_),
    .B(_12617_),
    .Y(_12618_));
 sg13g2_a21oi_1 _19623_ (.A1(net763),
    .A2(net49),
    .Y(_00423_),
    .B1(_12618_));
 sg13g2_mux2_1 _19624_ (.A0(\cpu.dcache.r_data[3][23] ),
    .A1(net1015),
    .S(_12611_),
    .X(_12619_));
 sg13g2_nor2_1 _19625_ (.A(_12595_),
    .B(_12619_),
    .Y(_12620_));
 sg13g2_a21oi_1 _19626_ (.A1(net762),
    .A2(net49),
    .Y(_00424_),
    .B1(_12620_));
 sg13g2_nor2_1 _19627_ (.A(net426),
    .B(_12404_),
    .Y(_12621_));
 sg13g2_buf_2 _19628_ (.A(_12621_),
    .X(_12622_));
 sg13g2_buf_1 _19629_ (.A(_12622_),
    .X(_12623_));
 sg13g2_nor2_1 _19630_ (.A(_12565_),
    .B(_12131_),
    .Y(_12624_));
 sg13g2_buf_1 _19631_ (.A(_12624_),
    .X(_12625_));
 sg13g2_nor2b_1 _19632_ (.A(net382),
    .B_N(\cpu.dcache.r_data[3][24] ),
    .Y(_12626_));
 sg13g2_a21oi_1 _19633_ (.A1(_12450_),
    .A2(net382),
    .Y(_12627_),
    .B1(_12626_));
 sg13g2_nand2_1 _19634_ (.Y(_12628_),
    .A(net431),
    .B(net48));
 sg13g2_o21ai_1 _19635_ (.B1(_12628_),
    .Y(_00425_),
    .A1(net48),
    .A2(_12627_));
 sg13g2_nor2b_1 _19636_ (.A(net382),
    .B_N(\cpu.dcache.r_data[3][25] ),
    .Y(_12629_));
 sg13g2_a21oi_1 _19637_ (.A1(net1018),
    .A2(net382),
    .Y(_12630_),
    .B1(_12629_));
 sg13g2_nand2_1 _19638_ (.Y(_12631_),
    .A(net430),
    .B(net48));
 sg13g2_o21ai_1 _19639_ (.B1(_12631_),
    .Y(_00426_),
    .A1(net48),
    .A2(_12630_));
 sg13g2_buf_1 _19640_ (.A(_12167_),
    .X(_12632_));
 sg13g2_nor2b_1 _19641_ (.A(net382),
    .B_N(\cpu.dcache.r_data[3][26] ),
    .Y(_12633_));
 sg13g2_a21oi_1 _19642_ (.A1(net1010),
    .A2(net382),
    .Y(_12634_),
    .B1(_12633_));
 sg13g2_nand2_1 _19643_ (.Y(_12635_),
    .A(net433),
    .B(_12622_));
 sg13g2_o21ai_1 _19644_ (.B1(_12635_),
    .Y(_00427_),
    .A1(_12623_),
    .A2(_12634_));
 sg13g2_nor2b_1 _19645_ (.A(net382),
    .B_N(\cpu.dcache.r_data[3][27] ),
    .Y(_12636_));
 sg13g2_a21oi_1 _19646_ (.A1(_12434_),
    .A2(net382),
    .Y(_12637_),
    .B1(_12636_));
 sg13g2_nand2_1 _19647_ (.Y(_12638_),
    .A(net429),
    .B(_12622_));
 sg13g2_o21ai_1 _19648_ (.B1(_12638_),
    .Y(_00428_),
    .A1(_12623_),
    .A2(_12637_));
 sg13g2_nor2_2 _19649_ (.A(net426),
    .B(_12298_),
    .Y(_12639_));
 sg13g2_mux2_1 _19650_ (.A0(\cpu.dcache.r_data[3][28] ),
    .A1(_12422_),
    .S(_12639_),
    .X(_12640_));
 sg13g2_nor2_1 _19651_ (.A(_12622_),
    .B(_12640_),
    .Y(_12641_));
 sg13g2_a21oi_1 _19652_ (.A1(net428),
    .A2(net48),
    .Y(_00429_),
    .B1(_12641_));
 sg13g2_mux2_1 _19653_ (.A0(\cpu.dcache.r_data[3][29] ),
    .A1(net1013),
    .S(_12639_),
    .X(_12642_));
 sg13g2_nor2_1 _19654_ (.A(_12622_),
    .B(_12642_),
    .Y(_12643_));
 sg13g2_a21oi_1 _19655_ (.A1(net427),
    .A2(net48),
    .Y(_00430_),
    .B1(_12643_));
 sg13g2_mux2_1 _19656_ (.A0(\cpu.dcache.r_data[3][2] ),
    .A1(_12509_),
    .S(_12571_),
    .X(_12644_));
 sg13g2_nor2_1 _19657_ (.A(_12568_),
    .B(_12644_),
    .Y(_12645_));
 sg13g2_a21oi_1 _19658_ (.A1(net765),
    .A2(_12569_),
    .Y(_00431_),
    .B1(_12645_));
 sg13g2_mux2_1 _19659_ (.A0(\cpu.dcache.r_data[3][30] ),
    .A1(net1012),
    .S(_12639_),
    .X(_12646_));
 sg13g2_nor2_1 _19660_ (.A(_12622_),
    .B(_12646_),
    .Y(_12647_));
 sg13g2_a21oi_1 _19661_ (.A1(net384),
    .A2(net48),
    .Y(_00432_),
    .B1(_12647_));
 sg13g2_mux2_1 _19662_ (.A0(\cpu.dcache.r_data[3][31] ),
    .A1(_12447_),
    .S(_12639_),
    .X(_12648_));
 sg13g2_nor2_1 _19663_ (.A(_12622_),
    .B(_12648_),
    .Y(_12649_));
 sg13g2_a21oi_1 _19664_ (.A1(net383),
    .A2(net48),
    .Y(_00433_),
    .B1(_12649_));
 sg13g2_nor2b_1 _19665_ (.A(_12571_),
    .B_N(\cpu.dcache.r_data[3][3] ),
    .Y(_12650_));
 sg13g2_a21oi_1 _19666_ (.A1(net1016),
    .A2(_12571_),
    .Y(_12651_),
    .B1(_12650_));
 sg13g2_buf_1 _19667_ (.A(_09992_),
    .X(_12652_));
 sg13g2_nand2_1 _19668_ (.Y(_12653_),
    .A(net1009),
    .B(net51));
 sg13g2_o21ai_1 _19669_ (.B1(_12653_),
    .Y(_00434_),
    .A1(net51),
    .A2(_12651_));
 sg13g2_nor2_1 _19670_ (.A(_12565_),
    .B(_12320_),
    .Y(_12654_));
 sg13g2_buf_2 _19671_ (.A(_12654_),
    .X(_12655_));
 sg13g2_nor2b_1 _19672_ (.A(_12655_),
    .B_N(\cpu.dcache.r_data[3][4] ),
    .Y(_12656_));
 sg13g2_a21oi_1 _19673_ (.A1(net1014),
    .A2(_12655_),
    .Y(_12657_),
    .B1(_12656_));
 sg13g2_nand2_1 _19674_ (.Y(_12658_),
    .A(net1011),
    .B(net51));
 sg13g2_o21ai_1 _19675_ (.B1(_12658_),
    .Y(_00435_),
    .A1(net51),
    .A2(_12657_));
 sg13g2_mux2_1 _19676_ (.A0(\cpu.dcache.r_data[3][5] ),
    .A1(net1013),
    .S(_12655_),
    .X(_12659_));
 sg13g2_nor2_1 _19677_ (.A(_12568_),
    .B(_12659_),
    .Y(_12660_));
 sg13g2_a21oi_1 _19678_ (.A1(net764),
    .A2(net51),
    .Y(_00436_),
    .B1(_12660_));
 sg13g2_mux2_1 _19679_ (.A0(\cpu.dcache.r_data[3][6] ),
    .A1(net1012),
    .S(_12655_),
    .X(_12661_));
 sg13g2_nor2_1 _19680_ (.A(_12568_),
    .B(_12661_),
    .Y(_12662_));
 sg13g2_a21oi_1 _19681_ (.A1(net763),
    .A2(_12569_),
    .Y(_00437_),
    .B1(_12662_));
 sg13g2_mux2_1 _19682_ (.A0(\cpu.dcache.r_data[3][7] ),
    .A1(net1015),
    .S(_12655_),
    .X(_12663_));
 sg13g2_nor2_1 _19683_ (.A(_12568_),
    .B(_12663_),
    .Y(_12664_));
 sg13g2_a21oi_1 _19684_ (.A1(net762),
    .A2(net51),
    .Y(_00438_),
    .B1(_12664_));
 sg13g2_nor2b_1 _19685_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[3][8] ),
    .Y(_12665_));
 sg13g2_a21oi_1 _19686_ (.A1(_12450_),
    .A2(_12578_),
    .Y(_12666_),
    .B1(_12665_));
 sg13g2_nand2_1 _19687_ (.Y(_12667_),
    .A(net431),
    .B(_12575_));
 sg13g2_o21ai_1 _19688_ (.B1(_12667_),
    .Y(_00439_),
    .A1(_12576_),
    .A2(_12666_));
 sg13g2_buf_1 _19689_ (.A(_12303_),
    .X(_12668_));
 sg13g2_nor2b_1 _19690_ (.A(_12578_),
    .B_N(\cpu.dcache.r_data[3][9] ),
    .Y(_12669_));
 sg13g2_a21oi_1 _19691_ (.A1(net1008),
    .A2(_12578_),
    .Y(_12670_),
    .B1(_12669_));
 sg13g2_nand2_1 _19692_ (.Y(_12671_),
    .A(net430),
    .B(_12575_));
 sg13g2_o21ai_1 _19693_ (.B1(_12671_),
    .Y(_00440_),
    .A1(net50),
    .A2(_12670_));
 sg13g2_buf_1 _19694_ (.A(_10031_),
    .X(_12672_));
 sg13g2_nor2_1 _19695_ (.A(_12672_),
    .B(_12342_),
    .Y(_12673_));
 sg13g2_buf_2 _19696_ (.A(_12673_),
    .X(_12674_));
 sg13g2_buf_1 _19697_ (.A(_12674_),
    .X(_12675_));
 sg13g2_nor2_1 _19698_ (.A(_12672_),
    .B(_12155_),
    .Y(_12676_));
 sg13g2_buf_2 _19699_ (.A(_12676_),
    .X(_12677_));
 sg13g2_mux2_1 _19700_ (.A0(\cpu.dcache.r_data[4][0] ),
    .A1(net1017),
    .S(_12677_),
    .X(_12678_));
 sg13g2_nor2_1 _19701_ (.A(_12674_),
    .B(_12678_),
    .Y(_12679_));
 sg13g2_a21oi_1 _19702_ (.A1(_09971_),
    .A2(net47),
    .Y(_00441_),
    .B1(_12679_));
 sg13g2_nor2_1 _19703_ (.A(net484),
    .B(_12352_),
    .Y(_12680_));
 sg13g2_buf_2 _19704_ (.A(_12680_),
    .X(_12681_));
 sg13g2_buf_1 _19705_ (.A(_12681_),
    .X(_12682_));
 sg13g2_nor2_1 _19706_ (.A(net484),
    .B(_12170_),
    .Y(_12683_));
 sg13g2_buf_2 _19707_ (.A(_12683_),
    .X(_12684_));
 sg13g2_nor2b_1 _19708_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_12685_));
 sg13g2_a21oi_1 _19709_ (.A1(net1010),
    .A2(_12684_),
    .Y(_12686_),
    .B1(_12685_));
 sg13g2_nand2_1 _19710_ (.Y(_12687_),
    .A(net433),
    .B(net46));
 sg13g2_o21ai_1 _19711_ (.B1(_12687_),
    .Y(_00442_),
    .A1(net46),
    .A2(_12686_));
 sg13g2_nor2b_1 _19712_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[4][11] ),
    .Y(_12688_));
 sg13g2_a21oi_1 _19713_ (.A1(_12434_),
    .A2(_12684_),
    .Y(_12689_),
    .B1(_12688_));
 sg13g2_nand2_1 _19714_ (.Y(_12690_),
    .A(net429),
    .B(net46));
 sg13g2_o21ai_1 _19715_ (.B1(_12690_),
    .Y(_00443_),
    .A1(_12682_),
    .A2(_12689_));
 sg13g2_buf_1 _19716_ (.A(_12145_),
    .X(_12691_));
 sg13g2_nor2_2 _19717_ (.A(net484),
    .B(_12198_),
    .Y(_12692_));
 sg13g2_mux2_1 _19718_ (.A0(\cpu.dcache.r_data[4][12] ),
    .A1(net1104),
    .S(_12692_),
    .X(_12693_));
 sg13g2_nor2_1 _19719_ (.A(_12681_),
    .B(_12693_),
    .Y(_12694_));
 sg13g2_a21oi_1 _19720_ (.A1(net428),
    .A2(net46),
    .Y(_00444_),
    .B1(_12694_));
 sg13g2_buf_1 _19721_ (.A(net1105),
    .X(_12695_));
 sg13g2_mux2_1 _19722_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(_12695_),
    .S(_12692_),
    .X(_12696_));
 sg13g2_nor2_1 _19723_ (.A(_12681_),
    .B(_12696_),
    .Y(_12697_));
 sg13g2_a21oi_1 _19724_ (.A1(net427),
    .A2(net46),
    .Y(_00445_),
    .B1(_12697_));
 sg13g2_buf_1 _19725_ (.A(net1111),
    .X(_12698_));
 sg13g2_mux2_1 _19726_ (.A0(\cpu.dcache.r_data[4][14] ),
    .A1(_12698_),
    .S(_12692_),
    .X(_12699_));
 sg13g2_nor2_1 _19727_ (.A(_12681_),
    .B(_12699_),
    .Y(_12700_));
 sg13g2_a21oi_1 _19728_ (.A1(net384),
    .A2(net46),
    .Y(_00446_),
    .B1(_12700_));
 sg13g2_mux2_1 _19729_ (.A0(\cpu.dcache.r_data[4][15] ),
    .A1(_12447_),
    .S(_12692_),
    .X(_12701_));
 sg13g2_nor2_1 _19730_ (.A(_12681_),
    .B(_12701_),
    .Y(_12702_));
 sg13g2_a21oi_1 _19731_ (.A1(net383),
    .A2(net46),
    .Y(_00447_),
    .B1(_12702_));
 sg13g2_buf_1 _19732_ (.A(_09970_),
    .X(_12703_));
 sg13g2_nor2_1 _19733_ (.A(net484),
    .B(_12375_),
    .Y(_12704_));
 sg13g2_buf_1 _19734_ (.A(_12704_),
    .X(_12705_));
 sg13g2_buf_1 _19735_ (.A(_12705_),
    .X(_12706_));
 sg13g2_nor2_1 _19736_ (.A(net484),
    .B(_12230_),
    .Y(_12707_));
 sg13g2_buf_1 _19737_ (.A(_12707_),
    .X(_12708_));
 sg13g2_mux2_1 _19738_ (.A0(\cpu.dcache.r_data[4][16] ),
    .A1(net1104),
    .S(_12708_),
    .X(_12709_));
 sg13g2_nor2_1 _19739_ (.A(_12705_),
    .B(_12709_),
    .Y(_12710_));
 sg13g2_a21oi_1 _19740_ (.A1(net761),
    .A2(net45),
    .Y(_00448_),
    .B1(_12710_));
 sg13g2_mux2_1 _19741_ (.A0(\cpu.dcache.r_data[4][17] ),
    .A1(net1007),
    .S(_12708_),
    .X(_12711_));
 sg13g2_nor2_1 _19742_ (.A(_12705_),
    .B(_12711_),
    .Y(_12712_));
 sg13g2_a21oi_1 _19743_ (.A1(net766),
    .A2(net45),
    .Y(_00449_),
    .B1(_12712_));
 sg13g2_mux2_1 _19744_ (.A0(\cpu.dcache.r_data[4][18] ),
    .A1(net1006),
    .S(_12708_),
    .X(_12713_));
 sg13g2_nor2_1 _19745_ (.A(_12705_),
    .B(_12713_),
    .Y(_12714_));
 sg13g2_a21oi_1 _19746_ (.A1(net765),
    .A2(net45),
    .Y(_00450_),
    .B1(_12714_));
 sg13g2_buf_1 _19747_ (.A(_12184_),
    .X(_12715_));
 sg13g2_nor2b_1 _19748_ (.A(_12708_),
    .B_N(\cpu.dcache.r_data[4][19] ),
    .Y(_12716_));
 sg13g2_a21oi_1 _19749_ (.A1(net1005),
    .A2(_12708_),
    .Y(_12717_),
    .B1(_12716_));
 sg13g2_nand2_1 _19750_ (.Y(_12718_),
    .A(net1009),
    .B(net45));
 sg13g2_o21ai_1 _19751_ (.B1(_12718_),
    .Y(_00451_),
    .A1(net45),
    .A2(_12717_));
 sg13g2_mux2_1 _19752_ (.A0(\cpu.dcache.r_data[4][1] ),
    .A1(net1007),
    .S(_12677_),
    .X(_12719_));
 sg13g2_nor2_1 _19753_ (.A(_12674_),
    .B(_12719_),
    .Y(_12720_));
 sg13g2_a21oi_1 _19754_ (.A1(_12237_),
    .A2(net47),
    .Y(_00452_),
    .B1(_12720_));
 sg13g2_nor2_1 _19755_ (.A(_10031_),
    .B(_12254_),
    .Y(_12721_));
 sg13g2_buf_2 _19756_ (.A(_12721_),
    .X(_12722_));
 sg13g2_nor2b_1 _19757_ (.A(_12722_),
    .B_N(\cpu.dcache.r_data[4][20] ),
    .Y(_12723_));
 sg13g2_a21oi_1 _19758_ (.A1(net1014),
    .A2(_12722_),
    .Y(_12724_),
    .B1(_12723_));
 sg13g2_nand2_1 _19759_ (.Y(_12725_),
    .A(net1011),
    .B(_12706_));
 sg13g2_o21ai_1 _19760_ (.B1(_12725_),
    .Y(_00453_),
    .A1(net45),
    .A2(_12724_));
 sg13g2_mux2_1 _19761_ (.A0(\cpu.dcache.r_data[4][21] ),
    .A1(net1007),
    .S(_12722_),
    .X(_12726_));
 sg13g2_nor2_1 _19762_ (.A(_12705_),
    .B(_12726_),
    .Y(_12727_));
 sg13g2_a21oi_1 _19763_ (.A1(net764),
    .A2(net45),
    .Y(_00454_),
    .B1(_12727_));
 sg13g2_mux2_1 _19764_ (.A0(\cpu.dcache.r_data[4][22] ),
    .A1(net1006),
    .S(_12722_),
    .X(_12728_));
 sg13g2_nor2_1 _19765_ (.A(_12705_),
    .B(_12728_),
    .Y(_12729_));
 sg13g2_a21oi_1 _19766_ (.A1(net763),
    .A2(net45),
    .Y(_00455_),
    .B1(_12729_));
 sg13g2_buf_1 _19767_ (.A(_12183_),
    .X(_12730_));
 sg13g2_mux2_1 _19768_ (.A0(\cpu.dcache.r_data[4][23] ),
    .A1(net1103),
    .S(_12722_),
    .X(_12731_));
 sg13g2_nor2_1 _19769_ (.A(_12705_),
    .B(_12731_),
    .Y(_12732_));
 sg13g2_a21oi_1 _19770_ (.A1(net762),
    .A2(_12706_),
    .Y(_00456_),
    .B1(_12732_));
 sg13g2_nand2_1 _19771_ (.Y(_12733_),
    .A(net441),
    .B(_12274_));
 sg13g2_buf_1 _19772_ (.A(_12733_),
    .X(_12734_));
 sg13g2_mux2_1 _19773_ (.A0(_12146_),
    .A1(\cpu.dcache.r_data[4][24] ),
    .S(net346),
    .X(_12735_));
 sg13g2_nor2_1 _19774_ (.A(net484),
    .B(_12404_),
    .Y(_12736_));
 sg13g2_buf_2 _19775_ (.A(_12736_),
    .X(_12737_));
 sg13g2_mux2_1 _19776_ (.A0(_12735_),
    .A1(net431),
    .S(net72),
    .X(_00457_));
 sg13g2_mux2_1 _19777_ (.A0(net1109),
    .A1(\cpu.dcache.r_data[4][25] ),
    .S(net346),
    .X(_12738_));
 sg13g2_mux2_1 _19778_ (.A0(_12738_),
    .A1(net430),
    .S(net72),
    .X(_00458_));
 sg13g2_mux2_1 _19779_ (.A0(net1108),
    .A1(\cpu.dcache.r_data[4][26] ),
    .S(net346),
    .X(_12739_));
 sg13g2_mux2_1 _19780_ (.A0(_12739_),
    .A1(_12181_),
    .S(_12737_),
    .X(_00459_));
 sg13g2_mux2_1 _19781_ (.A0(_12221_),
    .A1(\cpu.dcache.r_data[4][27] ),
    .S(net346),
    .X(_12740_));
 sg13g2_mux2_1 _19782_ (.A0(_12740_),
    .A1(net429),
    .S(_12737_),
    .X(_00460_));
 sg13g2_nor2_2 _19783_ (.A(net484),
    .B(_12298_),
    .Y(_12741_));
 sg13g2_mux2_1 _19784_ (.A0(\cpu.dcache.r_data[4][28] ),
    .A1(net1104),
    .S(_12741_),
    .X(_12742_));
 sg13g2_nor2_1 _19785_ (.A(net72),
    .B(_12742_),
    .Y(_12743_));
 sg13g2_a21oi_1 _19786_ (.A1(net428),
    .A2(net72),
    .Y(_00461_),
    .B1(_12743_));
 sg13g2_mux2_1 _19787_ (.A0(\cpu.dcache.r_data[4][29] ),
    .A1(_12695_),
    .S(_12741_),
    .X(_12744_));
 sg13g2_nor2_1 _19788_ (.A(net72),
    .B(_12744_),
    .Y(_12745_));
 sg13g2_a21oi_1 _19789_ (.A1(net427),
    .A2(net72),
    .Y(_00462_),
    .B1(_12745_));
 sg13g2_mux2_1 _19790_ (.A0(\cpu.dcache.r_data[4][2] ),
    .A1(net1006),
    .S(_12677_),
    .X(_12746_));
 sg13g2_nor2_1 _19791_ (.A(_12674_),
    .B(_12746_),
    .Y(_12747_));
 sg13g2_a21oi_1 _19792_ (.A1(_12241_),
    .A2(net47),
    .Y(_00463_),
    .B1(_12747_));
 sg13g2_mux2_1 _19793_ (.A0(\cpu.dcache.r_data[4][30] ),
    .A1(net1006),
    .S(_12741_),
    .X(_12748_));
 sg13g2_nor2_1 _19794_ (.A(_12736_),
    .B(_12748_),
    .Y(_12749_));
 sg13g2_a21oi_1 _19795_ (.A1(net384),
    .A2(net72),
    .Y(_00464_),
    .B1(_12749_));
 sg13g2_mux2_1 _19796_ (.A0(\cpu.dcache.r_data[4][31] ),
    .A1(_12730_),
    .S(_12741_),
    .X(_12750_));
 sg13g2_nor2_1 _19797_ (.A(_12736_),
    .B(_12750_),
    .Y(_12751_));
 sg13g2_a21oi_1 _19798_ (.A1(net383),
    .A2(net72),
    .Y(_00465_),
    .B1(_12751_));
 sg13g2_nor2b_1 _19799_ (.A(_12677_),
    .B_N(\cpu.dcache.r_data[4][3] ),
    .Y(_12752_));
 sg13g2_a21oi_1 _19800_ (.A1(net1005),
    .A2(_12677_),
    .Y(_02672_),
    .B1(_12752_));
 sg13g2_nand2_1 _19801_ (.Y(_02673_),
    .A(_12652_),
    .B(net47));
 sg13g2_o21ai_1 _19802_ (.B1(_02673_),
    .Y(_00466_),
    .A1(_12675_),
    .A2(_02672_));
 sg13g2_buf_1 _19803_ (.A(net1106),
    .X(_02674_));
 sg13g2_nor2_1 _19804_ (.A(_10031_),
    .B(_12320_),
    .Y(_02675_));
 sg13g2_buf_2 _19805_ (.A(_02675_),
    .X(_02676_));
 sg13g2_nor2b_1 _19806_ (.A(_02676_),
    .B_N(\cpu.dcache.r_data[4][4] ),
    .Y(_02677_));
 sg13g2_a21oi_1 _19807_ (.A1(net1004),
    .A2(_02676_),
    .Y(_02678_),
    .B1(_02677_));
 sg13g2_nand2_1 _19808_ (.Y(_02679_),
    .A(net1011),
    .B(net47));
 sg13g2_o21ai_1 _19809_ (.B1(_02679_),
    .Y(_00467_),
    .A1(net47),
    .A2(_02678_));
 sg13g2_mux2_1 _19810_ (.A0(\cpu.dcache.r_data[4][5] ),
    .A1(net1007),
    .S(_02676_),
    .X(_02680_));
 sg13g2_nor2_1 _19811_ (.A(_12674_),
    .B(_02680_),
    .Y(_02681_));
 sg13g2_a21oi_1 _19812_ (.A1(net764),
    .A2(net47),
    .Y(_00468_),
    .B1(_02681_));
 sg13g2_mux2_1 _19813_ (.A0(\cpu.dcache.r_data[4][6] ),
    .A1(net1006),
    .S(_02676_),
    .X(_02682_));
 sg13g2_nor2_1 _19814_ (.A(_12674_),
    .B(_02682_),
    .Y(_02683_));
 sg13g2_a21oi_1 _19815_ (.A1(_12266_),
    .A2(_12675_),
    .Y(_00469_),
    .B1(_02683_));
 sg13g2_mux2_1 _19816_ (.A0(\cpu.dcache.r_data[4][7] ),
    .A1(net1103),
    .S(_02676_),
    .X(_02684_));
 sg13g2_nor2_1 _19817_ (.A(_12674_),
    .B(_02684_),
    .Y(_02685_));
 sg13g2_a21oi_1 _19818_ (.A1(net762),
    .A2(net47),
    .Y(_00470_),
    .B1(_02685_));
 sg13g2_nor2b_1 _19819_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[4][8] ),
    .Y(_02686_));
 sg13g2_a21oi_1 _19820_ (.A1(net1004),
    .A2(_12684_),
    .Y(_02687_),
    .B1(_02686_));
 sg13g2_nand2_1 _19821_ (.Y(_02688_),
    .A(net431),
    .B(_12681_));
 sg13g2_o21ai_1 _19822_ (.B1(_02688_),
    .Y(_00471_),
    .A1(_12682_),
    .A2(_02687_));
 sg13g2_nor2b_1 _19823_ (.A(_12684_),
    .B_N(\cpu.dcache.r_data[4][9] ),
    .Y(_02689_));
 sg13g2_a21oi_1 _19824_ (.A1(net1008),
    .A2(_12684_),
    .Y(_02690_),
    .B1(_02689_));
 sg13g2_nand2_1 _19825_ (.Y(_02691_),
    .A(net430),
    .B(_12681_));
 sg13g2_o21ai_1 _19826_ (.B1(_02691_),
    .Y(_00472_),
    .A1(net46),
    .A2(_02690_));
 sg13g2_buf_1 _19827_ (.A(_09547_),
    .X(_02692_));
 sg13g2_nor2_1 _19828_ (.A(net760),
    .B(_12342_),
    .Y(_02693_));
 sg13g2_buf_1 _19829_ (.A(_02693_),
    .X(_02694_));
 sg13g2_buf_1 _19830_ (.A(_02694_),
    .X(_02695_));
 sg13g2_nor2_1 _19831_ (.A(net760),
    .B(_12155_),
    .Y(_02696_));
 sg13g2_buf_2 _19832_ (.A(_02696_),
    .X(_02697_));
 sg13g2_mux2_1 _19833_ (.A0(\cpu.dcache.r_data[5][0] ),
    .A1(net1104),
    .S(_02697_),
    .X(_02698_));
 sg13g2_nor2_1 _19834_ (.A(_02694_),
    .B(_02698_),
    .Y(_02699_));
 sg13g2_a21oi_1 _19835_ (.A1(net761),
    .A2(net44),
    .Y(_00473_),
    .B1(_02699_));
 sg13g2_nor2_1 _19836_ (.A(net760),
    .B(_12352_),
    .Y(_02700_));
 sg13g2_buf_2 _19837_ (.A(_02700_),
    .X(_02701_));
 sg13g2_buf_1 _19838_ (.A(_02701_),
    .X(_02702_));
 sg13g2_nor2_1 _19839_ (.A(net760),
    .B(_12170_),
    .Y(_02703_));
 sg13g2_buf_2 _19840_ (.A(_02703_),
    .X(_02704_));
 sg13g2_nor2b_1 _19841_ (.A(_02704_),
    .B_N(\cpu.dcache.r_data[5][10] ),
    .Y(_02705_));
 sg13g2_a21oi_1 _19842_ (.A1(net1010),
    .A2(_02704_),
    .Y(_02706_),
    .B1(_02705_));
 sg13g2_nand2_1 _19843_ (.Y(_02707_),
    .A(_12180_),
    .B(net43));
 sg13g2_o21ai_1 _19844_ (.B1(_02707_),
    .Y(_00474_),
    .A1(net43),
    .A2(_02706_));
 sg13g2_nor2b_1 _19845_ (.A(_02704_),
    .B_N(\cpu.dcache.r_data[5][11] ),
    .Y(_02708_));
 sg13g2_a21oi_1 _19846_ (.A1(net1005),
    .A2(_02704_),
    .Y(_02709_),
    .B1(_02708_));
 sg13g2_nand2_1 _19847_ (.Y(_02710_),
    .A(net429),
    .B(net43));
 sg13g2_o21ai_1 _19848_ (.B1(_02710_),
    .Y(_00475_),
    .A1(net43),
    .A2(_02709_));
 sg13g2_nor2_2 _19849_ (.A(net760),
    .B(_12198_),
    .Y(_02711_));
 sg13g2_mux2_1 _19850_ (.A0(\cpu.dcache.r_data[5][12] ),
    .A1(net1104),
    .S(_02711_),
    .X(_02712_));
 sg13g2_nor2_1 _19851_ (.A(_02701_),
    .B(_02712_),
    .Y(_02713_));
 sg13g2_a21oi_1 _19852_ (.A1(_12295_),
    .A2(net43),
    .Y(_00476_),
    .B1(_02713_));
 sg13g2_mux2_1 _19853_ (.A0(\cpu.dcache.r_data[5][13] ),
    .A1(net1007),
    .S(_02711_),
    .X(_02714_));
 sg13g2_nor2_1 _19854_ (.A(_02701_),
    .B(_02714_),
    .Y(_02715_));
 sg13g2_a21oi_1 _19855_ (.A1(net427),
    .A2(net43),
    .Y(_00477_),
    .B1(_02715_));
 sg13g2_mux2_1 _19856_ (.A0(\cpu.dcache.r_data[5][14] ),
    .A1(_12698_),
    .S(_02711_),
    .X(_02716_));
 sg13g2_nor2_1 _19857_ (.A(_02701_),
    .B(_02716_),
    .Y(_02717_));
 sg13g2_a21oi_1 _19858_ (.A1(_12309_),
    .A2(net43),
    .Y(_00478_),
    .B1(_02717_));
 sg13g2_mux2_1 _19859_ (.A0(\cpu.dcache.r_data[5][15] ),
    .A1(_12730_),
    .S(_02711_),
    .X(_02718_));
 sg13g2_nor2_1 _19860_ (.A(_02701_),
    .B(_02718_),
    .Y(_02719_));
 sg13g2_a21oi_1 _19861_ (.A1(net383),
    .A2(net43),
    .Y(_00479_),
    .B1(_02719_));
 sg13g2_nor2_1 _19862_ (.A(net760),
    .B(_12375_),
    .Y(_02720_));
 sg13g2_buf_1 _19863_ (.A(_02720_),
    .X(_02721_));
 sg13g2_buf_1 _19864_ (.A(_02721_),
    .X(_02722_));
 sg13g2_nor2_1 _19865_ (.A(net924),
    .B(_12230_),
    .Y(_02723_));
 sg13g2_buf_2 _19866_ (.A(_02723_),
    .X(_02724_));
 sg13g2_mux2_1 _19867_ (.A0(\cpu.dcache.r_data[5][16] ),
    .A1(net1104),
    .S(_02724_),
    .X(_02725_));
 sg13g2_nor2_1 _19868_ (.A(_02721_),
    .B(_02725_),
    .Y(_02726_));
 sg13g2_a21oi_1 _19869_ (.A1(net761),
    .A2(net42),
    .Y(_00480_),
    .B1(_02726_));
 sg13g2_buf_1 _19870_ (.A(_12236_),
    .X(_02727_));
 sg13g2_mux2_1 _19871_ (.A0(\cpu.dcache.r_data[5][17] ),
    .A1(net1007),
    .S(_02724_),
    .X(_02728_));
 sg13g2_nor2_1 _19872_ (.A(_02721_),
    .B(_02728_),
    .Y(_02729_));
 sg13g2_a21oi_1 _19873_ (.A1(net759),
    .A2(net42),
    .Y(_00481_),
    .B1(_02729_));
 sg13g2_buf_1 _19874_ (.A(net896),
    .X(_02730_));
 sg13g2_mux2_1 _19875_ (.A0(\cpu.dcache.r_data[5][18] ),
    .A1(net1006),
    .S(_02724_),
    .X(_02731_));
 sg13g2_nor2_1 _19876_ (.A(_02721_),
    .B(_02731_),
    .Y(_02732_));
 sg13g2_a21oi_1 _19877_ (.A1(net758),
    .A2(net42),
    .Y(_00482_),
    .B1(_02732_));
 sg13g2_nor2b_1 _19878_ (.A(_02724_),
    .B_N(\cpu.dcache.r_data[5][19] ),
    .Y(_02733_));
 sg13g2_a21oi_1 _19879_ (.A1(net1005),
    .A2(_02724_),
    .Y(_02734_),
    .B1(_02733_));
 sg13g2_nand2_1 _19880_ (.Y(_02735_),
    .A(net1009),
    .B(net42));
 sg13g2_o21ai_1 _19881_ (.B1(_02735_),
    .Y(_00483_),
    .A1(net42),
    .A2(_02734_));
 sg13g2_mux2_1 _19882_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(net1007),
    .S(_02697_),
    .X(_02736_));
 sg13g2_nor2_1 _19883_ (.A(_02694_),
    .B(_02736_),
    .Y(_02737_));
 sg13g2_a21oi_1 _19884_ (.A1(net759),
    .A2(net44),
    .Y(_00484_),
    .B1(_02737_));
 sg13g2_nor2_1 _19885_ (.A(net924),
    .B(_12254_),
    .Y(_02738_));
 sg13g2_buf_2 _19886_ (.A(_02738_),
    .X(_02739_));
 sg13g2_nor2b_1 _19887_ (.A(_02739_),
    .B_N(\cpu.dcache.r_data[5][20] ),
    .Y(_02740_));
 sg13g2_a21oi_1 _19888_ (.A1(net1004),
    .A2(_02739_),
    .Y(_02741_),
    .B1(_02740_));
 sg13g2_nand2_1 _19889_ (.Y(_02742_),
    .A(net1011),
    .B(net42));
 sg13g2_o21ai_1 _19890_ (.B1(_02742_),
    .Y(_00485_),
    .A1(_02722_),
    .A2(_02741_));
 sg13g2_buf_1 _19891_ (.A(_12202_),
    .X(_02743_));
 sg13g2_mux2_1 _19892_ (.A0(\cpu.dcache.r_data[5][21] ),
    .A1(net1007),
    .S(_02739_),
    .X(_02744_));
 sg13g2_nor2_1 _19893_ (.A(_02721_),
    .B(_02744_),
    .Y(_02745_));
 sg13g2_a21oi_1 _19894_ (.A1(net892),
    .A2(net42),
    .Y(_00486_),
    .B1(_02745_));
 sg13g2_buf_1 _19895_ (.A(net894),
    .X(_02746_));
 sg13g2_mux2_1 _19896_ (.A0(\cpu.dcache.r_data[5][22] ),
    .A1(net1006),
    .S(_02739_),
    .X(_02747_));
 sg13g2_nor2_1 _19897_ (.A(_02721_),
    .B(_02747_),
    .Y(_02748_));
 sg13g2_a21oi_1 _19898_ (.A1(net757),
    .A2(net42),
    .Y(_00487_),
    .B1(_02748_));
 sg13g2_buf_1 _19899_ (.A(_12217_),
    .X(_02749_));
 sg13g2_mux2_1 _19900_ (.A0(\cpu.dcache.r_data[5][23] ),
    .A1(net1103),
    .S(_02739_),
    .X(_02750_));
 sg13g2_nor2_1 _19901_ (.A(_02721_),
    .B(_02750_),
    .Y(_02751_));
 sg13g2_a21oi_1 _19902_ (.A1(net891),
    .A2(_02722_),
    .Y(_00488_),
    .B1(_02751_));
 sg13g2_nor2_1 _19903_ (.A(_02692_),
    .B(_12404_),
    .Y(_02752_));
 sg13g2_buf_2 _19904_ (.A(_02752_),
    .X(_02753_));
 sg13g2_buf_1 _19905_ (.A(_02753_),
    .X(_02754_));
 sg13g2_nor2_1 _19906_ (.A(net760),
    .B(_12131_),
    .Y(_02755_));
 sg13g2_buf_1 _19907_ (.A(_02755_),
    .X(_02756_));
 sg13g2_nor2b_1 _19908_ (.A(_02756_),
    .B_N(\cpu.dcache.r_data[5][24] ),
    .Y(_02757_));
 sg13g2_a21oi_1 _19909_ (.A1(net1004),
    .A2(_02756_),
    .Y(_02758_),
    .B1(_02757_));
 sg13g2_nand2_1 _19910_ (.Y(_02759_),
    .A(net431),
    .B(net41));
 sg13g2_o21ai_1 _19911_ (.B1(_02759_),
    .Y(_00489_),
    .A1(net41),
    .A2(_02758_));
 sg13g2_nor2b_1 _19912_ (.A(net550),
    .B_N(\cpu.dcache.r_data[5][25] ),
    .Y(_02760_));
 sg13g2_a21oi_1 _19913_ (.A1(net1008),
    .A2(net550),
    .Y(_02761_),
    .B1(_02760_));
 sg13g2_nand2_1 _19914_ (.Y(_02762_),
    .A(net430),
    .B(net41));
 sg13g2_o21ai_1 _19915_ (.B1(_02762_),
    .Y(_00490_),
    .A1(_02754_),
    .A2(_02761_));
 sg13g2_nor2b_1 _19916_ (.A(net550),
    .B_N(\cpu.dcache.r_data[5][26] ),
    .Y(_02763_));
 sg13g2_a21oi_1 _19917_ (.A1(net1010),
    .A2(net550),
    .Y(_02764_),
    .B1(_02763_));
 sg13g2_nand2_1 _19918_ (.Y(_02765_),
    .A(_12180_),
    .B(_02753_));
 sg13g2_o21ai_1 _19919_ (.B1(_02765_),
    .Y(_00491_),
    .A1(net41),
    .A2(_02764_));
 sg13g2_nor2b_1 _19920_ (.A(net550),
    .B_N(\cpu.dcache.r_data[5][27] ),
    .Y(_02766_));
 sg13g2_a21oi_1 _19921_ (.A1(net1005),
    .A2(net550),
    .Y(_02767_),
    .B1(_02766_));
 sg13g2_nand2_1 _19922_ (.Y(_02768_),
    .A(_12189_),
    .B(_02753_));
 sg13g2_o21ai_1 _19923_ (.B1(_02768_),
    .Y(_00492_),
    .A1(_02754_),
    .A2(_02767_));
 sg13g2_nor2_2 _19924_ (.A(_02692_),
    .B(_12298_),
    .Y(_02769_));
 sg13g2_mux2_1 _19925_ (.A0(\cpu.dcache.r_data[5][28] ),
    .A1(_12691_),
    .S(_02769_),
    .X(_02770_));
 sg13g2_nor2_1 _19926_ (.A(_02753_),
    .B(_02770_),
    .Y(_02771_));
 sg13g2_a21oi_1 _19927_ (.A1(_12194_),
    .A2(net41),
    .Y(_00493_),
    .B1(_02771_));
 sg13g2_buf_1 _19928_ (.A(_12206_),
    .X(_02772_));
 sg13g2_mux2_1 _19929_ (.A0(\cpu.dcache.r_data[5][29] ),
    .A1(net1102),
    .S(_02769_),
    .X(_02773_));
 sg13g2_nor2_1 _19930_ (.A(_02753_),
    .B(_02773_),
    .Y(_02774_));
 sg13g2_a21oi_1 _19931_ (.A1(_12205_),
    .A2(net41),
    .Y(_00494_),
    .B1(_02774_));
 sg13g2_mux2_1 _19932_ (.A0(\cpu.dcache.r_data[5][2] ),
    .A1(net1006),
    .S(_02697_),
    .X(_02775_));
 sg13g2_nor2_1 _19933_ (.A(_02694_),
    .B(_02775_),
    .Y(_02776_));
 sg13g2_a21oi_1 _19934_ (.A1(net758),
    .A2(net44),
    .Y(_00495_),
    .B1(_02776_));
 sg13g2_buf_1 _19935_ (.A(_12166_),
    .X(_02777_));
 sg13g2_mux2_1 _19936_ (.A0(\cpu.dcache.r_data[5][30] ),
    .A1(net1101),
    .S(_02769_),
    .X(_02778_));
 sg13g2_nor2_1 _19937_ (.A(_02753_),
    .B(_02778_),
    .Y(_02779_));
 sg13g2_a21oi_1 _19938_ (.A1(_12213_),
    .A2(net41),
    .Y(_00496_),
    .B1(_02779_));
 sg13g2_mux2_1 _19939_ (.A0(\cpu.dcache.r_data[5][31] ),
    .A1(net1103),
    .S(_02769_),
    .X(_02780_));
 sg13g2_nor2_1 _19940_ (.A(_02753_),
    .B(_02780_),
    .Y(_02781_));
 sg13g2_a21oi_1 _19941_ (.A1(_12220_),
    .A2(net41),
    .Y(_00497_),
    .B1(_02781_));
 sg13g2_nor2b_1 _19942_ (.A(_02697_),
    .B_N(\cpu.dcache.r_data[5][3] ),
    .Y(_02782_));
 sg13g2_a21oi_1 _19943_ (.A1(net1005),
    .A2(_02697_),
    .Y(_02783_),
    .B1(_02782_));
 sg13g2_nand2_1 _19944_ (.Y(_02784_),
    .A(net1009),
    .B(net44));
 sg13g2_o21ai_1 _19945_ (.B1(_02784_),
    .Y(_00498_),
    .A1(net44),
    .A2(_02783_));
 sg13g2_nor2_1 _19946_ (.A(net924),
    .B(_12320_),
    .Y(_02785_));
 sg13g2_buf_2 _19947_ (.A(_02785_),
    .X(_02786_));
 sg13g2_nor2b_1 _19948_ (.A(_02786_),
    .B_N(\cpu.dcache.r_data[5][4] ),
    .Y(_02787_));
 sg13g2_a21oi_1 _19949_ (.A1(net1004),
    .A2(_02786_),
    .Y(_02788_),
    .B1(_02787_));
 sg13g2_nand2_1 _19950_ (.Y(_02789_),
    .A(net1011),
    .B(net44));
 sg13g2_o21ai_1 _19951_ (.B1(_02789_),
    .Y(_00499_),
    .A1(net44),
    .A2(_02788_));
 sg13g2_mux2_1 _19952_ (.A0(\cpu.dcache.r_data[5][5] ),
    .A1(net1102),
    .S(_02786_),
    .X(_02790_));
 sg13g2_nor2_1 _19953_ (.A(_02694_),
    .B(_02790_),
    .Y(_02791_));
 sg13g2_a21oi_1 _19954_ (.A1(net892),
    .A2(net44),
    .Y(_00500_),
    .B1(_02791_));
 sg13g2_mux2_1 _19955_ (.A0(\cpu.dcache.r_data[5][6] ),
    .A1(net1101),
    .S(_02786_),
    .X(_02792_));
 sg13g2_nor2_1 _19956_ (.A(_02694_),
    .B(_02792_),
    .Y(_02793_));
 sg13g2_a21oi_1 _19957_ (.A1(net757),
    .A2(_02695_),
    .Y(_00501_),
    .B1(_02793_));
 sg13g2_mux2_1 _19958_ (.A0(\cpu.dcache.r_data[5][7] ),
    .A1(net1103),
    .S(_02786_),
    .X(_02794_));
 sg13g2_nor2_1 _19959_ (.A(_02694_),
    .B(_02794_),
    .Y(_02795_));
 sg13g2_a21oi_1 _19960_ (.A1(net891),
    .A2(_02695_),
    .Y(_00502_),
    .B1(_02795_));
 sg13g2_nor2b_1 _19961_ (.A(_02704_),
    .B_N(\cpu.dcache.r_data[5][8] ),
    .Y(_02796_));
 sg13g2_a21oi_1 _19962_ (.A1(net1004),
    .A2(_02704_),
    .Y(_02797_),
    .B1(_02796_));
 sg13g2_nand2_1 _19963_ (.Y(_02798_),
    .A(_12281_),
    .B(_02701_));
 sg13g2_o21ai_1 _19964_ (.B1(_02798_),
    .Y(_00503_),
    .A1(_02702_),
    .A2(_02797_));
 sg13g2_nor2b_1 _19965_ (.A(_02704_),
    .B_N(\cpu.dcache.r_data[5][9] ),
    .Y(_02799_));
 sg13g2_a21oi_1 _19966_ (.A1(net1008),
    .A2(_02704_),
    .Y(_02800_),
    .B1(_02799_));
 sg13g2_nand2_1 _19967_ (.Y(_02801_),
    .A(_12290_),
    .B(_02701_));
 sg13g2_o21ai_1 _19968_ (.B1(_02801_),
    .Y(_00504_),
    .A1(_02702_),
    .A2(_02800_));
 sg13g2_buf_1 _19969_ (.A(_09556_),
    .X(_02802_));
 sg13g2_nor2_1 _19970_ (.A(net756),
    .B(_12342_),
    .Y(_02803_));
 sg13g2_buf_1 _19971_ (.A(_02803_),
    .X(_02804_));
 sg13g2_buf_1 _19972_ (.A(_02804_),
    .X(_02805_));
 sg13g2_nor2_1 _19973_ (.A(net756),
    .B(_12155_),
    .Y(_02806_));
 sg13g2_buf_1 _19974_ (.A(_02806_),
    .X(_02807_));
 sg13g2_mux2_1 _19975_ (.A0(\cpu.dcache.r_data[6][0] ),
    .A1(net1104),
    .S(_02807_),
    .X(_02808_));
 sg13g2_nor2_1 _19976_ (.A(_02804_),
    .B(_02808_),
    .Y(_02809_));
 sg13g2_a21oi_1 _19977_ (.A1(net761),
    .A2(net40),
    .Y(_00505_),
    .B1(_02809_));
 sg13g2_nor2_1 _19978_ (.A(net756),
    .B(_12352_),
    .Y(_02810_));
 sg13g2_buf_2 _19979_ (.A(_02810_),
    .X(_02811_));
 sg13g2_buf_1 _19980_ (.A(_02811_),
    .X(_02812_));
 sg13g2_nor2_1 _19981_ (.A(net756),
    .B(_12170_),
    .Y(_02813_));
 sg13g2_buf_2 _19982_ (.A(_02813_),
    .X(_02814_));
 sg13g2_nor2b_1 _19983_ (.A(_02814_),
    .B_N(\cpu.dcache.r_data[6][10] ),
    .Y(_02815_));
 sg13g2_a21oi_1 _19984_ (.A1(net1010),
    .A2(_02814_),
    .Y(_02816_),
    .B1(_02815_));
 sg13g2_nand2_1 _19985_ (.Y(_02817_),
    .A(_12180_),
    .B(net39));
 sg13g2_o21ai_1 _19986_ (.B1(_02817_),
    .Y(_00506_),
    .A1(_02812_),
    .A2(_02816_));
 sg13g2_nor2b_1 _19987_ (.A(_02814_),
    .B_N(\cpu.dcache.r_data[6][11] ),
    .Y(_02818_));
 sg13g2_a21oi_1 _19988_ (.A1(_12715_),
    .A2(_02814_),
    .Y(_02819_),
    .B1(_02818_));
 sg13g2_nand2_1 _19989_ (.Y(_02820_),
    .A(_12189_),
    .B(net39));
 sg13g2_o21ai_1 _19990_ (.B1(_02820_),
    .Y(_00507_),
    .A1(net39),
    .A2(_02819_));
 sg13g2_nor2_2 _19991_ (.A(net756),
    .B(_12198_),
    .Y(_02821_));
 sg13g2_mux2_1 _19992_ (.A0(\cpu.dcache.r_data[6][12] ),
    .A1(_12691_),
    .S(_02821_),
    .X(_02822_));
 sg13g2_nor2_1 _19993_ (.A(_02811_),
    .B(_02822_),
    .Y(_02823_));
 sg13g2_a21oi_1 _19994_ (.A1(_12194_),
    .A2(net39),
    .Y(_00508_),
    .B1(_02823_));
 sg13g2_mux2_1 _19995_ (.A0(\cpu.dcache.r_data[6][13] ),
    .A1(net1102),
    .S(_02821_),
    .X(_02824_));
 sg13g2_nor2_1 _19996_ (.A(_02811_),
    .B(_02824_),
    .Y(_02825_));
 sg13g2_a21oi_1 _19997_ (.A1(_12205_),
    .A2(net39),
    .Y(_00509_),
    .B1(_02825_));
 sg13g2_mux2_1 _19998_ (.A0(\cpu.dcache.r_data[6][14] ),
    .A1(net1101),
    .S(_02821_),
    .X(_02826_));
 sg13g2_nor2_1 _19999_ (.A(_02811_),
    .B(_02826_),
    .Y(_02827_));
 sg13g2_a21oi_1 _20000_ (.A1(_12213_),
    .A2(net39),
    .Y(_00510_),
    .B1(_02827_));
 sg13g2_mux2_1 _20001_ (.A0(\cpu.dcache.r_data[6][15] ),
    .A1(net1103),
    .S(_02821_),
    .X(_02828_));
 sg13g2_nor2_1 _20002_ (.A(_02811_),
    .B(_02828_),
    .Y(_02829_));
 sg13g2_a21oi_1 _20003_ (.A1(_12220_),
    .A2(net39),
    .Y(_00511_),
    .B1(_02829_));
 sg13g2_nor2_1 _20004_ (.A(net756),
    .B(_12375_),
    .Y(_02830_));
 sg13g2_buf_1 _20005_ (.A(_02830_),
    .X(_02831_));
 sg13g2_buf_1 _20006_ (.A(_02831_),
    .X(_02832_));
 sg13g2_nor2_1 _20007_ (.A(_09556_),
    .B(_12230_),
    .Y(_02833_));
 sg13g2_buf_2 _20008_ (.A(_02833_),
    .X(_02834_));
 sg13g2_mux2_1 _20009_ (.A0(\cpu.dcache.r_data[6][16] ),
    .A1(net1104),
    .S(_02834_),
    .X(_02835_));
 sg13g2_nor2_1 _20010_ (.A(_02831_),
    .B(_02835_),
    .Y(_02836_));
 sg13g2_a21oi_1 _20011_ (.A1(net761),
    .A2(net38),
    .Y(_00512_),
    .B1(_02836_));
 sg13g2_mux2_1 _20012_ (.A0(\cpu.dcache.r_data[6][17] ),
    .A1(net1102),
    .S(_02834_),
    .X(_02837_));
 sg13g2_nor2_1 _20013_ (.A(_02831_),
    .B(_02837_),
    .Y(_02838_));
 sg13g2_a21oi_1 _20014_ (.A1(net759),
    .A2(net38),
    .Y(_00513_),
    .B1(_02838_));
 sg13g2_mux2_1 _20015_ (.A0(\cpu.dcache.r_data[6][18] ),
    .A1(net1101),
    .S(_02834_),
    .X(_02839_));
 sg13g2_nor2_1 _20016_ (.A(_02831_),
    .B(_02839_),
    .Y(_02840_));
 sg13g2_a21oi_1 _20017_ (.A1(net758),
    .A2(net38),
    .Y(_00514_),
    .B1(_02840_));
 sg13g2_nor2b_1 _20018_ (.A(_02834_),
    .B_N(\cpu.dcache.r_data[6][19] ),
    .Y(_02841_));
 sg13g2_a21oi_1 _20019_ (.A1(net1005),
    .A2(_02834_),
    .Y(_02842_),
    .B1(_02841_));
 sg13g2_nand2_1 _20020_ (.Y(_02843_),
    .A(net1009),
    .B(net38));
 sg13g2_o21ai_1 _20021_ (.B1(_02843_),
    .Y(_00515_),
    .A1(net38),
    .A2(_02842_));
 sg13g2_mux2_1 _20022_ (.A0(\cpu.dcache.r_data[6][1] ),
    .A1(net1102),
    .S(_02807_),
    .X(_02844_));
 sg13g2_nor2_1 _20023_ (.A(_02804_),
    .B(_02844_),
    .Y(_02845_));
 sg13g2_a21oi_1 _20024_ (.A1(net759),
    .A2(net40),
    .Y(_00516_),
    .B1(_02845_));
 sg13g2_nor2_1 _20025_ (.A(_09556_),
    .B(_12254_),
    .Y(_02846_));
 sg13g2_buf_1 _20026_ (.A(_02846_),
    .X(_02847_));
 sg13g2_nor2b_1 _20027_ (.A(_02847_),
    .B_N(\cpu.dcache.r_data[6][20] ),
    .Y(_02848_));
 sg13g2_a21oi_1 _20028_ (.A1(net1004),
    .A2(_02847_),
    .Y(_02849_),
    .B1(_02848_));
 sg13g2_nand2_1 _20029_ (.Y(_02850_),
    .A(net1011),
    .B(_02832_));
 sg13g2_o21ai_1 _20030_ (.B1(_02850_),
    .Y(_00517_),
    .A1(_02832_),
    .A2(_02849_));
 sg13g2_mux2_1 _20031_ (.A0(\cpu.dcache.r_data[6][21] ),
    .A1(net1102),
    .S(_02847_),
    .X(_02851_));
 sg13g2_nor2_1 _20032_ (.A(_02831_),
    .B(_02851_),
    .Y(_02852_));
 sg13g2_a21oi_1 _20033_ (.A1(net892),
    .A2(net38),
    .Y(_00518_),
    .B1(_02852_));
 sg13g2_mux2_1 _20034_ (.A0(\cpu.dcache.r_data[6][22] ),
    .A1(net1101),
    .S(_02847_),
    .X(_02853_));
 sg13g2_nor2_1 _20035_ (.A(_02831_),
    .B(_02853_),
    .Y(_02854_));
 sg13g2_a21oi_1 _20036_ (.A1(net757),
    .A2(net38),
    .Y(_00519_),
    .B1(_02854_));
 sg13g2_mux2_1 _20037_ (.A0(\cpu.dcache.r_data[6][23] ),
    .A1(net1103),
    .S(_02847_),
    .X(_02855_));
 sg13g2_nor2_1 _20038_ (.A(_02831_),
    .B(_02855_),
    .Y(_02856_));
 sg13g2_a21oi_1 _20039_ (.A1(net891),
    .A2(net38),
    .Y(_00520_),
    .B1(_02856_));
 sg13g2_nor2_1 _20040_ (.A(_02802_),
    .B(_12404_),
    .Y(_02857_));
 sg13g2_buf_2 _20041_ (.A(_02857_),
    .X(_02858_));
 sg13g2_buf_1 _20042_ (.A(_02858_),
    .X(_02859_));
 sg13g2_nor2_1 _20043_ (.A(net756),
    .B(_12131_),
    .Y(_02860_));
 sg13g2_buf_1 _20044_ (.A(_02860_),
    .X(_02861_));
 sg13g2_nor2b_1 _20045_ (.A(_02861_),
    .B_N(\cpu.dcache.r_data[6][24] ),
    .Y(_02862_));
 sg13g2_a21oi_1 _20046_ (.A1(_02674_),
    .A2(net549),
    .Y(_02863_),
    .B1(_02862_));
 sg13g2_nand2_1 _20047_ (.Y(_02864_),
    .A(_12281_),
    .B(net37));
 sg13g2_o21ai_1 _20048_ (.B1(_02864_),
    .Y(_00521_),
    .A1(net37),
    .A2(_02863_));
 sg13g2_nor2b_1 _20049_ (.A(net549),
    .B_N(\cpu.dcache.r_data[6][25] ),
    .Y(_02865_));
 sg13g2_a21oi_1 _20050_ (.A1(net1008),
    .A2(net549),
    .Y(_02866_),
    .B1(_02865_));
 sg13g2_nand2_1 _20051_ (.Y(_02867_),
    .A(_12290_),
    .B(net37));
 sg13g2_o21ai_1 _20052_ (.B1(_02867_),
    .Y(_00522_),
    .A1(_02859_),
    .A2(_02866_));
 sg13g2_nor2b_1 _20053_ (.A(net549),
    .B_N(\cpu.dcache.r_data[6][26] ),
    .Y(_02868_));
 sg13g2_a21oi_1 _20054_ (.A1(net1010),
    .A2(net549),
    .Y(_02869_),
    .B1(_02868_));
 sg13g2_nand2_1 _20055_ (.Y(_02870_),
    .A(_12180_),
    .B(_02858_));
 sg13g2_o21ai_1 _20056_ (.B1(_02870_),
    .Y(_00523_),
    .A1(net37),
    .A2(_02869_));
 sg13g2_nor2b_1 _20057_ (.A(net549),
    .B_N(\cpu.dcache.r_data[6][27] ),
    .Y(_02871_));
 sg13g2_a21oi_1 _20058_ (.A1(_12715_),
    .A2(net549),
    .Y(_02872_),
    .B1(_02871_));
 sg13g2_nand2_1 _20059_ (.Y(_02873_),
    .A(_12189_),
    .B(_02858_));
 sg13g2_o21ai_1 _20060_ (.B1(_02873_),
    .Y(_00524_),
    .A1(_02859_),
    .A2(_02872_));
 sg13g2_nor2_2 _20061_ (.A(_02802_),
    .B(_12298_),
    .Y(_02874_));
 sg13g2_mux2_1 _20062_ (.A0(\cpu.dcache.r_data[6][28] ),
    .A1(_12250_),
    .S(_02874_),
    .X(_02875_));
 sg13g2_nor2_1 _20063_ (.A(_02858_),
    .B(_02875_),
    .Y(_02876_));
 sg13g2_a21oi_1 _20064_ (.A1(_12194_),
    .A2(net37),
    .Y(_00525_),
    .B1(_02876_));
 sg13g2_mux2_1 _20065_ (.A0(\cpu.dcache.r_data[6][29] ),
    .A1(_02772_),
    .S(_02874_),
    .X(_02877_));
 sg13g2_nor2_1 _20066_ (.A(_02858_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_a21oi_1 _20067_ (.A1(_12205_),
    .A2(net37),
    .Y(_00526_),
    .B1(_02878_));
 sg13g2_mux2_1 _20068_ (.A0(\cpu.dcache.r_data[6][2] ),
    .A1(net1101),
    .S(_02807_),
    .X(_02879_));
 sg13g2_nor2_1 _20069_ (.A(_02804_),
    .B(_02879_),
    .Y(_02880_));
 sg13g2_a21oi_1 _20070_ (.A1(net758),
    .A2(net40),
    .Y(_00527_),
    .B1(_02880_));
 sg13g2_mux2_1 _20071_ (.A0(\cpu.dcache.r_data[6][30] ),
    .A1(_02777_),
    .S(_02874_),
    .X(_02881_));
 sg13g2_nor2_1 _20072_ (.A(_02858_),
    .B(_02881_),
    .Y(_02882_));
 sg13g2_a21oi_1 _20073_ (.A1(_12213_),
    .A2(net37),
    .Y(_00528_),
    .B1(_02882_));
 sg13g2_mux2_1 _20074_ (.A0(\cpu.dcache.r_data[6][31] ),
    .A1(net1103),
    .S(_02874_),
    .X(_02883_));
 sg13g2_nor2_1 _20075_ (.A(_02858_),
    .B(_02883_),
    .Y(_02884_));
 sg13g2_a21oi_1 _20076_ (.A1(_12220_),
    .A2(net37),
    .Y(_00529_),
    .B1(_02884_));
 sg13g2_nor2b_1 _20077_ (.A(_02807_),
    .B_N(\cpu.dcache.r_data[6][3] ),
    .Y(_02885_));
 sg13g2_a21oi_1 _20078_ (.A1(net1005),
    .A2(_02807_),
    .Y(_02886_),
    .B1(_02885_));
 sg13g2_nand2_1 _20079_ (.Y(_02887_),
    .A(net1009),
    .B(net40));
 sg13g2_o21ai_1 _20080_ (.B1(_02887_),
    .Y(_00530_),
    .A1(net40),
    .A2(_02886_));
 sg13g2_nor2_1 _20081_ (.A(_09556_),
    .B(_12320_),
    .Y(_02888_));
 sg13g2_buf_2 _20082_ (.A(_02888_),
    .X(_02889_));
 sg13g2_nor2b_1 _20083_ (.A(_02889_),
    .B_N(\cpu.dcache.r_data[6][4] ),
    .Y(_02890_));
 sg13g2_a21oi_1 _20084_ (.A1(net1004),
    .A2(_02889_),
    .Y(_02891_),
    .B1(_02890_));
 sg13g2_nand2_1 _20085_ (.Y(_02892_),
    .A(_12549_),
    .B(net40));
 sg13g2_o21ai_1 _20086_ (.B1(_02892_),
    .Y(_00531_),
    .A1(net40),
    .A2(_02891_));
 sg13g2_mux2_1 _20087_ (.A0(\cpu.dcache.r_data[6][5] ),
    .A1(net1102),
    .S(_02889_),
    .X(_02893_));
 sg13g2_nor2_1 _20088_ (.A(_02804_),
    .B(_02893_),
    .Y(_02894_));
 sg13g2_a21oi_1 _20089_ (.A1(net892),
    .A2(_02805_),
    .Y(_00532_),
    .B1(_02894_));
 sg13g2_mux2_1 _20090_ (.A0(\cpu.dcache.r_data[6][6] ),
    .A1(net1101),
    .S(_02889_),
    .X(_02895_));
 sg13g2_nor2_1 _20091_ (.A(_02804_),
    .B(_02895_),
    .Y(_02896_));
 sg13g2_a21oi_1 _20092_ (.A1(net757),
    .A2(_02805_),
    .Y(_00533_),
    .B1(_02896_));
 sg13g2_mux2_1 _20093_ (.A0(\cpu.dcache.r_data[6][7] ),
    .A1(net1110),
    .S(_02889_),
    .X(_02897_));
 sg13g2_nor2_1 _20094_ (.A(_02804_),
    .B(_02897_),
    .Y(_02898_));
 sg13g2_a21oi_1 _20095_ (.A1(net891),
    .A2(net40),
    .Y(_00534_),
    .B1(_02898_));
 sg13g2_nor2b_1 _20096_ (.A(_02814_),
    .B_N(\cpu.dcache.r_data[6][8] ),
    .Y(_02899_));
 sg13g2_a21oi_1 _20097_ (.A1(_02674_),
    .A2(_02814_),
    .Y(_02900_),
    .B1(_02899_));
 sg13g2_nand2_1 _20098_ (.Y(_02901_),
    .A(_12281_),
    .B(_02811_));
 sg13g2_o21ai_1 _20099_ (.B1(_02901_),
    .Y(_00535_),
    .A1(net39),
    .A2(_02900_));
 sg13g2_nor2b_1 _20100_ (.A(_02814_),
    .B_N(\cpu.dcache.r_data[6][9] ),
    .Y(_02902_));
 sg13g2_a21oi_1 _20101_ (.A1(net1008),
    .A2(_02814_),
    .Y(_02903_),
    .B1(_02902_));
 sg13g2_nand2_1 _20102_ (.Y(_02904_),
    .A(_12290_),
    .B(_02811_));
 sg13g2_o21ai_1 _20103_ (.B1(_02904_),
    .Y(_00536_),
    .A1(_02812_),
    .A2(_02903_));
 sg13g2_buf_1 _20104_ (.A(_09892_),
    .X(_02905_));
 sg13g2_nor2_1 _20105_ (.A(net381),
    .B(_12342_),
    .Y(_02906_));
 sg13g2_buf_1 _20106_ (.A(_02906_),
    .X(_02907_));
 sg13g2_buf_1 _20107_ (.A(_02907_),
    .X(_02908_));
 sg13g2_nor2_1 _20108_ (.A(net381),
    .B(_12155_),
    .Y(_02909_));
 sg13g2_buf_2 _20109_ (.A(_02909_),
    .X(_02910_));
 sg13g2_mux2_1 _20110_ (.A0(\cpu.dcache.r_data[7][0] ),
    .A1(net1106),
    .S(_02910_),
    .X(_02911_));
 sg13g2_nor2_1 _20111_ (.A(_02907_),
    .B(_02911_),
    .Y(_02912_));
 sg13g2_a21oi_1 _20112_ (.A1(net761),
    .A2(_02908_),
    .Y(_00537_),
    .B1(_02912_));
 sg13g2_nor2_1 _20113_ (.A(net381),
    .B(_12352_),
    .Y(_02913_));
 sg13g2_buf_2 _20114_ (.A(_02913_),
    .X(_02914_));
 sg13g2_buf_1 _20115_ (.A(_02914_),
    .X(_02915_));
 sg13g2_nor2_1 _20116_ (.A(_02905_),
    .B(_12170_),
    .Y(_02916_));
 sg13g2_buf_2 _20117_ (.A(_02916_),
    .X(_02917_));
 sg13g2_nor2b_1 _20118_ (.A(_02917_),
    .B_N(\cpu.dcache.r_data[7][10] ),
    .Y(_02918_));
 sg13g2_a21oi_1 _20119_ (.A1(net1010),
    .A2(_02917_),
    .Y(_02919_),
    .B1(_02918_));
 sg13g2_nand2_1 _20120_ (.Y(_02920_),
    .A(_12180_),
    .B(net35));
 sg13g2_o21ai_1 _20121_ (.B1(_02920_),
    .Y(_00538_),
    .A1(net35),
    .A2(_02919_));
 sg13g2_buf_2 _20122_ (.A(net1110),
    .X(_02921_));
 sg13g2_nor2b_1 _20123_ (.A(_02917_),
    .B_N(\cpu.dcache.r_data[7][11] ),
    .Y(_02922_));
 sg13g2_a21oi_1 _20124_ (.A1(net1003),
    .A2(_02917_),
    .Y(_02923_),
    .B1(_02922_));
 sg13g2_nand2_1 _20125_ (.Y(_02924_),
    .A(_12189_),
    .B(net35));
 sg13g2_o21ai_1 _20126_ (.B1(_02924_),
    .Y(_00539_),
    .A1(net35),
    .A2(_02923_));
 sg13g2_nor2_2 _20127_ (.A(net381),
    .B(_12198_),
    .Y(_02925_));
 sg13g2_mux2_1 _20128_ (.A0(\cpu.dcache.r_data[7][12] ),
    .A1(net1106),
    .S(_02925_),
    .X(_02926_));
 sg13g2_nor2_1 _20129_ (.A(_02914_),
    .B(_02926_),
    .Y(_02927_));
 sg13g2_a21oi_1 _20130_ (.A1(_12194_),
    .A2(net35),
    .Y(_00540_),
    .B1(_02927_));
 sg13g2_mux2_1 _20131_ (.A0(\cpu.dcache.r_data[7][13] ),
    .A1(_02772_),
    .S(_02925_),
    .X(_02928_));
 sg13g2_nor2_1 _20132_ (.A(_02914_),
    .B(_02928_),
    .Y(_02929_));
 sg13g2_a21oi_1 _20133_ (.A1(_12205_),
    .A2(net35),
    .Y(_00541_),
    .B1(_02929_));
 sg13g2_mux2_1 _20134_ (.A0(\cpu.dcache.r_data[7][14] ),
    .A1(_02777_),
    .S(_02925_),
    .X(_02930_));
 sg13g2_nor2_1 _20135_ (.A(_02914_),
    .B(_02930_),
    .Y(_02931_));
 sg13g2_a21oi_1 _20136_ (.A1(_12213_),
    .A2(net35),
    .Y(_00542_),
    .B1(_02931_));
 sg13g2_mux2_1 _20137_ (.A0(\cpu.dcache.r_data[7][15] ),
    .A1(net1110),
    .S(_02925_),
    .X(_02932_));
 sg13g2_nor2_1 _20138_ (.A(_02914_),
    .B(_02932_),
    .Y(_02933_));
 sg13g2_a21oi_1 _20139_ (.A1(_12220_),
    .A2(net35),
    .Y(_00543_),
    .B1(_02933_));
 sg13g2_nor2_1 _20140_ (.A(net381),
    .B(_12375_),
    .Y(_02934_));
 sg13g2_buf_1 _20141_ (.A(_02934_),
    .X(_02935_));
 sg13g2_buf_1 _20142_ (.A(_02935_),
    .X(_02936_));
 sg13g2_nor2_1 _20143_ (.A(net381),
    .B(_12230_),
    .Y(_02937_));
 sg13g2_buf_2 _20144_ (.A(_02937_),
    .X(_02938_));
 sg13g2_mux2_1 _20145_ (.A0(\cpu.dcache.r_data[7][16] ),
    .A1(net1106),
    .S(_02938_),
    .X(_02939_));
 sg13g2_nor2_1 _20146_ (.A(_02935_),
    .B(_02939_),
    .Y(_02940_));
 sg13g2_a21oi_1 _20147_ (.A1(net761),
    .A2(net34),
    .Y(_00544_),
    .B1(_02940_));
 sg13g2_mux2_1 _20148_ (.A0(\cpu.dcache.r_data[7][17] ),
    .A1(net1102),
    .S(_02938_),
    .X(_02941_));
 sg13g2_nor2_1 _20149_ (.A(_02935_),
    .B(_02941_),
    .Y(_02942_));
 sg13g2_a21oi_1 _20150_ (.A1(net759),
    .A2(net34),
    .Y(_00545_),
    .B1(_02942_));
 sg13g2_mux2_1 _20151_ (.A0(\cpu.dcache.r_data[7][18] ),
    .A1(net1101),
    .S(_02938_),
    .X(_02943_));
 sg13g2_nor2_1 _20152_ (.A(_02935_),
    .B(_02943_),
    .Y(_02944_));
 sg13g2_a21oi_1 _20153_ (.A1(net758),
    .A2(net34),
    .Y(_00546_),
    .B1(_02944_));
 sg13g2_nor2b_1 _20154_ (.A(_02938_),
    .B_N(\cpu.dcache.r_data[7][19] ),
    .Y(_02945_));
 sg13g2_a21oi_1 _20155_ (.A1(net1003),
    .A2(_02938_),
    .Y(_02946_),
    .B1(_02945_));
 sg13g2_nand2_1 _20156_ (.Y(_02947_),
    .A(net1009),
    .B(net34));
 sg13g2_o21ai_1 _20157_ (.B1(_02947_),
    .Y(_00547_),
    .A1(net34),
    .A2(_02946_));
 sg13g2_mux2_1 _20158_ (.A0(\cpu.dcache.r_data[7][1] ),
    .A1(net1105),
    .S(_02910_),
    .X(_02948_));
 sg13g2_nor2_1 _20159_ (.A(_02907_),
    .B(_02948_),
    .Y(_02949_));
 sg13g2_a21oi_1 _20160_ (.A1(net759),
    .A2(net36),
    .Y(_00548_),
    .B1(_02949_));
 sg13g2_buf_2 _20161_ (.A(net1106),
    .X(_02950_));
 sg13g2_nor2_1 _20162_ (.A(_09892_),
    .B(_12254_),
    .Y(_02951_));
 sg13g2_buf_2 _20163_ (.A(_02951_),
    .X(_02952_));
 sg13g2_nor2b_1 _20164_ (.A(_02952_),
    .B_N(\cpu.dcache.r_data[7][20] ),
    .Y(_02953_));
 sg13g2_a21oi_1 _20165_ (.A1(net1002),
    .A2(_02952_),
    .Y(_02954_),
    .B1(_02953_));
 sg13g2_nand2_1 _20166_ (.Y(_02955_),
    .A(_12549_),
    .B(net34));
 sg13g2_o21ai_1 _20167_ (.B1(_02955_),
    .Y(_00549_),
    .A1(net34),
    .A2(_02954_));
 sg13g2_mux2_1 _20168_ (.A0(\cpu.dcache.r_data[7][21] ),
    .A1(net1105),
    .S(_02952_),
    .X(_02956_));
 sg13g2_nor2_1 _20169_ (.A(_02935_),
    .B(_02956_),
    .Y(_02957_));
 sg13g2_a21oi_1 _20170_ (.A1(net892),
    .A2(_02936_),
    .Y(_00550_),
    .B1(_02957_));
 sg13g2_mux2_1 _20171_ (.A0(\cpu.dcache.r_data[7][22] ),
    .A1(net1111),
    .S(_02952_),
    .X(_02958_));
 sg13g2_nor2_1 _20172_ (.A(_02935_),
    .B(_02958_),
    .Y(_02959_));
 sg13g2_a21oi_1 _20173_ (.A1(net757),
    .A2(_02936_),
    .Y(_00551_),
    .B1(_02959_));
 sg13g2_mux2_1 _20174_ (.A0(\cpu.dcache.r_data[7][23] ),
    .A1(net1110),
    .S(_02952_),
    .X(_02960_));
 sg13g2_nor2_1 _20175_ (.A(_02935_),
    .B(_02960_),
    .Y(_02961_));
 sg13g2_a21oi_1 _20176_ (.A1(net891),
    .A2(net34),
    .Y(_00552_),
    .B1(_02961_));
 sg13g2_nor2_1 _20177_ (.A(_02905_),
    .B(_12404_),
    .Y(_02962_));
 sg13g2_buf_2 _20178_ (.A(_02962_),
    .X(_02963_));
 sg13g2_buf_1 _20179_ (.A(_02963_),
    .X(_02964_));
 sg13g2_nor2_1 _20180_ (.A(_09892_),
    .B(_12131_),
    .Y(_02965_));
 sg13g2_buf_1 _20181_ (.A(_02965_),
    .X(_02966_));
 sg13g2_nor2b_1 _20182_ (.A(net345),
    .B_N(\cpu.dcache.r_data[7][24] ),
    .Y(_02967_));
 sg13g2_a21oi_1 _20183_ (.A1(net1002),
    .A2(net345),
    .Y(_02968_),
    .B1(_02967_));
 sg13g2_nand2_1 _20184_ (.Y(_02969_),
    .A(_12281_),
    .B(net33));
 sg13g2_o21ai_1 _20185_ (.B1(_02969_),
    .Y(_00553_),
    .A1(net33),
    .A2(_02968_));
 sg13g2_nor2b_1 _20186_ (.A(net345),
    .B_N(\cpu.dcache.r_data[7][25] ),
    .Y(_02970_));
 sg13g2_a21oi_1 _20187_ (.A1(net1008),
    .A2(net345),
    .Y(_02971_),
    .B1(_02970_));
 sg13g2_nand2_1 _20188_ (.Y(_02972_),
    .A(_12290_),
    .B(net33));
 sg13g2_o21ai_1 _20189_ (.B1(_02972_),
    .Y(_00554_),
    .A1(net33),
    .A2(_02971_));
 sg13g2_nor2b_1 _20190_ (.A(net345),
    .B_N(\cpu.dcache.r_data[7][26] ),
    .Y(_02973_));
 sg13g2_a21oi_1 _20191_ (.A1(net1010),
    .A2(net345),
    .Y(_02974_),
    .B1(_02973_));
 sg13g2_nand2_1 _20192_ (.Y(_02975_),
    .A(_12180_),
    .B(_02963_));
 sg13g2_o21ai_1 _20193_ (.B1(_02975_),
    .Y(_00555_),
    .A1(_02964_),
    .A2(_02974_));
 sg13g2_nor2b_1 _20194_ (.A(net345),
    .B_N(\cpu.dcache.r_data[7][27] ),
    .Y(_02976_));
 sg13g2_a21oi_1 _20195_ (.A1(net1003),
    .A2(net345),
    .Y(_02977_),
    .B1(_02976_));
 sg13g2_nand2_1 _20196_ (.Y(_02978_),
    .A(_12189_),
    .B(_02963_));
 sg13g2_o21ai_1 _20197_ (.B1(_02978_),
    .Y(_00556_),
    .A1(_02964_),
    .A2(_02977_));
 sg13g2_nor2_2 _20198_ (.A(net381),
    .B(_12298_),
    .Y(_02979_));
 sg13g2_mux2_1 _20199_ (.A0(\cpu.dcache.r_data[7][28] ),
    .A1(net1106),
    .S(_02979_),
    .X(_02980_));
 sg13g2_nor2_1 _20200_ (.A(_02963_),
    .B(_02980_),
    .Y(_02981_));
 sg13g2_a21oi_1 _20201_ (.A1(_12194_),
    .A2(net33),
    .Y(_00557_),
    .B1(_02981_));
 sg13g2_mux2_1 _20202_ (.A0(\cpu.dcache.r_data[7][29] ),
    .A1(net1105),
    .S(_02979_),
    .X(_02982_));
 sg13g2_nor2_1 _20203_ (.A(_02963_),
    .B(_02982_),
    .Y(_02983_));
 sg13g2_a21oi_1 _20204_ (.A1(_12205_),
    .A2(net33),
    .Y(_00558_),
    .B1(_02983_));
 sg13g2_mux2_1 _20205_ (.A0(\cpu.dcache.r_data[7][2] ),
    .A1(net1111),
    .S(_02910_),
    .X(_02984_));
 sg13g2_nor2_1 _20206_ (.A(_02907_),
    .B(_02984_),
    .Y(_02985_));
 sg13g2_a21oi_1 _20207_ (.A1(net758),
    .A2(net36),
    .Y(_00559_),
    .B1(_02985_));
 sg13g2_mux2_1 _20208_ (.A0(\cpu.dcache.r_data[7][30] ),
    .A1(net1111),
    .S(_02979_),
    .X(_02986_));
 sg13g2_nor2_1 _20209_ (.A(_02963_),
    .B(_02986_),
    .Y(_02987_));
 sg13g2_a21oi_1 _20210_ (.A1(_12213_),
    .A2(net33),
    .Y(_00560_),
    .B1(_02987_));
 sg13g2_mux2_1 _20211_ (.A0(\cpu.dcache.r_data[7][31] ),
    .A1(net1110),
    .S(_02979_),
    .X(_02988_));
 sg13g2_nor2_1 _20212_ (.A(_02963_),
    .B(_02988_),
    .Y(_02989_));
 sg13g2_a21oi_1 _20213_ (.A1(_12220_),
    .A2(net33),
    .Y(_00561_),
    .B1(_02989_));
 sg13g2_nor2b_1 _20214_ (.A(_02910_),
    .B_N(\cpu.dcache.r_data[7][3] ),
    .Y(_02990_));
 sg13g2_a21oi_1 _20215_ (.A1(net1003),
    .A2(_02910_),
    .Y(_02991_),
    .B1(_02990_));
 sg13g2_nand2_1 _20216_ (.Y(_02992_),
    .A(_12652_),
    .B(net36));
 sg13g2_o21ai_1 _20217_ (.B1(_02992_),
    .Y(_00562_),
    .A1(net36),
    .A2(_02991_));
 sg13g2_nor2_1 _20218_ (.A(_09892_),
    .B(_12320_),
    .Y(_02993_));
 sg13g2_buf_2 _20219_ (.A(_02993_),
    .X(_02994_));
 sg13g2_nor2b_1 _20220_ (.A(_02994_),
    .B_N(\cpu.dcache.r_data[7][4] ),
    .Y(_02995_));
 sg13g2_a21oi_1 _20221_ (.A1(net1002),
    .A2(_02994_),
    .Y(_02996_),
    .B1(_02995_));
 sg13g2_nand2_1 _20222_ (.Y(_02997_),
    .A(net1057),
    .B(_02908_));
 sg13g2_o21ai_1 _20223_ (.B1(_02997_),
    .Y(_00563_),
    .A1(net36),
    .A2(_02996_));
 sg13g2_mux2_1 _20224_ (.A0(\cpu.dcache.r_data[7][5] ),
    .A1(net1105),
    .S(_02994_),
    .X(_02998_));
 sg13g2_nor2_1 _20225_ (.A(_02907_),
    .B(_02998_),
    .Y(_02999_));
 sg13g2_a21oi_1 _20226_ (.A1(net892),
    .A2(net36),
    .Y(_00564_),
    .B1(_02999_));
 sg13g2_mux2_1 _20227_ (.A0(\cpu.dcache.r_data[7][6] ),
    .A1(net1111),
    .S(_02994_),
    .X(_03000_));
 sg13g2_nor2_1 _20228_ (.A(_02907_),
    .B(_03000_),
    .Y(_03001_));
 sg13g2_a21oi_1 _20229_ (.A1(net757),
    .A2(net36),
    .Y(_00565_),
    .B1(_03001_));
 sg13g2_mux2_1 _20230_ (.A0(\cpu.dcache.r_data[7][7] ),
    .A1(net1110),
    .S(_02994_),
    .X(_03002_));
 sg13g2_nor2_1 _20231_ (.A(_02907_),
    .B(_03002_),
    .Y(_03003_));
 sg13g2_a21oi_1 _20232_ (.A1(net891),
    .A2(net36),
    .Y(_00566_),
    .B1(_03003_));
 sg13g2_nor2b_1 _20233_ (.A(_02917_),
    .B_N(\cpu.dcache.r_data[7][8] ),
    .Y(_03004_));
 sg13g2_a21oi_1 _20234_ (.A1(net1002),
    .A2(_02917_),
    .Y(_03005_),
    .B1(_03004_));
 sg13g2_nand2_1 _20235_ (.Y(_03006_),
    .A(_12281_),
    .B(_02914_));
 sg13g2_o21ai_1 _20236_ (.B1(_03006_),
    .Y(_00567_),
    .A1(_02915_),
    .A2(_03005_));
 sg13g2_nor2b_1 _20237_ (.A(_02917_),
    .B_N(\cpu.dcache.r_data[7][9] ),
    .Y(_03007_));
 sg13g2_a21oi_1 _20238_ (.A1(net1008),
    .A2(_02917_),
    .Y(_03008_),
    .B1(_03007_));
 sg13g2_nand2_1 _20239_ (.Y(_03009_),
    .A(_12290_),
    .B(_02914_));
 sg13g2_o21ai_1 _20240_ (.B1(_03009_),
    .Y(_00568_),
    .A1(_02915_),
    .A2(_03008_));
 sg13g2_and2_1 _20241_ (.A(_11634_),
    .B(_12124_),
    .X(_03010_));
 sg13g2_buf_1 _20242_ (.A(net1166),
    .X(_03011_));
 sg13g2_buf_1 _20243_ (.A(\cpu.d_rstrobe_d ),
    .X(_03012_));
 sg13g2_nand2b_1 _20244_ (.Y(_03013_),
    .B(_12148_),
    .A_N(_03012_));
 sg13g2_nor4_1 _20245_ (.A(net1001),
    .B(_09303_),
    .C(_08355_),
    .D(_03013_),
    .Y(_03014_));
 sg13g2_or2_1 _20246_ (.X(_03015_),
    .B(_03014_),
    .A(_03010_));
 sg13g2_buf_2 _20247_ (.A(_03015_),
    .X(_03016_));
 sg13g2_nand2b_1 _20248_ (.Y(_03017_),
    .B(_03012_),
    .A_N(net1029));
 sg13g2_nand2_1 _20249_ (.Y(_03018_),
    .A(_12296_),
    .B(_12129_));
 sg13g2_a21oi_1 _20250_ (.A1(_03013_),
    .A2(_03017_),
    .Y(_03019_),
    .B1(_03018_));
 sg13g2_or2_1 _20251_ (.X(_03020_),
    .B(_03010_),
    .A(_03019_));
 sg13g2_buf_2 _20252_ (.A(_03020_),
    .X(_03021_));
 sg13g2_nor2b_1 _20253_ (.A(_12147_),
    .B_N(_03021_),
    .Y(_03022_));
 sg13g2_mux2_1 _20254_ (.A0(\cpu.dcache.r_dirty[0] ),
    .A1(_03016_),
    .S(_03022_),
    .X(_00569_));
 sg13g2_buf_1 _20255_ (.A(net643),
    .X(_03023_));
 sg13g2_buf_1 _20256_ (.A(net548),
    .X(_03024_));
 sg13g2_buf_1 _20257_ (.A(net483),
    .X(_03025_));
 sg13g2_nand2_1 _20258_ (.Y(_03026_),
    .A(_03025_),
    .B(_03021_));
 sg13g2_mux2_1 _20259_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[1] ),
    .S(_03026_),
    .X(_00570_));
 sg13g2_buf_1 _20260_ (.A(net641),
    .X(_03027_));
 sg13g2_buf_1 _20261_ (.A(net547),
    .X(_03028_));
 sg13g2_buf_1 _20262_ (.A(net482),
    .X(_03029_));
 sg13g2_nand2_1 _20263_ (.Y(_03030_),
    .A(_03029_),
    .B(_03021_));
 sg13g2_mux2_1 _20264_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[2] ),
    .S(_03030_),
    .X(_00571_));
 sg13g2_buf_1 _20265_ (.A(_09360_),
    .X(_03031_));
 sg13g2_buf_1 _20266_ (.A(net546),
    .X(_03032_));
 sg13g2_buf_1 _20267_ (.A(net481),
    .X(_03033_));
 sg13g2_nand2_1 _20268_ (.Y(_03034_),
    .A(_03033_),
    .B(_03021_));
 sg13g2_mux2_1 _20269_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[3] ),
    .S(_03034_),
    .X(_00572_));
 sg13g2_nand2_1 _20270_ (.Y(_03035_),
    .A(_10019_),
    .B(_03021_));
 sg13g2_mux2_1 _20271_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[4] ),
    .S(_03035_),
    .X(_00573_));
 sg13g2_buf_1 _20272_ (.A(net639),
    .X(_03036_));
 sg13g2_buf_1 _20273_ (.A(net545),
    .X(_03037_));
 sg13g2_buf_1 _20274_ (.A(net480),
    .X(_03038_));
 sg13g2_nand2_1 _20275_ (.Y(_03039_),
    .A(_03038_),
    .B(_03021_));
 sg13g2_mux2_1 _20276_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[5] ),
    .S(_03039_),
    .X(_00574_));
 sg13g2_buf_1 _20277_ (.A(net644),
    .X(_03040_));
 sg13g2_buf_1 _20278_ (.A(net544),
    .X(_03041_));
 sg13g2_buf_1 _20279_ (.A(net479),
    .X(_03042_));
 sg13g2_buf_1 _20280_ (.A(net421),
    .X(_03043_));
 sg13g2_nand2_1 _20281_ (.Y(_03044_),
    .A(_03043_),
    .B(_03021_));
 sg13g2_mux2_1 _20282_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[6] ),
    .S(_03044_),
    .X(_00575_));
 sg13g2_buf_1 _20283_ (.A(net703),
    .X(_03045_));
 sg13g2_buf_1 _20284_ (.A(net621),
    .X(_03046_));
 sg13g2_buf_1 _20285_ (.A(net543),
    .X(_03047_));
 sg13g2_buf_1 _20286_ (.A(net478),
    .X(_03048_));
 sg13g2_nand2_1 _20287_ (.Y(_03049_),
    .A(_03048_),
    .B(_03021_));
 sg13g2_mux2_1 _20288_ (.A0(_03016_),
    .A1(\cpu.dcache.r_dirty[7] ),
    .S(_03049_),
    .X(_00576_));
 sg13g2_buf_1 _20289_ (.A(_12074_),
    .X(_03050_));
 sg13g2_buf_1 _20290_ (.A(net755),
    .X(_03051_));
 sg13g2_buf_1 _20291_ (.A(net432),
    .X(_03052_));
 sg13g2_buf_1 _20292_ (.A(_12276_),
    .X(_03053_));
 sg13g2_nand2_1 _20293_ (.Y(_03054_),
    .A(\cpu.dcache.r_tag[0][5] ),
    .B(_03053_));
 sg13g2_o21ai_1 _20294_ (.B1(_03054_),
    .Y(_00580_),
    .A1(net674),
    .A2(net379));
 sg13g2_mux2_1 _20295_ (.A0(net442),
    .A1(\cpu.dcache.r_tag[0][15] ),
    .S(_03052_),
    .X(_00581_));
 sg13g2_mux2_1 _20296_ (.A0(net390),
    .A1(\cpu.dcache.r_tag[0][16] ),
    .S(net379),
    .X(_00582_));
 sg13g2_mux2_1 _20297_ (.A0(net391),
    .A1(\cpu.dcache.r_tag[0][17] ),
    .S(_03052_),
    .X(_00583_));
 sg13g2_mux2_1 _20298_ (.A0(net445),
    .A1(\cpu.dcache.r_tag[0][18] ),
    .S(net379),
    .X(_00584_));
 sg13g2_mux2_1 _20299_ (.A0(net389),
    .A1(\cpu.dcache.r_tag[0][19] ),
    .S(net379),
    .X(_00585_));
 sg13g2_mux2_1 _20300_ (.A0(net444),
    .A1(\cpu.dcache.r_tag[0][20] ),
    .S(_03053_),
    .X(_00586_));
 sg13g2_mux2_1 _20301_ (.A0(net387),
    .A1(\cpu.dcache.r_tag[0][21] ),
    .S(net419),
    .X(_00587_));
 sg13g2_mux2_1 _20302_ (.A0(net443),
    .A1(\cpu.dcache.r_tag[0][22] ),
    .S(net419),
    .X(_00588_));
 sg13g2_nand2_1 _20303_ (.Y(_03055_),
    .A(\cpu.dcache.r_tag[0][23] ),
    .B(net432));
 sg13g2_o21ai_1 _20304_ (.B1(_03055_),
    .Y(_00589_),
    .A1(_09789_),
    .A2(net379));
 sg13g2_buf_2 _20305_ (.A(_09164_),
    .X(_03056_));
 sg13g2_buf_1 _20306_ (.A(net1000),
    .X(_03057_));
 sg13g2_buf_1 _20307_ (.A(net890),
    .X(_03058_));
 sg13g2_mux2_1 _20308_ (.A0(net754),
    .A1(\cpu.dcache.r_tag[0][6] ),
    .S(net419),
    .X(_00590_));
 sg13g2_buf_1 _20309_ (.A(_09167_),
    .X(_03059_));
 sg13g2_buf_1 _20310_ (.A(_03059_),
    .X(_03060_));
 sg13g2_nand2_1 _20311_ (.Y(_03061_),
    .A(\cpu.dcache.r_tag[0][7] ),
    .B(net432));
 sg13g2_o21ai_1 _20312_ (.B1(_03061_),
    .Y(_00591_),
    .A1(net753),
    .A2(net379));
 sg13g2_buf_1 _20313_ (.A(_10920_),
    .X(_03062_));
 sg13g2_buf_1 _20314_ (.A(net888),
    .X(_03063_));
 sg13g2_nand2_1 _20315_ (.Y(_03064_),
    .A(\cpu.dcache.r_tag[0][8] ),
    .B(_12277_));
 sg13g2_o21ai_1 _20316_ (.B1(_03064_),
    .Y(_00592_),
    .A1(net752),
    .A2(net379));
 sg13g2_buf_1 _20317_ (.A(_10876_),
    .X(_03065_));
 sg13g2_buf_1 _20318_ (.A(net887),
    .X(_03066_));
 sg13g2_nand2_1 _20319_ (.Y(_03067_),
    .A(\cpu.dcache.r_tag[0][9] ),
    .B(_12277_));
 sg13g2_o21ai_1 _20320_ (.B1(_03067_),
    .Y(_00593_),
    .A1(net751),
    .A2(net379));
 sg13g2_buf_1 _20321_ (.A(net1143),
    .X(_03068_));
 sg13g2_buf_1 _20322_ (.A(net999),
    .X(_03069_));
 sg13g2_mux2_1 _20323_ (.A0(net886),
    .A1(\cpu.dcache.r_tag[0][10] ),
    .S(net419),
    .X(_00594_));
 sg13g2_buf_1 _20324_ (.A(net1135),
    .X(_03070_));
 sg13g2_buf_1 _20325_ (.A(net998),
    .X(_03071_));
 sg13g2_mux2_1 _20326_ (.A0(net885),
    .A1(\cpu.dcache.r_tag[0][11] ),
    .S(net419),
    .X(_00595_));
 sg13g2_mux2_1 _20327_ (.A0(net351),
    .A1(\cpu.dcache.r_tag[0][12] ),
    .S(net419),
    .X(_00596_));
 sg13g2_mux2_1 _20328_ (.A0(net388),
    .A1(\cpu.dcache.r_tag[0][13] ),
    .S(net419),
    .X(_00597_));
 sg13g2_mux2_1 _20329_ (.A0(net446),
    .A1(\cpu.dcache.r_tag[0][14] ),
    .S(net419),
    .X(_00598_));
 sg13g2_buf_2 _20330_ (.A(net678),
    .X(_03072_));
 sg13g2_buf_1 _20331_ (.A(net620),
    .X(_03073_));
 sg13g2_buf_1 _20332_ (.A(_12409_),
    .X(_03074_));
 sg13g2_mux2_1 _20333_ (.A0(\cpu.dcache.r_tag[1][5] ),
    .A1(net542),
    .S(net477),
    .X(_00599_));
 sg13g2_mux2_1 _20334_ (.A0(\cpu.dcache.r_tag[1][15] ),
    .A1(net442),
    .S(net477),
    .X(_00600_));
 sg13g2_mux2_1 _20335_ (.A0(\cpu.dcache.r_tag[1][16] ),
    .A1(net390),
    .S(net477),
    .X(_00601_));
 sg13g2_mux2_1 _20336_ (.A0(\cpu.dcache.r_tag[1][17] ),
    .A1(net391),
    .S(net477),
    .X(_00602_));
 sg13g2_mux2_1 _20337_ (.A0(\cpu.dcache.r_tag[1][18] ),
    .A1(net445),
    .S(net477),
    .X(_00603_));
 sg13g2_mux2_1 _20338_ (.A0(\cpu.dcache.r_tag[1][19] ),
    .A1(net389),
    .S(net477),
    .X(_00604_));
 sg13g2_mux2_1 _20339_ (.A0(\cpu.dcache.r_tag[1][20] ),
    .A1(net444),
    .S(_03074_),
    .X(_00605_));
 sg13g2_mux2_1 _20340_ (.A0(\cpu.dcache.r_tag[1][21] ),
    .A1(net387),
    .S(net477),
    .X(_00606_));
 sg13g2_mux2_1 _20341_ (.A0(\cpu.dcache.r_tag[1][22] ),
    .A1(net443),
    .S(_03074_),
    .X(_00607_));
 sg13g2_mux2_1 _20342_ (.A0(\cpu.dcache.r_tag[1][23] ),
    .A1(_09614_),
    .S(net477),
    .X(_00608_));
 sg13g2_buf_1 _20343_ (.A(net890),
    .X(_03075_));
 sg13g2_buf_1 _20344_ (.A(_12409_),
    .X(_03076_));
 sg13g2_mux2_1 _20345_ (.A0(\cpu.dcache.r_tag[1][6] ),
    .A1(net750),
    .S(net476),
    .X(_00609_));
 sg13g2_buf_2 _20346_ (.A(net1154),
    .X(_03077_));
 sg13g2_buf_1 _20347_ (.A(net997),
    .X(_03078_));
 sg13g2_mux2_1 _20348_ (.A0(\cpu.dcache.r_tag[1][7] ),
    .A1(net884),
    .S(net476),
    .X(_00610_));
 sg13g2_buf_1 _20349_ (.A(_09165_),
    .X(_03079_));
 sg13g2_buf_1 _20350_ (.A(net996),
    .X(_03080_));
 sg13g2_mux2_1 _20351_ (.A0(\cpu.dcache.r_tag[1][8] ),
    .A1(net883),
    .S(net476),
    .X(_00611_));
 sg13g2_buf_1 _20352_ (.A(_10234_),
    .X(_03081_));
 sg13g2_buf_1 _20353_ (.A(net995),
    .X(_03082_));
 sg13g2_mux2_1 _20354_ (.A0(\cpu.dcache.r_tag[1][9] ),
    .A1(net882),
    .S(net476),
    .X(_00612_));
 sg13g2_buf_1 _20355_ (.A(net999),
    .X(_03083_));
 sg13g2_mux2_1 _20356_ (.A0(\cpu.dcache.r_tag[1][10] ),
    .A1(net881),
    .S(_03076_),
    .X(_00613_));
 sg13g2_buf_1 _20357_ (.A(net998),
    .X(_03084_));
 sg13g2_mux2_1 _20358_ (.A0(\cpu.dcache.r_tag[1][11] ),
    .A1(net880),
    .S(_03076_),
    .X(_00614_));
 sg13g2_mux2_1 _20359_ (.A0(\cpu.dcache.r_tag[1][12] ),
    .A1(net351),
    .S(net476),
    .X(_00615_));
 sg13g2_mux2_1 _20360_ (.A0(\cpu.dcache.r_tag[1][13] ),
    .A1(net388),
    .S(net476),
    .X(_00616_));
 sg13g2_mux2_1 _20361_ (.A0(\cpu.dcache.r_tag[1][14] ),
    .A1(net446),
    .S(net476),
    .X(_00617_));
 sg13g2_buf_1 _20362_ (.A(_12518_),
    .X(_03085_));
 sg13g2_mux2_1 _20363_ (.A0(\cpu.dcache.r_tag[2][5] ),
    .A1(net542),
    .S(net475),
    .X(_00618_));
 sg13g2_mux2_1 _20364_ (.A0(\cpu.dcache.r_tag[2][15] ),
    .A1(net442),
    .S(net475),
    .X(_00619_));
 sg13g2_mux2_1 _20365_ (.A0(\cpu.dcache.r_tag[2][16] ),
    .A1(net390),
    .S(net475),
    .X(_00620_));
 sg13g2_mux2_1 _20366_ (.A0(\cpu.dcache.r_tag[2][17] ),
    .A1(net391),
    .S(net475),
    .X(_00621_));
 sg13g2_mux2_1 _20367_ (.A0(\cpu.dcache.r_tag[2][18] ),
    .A1(net445),
    .S(net475),
    .X(_00622_));
 sg13g2_mux2_1 _20368_ (.A0(\cpu.dcache.r_tag[2][19] ),
    .A1(net389),
    .S(net475),
    .X(_00623_));
 sg13g2_mux2_1 _20369_ (.A0(\cpu.dcache.r_tag[2][20] ),
    .A1(net444),
    .S(_03085_),
    .X(_00624_));
 sg13g2_mux2_1 _20370_ (.A0(\cpu.dcache.r_tag[2][21] ),
    .A1(net387),
    .S(net475),
    .X(_00625_));
 sg13g2_mux2_1 _20371_ (.A0(\cpu.dcache.r_tag[2][22] ),
    .A1(net443),
    .S(_03085_),
    .X(_00626_));
 sg13g2_buf_1 _20372_ (.A(_12517_),
    .X(_03086_));
 sg13g2_mux2_1 _20373_ (.A0(\cpu.dcache.r_tag[2][23] ),
    .A1(_09614_),
    .S(_03086_),
    .X(_00627_));
 sg13g2_mux2_1 _20374_ (.A0(\cpu.dcache.r_tag[2][6] ),
    .A1(net750),
    .S(_03086_),
    .X(_00628_));
 sg13g2_nand2_1 _20375_ (.Y(_03087_),
    .A(net997),
    .B(net541));
 sg13g2_o21ai_1 _20376_ (.B1(_03087_),
    .Y(_00629_),
    .A1(_09550_),
    .A2(net475));
 sg13g2_mux2_1 _20377_ (.A0(\cpu.dcache.r_tag[2][8] ),
    .A1(net883),
    .S(net541),
    .X(_00630_));
 sg13g2_mux2_1 _20378_ (.A0(\cpu.dcache.r_tag[2][9] ),
    .A1(net882),
    .S(net541),
    .X(_00631_));
 sg13g2_mux2_1 _20379_ (.A0(\cpu.dcache.r_tag[2][10] ),
    .A1(net881),
    .S(net541),
    .X(_00632_));
 sg13g2_mux2_1 _20380_ (.A0(\cpu.dcache.r_tag[2][11] ),
    .A1(net880),
    .S(net541),
    .X(_00633_));
 sg13g2_mux2_1 _20381_ (.A0(\cpu.dcache.r_tag[2][12] ),
    .A1(net351),
    .S(net541),
    .X(_00634_));
 sg13g2_mux2_1 _20382_ (.A0(\cpu.dcache.r_tag[2][13] ),
    .A1(net388),
    .S(net541),
    .X(_00635_));
 sg13g2_mux2_1 _20383_ (.A0(\cpu.dcache.r_tag[2][14] ),
    .A1(net446),
    .S(net541),
    .X(_00636_));
 sg13g2_buf_1 _20384_ (.A(_12625_),
    .X(_03088_));
 sg13g2_mux2_1 _20385_ (.A0(\cpu.dcache.r_tag[3][5] ),
    .A1(net542),
    .S(net344),
    .X(_00637_));
 sg13g2_mux2_1 _20386_ (.A0(\cpu.dcache.r_tag[3][15] ),
    .A1(_09727_),
    .S(net344),
    .X(_00638_));
 sg13g2_mux2_1 _20387_ (.A0(\cpu.dcache.r_tag[3][16] ),
    .A1(net390),
    .S(net344),
    .X(_00639_));
 sg13g2_mux2_1 _20388_ (.A0(\cpu.dcache.r_tag[3][17] ),
    .A1(net391),
    .S(net344),
    .X(_00640_));
 sg13g2_mux2_1 _20389_ (.A0(\cpu.dcache.r_tag[3][18] ),
    .A1(net445),
    .S(net344),
    .X(_00641_));
 sg13g2_mux2_1 _20390_ (.A0(\cpu.dcache.r_tag[3][19] ),
    .A1(net389),
    .S(net344),
    .X(_00642_));
 sg13g2_mux2_1 _20391_ (.A0(\cpu.dcache.r_tag[3][20] ),
    .A1(_09680_),
    .S(_03088_),
    .X(_00643_));
 sg13g2_mux2_1 _20392_ (.A0(\cpu.dcache.r_tag[3][21] ),
    .A1(net387),
    .S(net344),
    .X(_00644_));
 sg13g2_mux2_1 _20393_ (.A0(\cpu.dcache.r_tag[3][22] ),
    .A1(net443),
    .S(_03088_),
    .X(_00645_));
 sg13g2_mux2_1 _20394_ (.A0(\cpu.dcache.r_tag[3][23] ),
    .A1(_09614_),
    .S(net344),
    .X(_00646_));
 sg13g2_buf_1 _20395_ (.A(_12625_),
    .X(_03089_));
 sg13g2_mux2_1 _20396_ (.A0(\cpu.dcache.r_tag[3][6] ),
    .A1(net750),
    .S(_03089_),
    .X(_00647_));
 sg13g2_mux2_1 _20397_ (.A0(\cpu.dcache.r_tag[3][7] ),
    .A1(net884),
    .S(net343),
    .X(_00648_));
 sg13g2_mux2_1 _20398_ (.A0(\cpu.dcache.r_tag[3][8] ),
    .A1(net883),
    .S(net343),
    .X(_00649_));
 sg13g2_mux2_1 _20399_ (.A0(\cpu.dcache.r_tag[3][9] ),
    .A1(net882),
    .S(net343),
    .X(_00650_));
 sg13g2_mux2_1 _20400_ (.A0(\cpu.dcache.r_tag[3][10] ),
    .A1(net881),
    .S(_03089_),
    .X(_00651_));
 sg13g2_mux2_1 _20401_ (.A0(\cpu.dcache.r_tag[3][11] ),
    .A1(net880),
    .S(net343),
    .X(_00652_));
 sg13g2_mux2_1 _20402_ (.A0(\cpu.dcache.r_tag[3][12] ),
    .A1(net351),
    .S(net343),
    .X(_00653_));
 sg13g2_mux2_1 _20403_ (.A0(\cpu.dcache.r_tag[3][13] ),
    .A1(net388),
    .S(net343),
    .X(_00654_));
 sg13g2_mux2_1 _20404_ (.A0(\cpu.dcache.r_tag[3][14] ),
    .A1(net446),
    .S(net343),
    .X(_00655_));
 sg13g2_buf_1 _20405_ (.A(net346),
    .X(_03090_));
 sg13g2_buf_1 _20406_ (.A(net346),
    .X(_03091_));
 sg13g2_nand2_1 _20407_ (.Y(_03092_),
    .A(\cpu.dcache.r_tag[4][5] ),
    .B(net297));
 sg13g2_o21ai_1 _20408_ (.B1(_03092_),
    .Y(_00656_),
    .A1(net674),
    .A2(net298));
 sg13g2_mux2_1 _20409_ (.A0(_09727_),
    .A1(\cpu.dcache.r_tag[4][15] ),
    .S(_03090_),
    .X(_00657_));
 sg13g2_mux2_1 _20410_ (.A0(net390),
    .A1(\cpu.dcache.r_tag[4][16] ),
    .S(net298),
    .X(_00658_));
 sg13g2_mux2_1 _20411_ (.A0(net391),
    .A1(\cpu.dcache.r_tag[4][17] ),
    .S(_03090_),
    .X(_00659_));
 sg13g2_mux2_1 _20412_ (.A0(_09658_),
    .A1(\cpu.dcache.r_tag[4][18] ),
    .S(net298),
    .X(_00660_));
 sg13g2_mux2_1 _20413_ (.A0(net389),
    .A1(\cpu.dcache.r_tag[4][19] ),
    .S(net298),
    .X(_00661_));
 sg13g2_mux2_1 _20414_ (.A0(net444),
    .A1(\cpu.dcache.r_tag[4][20] ),
    .S(_03091_),
    .X(_00662_));
 sg13g2_mux2_1 _20415_ (.A0(net387),
    .A1(\cpu.dcache.r_tag[4][21] ),
    .S(net297),
    .X(_00663_));
 sg13g2_mux2_1 _20416_ (.A0(net443),
    .A1(\cpu.dcache.r_tag[4][22] ),
    .S(_03091_),
    .X(_00664_));
 sg13g2_nand2_1 _20417_ (.Y(_03093_),
    .A(\cpu.dcache.r_tag[4][23] ),
    .B(net346));
 sg13g2_o21ai_1 _20418_ (.B1(_03093_),
    .Y(_00665_),
    .A1(_09789_),
    .A2(net298));
 sg13g2_mux2_1 _20419_ (.A0(net754),
    .A1(\cpu.dcache.r_tag[4][6] ),
    .S(net297),
    .X(_00666_));
 sg13g2_nand2_1 _20420_ (.Y(_03094_),
    .A(\cpu.dcache.r_tag[4][7] ),
    .B(net346));
 sg13g2_o21ai_1 _20421_ (.B1(_03094_),
    .Y(_00667_),
    .A1(net753),
    .A2(net298));
 sg13g2_nand2_1 _20422_ (.Y(_03095_),
    .A(\cpu.dcache.r_tag[4][8] ),
    .B(_12734_));
 sg13g2_o21ai_1 _20423_ (.B1(_03095_),
    .Y(_00668_),
    .A1(net752),
    .A2(net298));
 sg13g2_nand2_1 _20424_ (.Y(_03096_),
    .A(\cpu.dcache.r_tag[4][9] ),
    .B(_12734_));
 sg13g2_o21ai_1 _20425_ (.B1(_03096_),
    .Y(_00669_),
    .A1(net751),
    .A2(net298));
 sg13g2_mux2_1 _20426_ (.A0(net886),
    .A1(\cpu.dcache.r_tag[4][10] ),
    .S(net297),
    .X(_00670_));
 sg13g2_mux2_1 _20427_ (.A0(net885),
    .A1(\cpu.dcache.r_tag[4][11] ),
    .S(net297),
    .X(_00671_));
 sg13g2_mux2_1 _20428_ (.A0(net351),
    .A1(\cpu.dcache.r_tag[4][12] ),
    .S(net297),
    .X(_00672_));
 sg13g2_mux2_1 _20429_ (.A0(net388),
    .A1(\cpu.dcache.r_tag[4][13] ),
    .S(net297),
    .X(_00673_));
 sg13g2_mux2_1 _20430_ (.A0(net446),
    .A1(\cpu.dcache.r_tag[4][14] ),
    .S(net297),
    .X(_00674_));
 sg13g2_buf_1 _20431_ (.A(net550),
    .X(_03097_));
 sg13g2_mux2_1 _20432_ (.A0(\cpu.dcache.r_tag[5][5] ),
    .A1(net542),
    .S(net474),
    .X(_00675_));
 sg13g2_mux2_1 _20433_ (.A0(\cpu.dcache.r_tag[5][15] ),
    .A1(net442),
    .S(net474),
    .X(_00676_));
 sg13g2_mux2_1 _20434_ (.A0(\cpu.dcache.r_tag[5][16] ),
    .A1(_09387_),
    .S(net474),
    .X(_00677_));
 sg13g2_mux2_1 _20435_ (.A0(\cpu.dcache.r_tag[5][17] ),
    .A1(_09331_),
    .S(net474),
    .X(_00678_));
 sg13g2_mux2_1 _20436_ (.A0(\cpu.dcache.r_tag[5][18] ),
    .A1(net445),
    .S(net474),
    .X(_00679_));
 sg13g2_mux2_1 _20437_ (.A0(\cpu.dcache.r_tag[5][19] ),
    .A1(net389),
    .S(net474),
    .X(_00680_));
 sg13g2_mux2_1 _20438_ (.A0(\cpu.dcache.r_tag[5][20] ),
    .A1(net444),
    .S(_03097_),
    .X(_00681_));
 sg13g2_mux2_1 _20439_ (.A0(\cpu.dcache.r_tag[5][21] ),
    .A1(net387),
    .S(net474),
    .X(_00682_));
 sg13g2_mux2_1 _20440_ (.A0(\cpu.dcache.r_tag[5][22] ),
    .A1(net443),
    .S(_03097_),
    .X(_00683_));
 sg13g2_buf_1 _20441_ (.A(_02755_),
    .X(_03098_));
 sg13g2_mux2_1 _20442_ (.A0(\cpu.dcache.r_tag[5][23] ),
    .A1(_09614_),
    .S(net540),
    .X(_00684_));
 sg13g2_mux2_1 _20443_ (.A0(\cpu.dcache.r_tag[5][6] ),
    .A1(net750),
    .S(net540),
    .X(_00685_));
 sg13g2_nand2_1 _20444_ (.Y(_03099_),
    .A(net997),
    .B(net540));
 sg13g2_o21ai_1 _20445_ (.B1(_03099_),
    .Y(_00686_),
    .A1(_09545_),
    .A2(net474));
 sg13g2_mux2_1 _20446_ (.A0(\cpu.dcache.r_tag[5][8] ),
    .A1(net883),
    .S(_03098_),
    .X(_00687_));
 sg13g2_mux2_1 _20447_ (.A0(\cpu.dcache.r_tag[5][9] ),
    .A1(net882),
    .S(_03098_),
    .X(_00688_));
 sg13g2_mux2_1 _20448_ (.A0(\cpu.dcache.r_tag[5][10] ),
    .A1(net881),
    .S(net540),
    .X(_00689_));
 sg13g2_mux2_1 _20449_ (.A0(\cpu.dcache.r_tag[5][11] ),
    .A1(net880),
    .S(net540),
    .X(_00690_));
 sg13g2_mux2_1 _20450_ (.A0(\cpu.dcache.r_tag[5][12] ),
    .A1(net351),
    .S(net540),
    .X(_00691_));
 sg13g2_mux2_1 _20451_ (.A0(\cpu.dcache.r_tag[5][13] ),
    .A1(net388),
    .S(net540),
    .X(_00692_));
 sg13g2_mux2_1 _20452_ (.A0(\cpu.dcache.r_tag[5][14] ),
    .A1(net446),
    .S(net540),
    .X(_00693_));
 sg13g2_buf_1 _20453_ (.A(net549),
    .X(_03100_));
 sg13g2_mux2_1 _20454_ (.A0(\cpu.dcache.r_tag[6][5] ),
    .A1(net542),
    .S(net473),
    .X(_00694_));
 sg13g2_mux2_1 _20455_ (.A0(\cpu.dcache.r_tag[6][15] ),
    .A1(net442),
    .S(net473),
    .X(_00695_));
 sg13g2_mux2_1 _20456_ (.A0(\cpu.dcache.r_tag[6][16] ),
    .A1(_09387_),
    .S(net473),
    .X(_00696_));
 sg13g2_mux2_1 _20457_ (.A0(\cpu.dcache.r_tag[6][17] ),
    .A1(_09331_),
    .S(net473),
    .X(_00697_));
 sg13g2_mux2_1 _20458_ (.A0(\cpu.dcache.r_tag[6][18] ),
    .A1(net445),
    .S(net473),
    .X(_00698_));
 sg13g2_mux2_1 _20459_ (.A0(\cpu.dcache.r_tag[6][19] ),
    .A1(net389),
    .S(net473),
    .X(_00699_));
 sg13g2_mux2_1 _20460_ (.A0(\cpu.dcache.r_tag[6][20] ),
    .A1(net444),
    .S(_03100_),
    .X(_00700_));
 sg13g2_mux2_1 _20461_ (.A0(\cpu.dcache.r_tag[6][21] ),
    .A1(net387),
    .S(net473),
    .X(_00701_));
 sg13g2_mux2_1 _20462_ (.A0(\cpu.dcache.r_tag[6][22] ),
    .A1(net443),
    .S(_03100_),
    .X(_00702_));
 sg13g2_buf_1 _20463_ (.A(_02860_),
    .X(_03101_));
 sg13g2_mux2_1 _20464_ (.A0(\cpu.dcache.r_tag[6][23] ),
    .A1(_09614_),
    .S(_03101_),
    .X(_00703_));
 sg13g2_buf_1 _20465_ (.A(net890),
    .X(_03102_));
 sg13g2_mux2_1 _20466_ (.A0(\cpu.dcache.r_tag[6][6] ),
    .A1(net749),
    .S(net539),
    .X(_00704_));
 sg13g2_nand2_1 _20467_ (.Y(_03103_),
    .A(net997),
    .B(net539));
 sg13g2_o21ai_1 _20468_ (.B1(_03103_),
    .Y(_00705_),
    .A1(_09554_),
    .A2(net473));
 sg13g2_mux2_1 _20469_ (.A0(\cpu.dcache.r_tag[6][8] ),
    .A1(net883),
    .S(net539),
    .X(_00706_));
 sg13g2_mux2_1 _20470_ (.A0(\cpu.dcache.r_tag[6][9] ),
    .A1(net882),
    .S(net539),
    .X(_00707_));
 sg13g2_buf_1 _20471_ (.A(net999),
    .X(_03104_));
 sg13g2_mux2_1 _20472_ (.A0(\cpu.dcache.r_tag[6][10] ),
    .A1(net879),
    .S(_03101_),
    .X(_00708_));
 sg13g2_buf_1 _20473_ (.A(net998),
    .X(_03105_));
 sg13g2_mux2_1 _20474_ (.A0(\cpu.dcache.r_tag[6][11] ),
    .A1(net878),
    .S(net539),
    .X(_00709_));
 sg13g2_mux2_1 _20475_ (.A0(\cpu.dcache.r_tag[6][12] ),
    .A1(net351),
    .S(net539),
    .X(_00710_));
 sg13g2_mux2_1 _20476_ (.A0(\cpu.dcache.r_tag[6][13] ),
    .A1(net388),
    .S(net539),
    .X(_00711_));
 sg13g2_mux2_1 _20477_ (.A0(\cpu.dcache.r_tag[6][14] ),
    .A1(net446),
    .S(net539),
    .X(_00712_));
 sg13g2_buf_1 _20478_ (.A(_02966_),
    .X(_03106_));
 sg13g2_mux2_1 _20479_ (.A0(\cpu.dcache.r_tag[7][5] ),
    .A1(net542),
    .S(net296),
    .X(_00713_));
 sg13g2_mux2_1 _20480_ (.A0(\cpu.dcache.r_tag[7][15] ),
    .A1(net442),
    .S(net296),
    .X(_00714_));
 sg13g2_mux2_1 _20481_ (.A0(\cpu.dcache.r_tag[7][16] ),
    .A1(net390),
    .S(net296),
    .X(_00715_));
 sg13g2_mux2_1 _20482_ (.A0(\cpu.dcache.r_tag[7][17] ),
    .A1(net391),
    .S(net296),
    .X(_00716_));
 sg13g2_mux2_1 _20483_ (.A0(\cpu.dcache.r_tag[7][18] ),
    .A1(_09658_),
    .S(net296),
    .X(_00717_));
 sg13g2_mux2_1 _20484_ (.A0(\cpu.dcache.r_tag[7][19] ),
    .A1(net389),
    .S(net296),
    .X(_00718_));
 sg13g2_mux2_1 _20485_ (.A0(\cpu.dcache.r_tag[7][20] ),
    .A1(net444),
    .S(_03106_),
    .X(_00719_));
 sg13g2_mux2_1 _20486_ (.A0(\cpu.dcache.r_tag[7][21] ),
    .A1(_09635_),
    .S(net296),
    .X(_00720_));
 sg13g2_mux2_1 _20487_ (.A0(\cpu.dcache.r_tag[7][22] ),
    .A1(net443),
    .S(_03106_),
    .X(_00721_));
 sg13g2_mux2_1 _20488_ (.A0(\cpu.dcache.r_tag[7][23] ),
    .A1(_09614_),
    .S(net296),
    .X(_00722_));
 sg13g2_buf_1 _20489_ (.A(_02966_),
    .X(_03107_));
 sg13g2_mux2_1 _20490_ (.A0(\cpu.dcache.r_tag[7][6] ),
    .A1(net749),
    .S(net295),
    .X(_00723_));
 sg13g2_mux2_1 _20491_ (.A0(\cpu.dcache.r_tag[7][7] ),
    .A1(net884),
    .S(net295),
    .X(_00724_));
 sg13g2_mux2_1 _20492_ (.A0(\cpu.dcache.r_tag[7][8] ),
    .A1(net883),
    .S(net295),
    .X(_00725_));
 sg13g2_mux2_1 _20493_ (.A0(\cpu.dcache.r_tag[7][9] ),
    .A1(net882),
    .S(net295),
    .X(_00726_));
 sg13g2_mux2_1 _20494_ (.A0(\cpu.dcache.r_tag[7][10] ),
    .A1(net879),
    .S(_03107_),
    .X(_00727_));
 sg13g2_mux2_1 _20495_ (.A0(\cpu.dcache.r_tag[7][11] ),
    .A1(net878),
    .S(_03107_),
    .X(_00728_));
 sg13g2_mux2_1 _20496_ (.A0(\cpu.dcache.r_tag[7][12] ),
    .A1(net351),
    .S(net295),
    .X(_00729_));
 sg13g2_mux2_1 _20497_ (.A0(\cpu.dcache.r_tag[7][13] ),
    .A1(net388),
    .S(net295),
    .X(_00730_));
 sg13g2_mux2_1 _20498_ (.A0(\cpu.dcache.r_tag[7][14] ),
    .A1(net446),
    .S(net295),
    .X(_00731_));
 sg13g2_buf_1 _20499_ (.A(_09840_),
    .X(_03108_));
 sg13g2_nor2_1 _20500_ (.A(net174),
    .B(net210),
    .Y(_03109_));
 sg13g2_buf_1 _20501_ (.A(_03109_),
    .X(_03110_));
 sg13g2_buf_1 _20502_ (.A(_03110_),
    .X(_03111_));
 sg13g2_buf_1 _20503_ (.A(_09834_),
    .X(_03112_));
 sg13g2_nor2_1 _20504_ (.A(net222),
    .B(net263),
    .Y(_03113_));
 sg13g2_buf_1 _20505_ (.A(_03113_),
    .X(_03114_));
 sg13g2_a21oi_1 _20506_ (.A1(net819),
    .A2(_08956_),
    .Y(_03115_),
    .B1(_08967_));
 sg13g2_buf_1 _20507_ (.A(_03115_),
    .X(_03116_));
 sg13g2_nor2_2 _20508_ (.A(_08931_),
    .B(net251),
    .Y(_03117_));
 sg13g2_a21oi_1 _20509_ (.A1(net236),
    .A2(net173),
    .Y(_03118_),
    .B1(_03117_));
 sg13g2_nor2_1 _20510_ (.A(net186),
    .B(_03118_),
    .Y(_03119_));
 sg13g2_a21oi_1 _20511_ (.A1(net187),
    .A2(net89),
    .Y(_03120_),
    .B1(_03119_));
 sg13g2_nand2_1 _20512_ (.Y(_03121_),
    .A(net1038),
    .B(_09101_));
 sg13g2_o21ai_1 _20513_ (.B1(_03121_),
    .Y(_00740_),
    .A1(net93),
    .A2(_03120_));
 sg13g2_buf_1 _20514_ (.A(net263),
    .X(_03122_));
 sg13g2_buf_1 _20515_ (.A(net221),
    .X(_03123_));
 sg13g2_inv_1 _20516_ (.Y(_03124_),
    .A(_09073_));
 sg13g2_buf_1 _20517_ (.A(_03124_),
    .X(_03125_));
 sg13g2_a22oi_1 _20518_ (.Y(_03126_),
    .B1(net294),
    .B2(net186),
    .A2(net209),
    .A1(net222));
 sg13g2_buf_1 _20519_ (.A(_08931_),
    .X(_03127_));
 sg13g2_buf_1 _20520_ (.A(net220),
    .X(_03128_));
 sg13g2_nand2_1 _20521_ (.Y(_03129_),
    .A(net197),
    .B(net158));
 sg13g2_o21ai_1 _20522_ (.B1(_03129_),
    .Y(_03130_),
    .A1(net198),
    .A2(_03126_));
 sg13g2_buf_1 _20523_ (.A(net251),
    .X(_03131_));
 sg13g2_buf_1 _20524_ (.A(_09821_),
    .X(_03132_));
 sg13g2_nor2_1 _20525_ (.A(net196),
    .B(net186),
    .Y(_03133_));
 sg13g2_nor2_1 _20526_ (.A(net219),
    .B(_03133_),
    .Y(_03134_));
 sg13g2_buf_1 _20527_ (.A(_08948_),
    .X(_03135_));
 sg13g2_buf_1 _20528_ (.A(net250),
    .X(_03136_));
 sg13g2_buf_1 _20529_ (.A(net218),
    .X(_03137_));
 sg13g2_o21ai_1 _20530_ (.B1(net195),
    .Y(_03138_),
    .A1(_03110_),
    .A2(_03134_));
 sg13g2_nor2b_1 _20531_ (.A(_03130_),
    .B_N(_03138_),
    .Y(_03139_));
 sg13g2_buf_1 _20532_ (.A(_08374_),
    .X(_03140_));
 sg13g2_buf_1 _20533_ (.A(net994),
    .X(_03141_));
 sg13g2_buf_1 _20534_ (.A(net877),
    .X(_03142_));
 sg13g2_nand2_1 _20535_ (.Y(_03143_),
    .A(_03142_),
    .B(net112));
 sg13g2_o21ai_1 _20536_ (.B1(_03143_),
    .Y(_00741_),
    .A1(net93),
    .A2(_03139_));
 sg13g2_nand2_1 _20537_ (.Y(_03144_),
    .A(_09840_),
    .B(net210));
 sg13g2_buf_1 _20538_ (.A(_03144_),
    .X(_03145_));
 sg13g2_nand2_1 _20539_ (.Y(_03146_),
    .A(net196),
    .B(net263));
 sg13g2_buf_1 _20540_ (.A(_03146_),
    .X(_03147_));
 sg13g2_nor3_1 _20541_ (.A(net113),
    .B(net145),
    .C(net144),
    .Y(_03148_));
 sg13g2_a21o_1 _20542_ (.A2(net92),
    .A1(\cpu.cond[1] ),
    .B1(_03148_),
    .X(_00742_));
 sg13g2_a22oi_1 _20543_ (.Y(_03149_),
    .B1(net89),
    .B2(net219),
    .A2(net144),
    .A1(net158));
 sg13g2_nand2_1 _20544_ (.Y(_03150_),
    .A(\cpu.cond[2] ),
    .B(net112));
 sg13g2_o21ai_1 _20545_ (.B1(_03150_),
    .Y(_00743_),
    .A1(net93),
    .A2(_03149_));
 sg13g2_nor4_1 _20546_ (.A(net156),
    .B(net145),
    .C(_09088_),
    .D(_09090_),
    .Y(_03151_));
 sg13g2_mux2_1 _20547_ (.A0(_03151_),
    .A1(_09277_),
    .S(net94),
    .X(_00744_));
 sg13g2_nand2_1 _20548_ (.Y(_03152_),
    .A(_09077_),
    .B(_09838_));
 sg13g2_nor2_1 _20549_ (.A(_00167_),
    .B(net734),
    .Y(_03153_));
 sg13g2_mux2_1 _20550_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(\cpu.icache.r_data[7][24] ),
    .S(net936),
    .X(_03154_));
 sg13g2_a22oi_1 _20551_ (.Y(_03155_),
    .B1(_03154_),
    .B2(net1077),
    .A2(_08891_),
    .A1(\cpu.icache.r_data[6][24] ));
 sg13g2_nor2_1 _20552_ (.A(net824),
    .B(_03155_),
    .Y(_03156_));
 sg13g2_a22oi_1 _20553_ (.Y(_03157_),
    .B1(_08593_),
    .B2(\cpu.icache.r_data[4][24] ),
    .A2(_08527_),
    .A1(\cpu.icache.r_data[3][24] ));
 sg13g2_a22oi_1 _20554_ (.Y(_03158_),
    .B1(net654),
    .B2(\cpu.icache.r_data[2][24] ),
    .A2(net655),
    .A1(\cpu.icache.r_data[1][24] ));
 sg13g2_nand2_1 _20555_ (.Y(_03159_),
    .A(_03157_),
    .B(_03158_));
 sg13g2_nor3_1 _20556_ (.A(_03153_),
    .B(_03156_),
    .C(_03159_),
    .Y(_03160_));
 sg13g2_nand2_1 _20557_ (.Y(_03161_),
    .A(_00166_),
    .B(net720));
 sg13g2_a22oi_1 _20558_ (.Y(_03162_),
    .B1(_08531_),
    .B2(\cpu.icache.r_data[5][8] ),
    .A2(_08477_),
    .A1(\cpu.icache.r_data[1][8] ));
 sg13g2_a22oi_1 _20559_ (.Y(_03163_),
    .B1(_08592_),
    .B2(\cpu.icache.r_data[4][8] ),
    .A2(_08486_),
    .A1(\cpu.icache.r_data[2][8] ));
 sg13g2_mux2_1 _20560_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(\cpu.icache.r_data[3][8] ),
    .S(net1079),
    .X(_03164_));
 sg13g2_a22oi_1 _20561_ (.Y(_03165_),
    .B1(_03164_),
    .B2(_08470_),
    .A2(_08481_),
    .A1(\cpu.icache.r_data[6][8] ));
 sg13g2_nand2b_1 _20562_ (.Y(_03166_),
    .B(net828),
    .A_N(_03165_));
 sg13g2_nand4_1 _20563_ (.B(_03162_),
    .C(_03163_),
    .A(net734),
    .Y(_03167_),
    .D(_03166_));
 sg13g2_a21oi_1 _20564_ (.A1(_03161_),
    .A2(_03167_),
    .Y(_03168_),
    .B1(net1074));
 sg13g2_a21oi_1 _20565_ (.A1(net1074),
    .A2(_03160_),
    .Y(_03169_),
    .B1(_03168_));
 sg13g2_buf_1 _20566_ (.A(_03169_),
    .X(_03170_));
 sg13g2_inv_1 _20567_ (.Y(_03171_),
    .A(_00168_));
 sg13g2_a22oi_1 _20568_ (.Y(_03172_),
    .B1(_08531_),
    .B2(\cpu.icache.r_data[5][9] ),
    .A2(_08513_),
    .A1(\cpu.icache.r_data[1][9] ));
 sg13g2_a22oi_1 _20569_ (.Y(_03173_),
    .B1(_08528_),
    .B2(\cpu.icache.r_data[3][9] ),
    .A2(_08518_),
    .A1(\cpu.icache.r_data[2][9] ));
 sg13g2_mux2_1 _20570_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(net1078),
    .X(_03174_));
 sg13g2_a22oi_1 _20571_ (.Y(_03175_),
    .B1(_03174_),
    .B2(net941),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][9] ));
 sg13g2_or2_1 _20572_ (.X(_03176_),
    .B(_03175_),
    .A(net938));
 sg13g2_nand4_1 _20573_ (.B(_03172_),
    .C(_03173_),
    .A(net734),
    .Y(_03177_),
    .D(_03176_));
 sg13g2_o21ai_1 _20574_ (.B1(_03177_),
    .Y(_03178_),
    .A1(_03171_),
    .A2(net658));
 sg13g2_nor2_1 _20575_ (.A(_00169_),
    .B(net734),
    .Y(_03179_));
 sg13g2_mux2_1 _20576_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(net936),
    .X(_03180_));
 sg13g2_a22oi_1 _20577_ (.Y(_03181_),
    .B1(_03180_),
    .B2(net820),
    .A2(_08597_),
    .A1(\cpu.icache.r_data[7][25] ));
 sg13g2_nor2_1 _20578_ (.A(net824),
    .B(_03181_),
    .Y(_03182_));
 sg13g2_a22oi_1 _20579_ (.Y(_03183_),
    .B1(_08531_),
    .B2(\cpu.icache.r_data[5][25] ),
    .A2(_08513_),
    .A1(\cpu.icache.r_data[1][25] ));
 sg13g2_a22oi_1 _20580_ (.Y(_03184_),
    .B1(_08528_),
    .B2(\cpu.icache.r_data[3][25] ),
    .A2(_08518_),
    .A1(\cpu.icache.r_data[2][25] ));
 sg13g2_nand2_1 _20581_ (.Y(_03185_),
    .A(_03183_),
    .B(_03184_));
 sg13g2_nor4_1 _20582_ (.A(net934),
    .B(_03179_),
    .C(_03182_),
    .D(_03185_),
    .Y(_03186_));
 sg13g2_a21oi_1 _20583_ (.A1(_08958_),
    .A2(_03178_),
    .Y(_03187_),
    .B1(_03186_));
 sg13g2_buf_2 _20584_ (.A(_03187_),
    .X(_03188_));
 sg13g2_nor2_1 _20585_ (.A(_00165_),
    .B(_08458_),
    .Y(_03189_));
 sg13g2_mux2_1 _20586_ (.A0(\cpu.icache.r_data[5][23] ),
    .A1(\cpu.icache.r_data[7][23] ),
    .S(net944),
    .X(_03190_));
 sg13g2_a22oi_1 _20587_ (.Y(_03191_),
    .B1(_03190_),
    .B2(net942),
    .A2(_08891_),
    .A1(\cpu.icache.r_data[6][23] ));
 sg13g2_nor2_1 _20588_ (.A(net719),
    .B(_03191_),
    .Y(_03192_));
 sg13g2_a22oi_1 _20589_ (.Y(_03193_),
    .B1(_08593_),
    .B2(\cpu.icache.r_data[4][23] ),
    .A2(net572),
    .A1(\cpu.icache.r_data[3][23] ));
 sg13g2_a22oi_1 _20590_ (.Y(_03194_),
    .B1(_08519_),
    .B2(\cpu.icache.r_data[2][23] ),
    .A2(net574),
    .A1(\cpu.icache.r_data[1][23] ));
 sg13g2_nand2_1 _20591_ (.Y(_03195_),
    .A(_03193_),
    .B(_03194_));
 sg13g2_nor3_1 _20592_ (.A(_03189_),
    .B(_03192_),
    .C(_03195_),
    .Y(_03196_));
 sg13g2_nand2_1 _20593_ (.Y(_03197_),
    .A(_00164_),
    .B(net650));
 sg13g2_a22oi_1 _20594_ (.Y(_03198_),
    .B1(_08567_),
    .B2(\cpu.icache.r_data[6][7] ),
    .A2(net656),
    .A1(\cpu.icache.r_data[2][7] ));
 sg13g2_a22oi_1 _20595_ (.Y(_03199_),
    .B1(net572),
    .B2(\cpu.icache.r_data[3][7] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_data[1][7] ));
 sg13g2_mux2_1 _20596_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(\cpu.icache.r_data[7][7] ),
    .S(net936),
    .X(_03200_));
 sg13g2_a22oi_1 _20597_ (.Y(_03201_),
    .B1(_03200_),
    .B2(_08470_),
    .A2(_08572_),
    .A1(\cpu.icache.r_data[4][7] ));
 sg13g2_or2_1 _20598_ (.X(_03202_),
    .B(_03201_),
    .A(_08570_));
 sg13g2_nand4_1 _20599_ (.B(_03198_),
    .C(_03199_),
    .A(net659),
    .Y(_03203_),
    .D(_03202_));
 sg13g2_a21oi_1 _20600_ (.A1(_03197_),
    .A2(_03203_),
    .Y(_03204_),
    .B1(net1074));
 sg13g2_a21oi_1 _20601_ (.A1(net935),
    .A2(_03196_),
    .Y(_03205_),
    .B1(_03204_));
 sg13g2_nor3_1 _20602_ (.A(net342),
    .B(_03188_),
    .C(_03205_),
    .Y(_03206_));
 sg13g2_nor2_1 _20603_ (.A(_03124_),
    .B(_09816_),
    .Y(_03207_));
 sg13g2_and2_1 _20604_ (.A(_03206_),
    .B(_03207_),
    .X(_03208_));
 sg13g2_buf_1 _20605_ (.A(_03208_),
    .X(_03209_));
 sg13g2_inv_1 _20606_ (.Y(_03210_),
    .A(_03209_));
 sg13g2_inv_1 _20607_ (.Y(_03211_),
    .A(_00174_));
 sg13g2_a22oi_1 _20608_ (.Y(_03212_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][4] ),
    .A2(_08915_),
    .A1(\cpu.icache.r_data[1][4] ));
 sg13g2_buf_1 _20609_ (.A(_08529_),
    .X(_03213_));
 sg13g2_a22oi_1 _20610_ (.Y(_03214_),
    .B1(net472),
    .B2(\cpu.icache.r_data[3][4] ),
    .A2(_08916_),
    .A1(\cpu.icache.r_data[2][4] ));
 sg13g2_mux2_1 _20611_ (.A0(\cpu.icache.r_data[4][4] ),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(net828),
    .X(_03215_));
 sg13g2_a22oi_1 _20612_ (.Y(_03216_),
    .B1(_03215_),
    .B2(net820),
    .A2(net822),
    .A1(\cpu.icache.r_data[7][4] ));
 sg13g2_or2_1 _20613_ (.X(_03217_),
    .B(_03216_),
    .A(net719));
 sg13g2_nand4_1 _20614_ (.B(_03212_),
    .C(_03214_),
    .A(net497),
    .Y(_03218_),
    .D(_03217_));
 sg13g2_o21ai_1 _20615_ (.B1(_03218_),
    .Y(_03219_),
    .A1(_03211_),
    .A2(net497));
 sg13g2_nor2_1 _20616_ (.A(_00175_),
    .B(net497),
    .Y(_03220_));
 sg13g2_mux2_1 _20617_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(net824),
    .X(_03221_));
 sg13g2_a22oi_1 _20618_ (.Y(_03222_),
    .B1(_03221_),
    .B2(_08912_),
    .A2(net830),
    .A1(\cpu.icache.r_data[6][20] ));
 sg13g2_nand2b_1 _20619_ (.Y(_03223_),
    .B(_08814_),
    .A_N(_03222_));
 sg13g2_a22oi_1 _20620_ (.Y(_03224_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][20] ),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][20] ));
 sg13g2_a22oi_1 _20621_ (.Y(_03225_),
    .B1(net726),
    .B2(\cpu.icache.r_data[4][20] ),
    .A2(net494),
    .A1(\cpu.icache.r_data[2][20] ));
 sg13g2_nand3_1 _20622_ (.B(_03224_),
    .C(_03225_),
    .A(_03223_),
    .Y(_03226_));
 sg13g2_o21ai_1 _20623_ (.B1(net935),
    .Y(_03227_),
    .A1(_03220_),
    .A2(_03226_));
 sg13g2_o21ai_1 _20624_ (.B1(_03227_),
    .Y(_03228_),
    .A1(net819),
    .A2(_03219_));
 sg13g2_buf_1 _20625_ (.A(_03228_),
    .X(_03229_));
 sg13g2_buf_1 _20626_ (.A(_03229_),
    .X(_03230_));
 sg13g2_nor4_1 _20627_ (.A(_09090_),
    .B(_03152_),
    .C(_03210_),
    .D(net217),
    .Y(_03231_));
 sg13g2_mux2_1 _20628_ (.A0(_03231_),
    .A1(\cpu.dec.do_flush_all ),
    .S(net94),
    .X(_00745_));
 sg13g2_nor3_2 _20629_ (.A(net220),
    .B(net222),
    .C(net221),
    .Y(_03232_));
 sg13g2_nand2_1 _20630_ (.Y(_03233_),
    .A(_09077_),
    .B(_03232_));
 sg13g2_nand2_1 _20631_ (.Y(_03234_),
    .A(\cpu.dec.do_flush_write ),
    .B(net112));
 sg13g2_o21ai_1 _20632_ (.B1(_03234_),
    .Y(_00746_),
    .A1(net93),
    .A2(_03233_));
 sg13g2_inv_1 _20633_ (.Y(_03235_),
    .A(_00170_));
 sg13g2_a22oi_1 _20634_ (.Y(_03236_),
    .B1(net571),
    .B2(\cpu.icache.r_data[5][2] ),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][2] ));
 sg13g2_a22oi_1 _20635_ (.Y(_03237_),
    .B1(net472),
    .B2(\cpu.icache.r_data[3][2] ),
    .A2(net494),
    .A1(\cpu.icache.r_data[2][2] ));
 sg13g2_mux2_1 _20636_ (.A0(\cpu.icache.r_data[4][2] ),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_08464_),
    .X(_03238_));
 sg13g2_a22oi_1 _20637_ (.Y(_03239_),
    .B1(_03238_),
    .B2(net820),
    .A2(net822),
    .A1(\cpu.icache.r_data[7][2] ));
 sg13g2_or2_1 _20638_ (.X(_03240_),
    .B(_03239_),
    .A(_08888_));
 sg13g2_nand4_1 _20639_ (.B(_03236_),
    .C(_03237_),
    .A(net497),
    .Y(_03241_),
    .D(_03240_));
 sg13g2_o21ai_1 _20640_ (.B1(_03241_),
    .Y(_03242_),
    .A1(_03235_),
    .A2(net497));
 sg13g2_nor2_1 _20641_ (.A(_00171_),
    .B(net497),
    .Y(_03243_));
 sg13g2_mux2_1 _20642_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(net824),
    .X(_03244_));
 sg13g2_a22oi_1 _20643_ (.Y(_03245_),
    .B1(_03244_),
    .B2(_08912_),
    .A2(net830),
    .A1(\cpu.icache.r_data[6][18] ));
 sg13g2_nand2b_1 _20644_ (.Y(_03246_),
    .B(_08814_),
    .A_N(_03245_));
 sg13g2_a22oi_1 _20645_ (.Y(_03247_),
    .B1(_08533_),
    .B2(\cpu.icache.r_data[5][18] ),
    .A2(net494),
    .A1(\cpu.icache.r_data[2][18] ));
 sg13g2_buf_1 _20646_ (.A(_08594_),
    .X(_03248_));
 sg13g2_a22oi_1 _20647_ (.Y(_03249_),
    .B1(net619),
    .B2(\cpu.icache.r_data[4][18] ),
    .A2(net495),
    .A1(\cpu.icache.r_data[1][18] ));
 sg13g2_nand3_1 _20648_ (.B(_03247_),
    .C(_03249_),
    .A(_03246_),
    .Y(_03250_));
 sg13g2_o21ai_1 _20649_ (.B1(_08972_),
    .Y(_03251_),
    .A1(_03243_),
    .A2(_03250_));
 sg13g2_o21ai_1 _20650_ (.B1(_03251_),
    .Y(_03252_),
    .A1(_08972_),
    .A2(_03242_));
 sg13g2_buf_1 _20651_ (.A(_03252_),
    .X(_03253_));
 sg13g2_buf_1 _20652_ (.A(_03253_),
    .X(_03254_));
 sg13g2_a22oi_1 _20653_ (.Y(_03255_),
    .B1(net155),
    .B2(net216),
    .A2(net187),
    .A1(net304));
 sg13g2_nand4_1 _20654_ (.B(net198),
    .C(net154),
    .A(net195),
    .Y(_03256_),
    .D(net217));
 sg13g2_o21ai_1 _20655_ (.B1(_03256_),
    .Y(_03257_),
    .A1(net145),
    .A2(_03255_));
 sg13g2_nor2_1 _20656_ (.A(net251),
    .B(net174),
    .Y(_03258_));
 sg13g2_nor2_1 _20657_ (.A(net250),
    .B(net186),
    .Y(_03259_));
 sg13g2_a22oi_1 _20658_ (.Y(_03260_),
    .B1(_03259_),
    .B2(net144),
    .A2(_03258_),
    .A1(net218));
 sg13g2_nor2_1 _20659_ (.A(net210),
    .B(_03260_),
    .Y(_03261_));
 sg13g2_buf_1 _20660_ (.A(net174),
    .X(_03262_));
 sg13g2_nor3_1 _20661_ (.A(net198),
    .B(net143),
    .C(net209),
    .Y(_03263_));
 sg13g2_o21ai_1 _20662_ (.B1(net304),
    .Y(_03264_),
    .A1(_03261_),
    .A2(_03263_));
 sg13g2_nor2b_1 _20663_ (.A(_03257_),
    .B_N(_03264_),
    .Y(_03265_));
 sg13g2_nand2_1 _20664_ (.Y(_03266_),
    .A(_11168_),
    .B(net112));
 sg13g2_o21ai_1 _20665_ (.B1(_03266_),
    .Y(_00747_),
    .A1(net93),
    .A2(_03265_));
 sg13g2_inv_1 _20666_ (.Y(_03267_),
    .A(\cpu.dec.imm[10] ));
 sg13g2_buf_1 _20667_ (.A(_09056_),
    .X(_03268_));
 sg13g2_nand2_1 _20668_ (.Y(_03269_),
    .A(net174),
    .B(net236));
 sg13g2_nand2b_1 _20669_ (.Y(_03270_),
    .B(_09077_),
    .A_N(_09837_));
 sg13g2_buf_1 _20670_ (.A(_03270_),
    .X(_03271_));
 sg13g2_nand2_1 _20671_ (.Y(_03272_),
    .A(_03269_),
    .B(_03271_));
 sg13g2_nand2_1 _20672_ (.Y(_03273_),
    .A(net294),
    .B(_03117_));
 sg13g2_buf_2 _20673_ (.A(_03273_),
    .X(_03274_));
 sg13g2_nand2_1 _20674_ (.Y(_03275_),
    .A(net220),
    .B(net221));
 sg13g2_nor2_1 _20675_ (.A(net222),
    .B(_03275_),
    .Y(_03276_));
 sg13g2_nand2_1 _20676_ (.Y(_03277_),
    .A(net217),
    .B(_03276_));
 sg13g2_o21ai_1 _20677_ (.B1(_03277_),
    .Y(_03278_),
    .A1(_03274_),
    .A2(_03271_));
 sg13g2_o21ai_1 _20678_ (.B1(net158),
    .Y(_03279_),
    .A1(_09836_),
    .A2(net217));
 sg13g2_buf_1 _20679_ (.A(_03279_),
    .X(_03280_));
 sg13g2_nand2_1 _20680_ (.Y(_03281_),
    .A(_09836_),
    .B(_03274_));
 sg13g2_a21oi_1 _20681_ (.A1(net173),
    .A2(net342),
    .Y(_03282_),
    .B1(_03281_));
 sg13g2_nor2_1 _20682_ (.A(_03280_),
    .B(_03282_),
    .Y(_03283_));
 sg13g2_a21oi_1 _20683_ (.A1(_03272_),
    .A2(_03278_),
    .Y(_03284_),
    .B1(_03283_));
 sg13g2_nor3_2 _20684_ (.A(_09821_),
    .B(net222),
    .C(net263),
    .Y(_03285_));
 sg13g2_mux2_1 _20685_ (.A0(_08971_),
    .A1(_03285_),
    .S(_09009_),
    .X(_03286_));
 sg13g2_and3_1 _20686_ (.X(_03287_),
    .A(_09826_),
    .B(net217),
    .C(_03286_));
 sg13g2_nor2_1 _20687_ (.A(_12041_),
    .B(_03287_),
    .Y(_03288_));
 sg13g2_buf_2 _20688_ (.A(_03288_),
    .X(_03289_));
 sg13g2_a22oi_1 _20689_ (.Y(_00748_),
    .B1(_03284_),
    .B2(_03289_),
    .A2(net88),
    .A1(_03267_));
 sg13g2_inv_1 _20690_ (.Y(_03290_),
    .A(\cpu.dec.imm[11] ));
 sg13g2_nor2_1 _20691_ (.A(net145),
    .B(net155),
    .Y(_03291_));
 sg13g2_buf_1 _20692_ (.A(_03291_),
    .X(_03292_));
 sg13g2_nor2_1 _20693_ (.A(_09821_),
    .B(net251),
    .Y(_03293_));
 sg13g2_buf_2 _20694_ (.A(_03293_),
    .X(_03294_));
 sg13g2_nand2_1 _20695_ (.Y(_03295_),
    .A(_08948_),
    .B(_03294_));
 sg13g2_buf_1 _20696_ (.A(_03295_),
    .X(_03296_));
 sg13g2_o21ai_1 _20697_ (.B1(_03274_),
    .Y(_03297_),
    .A1(_08885_),
    .A2(net108));
 sg13g2_o21ai_1 _20698_ (.B1(net218),
    .Y(_03298_),
    .A1(net354),
    .A2(_03294_));
 sg13g2_o21ai_1 _20699_ (.B1(net196),
    .Y(_03299_),
    .A1(_09823_),
    .A2(net354));
 sg13g2_nand2_1 _20700_ (.Y(_03300_),
    .A(_03298_),
    .B(_03299_));
 sg13g2_inv_1 _20701_ (.Y(_03301_),
    .A(net342));
 sg13g2_inv_1 _20702_ (.Y(_03302_),
    .A(net355));
 sg13g2_buf_1 _20703_ (.A(_03205_),
    .X(_03303_));
 sg13g2_or3_1 _20704_ (.A(_03302_),
    .B(_03188_),
    .C(net293),
    .X(_03304_));
 sg13g2_nor2_1 _20705_ (.A(_03301_),
    .B(_03304_),
    .Y(_03305_));
 sg13g2_buf_1 _20706_ (.A(_03305_),
    .X(_03306_));
 sg13g2_inv_1 _20707_ (.Y(_03307_),
    .A(_03229_));
 sg13g2_a21oi_1 _20708_ (.A1(_03307_),
    .A2(_03305_),
    .Y(_03308_),
    .B1(_03295_));
 sg13g2_buf_1 _20709_ (.A(_03308_),
    .X(_03309_));
 sg13g2_o21ai_1 _20710_ (.B1(_03309_),
    .Y(_03310_),
    .A1(net304),
    .A2(net194));
 sg13g2_a21oi_1 _20711_ (.A1(_03300_),
    .A2(_03310_),
    .Y(_03311_),
    .B1(_03280_));
 sg13g2_a21oi_1 _20712_ (.A1(_03292_),
    .A2(_03297_),
    .Y(_03312_),
    .B1(_03311_));
 sg13g2_a22oi_1 _20713_ (.Y(_00749_),
    .B1(_03289_),
    .B2(_03312_),
    .A2(net88),
    .A1(_03290_));
 sg13g2_o21ai_1 _20714_ (.B1(_03274_),
    .Y(_03313_),
    .A1(_08908_),
    .A2(net108));
 sg13g2_o21ai_1 _20715_ (.B1(_03309_),
    .Y(_03314_),
    .A1(net357),
    .A2(net194));
 sg13g2_a21oi_1 _20716_ (.A1(_03300_),
    .A2(_03314_),
    .Y(_03315_),
    .B1(_03280_));
 sg13g2_a21oi_1 _20717_ (.A1(_03292_),
    .A2(_03313_),
    .Y(_03316_),
    .B1(_03315_));
 sg13g2_a22oi_1 _20718_ (.Y(_00750_),
    .B1(_03289_),
    .B2(_03316_),
    .A2(net88),
    .A1(_11291_));
 sg13g2_a21oi_1 _20719_ (.A1(net144),
    .A2(net108),
    .Y(_03317_),
    .B1(net354));
 sg13g2_o21ai_1 _20720_ (.B1(_03309_),
    .Y(_03318_),
    .A1(net294),
    .A2(_03306_));
 sg13g2_a21oi_1 _20721_ (.A1(_03300_),
    .A2(_03318_),
    .Y(_03319_),
    .B1(_03280_));
 sg13g2_a21oi_1 _20722_ (.A1(_03292_),
    .A2(_03317_),
    .Y(_03320_),
    .B1(_03319_));
 sg13g2_a22oi_1 _20723_ (.Y(_00751_),
    .B1(_03289_),
    .B2(_03320_),
    .A2(net88),
    .A1(_11298_));
 sg13g2_inv_1 _20724_ (.Y(_03321_),
    .A(\cpu.dec.imm[14] ));
 sg13g2_o21ai_1 _20725_ (.B1(_03274_),
    .Y(_03322_),
    .A1(net356),
    .A2(net108));
 sg13g2_nand2_1 _20726_ (.Y(_03323_),
    .A(_03292_),
    .B(_03322_));
 sg13g2_o21ai_1 _20727_ (.B1(_03309_),
    .Y(_03324_),
    .A1(_09083_),
    .A2(_03306_));
 sg13g2_a21oi_1 _20728_ (.A1(_03300_),
    .A2(_03324_),
    .Y(_03325_),
    .B1(_03280_));
 sg13g2_nor3_1 _20729_ (.A(net146),
    .B(_03287_),
    .C(_03325_),
    .Y(_03326_));
 sg13g2_a22oi_1 _20730_ (.Y(_00752_),
    .B1(_03323_),
    .B2(_03326_),
    .A2(_03268_),
    .A1(_03321_));
 sg13g2_o21ai_1 _20731_ (.B1(_03274_),
    .Y(_03327_),
    .A1(_09083_),
    .A2(_03296_));
 sg13g2_nand2_1 _20732_ (.Y(_03328_),
    .A(_03292_),
    .B(_03327_));
 sg13g2_a22oi_1 _20733_ (.Y(_00753_),
    .B1(_03326_),
    .B2(_03328_),
    .A2(_03268_),
    .A1(_11335_));
 sg13g2_nor2_1 _20734_ (.A(net263),
    .B(net236),
    .Y(_03329_));
 sg13g2_xnor2_1 _20735_ (.Y(_03330_),
    .A(net250),
    .B(_03329_));
 sg13g2_inv_1 _20736_ (.Y(_03331_),
    .A(_03305_));
 sg13g2_nor3_1 _20737_ (.A(net251),
    .B(net210),
    .C(_03331_),
    .Y(_03332_));
 sg13g2_o21ai_1 _20738_ (.B1(net197),
    .Y(_03333_),
    .A1(_03330_),
    .A2(_03332_));
 sg13g2_nand3_1 _20739_ (.B(net143),
    .C(_03333_),
    .A(net156),
    .Y(_03334_));
 sg13g2_nand2_1 _20740_ (.Y(_03335_),
    .A(net222),
    .B(net210));
 sg13g2_nor2_1 _20741_ (.A(net196),
    .B(_03335_),
    .Y(_03336_));
 sg13g2_a21oi_1 _20742_ (.A1(net195),
    .A2(net209),
    .Y(_03337_),
    .B1(_03336_));
 sg13g2_o21ai_1 _20743_ (.B1(net144),
    .Y(_03338_),
    .A1(net198),
    .A2(_03337_));
 sg13g2_a22oi_1 _20744_ (.Y(_03339_),
    .B1(net726),
    .B2(\cpu.icache.r_data[4][3] ),
    .A2(_08519_),
    .A1(\cpu.icache.r_data[2][3] ));
 sg13g2_a22oi_1 _20745_ (.Y(_03340_),
    .B1(_08529_),
    .B2(\cpu.icache.r_data[3][3] ),
    .A2(_08514_),
    .A1(\cpu.icache.r_data[1][3] ));
 sg13g2_mux2_1 _20746_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(\cpu.icache.r_data[7][3] ),
    .S(net944),
    .X(_03341_));
 sg13g2_a22oi_1 _20747_ (.Y(_03342_),
    .B1(_03341_),
    .B2(_08471_),
    .A2(_08891_),
    .A1(\cpu.icache.r_data[6][3] ));
 sg13g2_or2_1 _20748_ (.X(_03343_),
    .B(_03342_),
    .A(_08570_));
 sg13g2_and4_1 _20749_ (.A(_08512_),
    .B(_03339_),
    .C(_03340_),
    .D(_03343_),
    .X(_03344_));
 sg13g2_a21oi_1 _20750_ (.A1(_00172_),
    .A2(_08736_),
    .Y(_03345_),
    .B1(_03344_));
 sg13g2_nor2_1 _20751_ (.A(_00173_),
    .B(_08461_),
    .Y(_03346_));
 sg13g2_mux2_1 _20752_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_08569_),
    .X(_03347_));
 sg13g2_a22oi_1 _20753_ (.Y(_03348_),
    .B1(_03347_),
    .B2(_08471_),
    .A2(net940),
    .A1(\cpu.icache.r_data[6][19] ));
 sg13g2_nand2b_1 _20754_ (.Y(_03349_),
    .B(net723),
    .A_N(_03348_));
 sg13g2_a22oi_1 _20755_ (.Y(_03350_),
    .B1(_08594_),
    .B2(\cpu.icache.r_data[4][19] ),
    .A2(_08479_),
    .A1(\cpu.icache.r_data[1][19] ));
 sg13g2_a22oi_1 _20756_ (.Y(_03351_),
    .B1(_08533_),
    .B2(\cpu.icache.r_data[5][19] ),
    .A2(_08488_),
    .A1(\cpu.icache.r_data[2][19] ));
 sg13g2_nand3_1 _20757_ (.B(_03350_),
    .C(_03351_),
    .A(_03349_),
    .Y(_03352_));
 sg13g2_or3_1 _20758_ (.A(_08958_),
    .B(_03346_),
    .C(_03352_),
    .X(_03353_));
 sg13g2_o21ai_1 _20759_ (.B1(_03353_),
    .Y(_03354_),
    .A1(net935),
    .A2(_03345_));
 sg13g2_buf_1 _20760_ (.A(_03354_),
    .X(_03355_));
 sg13g2_buf_1 _20761_ (.A(_03355_),
    .X(_03356_));
 sg13g2_nor2_1 _20762_ (.A(net186),
    .B(net249),
    .Y(_03357_));
 sg13g2_a221oi_1 _20763_ (.B2(_03357_),
    .C1(net146),
    .B1(_03338_),
    .A1(net357),
    .Y(_03358_),
    .A2(_03334_));
 sg13g2_a21oi_1 _20764_ (.A1(_10590_),
    .A2(net146),
    .Y(_00754_),
    .B1(_03358_));
 sg13g2_a21oi_1 _20765_ (.A1(_03122_),
    .A2(_03108_),
    .Y(_03359_),
    .B1(net236));
 sg13g2_inv_1 _20766_ (.Y(_03360_),
    .A(_03329_));
 sg13g2_nor2_1 _20767_ (.A(_03112_),
    .B(_03360_),
    .Y(_03361_));
 sg13g2_inv_1 _20768_ (.Y(_03362_),
    .A(_03361_));
 sg13g2_o21ai_1 _20769_ (.B1(_03362_),
    .Y(_03363_),
    .A1(_03137_),
    .A2(_03359_));
 sg13g2_a21oi_1 _20770_ (.A1(net197),
    .A2(_03363_),
    .Y(_03364_),
    .B1(net89));
 sg13g2_nand2b_1 _20771_ (.Y(_03365_),
    .B(_03152_),
    .A_N(_03119_));
 sg13g2_nand2_1 _20772_ (.Y(_03366_),
    .A(net221),
    .B(net154));
 sg13g2_nand4_1 _20773_ (.B(net158),
    .C(_03294_),
    .A(net218),
    .Y(_03367_),
    .D(net194));
 sg13g2_nand2_1 _20774_ (.Y(_03368_),
    .A(_03366_),
    .B(_03367_));
 sg13g2_nand2_2 _20775_ (.Y(_03369_),
    .A(_08991_),
    .B(net210));
 sg13g2_nor2_1 _20776_ (.A(_03369_),
    .B(_03285_),
    .Y(_03370_));
 sg13g2_a22oi_1 _20777_ (.Y(_03371_),
    .B1(_03370_),
    .B2(net219),
    .A2(net174),
    .A1(_08971_));
 sg13g2_nor2_1 _20778_ (.A(net249),
    .B(_03371_),
    .Y(_03372_));
 sg13g2_a221oi_1 _20779_ (.B2(net304),
    .C1(_03372_),
    .B1(_03368_),
    .A1(_03230_),
    .Y(_03373_),
    .A2(_03365_));
 sg13g2_o21ai_1 _20780_ (.B1(_03373_),
    .Y(_03374_),
    .A1(net355),
    .A2(_03364_));
 sg13g2_mux2_1 _20781_ (.A0(_03374_),
    .A1(_10551_),
    .S(_09094_),
    .X(_00755_));
 sg13g2_inv_1 _20782_ (.Y(_03375_),
    .A(_11221_));
 sg13g2_nand2_1 _20783_ (.Y(_03376_),
    .A(net158),
    .B(_09836_));
 sg13g2_nand2_1 _20784_ (.Y(_03377_),
    .A(net187),
    .B(net217));
 sg13g2_nand2_1 _20785_ (.Y(_03378_),
    .A(_03302_),
    .B(_03117_));
 sg13g2_a22oi_1 _20786_ (.Y(_03379_),
    .B1(_03377_),
    .B2(_03378_),
    .A2(_03271_),
    .A1(_03376_));
 sg13g2_nor2_1 _20787_ (.A(net145),
    .B(_09836_),
    .Y(_03380_));
 sg13g2_a22oi_1 _20788_ (.Y(_03381_),
    .B1(_03380_),
    .B2(net304),
    .A2(_03370_),
    .A1(net217));
 sg13g2_nand3_1 _20789_ (.B(net195),
    .C(net158),
    .A(net304),
    .Y(_03382_));
 sg13g2_a21oi_1 _20790_ (.A1(_03381_),
    .A2(_03382_),
    .Y(_03383_),
    .B1(net198));
 sg13g2_a22oi_1 _20791_ (.Y(_03384_),
    .B1(_03330_),
    .B2(net197),
    .A2(_03360_),
    .A1(net186));
 sg13g2_a21oi_1 _20792_ (.A1(_03367_),
    .A2(_03384_),
    .Y(_03385_),
    .B1(net356));
 sg13g2_nor4_1 _20793_ (.A(net146),
    .B(_03379_),
    .C(_03383_),
    .D(_03385_),
    .Y(_03386_));
 sg13g2_a21oi_1 _20794_ (.A1(_03375_),
    .A2(net146),
    .Y(_00756_),
    .B1(_03386_));
 sg13g2_nor2_1 _20795_ (.A(_03127_),
    .B(_03122_),
    .Y(_03387_));
 sg13g2_a21oi_1 _20796_ (.A1(net197),
    .A2(net209),
    .Y(_03388_),
    .B1(_03387_));
 sg13g2_o21ai_1 _20797_ (.B1(net143),
    .Y(_03389_),
    .A1(net195),
    .A2(_03388_));
 sg13g2_nand2_1 _20798_ (.Y(_03390_),
    .A(_03135_),
    .B(_09010_));
 sg13g2_or4_1 _20799_ (.A(net196),
    .B(_09073_),
    .C(_03331_),
    .D(_03390_),
    .X(_03391_));
 sg13g2_o21ai_1 _20800_ (.B1(_03391_),
    .Y(_03392_),
    .A1(net197),
    .A2(net356));
 sg13g2_o21ai_1 _20801_ (.B1(net219),
    .Y(_03393_),
    .A1(net356),
    .A2(_03390_));
 sg13g2_o21ai_1 _20802_ (.B1(_03393_),
    .Y(_03394_),
    .A1(net219),
    .A2(_03392_));
 sg13g2_a21oi_1 _20803_ (.A1(_03376_),
    .A2(_03271_),
    .Y(_03395_),
    .B1(_03394_));
 sg13g2_a21oi_1 _20804_ (.A1(net294),
    .A2(_03389_),
    .Y(_03396_),
    .B1(_03395_));
 sg13g2_buf_1 _20805_ (.A(_08859_),
    .X(_03397_));
 sg13g2_nand2_1 _20806_ (.Y(_03398_),
    .A(\cpu.dec.imm[4] ),
    .B(net107));
 sg13g2_o21ai_1 _20807_ (.B1(_03398_),
    .Y(_00757_),
    .A1(net93),
    .A2(_03396_));
 sg13g2_nor2_1 _20808_ (.A(net108),
    .B(net194),
    .Y(_03399_));
 sg13g2_nand3_1 _20809_ (.B(net174),
    .C(_03147_),
    .A(net156),
    .Y(_03400_));
 sg13g2_nand2_1 _20810_ (.Y(_03401_),
    .A(net210),
    .B(_03400_));
 sg13g2_o21ai_1 _20811_ (.B1(_03401_),
    .Y(_03402_),
    .A1(_03269_),
    .A2(_03399_));
 sg13g2_nor2_2 _20812_ (.A(net220),
    .B(_08948_),
    .Y(_03403_));
 sg13g2_a22oi_1 _20813_ (.Y(_03404_),
    .B1(net216),
    .B2(_03403_),
    .A2(_03136_),
    .A1(_08884_));
 sg13g2_nor2_1 _20814_ (.A(_03123_),
    .B(_03404_),
    .Y(_03405_));
 sg13g2_nor3_1 _20815_ (.A(_08885_),
    .B(net195),
    .C(_03387_),
    .Y(_03406_));
 sg13g2_or2_1 _20816_ (.X(_03407_),
    .B(_03406_),
    .A(_03405_));
 sg13g2_a22oi_1 _20817_ (.Y(_03408_),
    .B1(_03407_),
    .B2(net89),
    .A2(_03402_),
    .A1(net216));
 sg13g2_nand2_1 _20818_ (.Y(_03409_),
    .A(\cpu.dec.imm[5] ),
    .B(net107));
 sg13g2_o21ai_1 _20819_ (.B1(_03409_),
    .Y(_00758_),
    .A1(_09095_),
    .A2(_03408_));
 sg13g2_inv_1 _20820_ (.Y(_03410_),
    .A(_03355_));
 sg13g2_nand2_1 _20821_ (.Y(_03411_),
    .A(net251),
    .B(net293));
 sg13g2_nor2_1 _20822_ (.A(net187),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_a21oi_1 _20823_ (.A1(net187),
    .A2(_03410_),
    .Y(_03413_),
    .B1(_03412_));
 sg13g2_nand2_1 _20824_ (.Y(_03414_),
    .A(net250),
    .B(net154));
 sg13g2_o21ai_1 _20825_ (.B1(_03414_),
    .Y(_03415_),
    .A1(net250),
    .A2(_03269_));
 sg13g2_nand2_1 _20826_ (.Y(_03416_),
    .A(net197),
    .B(_03415_));
 sg13g2_a21oi_1 _20827_ (.A1(_03366_),
    .A2(_03416_),
    .Y(_03417_),
    .B1(net249));
 sg13g2_nor2_1 _20828_ (.A(net108),
    .B(net249),
    .Y(_03418_));
 sg13g2_a22oi_1 _20829_ (.Y(_03419_),
    .B1(net194),
    .B2(_03418_),
    .A2(net293),
    .A1(net173));
 sg13g2_nand3_1 _20830_ (.B(net174),
    .C(_03117_),
    .A(_08884_),
    .Y(_03420_));
 sg13g2_o21ai_1 _20831_ (.B1(_03420_),
    .Y(_03421_),
    .A1(_03376_),
    .A2(_03419_));
 sg13g2_nor3_1 _20832_ (.A(net89),
    .B(_03417_),
    .C(_03421_),
    .Y(_03422_));
 sg13g2_a21oi_1 _20833_ (.A1(net89),
    .A2(_03413_),
    .Y(_03423_),
    .B1(_03422_));
 sg13g2_mux2_1 _20834_ (.A0(_03423_),
    .A1(\cpu.dec.imm[6] ),
    .S(net94),
    .X(_00759_));
 sg13g2_inv_1 _20835_ (.Y(_03424_),
    .A(\cpu.dec.imm[7] ));
 sg13g2_nand2_1 _20836_ (.Y(_03425_),
    .A(net251),
    .B(_03110_));
 sg13g2_nor2_1 _20837_ (.A(net187),
    .B(_03425_),
    .Y(_03426_));
 sg13g2_a22oi_1 _20838_ (.Y(_03427_),
    .B1(net342),
    .B2(_03426_),
    .A2(_03119_),
    .A1(net357));
 sg13g2_a21oi_1 _20839_ (.A1(_03123_),
    .A2(net194),
    .Y(_03428_),
    .B1(_03112_));
 sg13g2_nor2_1 _20840_ (.A(_03129_),
    .B(_03428_),
    .Y(_03429_));
 sg13g2_nor2_1 _20841_ (.A(net195),
    .B(_03366_),
    .Y(_03430_));
 sg13g2_o21ai_1 _20842_ (.B1(net217),
    .Y(_03431_),
    .A1(_03429_),
    .A2(_03430_));
 sg13g2_and2_1 _20843_ (.A(_03427_),
    .B(_03431_),
    .X(_03432_));
 sg13g2_a22oi_1 _20844_ (.Y(_00760_),
    .B1(_03289_),
    .B2(_03432_),
    .A2(net88),
    .A1(_03424_));
 sg13g2_inv_1 _20845_ (.Y(_03433_),
    .A(\cpu.dec.imm[8] ));
 sg13g2_inv_1 _20846_ (.Y(_03434_),
    .A(_03253_));
 sg13g2_o21ai_1 _20847_ (.B1(_03274_),
    .Y(_03435_),
    .A1(_03434_),
    .A2(net108));
 sg13g2_o21ai_1 _20848_ (.B1(_03309_),
    .Y(_03436_),
    .A1(net216),
    .A2(net194));
 sg13g2_a21oi_1 _20849_ (.A1(net173),
    .A2(_03188_),
    .Y(_03437_),
    .B1(_03281_));
 sg13g2_a21oi_1 _20850_ (.A1(_03436_),
    .A2(_03437_),
    .Y(_03438_),
    .B1(_03280_));
 sg13g2_a221oi_1 _20851_ (.B2(_03292_),
    .C1(_03438_),
    .B1(_03435_),
    .A1(_03188_),
    .Y(_03439_),
    .A2(_03426_));
 sg13g2_a22oi_1 _20852_ (.Y(_00761_),
    .B1(_03289_),
    .B2(_03439_),
    .A2(net88),
    .A1(_03433_));
 sg13g2_inv_1 _20853_ (.Y(_03440_),
    .A(\cpu.dec.imm[9] ));
 sg13g2_o21ai_1 _20854_ (.B1(_03274_),
    .Y(_03441_),
    .A1(_03296_),
    .A2(net249));
 sg13g2_o21ai_1 _20855_ (.B1(_03309_),
    .Y(_03442_),
    .A1(net194),
    .A2(_03410_));
 sg13g2_a21oi_1 _20856_ (.A1(_03302_),
    .A2(net173),
    .Y(_03443_),
    .B1(_03281_));
 sg13g2_a21oi_1 _20857_ (.A1(_03442_),
    .A2(_03443_),
    .Y(_03444_),
    .B1(_03280_));
 sg13g2_a21oi_1 _20858_ (.A1(_03292_),
    .A2(_03441_),
    .Y(_03445_),
    .B1(_03444_));
 sg13g2_a22oi_1 _20859_ (.Y(_00762_),
    .B1(_03289_),
    .B2(_03445_),
    .A2(net88),
    .A1(_03440_));
 sg13g2_nor4_1 _20860_ (.A(_08560_),
    .B(_08908_),
    .C(_03152_),
    .D(_03210_),
    .Y(_03446_));
 sg13g2_buf_1 _20861_ (.A(\cpu.dec.do_inv_mmu ),
    .X(_03447_));
 sg13g2_mux2_1 _20862_ (.A0(_03446_),
    .A1(_03447_),
    .S(net94),
    .X(_00763_));
 sg13g2_xnor2_1 _20863_ (.Y(_03448_),
    .A(_08948_),
    .B(net263));
 sg13g2_nor3_1 _20864_ (.A(_03132_),
    .B(_03145_),
    .C(_03448_),
    .Y(_03449_));
 sg13g2_mux2_1 _20865_ (.A0(_03449_),
    .A1(\cpu.dec.io ),
    .S(net94),
    .X(_00764_));
 sg13g2_nor2_1 _20866_ (.A(_08884_),
    .B(_08907_),
    .Y(_03450_));
 sg13g2_nand4_1 _20867_ (.B(_03307_),
    .C(_03434_),
    .A(_03450_),
    .Y(_03451_),
    .D(_03356_));
 sg13g2_nor3_2 _20868_ (.A(net156),
    .B(_03369_),
    .C(_03451_),
    .Y(_03452_));
 sg13g2_mux2_1 _20869_ (.A0(_03452_),
    .A1(\cpu.dec.jmp ),
    .S(_09094_),
    .X(_00765_));
 sg13g2_a21oi_1 _20870_ (.A1(net143),
    .A2(_03335_),
    .Y(_03453_),
    .B1(_03275_));
 sg13g2_mux2_1 _20871_ (.A0(_03453_),
    .A1(_11616_),
    .S(net94),
    .X(_00766_));
 sg13g2_nor3_1 _20872_ (.A(_09056_),
    .B(net294),
    .C(_09080_),
    .Y(_03454_));
 sg13g2_a21o_1 _20873_ (.A2(net92),
    .A1(_09278_),
    .B1(_03454_),
    .X(_00767_));
 sg13g2_o21ai_1 _20874_ (.B1(_09097_),
    .Y(_03455_),
    .A1(_09083_),
    .A2(net294));
 sg13g2_nand3_1 _20875_ (.B(_09826_),
    .C(net354),
    .A(_03128_),
    .Y(_03456_));
 sg13g2_nand3_1 _20876_ (.B(net174),
    .C(_09052_),
    .A(_03132_),
    .Y(_03457_));
 sg13g2_nand4_1 _20877_ (.B(_09009_),
    .C(_03456_),
    .A(_09823_),
    .Y(_03458_),
    .D(_03457_));
 sg13g2_o21ai_1 _20878_ (.B1(_03458_),
    .Y(_03459_),
    .A1(_09013_),
    .A2(_03455_));
 sg13g2_nor2_1 _20879_ (.A(net107),
    .B(_03459_),
    .Y(_03460_));
 sg13g2_a21oi_1 _20880_ (.A1(_10228_),
    .A2(net88),
    .Y(_00768_),
    .B1(_03460_));
 sg13g2_nor2_1 _20881_ (.A(_03117_),
    .B(net173),
    .Y(_03461_));
 sg13g2_o21ai_1 _20882_ (.B1(_03461_),
    .Y(_03462_),
    .A1(net196),
    .A2(net216));
 sg13g2_o21ai_1 _20883_ (.B1(_03108_),
    .Y(_03463_),
    .A1(_03136_),
    .A2(_03411_));
 sg13g2_o21ai_1 _20884_ (.B1(_03128_),
    .Y(_03464_),
    .A1(net173),
    .A2(net293));
 sg13g2_nand2b_1 _20885_ (.Y(_03465_),
    .B(_03464_),
    .A_N(_03463_));
 sg13g2_inv_1 _20886_ (.Y(_03466_),
    .A(_03411_));
 sg13g2_nand2_1 _20887_ (.Y(_03467_),
    .A(net250),
    .B(_03303_));
 sg13g2_o21ai_1 _20888_ (.B1(_03467_),
    .Y(_03468_),
    .A1(net250),
    .A2(_03434_));
 sg13g2_a22oi_1 _20889_ (.Y(_03469_),
    .B1(_03468_),
    .B2(_03294_),
    .A2(_03466_),
    .A1(_03403_));
 sg13g2_nor2_1 _20890_ (.A(net145),
    .B(_03469_),
    .Y(_03470_));
 sg13g2_a221oi_1 _20891_ (.B2(net209),
    .C1(_03470_),
    .B1(_03465_),
    .A1(_03125_),
    .Y(_03471_),
    .A2(_03452_));
 sg13g2_a21oi_1 _20892_ (.A1(_09823_),
    .A2(_03451_),
    .Y(_03472_),
    .B1(net220));
 sg13g2_nor2_1 _20893_ (.A(_03369_),
    .B(_03472_),
    .Y(_03473_));
 sg13g2_nand2_1 _20894_ (.Y(_03474_),
    .A(net293),
    .B(_03473_));
 sg13g2_a221oi_1 _20895_ (.B2(_03474_),
    .C1(net113),
    .B1(_03471_),
    .A1(_03111_),
    .Y(_03475_),
    .A2(_03462_));
 sg13g2_a21o_1 _20896_ (.A2(net92),
    .A1(\cpu.dec.r_rd[0] ),
    .B1(_03475_),
    .X(_00769_));
 sg13g2_a21oi_1 _20897_ (.A1(net158),
    .A2(_03461_),
    .Y(_03476_),
    .B1(_03473_));
 sg13g2_nand2b_1 _20898_ (.Y(_03477_),
    .B(_03110_),
    .A_N(_03114_));
 sg13g2_nor2_1 _20899_ (.A(net196),
    .B(_03477_),
    .Y(_03478_));
 sg13g2_nand2_1 _20900_ (.Y(_03479_),
    .A(net221),
    .B(_03356_));
 sg13g2_a22oi_1 _20901_ (.Y(_03480_),
    .B1(_03479_),
    .B2(net220),
    .A2(net342),
    .A1(net251));
 sg13g2_nand3_1 _20902_ (.B(net342),
    .C(_03294_),
    .A(net218),
    .Y(_03481_));
 sg13g2_o21ai_1 _20903_ (.B1(_03481_),
    .Y(_03482_),
    .A1(net218),
    .A2(_03480_));
 sg13g2_and2_1 _20904_ (.A(_09077_),
    .B(_03482_),
    .X(_03483_));
 sg13g2_nand3_1 _20905_ (.B(_03209_),
    .C(_03229_),
    .A(_03450_),
    .Y(_03484_));
 sg13g2_nor3_1 _20906_ (.A(_03253_),
    .B(net249),
    .C(_03484_),
    .Y(_03485_));
 sg13g2_nand2b_1 _20907_ (.Y(_03486_),
    .B(net155),
    .A_N(_03485_));
 sg13g2_a22oi_1 _20908_ (.Y(_03487_),
    .B1(_03483_),
    .B2(_03486_),
    .A2(_03478_),
    .A1(_03410_));
 sg13g2_o21ai_1 _20909_ (.B1(_03487_),
    .Y(_03488_),
    .A1(_03301_),
    .A2(_03476_));
 sg13g2_mux2_1 _20910_ (.A0(_03488_),
    .A1(\cpu.dec.r_rd[1] ),
    .S(net94),
    .X(_00770_));
 sg13g2_inv_2 _20911_ (.Y(_03489_),
    .A(_03188_));
 sg13g2_nand2_1 _20912_ (.Y(_03490_),
    .A(_03135_),
    .B(_03188_));
 sg13g2_o21ai_1 _20913_ (.B1(_03490_),
    .Y(_03491_),
    .A1(net218),
    .A2(_03307_));
 sg13g2_nor2_1 _20914_ (.A(net221),
    .B(_03489_),
    .Y(_03492_));
 sg13g2_a22oi_1 _20915_ (.Y(_03493_),
    .B1(_03492_),
    .B2(_03403_),
    .A2(_03491_),
    .A1(_03294_));
 sg13g2_inv_1 _20916_ (.Y(_03494_),
    .A(_03493_));
 sg13g2_a22oi_1 _20917_ (.Y(_03495_),
    .B1(_03494_),
    .B2(_09077_),
    .A2(_03478_),
    .A1(_03230_));
 sg13g2_o21ai_1 _20918_ (.B1(_03495_),
    .Y(_03496_),
    .A1(_03489_),
    .A2(_03476_));
 sg13g2_mux2_1 _20919_ (.A0(_03496_),
    .A1(\cpu.dec.r_rd[2] ),
    .S(net112),
    .X(_00771_));
 sg13g2_nor4_2 _20920_ (.A(_08909_),
    .B(_03229_),
    .C(_03253_),
    .Y(_03497_),
    .D(_03410_));
 sg13g2_nor3_1 _20921_ (.A(_09075_),
    .B(_09050_),
    .C(_03497_),
    .Y(_03498_));
 sg13g2_o21ai_1 _20922_ (.B1(net219),
    .Y(_03499_),
    .A1(net143),
    .A2(_03498_));
 sg13g2_o21ai_1 _20923_ (.B1(net198),
    .Y(_03500_),
    .A1(net186),
    .A2(_03302_));
 sg13g2_a22oi_1 _20924_ (.Y(_03501_),
    .B1(_03258_),
    .B2(net355),
    .A2(_03133_),
    .A1(_03131_));
 sg13g2_nor2_1 _20925_ (.A(net209),
    .B(_03501_),
    .Y(_03502_));
 sg13g2_a221oi_1 _20926_ (.B2(_03137_),
    .C1(_03502_),
    .B1(_03500_),
    .A1(net196),
    .Y(_03503_),
    .A2(_03499_));
 sg13g2_mux2_1 _20927_ (.A0(_03503_),
    .A1(\cpu.dec.r_rd[3] ),
    .S(net112),
    .X(_00772_));
 sg13g2_nand2b_1 _20928_ (.Y(_03504_),
    .B(_03146_),
    .A_N(_09823_));
 sg13g2_o21ai_1 _20929_ (.B1(_08971_),
    .Y(_03505_),
    .A1(_03124_),
    .A2(_03497_));
 sg13g2_buf_1 _20930_ (.A(_03505_),
    .X(_03506_));
 sg13g2_o21ai_1 _20931_ (.B1(_03506_),
    .Y(_03507_),
    .A1(net221),
    .A2(_03403_));
 sg13g2_a22oi_1 _20932_ (.Y(_03508_),
    .B1(_03507_),
    .B2(net154),
    .A2(_03504_),
    .A1(net158));
 sg13g2_o21ai_1 _20933_ (.B1(_03508_),
    .Y(_03509_),
    .A1(_03271_),
    .A2(_03276_));
 sg13g2_a21oi_1 _20934_ (.A1(net293),
    .A2(_03509_),
    .Y(_03510_),
    .B1(net89));
 sg13g2_a21oi_1 _20935_ (.A1(_03425_),
    .A2(net293),
    .Y(_03511_),
    .B1(net187));
 sg13g2_nor3_1 _20936_ (.A(net146),
    .B(_03510_),
    .C(_03511_),
    .Y(_03512_));
 sg13g2_a21o_1 _20937_ (.A2(net92),
    .A1(_10733_),
    .B1(_03512_),
    .X(_00773_));
 sg13g2_a21oi_1 _20938_ (.A1(net187),
    .A2(_03506_),
    .Y(_03513_),
    .B1(_03301_));
 sg13g2_o21ai_1 _20939_ (.B1(net154),
    .Y(_03514_),
    .A1(net198),
    .A2(_03513_));
 sg13g2_o21ai_1 _20940_ (.B1(net220),
    .Y(_03515_),
    .A1(net222),
    .A2(_03304_));
 sg13g2_a21oi_1 _20941_ (.A1(net221),
    .A2(_03515_),
    .Y(_03516_),
    .B1(_09823_));
 sg13g2_o21ai_1 _20942_ (.B1(net143),
    .Y(_03517_),
    .A1(_03301_),
    .A2(_03516_));
 sg13g2_nor2_1 _20943_ (.A(net155),
    .B(_03170_),
    .Y(_03518_));
 sg13g2_nor3_1 _20944_ (.A(net145),
    .B(_03276_),
    .C(_03518_),
    .Y(_03519_));
 sg13g2_a21oi_1 _20945_ (.A1(net209),
    .A2(_03517_),
    .Y(_03520_),
    .B1(_03519_));
 sg13g2_o21ai_1 _20946_ (.B1(net156),
    .Y(_03521_),
    .A1(net219),
    .A2(_03170_));
 sg13g2_a221oi_1 _20947_ (.B2(_03111_),
    .C1(net113),
    .B1(_03521_),
    .A1(_03514_),
    .Y(_03522_),
    .A2(_03520_));
 sg13g2_a21o_1 _20948_ (.A2(net92),
    .A1(_10756_),
    .B1(_03522_),
    .X(_00774_));
 sg13g2_o21ai_1 _20949_ (.B1(_09077_),
    .Y(_03523_),
    .A1(net155),
    .A2(_03188_));
 sg13g2_o21ai_1 _20950_ (.B1(_03523_),
    .Y(_03524_),
    .A1(_03489_),
    .A2(_03508_));
 sg13g2_nor2_1 _20951_ (.A(net219),
    .B(_03489_),
    .Y(_03525_));
 sg13g2_a22oi_1 _20952_ (.Y(_03526_),
    .B1(_03525_),
    .B2(net89),
    .A2(_03524_),
    .A1(net108));
 sg13g2_nand2_1 _20953_ (.Y(_03527_),
    .A(_10744_),
    .B(net107));
 sg13g2_o21ai_1 _20954_ (.B1(_03527_),
    .Y(_00775_),
    .A1(net93),
    .A2(_03526_));
 sg13g2_or2_1 _20955_ (.X(_03528_),
    .B(_03506_),
    .A(net355));
 sg13g2_a21oi_1 _20956_ (.A1(_03403_),
    .A2(_03528_),
    .Y(_03529_),
    .B1(net236));
 sg13g2_nand2_1 _20957_ (.Y(_03530_),
    .A(net250),
    .B(_08991_));
 sg13g2_o21ai_1 _20958_ (.B1(_03530_),
    .Y(_03531_),
    .A1(net218),
    .A2(net145));
 sg13g2_a22oi_1 _20959_ (.Y(_03532_),
    .B1(_03531_),
    .B2(net197),
    .A2(net236),
    .A1(net195));
 sg13g2_o21ai_1 _20960_ (.B1(_03532_),
    .Y(_03533_),
    .A1(net143),
    .A2(_03529_));
 sg13g2_nor2_1 _20961_ (.A(net198),
    .B(_03533_),
    .Y(_03534_));
 sg13g2_a221oi_1 _20962_ (.B2(net154),
    .C1(_03131_),
    .B1(_03528_),
    .A1(_03133_),
    .Y(_03535_),
    .A2(_03335_));
 sg13g2_nor3_1 _20963_ (.A(_12042_),
    .B(_03534_),
    .C(_03535_),
    .Y(_03536_));
 sg13g2_a21oi_1 _20964_ (.A1(_10737_),
    .A2(net146),
    .Y(_00776_),
    .B1(_03536_));
 sg13g2_nand3_1 _20965_ (.B(_09051_),
    .C(net294),
    .A(net357),
    .Y(_03537_));
 sg13g2_a221oi_1 _20966_ (.B2(_08971_),
    .C1(_03145_),
    .B1(_03537_),
    .A1(_03127_),
    .Y(_03538_),
    .A2(net173));
 sg13g2_buf_1 _20967_ (.A(_03538_),
    .X(_03539_));
 sg13g2_nor2_2 _20968_ (.A(_03369_),
    .B(net144),
    .Y(_03540_));
 sg13g2_nand2b_1 _20969_ (.Y(_03541_),
    .B(_03540_),
    .A_N(net293));
 sg13g2_o21ai_1 _20970_ (.B1(_03541_),
    .Y(_03542_),
    .A1(net216),
    .A2(_03540_));
 sg13g2_nor3_1 _20971_ (.A(net113),
    .B(_03539_),
    .C(_03542_),
    .Y(_03543_));
 sg13g2_a21o_1 _20972_ (.A2(net92),
    .A1(_10383_),
    .B1(_03543_),
    .X(_00777_));
 sg13g2_nor3_1 _20973_ (.A(net249),
    .B(_03539_),
    .C(_03540_),
    .Y(_03544_));
 sg13g2_a21oi_1 _20974_ (.A1(net342),
    .A2(_03540_),
    .Y(_03545_),
    .B1(_03544_));
 sg13g2_nand2_1 _20975_ (.Y(_03546_),
    .A(_10250_),
    .B(net107));
 sg13g2_o21ai_1 _20976_ (.B1(_03546_),
    .Y(_00778_),
    .A1(net95),
    .A2(_03545_));
 sg13g2_o21ai_1 _20977_ (.B1(_03377_),
    .Y(_03547_),
    .A1(net144),
    .A2(_03489_));
 sg13g2_nor3_1 _20978_ (.A(_03307_),
    .B(_03539_),
    .C(_03540_),
    .Y(_03548_));
 sg13g2_a21oi_1 _20979_ (.A1(net154),
    .A2(_03547_),
    .Y(_03549_),
    .B1(_03548_));
 sg13g2_nand2_1 _20980_ (.Y(_03550_),
    .A(_10270_),
    .B(net107));
 sg13g2_o21ai_1 _20981_ (.B1(_03550_),
    .Y(_00779_),
    .A1(net95),
    .A2(_03549_));
 sg13g2_o21ai_1 _20982_ (.B1(net144),
    .Y(_03551_),
    .A1(net304),
    .A2(net156));
 sg13g2_and3_1 _20983_ (.X(_03552_),
    .A(net154),
    .B(_03378_),
    .C(_03551_));
 sg13g2_nor3_1 _20984_ (.A(net113),
    .B(_03539_),
    .C(_03552_),
    .Y(_03553_));
 sg13g2_a21o_1 _20985_ (.A2(net92),
    .A1(_10291_),
    .B1(_03553_),
    .X(_00780_));
 sg13g2_nor4_1 _20986_ (.A(_08860_),
    .B(net354),
    .C(_09079_),
    .D(_09090_),
    .Y(_03554_));
 sg13g2_a21o_1 _20987_ (.A2(_09820_),
    .A1(_10139_),
    .B1(_03554_),
    .X(_00781_));
 sg13g2_nor4_1 _20988_ (.A(net357),
    .B(_09013_),
    .C(_09052_),
    .D(net354),
    .Y(_03555_));
 sg13g2_mux2_1 _20989_ (.A0(_03555_),
    .A1(\cpu.dec.r_set_cc ),
    .S(net112),
    .X(_00782_));
 sg13g2_nor2_1 _20990_ (.A(net143),
    .B(_03147_),
    .Y(_03556_));
 sg13g2_a21oi_1 _20991_ (.A1(_03262_),
    .A2(_03361_),
    .Y(_03557_),
    .B1(_03556_));
 sg13g2_buf_1 _20992_ (.A(\cpu.dec.r_store ),
    .X(_03558_));
 sg13g2_nand2_1 _20993_ (.Y(_03559_),
    .A(_03558_),
    .B(_03397_));
 sg13g2_o21ai_1 _20994_ (.B1(_03559_),
    .Y(_00783_),
    .A1(net95),
    .A2(_03557_));
 sg13g2_nand2b_1 _20995_ (.Y(_03560_),
    .B(_03485_),
    .A_N(_03152_));
 sg13g2_nand2_1 _20996_ (.Y(_03561_),
    .A(\cpu.dec.r_swapsp ),
    .B(net107));
 sg13g2_o21ai_1 _20997_ (.B1(_03561_),
    .Y(_00784_),
    .A1(net95),
    .A2(_03560_));
 sg13g2_nand2_1 _20998_ (.Y(_03562_),
    .A(net216),
    .B(net249));
 sg13g2_nor4_1 _20999_ (.A(net114),
    .B(_03152_),
    .C(_03484_),
    .D(_03562_),
    .Y(_03563_));
 sg13g2_a21o_1 _21000_ (.A2(_09820_),
    .A1(\cpu.dec.r_sys_call ),
    .B1(_03563_),
    .X(_00785_));
 sg13g2_nand2_1 _21001_ (.Y(_03564_),
    .A(net342),
    .B(_03303_));
 sg13g2_xnor2_1 _21002_ (.Y(_03565_),
    .A(_03489_),
    .B(_03564_));
 sg13g2_nor3_1 _21003_ (.A(net1163),
    .B(_03302_),
    .C(_03565_),
    .Y(_03566_));
 sg13g2_a22oi_1 _21004_ (.Y(_03567_),
    .B1(_09097_),
    .B2(_08907_),
    .A2(net356),
    .A1(_08884_));
 sg13g2_nand3_1 _21005_ (.B(_09074_),
    .C(net216),
    .A(net356),
    .Y(_03568_));
 sg13g2_o21ai_1 _21006_ (.B1(_03568_),
    .Y(_03569_),
    .A1(_09074_),
    .A2(_03567_));
 sg13g2_a22oi_1 _21007_ (.Y(_03570_),
    .B1(_03569_),
    .B2(_09096_),
    .A2(_03566_),
    .A1(_03399_));
 sg13g2_buf_1 _21008_ (.A(_08301_),
    .X(_03571_));
 sg13g2_nor2_1 _21009_ (.A(net993),
    .B(_10402_),
    .Y(_03572_));
 sg13g2_o21ai_1 _21010_ (.B1(net220),
    .Y(_03573_),
    .A1(_03448_),
    .A2(_03572_));
 sg13g2_nor3_1 _21011_ (.A(net222),
    .B(_03116_),
    .C(_03566_),
    .Y(_03574_));
 sg13g2_nand3_1 _21012_ (.B(_03207_),
    .C(_03497_),
    .A(net993),
    .Y(_03575_));
 sg13g2_a22oi_1 _21013_ (.Y(_03576_),
    .B1(_03232_),
    .B2(_03575_),
    .A2(net356),
    .A1(_09823_));
 sg13g2_o21ai_1 _21014_ (.B1(_03576_),
    .Y(_03577_),
    .A1(_03573_),
    .A2(_03574_));
 sg13g2_nor2_1 _21015_ (.A(_08885_),
    .B(_03229_),
    .Y(_03578_));
 sg13g2_o21ai_1 _21016_ (.B1(_03209_),
    .Y(_03579_),
    .A1(net357),
    .A2(_03578_));
 sg13g2_nand2b_1 _21017_ (.Y(_03580_),
    .B(_03579_),
    .A_N(_03485_));
 sg13g2_nand3_1 _21018_ (.B(_09838_),
    .C(_03580_),
    .A(net993),
    .Y(_03581_));
 sg13g2_nand3_1 _21019_ (.B(_03577_),
    .C(_03581_),
    .A(_09077_),
    .Y(_03582_));
 sg13g2_o21ai_1 _21020_ (.B1(_03582_),
    .Y(_03583_),
    .A1(_03269_),
    .A2(_03570_));
 sg13g2_a21oi_1 _21021_ (.A1(_03116_),
    .A2(_03506_),
    .Y(_03584_),
    .B1(_03302_));
 sg13g2_nor2_1 _21022_ (.A(_03571_),
    .B(_03565_),
    .Y(_03585_));
 sg13g2_o21ai_1 _21023_ (.B1(_03585_),
    .Y(_03586_),
    .A1(_03285_),
    .A2(_03584_));
 sg13g2_o21ai_1 _21024_ (.B1(net155),
    .Y(_03587_),
    .A1(net294),
    .A2(_03254_));
 sg13g2_a21oi_1 _21025_ (.A1(_03450_),
    .A2(_03125_),
    .Y(_03588_),
    .B1(_03587_));
 sg13g2_nand2_1 _21026_ (.Y(_03589_),
    .A(_03254_),
    .B(_03410_));
 sg13g2_xnor2_1 _21027_ (.Y(_03590_),
    .A(_03307_),
    .B(_03589_));
 sg13g2_nor2_1 _21028_ (.A(net993),
    .B(_09073_),
    .Y(_03591_));
 sg13g2_a21oi_1 _21029_ (.A1(_08265_),
    .A2(_09073_),
    .Y(_03592_),
    .B1(_03591_));
 sg13g2_nor4_1 _21030_ (.A(_08884_),
    .B(_09825_),
    .C(_03590_),
    .D(_03592_),
    .Y(_03593_));
 sg13g2_nor4_1 _21031_ (.A(net209),
    .B(_03232_),
    .C(_03588_),
    .D(_03593_),
    .Y(_03594_));
 sg13g2_a21oi_1 _21032_ (.A1(_03586_),
    .A2(_03594_),
    .Y(_03595_),
    .B1(_03262_));
 sg13g2_nand3_1 _21033_ (.B(_03206_),
    .C(_03497_),
    .A(net155),
    .Y(_03596_));
 sg13g2_a21oi_1 _21034_ (.A1(_08885_),
    .A2(_03206_),
    .Y(_03597_),
    .B1(net156));
 sg13g2_nor2_1 _21035_ (.A(_03477_),
    .B(_03597_),
    .Y(_03598_));
 sg13g2_o21ai_1 _21036_ (.B1(_03598_),
    .Y(_03599_),
    .A1(_09816_),
    .A2(_03596_));
 sg13g2_o21ai_1 _21037_ (.B1(_03599_),
    .Y(_03600_),
    .A1(_03583_),
    .A2(_03595_));
 sg13g2_nand2_1 _21038_ (.Y(_03601_),
    .A(_09110_),
    .B(net107));
 sg13g2_o21ai_1 _21039_ (.B1(_03601_),
    .Y(_00786_),
    .A1(net146),
    .A2(_03600_));
 sg13g2_buf_1 _21040_ (.A(net1162),
    .X(_03602_));
 sg13g2_buf_1 _21041_ (.A(net992),
    .X(_03603_));
 sg13g2_nand2b_1 _21042_ (.Y(_03604_),
    .B(_10144_),
    .A_N(net1043));
 sg13g2_buf_1 _21043_ (.A(_03604_),
    .X(_03605_));
 sg13g2_nand3_1 _21044_ (.B(_11430_),
    .C(_10150_),
    .A(net1141),
    .Y(_03606_));
 sg13g2_buf_1 _21045_ (.A(_03606_),
    .X(_03607_));
 sg13g2_nor2_1 _21046_ (.A(_03605_),
    .B(_03607_),
    .Y(_03608_));
 sg13g2_buf_4 _21047_ (.X(_03609_),
    .A(_03608_));
 sg13g2_buf_1 _21048_ (.A(_03609_),
    .X(_03610_));
 sg13g2_mux2_1 _21049_ (.A0(\cpu.ex.r_10[0] ),
    .A1(net876),
    .S(net538),
    .X(_00791_));
 sg13g2_mux2_1 _21050_ (.A0(\cpu.ex.r_10[10] ),
    .A1(net879),
    .S(_03610_),
    .X(_00792_));
 sg13g2_mux2_1 _21051_ (.A0(\cpu.ex.r_10[11] ),
    .A1(net878),
    .S(net538),
    .X(_00793_));
 sg13g2_buf_1 _21052_ (.A(net627),
    .X(_03611_));
 sg13g2_nand2_1 _21053_ (.Y(_03612_),
    .A(net537),
    .B(_03609_));
 sg13g2_o21ai_1 _21054_ (.B1(_03612_),
    .Y(_00794_),
    .A1(_11281_),
    .A2(net538));
 sg13g2_buf_1 _21055_ (.A(net628),
    .X(_03613_));
 sg13g2_buf_1 _21056_ (.A(net536),
    .X(_03614_));
 sg13g2_mux2_1 _21057_ (.A0(\cpu.ex.r_10[13] ),
    .A1(net471),
    .S(net538),
    .X(_00795_));
 sg13g2_buf_1 _21058_ (.A(net698),
    .X(_03615_));
 sg13g2_buf_1 _21059_ (.A(net618),
    .X(_03616_));
 sg13g2_mux2_1 _21060_ (.A0(\cpu.ex.r_10[14] ),
    .A1(net535),
    .S(_03610_),
    .X(_00796_));
 sg13g2_buf_1 _21061_ (.A(_10730_),
    .X(_03617_));
 sg13g2_buf_1 _21062_ (.A(net617),
    .X(_03618_));
 sg13g2_mux2_1 _21063_ (.A0(\cpu.ex.r_10[15] ),
    .A1(net534),
    .S(net538),
    .X(_00797_));
 sg13g2_buf_1 _21064_ (.A(_10028_),
    .X(_03619_));
 sg13g2_mux2_1 _21065_ (.A0(\cpu.ex.r_10[1] ),
    .A1(net470),
    .S(net538),
    .X(_00798_));
 sg13g2_buf_2 _21066_ (.A(net622),
    .X(_03620_));
 sg13g2_buf_1 _21067_ (.A(net533),
    .X(_03621_));
 sg13g2_mux2_1 _21068_ (.A0(\cpu.ex.r_10[2] ),
    .A1(net469),
    .S(net538),
    .X(_00799_));
 sg13g2_buf_1 _21069_ (.A(_09193_),
    .X(_03622_));
 sg13g2_buf_1 _21070_ (.A(net418),
    .X(_03623_));
 sg13g2_mux2_1 _21071_ (.A0(\cpu.ex.r_10[3] ),
    .A1(net378),
    .S(net538),
    .X(_00800_));
 sg13g2_buf_2 _21072_ (.A(net677),
    .X(_03624_));
 sg13g2_buf_1 _21073_ (.A(net616),
    .X(_03625_));
 sg13g2_mux2_1 _21074_ (.A0(\cpu.ex.r_10[4] ),
    .A1(net532),
    .S(_03609_),
    .X(_00801_));
 sg13g2_mux2_1 _21075_ (.A0(\cpu.ex.r_10[5] ),
    .A1(_03073_),
    .S(_03609_),
    .X(_00802_));
 sg13g2_mux2_1 _21076_ (.A0(\cpu.ex.r_10[6] ),
    .A1(net749),
    .S(_03609_),
    .X(_00803_));
 sg13g2_mux2_1 _21077_ (.A0(\cpu.ex.r_10[7] ),
    .A1(net884),
    .S(_03609_),
    .X(_00804_));
 sg13g2_mux2_1 _21078_ (.A0(\cpu.ex.r_10[8] ),
    .A1(net883),
    .S(_03609_),
    .X(_00805_));
 sg13g2_mux2_1 _21079_ (.A0(\cpu.ex.r_10[9] ),
    .A1(net882),
    .S(_03609_),
    .X(_00806_));
 sg13g2_nor2_1 _21080_ (.A(_11449_),
    .B(_03607_),
    .Y(_03626_));
 sg13g2_buf_1 _21081_ (.A(_03626_),
    .X(_03627_));
 sg13g2_buf_1 _21082_ (.A(net615),
    .X(_03628_));
 sg13g2_mux2_1 _21083_ (.A0(\cpu.ex.r_11[0] ),
    .A1(net876),
    .S(net531),
    .X(_00807_));
 sg13g2_mux2_1 _21084_ (.A0(\cpu.ex.r_11[10] ),
    .A1(net879),
    .S(net531),
    .X(_00808_));
 sg13g2_mux2_1 _21085_ (.A0(\cpu.ex.r_11[11] ),
    .A1(net878),
    .S(_03628_),
    .X(_00809_));
 sg13g2_buf_1 _21086_ (.A(net537),
    .X(_03629_));
 sg13g2_mux2_1 _21087_ (.A0(\cpu.ex.r_11[12] ),
    .A1(net468),
    .S(net531),
    .X(_00810_));
 sg13g2_mux2_1 _21088_ (.A0(\cpu.ex.r_11[13] ),
    .A1(net471),
    .S(net531),
    .X(_00811_));
 sg13g2_nand2_1 _21089_ (.Y(_03630_),
    .A(net618),
    .B(net615));
 sg13g2_o21ai_1 _21090_ (.B1(_03630_),
    .Y(_00812_),
    .A1(_10670_),
    .A2(net531));
 sg13g2_mux2_1 _21091_ (.A0(\cpu.ex.r_11[15] ),
    .A1(net534),
    .S(net531),
    .X(_00813_));
 sg13g2_mux2_1 _21092_ (.A0(\cpu.ex.r_11[1] ),
    .A1(net470),
    .S(net531),
    .X(_00814_));
 sg13g2_mux2_1 _21093_ (.A0(\cpu.ex.r_11[2] ),
    .A1(net469),
    .S(net531),
    .X(_00815_));
 sg13g2_mux2_1 _21094_ (.A0(\cpu.ex.r_11[3] ),
    .A1(_03623_),
    .S(net615),
    .X(_00816_));
 sg13g2_mux2_1 _21095_ (.A0(\cpu.ex.r_11[4] ),
    .A1(net532),
    .S(net615),
    .X(_00817_));
 sg13g2_mux2_1 _21096_ (.A0(\cpu.ex.r_11[5] ),
    .A1(net542),
    .S(net615),
    .X(_00818_));
 sg13g2_nand2_1 _21097_ (.Y(_03631_),
    .A(net890),
    .B(_03627_));
 sg13g2_o21ai_1 _21098_ (.B1(_03631_),
    .Y(_00819_),
    .A1(_11143_),
    .A2(_03628_));
 sg13g2_mux2_1 _21099_ (.A0(\cpu.ex.r_11[7] ),
    .A1(net884),
    .S(net615),
    .X(_00820_));
 sg13g2_mux2_1 _21100_ (.A0(\cpu.ex.r_11[8] ),
    .A1(net883),
    .S(net615),
    .X(_00821_));
 sg13g2_mux2_1 _21101_ (.A0(\cpu.ex.r_11[9] ),
    .A1(net882),
    .S(net615),
    .X(_00822_));
 sg13g2_nand3_1 _21102_ (.B(_10148_),
    .C(_10150_),
    .A(net1141),
    .Y(_03632_));
 sg13g2_buf_1 _21103_ (.A(_03632_),
    .X(_03633_));
 sg13g2_nor3_1 _21104_ (.A(_10144_),
    .B(_10633_),
    .C(_03633_),
    .Y(_03634_));
 sg13g2_buf_2 _21105_ (.A(_03634_),
    .X(_03635_));
 sg13g2_buf_1 _21106_ (.A(_03635_),
    .X(_03636_));
 sg13g2_mux2_1 _21107_ (.A0(\cpu.ex.r_12[0] ),
    .A1(net876),
    .S(net614),
    .X(_00823_));
 sg13g2_mux2_1 _21108_ (.A0(\cpu.ex.r_12[10] ),
    .A1(net879),
    .S(_03636_),
    .X(_00824_));
 sg13g2_mux2_1 _21109_ (.A0(\cpu.ex.r_12[11] ),
    .A1(net878),
    .S(_03636_),
    .X(_00825_));
 sg13g2_mux2_1 _21110_ (.A0(\cpu.ex.r_12[12] ),
    .A1(net468),
    .S(net614),
    .X(_00826_));
 sg13g2_mux2_1 _21111_ (.A0(\cpu.ex.r_12[13] ),
    .A1(net471),
    .S(net614),
    .X(_00827_));
 sg13g2_mux2_1 _21112_ (.A0(\cpu.ex.r_12[14] ),
    .A1(net535),
    .S(net614),
    .X(_00828_));
 sg13g2_mux2_1 _21113_ (.A0(\cpu.ex.r_12[15] ),
    .A1(net534),
    .S(net614),
    .X(_00829_));
 sg13g2_mux2_1 _21114_ (.A0(\cpu.ex.r_12[1] ),
    .A1(net470),
    .S(net614),
    .X(_00830_));
 sg13g2_mux2_1 _21115_ (.A0(\cpu.ex.r_12[2] ),
    .A1(net469),
    .S(net614),
    .X(_00831_));
 sg13g2_mux2_1 _21116_ (.A0(\cpu.ex.r_12[3] ),
    .A1(_03623_),
    .S(net614),
    .X(_00832_));
 sg13g2_mux2_1 _21117_ (.A0(\cpu.ex.r_12[4] ),
    .A1(net532),
    .S(_03635_),
    .X(_00833_));
 sg13g2_mux2_1 _21118_ (.A0(\cpu.ex.r_12[5] ),
    .A1(_03073_),
    .S(_03635_),
    .X(_00834_));
 sg13g2_mux2_1 _21119_ (.A0(\cpu.ex.r_12[6] ),
    .A1(net749),
    .S(_03635_),
    .X(_00835_));
 sg13g2_mux2_1 _21120_ (.A0(\cpu.ex.r_12[7] ),
    .A1(net884),
    .S(_03635_),
    .X(_00836_));
 sg13g2_mux2_1 _21121_ (.A0(\cpu.ex.r_12[8] ),
    .A1(_03080_),
    .S(_03635_),
    .X(_00837_));
 sg13g2_mux2_1 _21122_ (.A0(\cpu.ex.r_12[9] ),
    .A1(_03082_),
    .S(_03635_),
    .X(_00838_));
 sg13g2_inv_1 _21123_ (.Y(_03637_),
    .A(net1142));
 sg13g2_nand2_1 _21124_ (.Y(_03638_),
    .A(_03637_),
    .B(net1043));
 sg13g2_nor2_1 _21125_ (.A(_03633_),
    .B(_03638_),
    .Y(_03639_));
 sg13g2_buf_2 _21126_ (.A(_03639_),
    .X(_03640_));
 sg13g2_buf_1 _21127_ (.A(_03640_),
    .X(_03641_));
 sg13g2_mux2_1 _21128_ (.A0(\cpu.ex.r_13[0] ),
    .A1(net876),
    .S(net613),
    .X(_00839_));
 sg13g2_mux2_1 _21129_ (.A0(\cpu.ex.r_13[10] ),
    .A1(net879),
    .S(_03641_),
    .X(_00840_));
 sg13g2_mux2_1 _21130_ (.A0(\cpu.ex.r_13[11] ),
    .A1(net878),
    .S(_03641_),
    .X(_00841_));
 sg13g2_mux2_1 _21131_ (.A0(\cpu.ex.r_13[12] ),
    .A1(_03629_),
    .S(net613),
    .X(_00842_));
 sg13g2_mux2_1 _21132_ (.A0(\cpu.ex.r_13[13] ),
    .A1(net471),
    .S(net613),
    .X(_00843_));
 sg13g2_mux2_1 _21133_ (.A0(\cpu.ex.r_13[14] ),
    .A1(net535),
    .S(net613),
    .X(_00844_));
 sg13g2_mux2_1 _21134_ (.A0(\cpu.ex.r_13[15] ),
    .A1(net534),
    .S(net613),
    .X(_00845_));
 sg13g2_mux2_1 _21135_ (.A0(\cpu.ex.r_13[1] ),
    .A1(net470),
    .S(net613),
    .X(_00846_));
 sg13g2_mux2_1 _21136_ (.A0(\cpu.ex.r_13[2] ),
    .A1(net469),
    .S(net613),
    .X(_00847_));
 sg13g2_mux2_1 _21137_ (.A0(\cpu.ex.r_13[3] ),
    .A1(net378),
    .S(net613),
    .X(_00848_));
 sg13g2_mux2_1 _21138_ (.A0(\cpu.ex.r_13[4] ),
    .A1(net532),
    .S(_03640_),
    .X(_00849_));
 sg13g2_buf_1 _21139_ (.A(_03072_),
    .X(_03642_));
 sg13g2_buf_1 _21140_ (.A(net530),
    .X(_03643_));
 sg13g2_mux2_1 _21141_ (.A0(\cpu.ex.r_13[5] ),
    .A1(net467),
    .S(_03640_),
    .X(_00850_));
 sg13g2_mux2_1 _21142_ (.A0(\cpu.ex.r_13[6] ),
    .A1(net749),
    .S(_03640_),
    .X(_00851_));
 sg13g2_mux2_1 _21143_ (.A0(\cpu.ex.r_13[7] ),
    .A1(net884),
    .S(_03640_),
    .X(_00852_));
 sg13g2_mux2_1 _21144_ (.A0(\cpu.ex.r_13[8] ),
    .A1(_03080_),
    .S(_03640_),
    .X(_00853_));
 sg13g2_mux2_1 _21145_ (.A0(\cpu.ex.r_13[9] ),
    .A1(_03082_),
    .S(_03640_),
    .X(_00854_));
 sg13g2_nor2_1 _21146_ (.A(_03605_),
    .B(_03633_),
    .Y(_03644_));
 sg13g2_buf_2 _21147_ (.A(_03644_),
    .X(_03645_));
 sg13g2_buf_1 _21148_ (.A(_03645_),
    .X(_03646_));
 sg13g2_mux2_1 _21149_ (.A0(\cpu.ex.r_14[0] ),
    .A1(net876),
    .S(net529),
    .X(_00855_));
 sg13g2_mux2_1 _21150_ (.A0(\cpu.ex.r_14[10] ),
    .A1(net879),
    .S(net529),
    .X(_00856_));
 sg13g2_mux2_1 _21151_ (.A0(\cpu.ex.r_14[11] ),
    .A1(net878),
    .S(net529),
    .X(_00857_));
 sg13g2_mux2_1 _21152_ (.A0(\cpu.ex.r_14[12] ),
    .A1(net468),
    .S(net529),
    .X(_00858_));
 sg13g2_mux2_1 _21153_ (.A0(\cpu.ex.r_14[13] ),
    .A1(_03614_),
    .S(net529),
    .X(_00859_));
 sg13g2_mux2_1 _21154_ (.A0(\cpu.ex.r_14[14] ),
    .A1(net535),
    .S(net529),
    .X(_00860_));
 sg13g2_mux2_1 _21155_ (.A0(\cpu.ex.r_14[15] ),
    .A1(_03618_),
    .S(net529),
    .X(_00861_));
 sg13g2_mux2_1 _21156_ (.A0(\cpu.ex.r_14[1] ),
    .A1(net470),
    .S(net529),
    .X(_00862_));
 sg13g2_mux2_1 _21157_ (.A0(\cpu.ex.r_14[2] ),
    .A1(_03621_),
    .S(_03646_),
    .X(_00863_));
 sg13g2_mux2_1 _21158_ (.A0(\cpu.ex.r_14[3] ),
    .A1(net378),
    .S(_03646_),
    .X(_00864_));
 sg13g2_mux2_1 _21159_ (.A0(\cpu.ex.r_14[4] ),
    .A1(_03625_),
    .S(_03645_),
    .X(_00865_));
 sg13g2_mux2_1 _21160_ (.A0(\cpu.ex.r_14[5] ),
    .A1(net467),
    .S(_03645_),
    .X(_00866_));
 sg13g2_mux2_1 _21161_ (.A0(\cpu.ex.r_14[6] ),
    .A1(net749),
    .S(_03645_),
    .X(_00867_));
 sg13g2_mux2_1 _21162_ (.A0(\cpu.ex.r_14[7] ),
    .A1(net884),
    .S(_03645_),
    .X(_00868_));
 sg13g2_buf_1 _21163_ (.A(_03079_),
    .X(_03647_));
 sg13g2_mux2_1 _21164_ (.A0(\cpu.ex.r_14[8] ),
    .A1(net875),
    .S(_03645_),
    .X(_00869_));
 sg13g2_buf_1 _21165_ (.A(net995),
    .X(_03648_));
 sg13g2_mux2_1 _21166_ (.A0(\cpu.ex.r_14[9] ),
    .A1(net874),
    .S(_03645_),
    .X(_00870_));
 sg13g2_nor2_1 _21167_ (.A(_11449_),
    .B(_03633_),
    .Y(_03649_));
 sg13g2_buf_2 _21168_ (.A(_03649_),
    .X(_03650_));
 sg13g2_buf_1 _21169_ (.A(_03650_),
    .X(_03651_));
 sg13g2_mux2_1 _21170_ (.A0(\cpu.ex.r_15[0] ),
    .A1(net876),
    .S(net612),
    .X(_00871_));
 sg13g2_mux2_1 _21171_ (.A0(\cpu.ex.r_15[10] ),
    .A1(net879),
    .S(_03651_),
    .X(_00872_));
 sg13g2_mux2_1 _21172_ (.A0(\cpu.ex.r_15[11] ),
    .A1(net878),
    .S(_03651_),
    .X(_00873_));
 sg13g2_mux2_1 _21173_ (.A0(\cpu.ex.r_15[12] ),
    .A1(net468),
    .S(net612),
    .X(_00874_));
 sg13g2_mux2_1 _21174_ (.A0(\cpu.ex.r_15[13] ),
    .A1(_03614_),
    .S(net612),
    .X(_00875_));
 sg13g2_mux2_1 _21175_ (.A0(\cpu.ex.r_15[14] ),
    .A1(_03616_),
    .S(net612),
    .X(_00876_));
 sg13g2_mux2_1 _21176_ (.A0(\cpu.ex.r_15[15] ),
    .A1(_03618_),
    .S(net612),
    .X(_00877_));
 sg13g2_mux2_1 _21177_ (.A0(\cpu.ex.r_15[1] ),
    .A1(net470),
    .S(net612),
    .X(_00878_));
 sg13g2_mux2_1 _21178_ (.A0(\cpu.ex.r_15[2] ),
    .A1(net469),
    .S(net612),
    .X(_00879_));
 sg13g2_mux2_1 _21179_ (.A0(\cpu.ex.r_15[3] ),
    .A1(net378),
    .S(net612),
    .X(_00880_));
 sg13g2_mux2_1 _21180_ (.A0(\cpu.ex.r_15[4] ),
    .A1(net532),
    .S(_03650_),
    .X(_00881_));
 sg13g2_mux2_1 _21181_ (.A0(\cpu.ex.r_15[5] ),
    .A1(net467),
    .S(_03650_),
    .X(_00882_));
 sg13g2_mux2_1 _21182_ (.A0(\cpu.ex.r_15[6] ),
    .A1(net749),
    .S(_03650_),
    .X(_00883_));
 sg13g2_mux2_1 _21183_ (.A0(\cpu.ex.r_15[7] ),
    .A1(_03078_),
    .S(_03650_),
    .X(_00884_));
 sg13g2_mux2_1 _21184_ (.A0(\cpu.ex.r_15[8] ),
    .A1(net875),
    .S(_03650_),
    .X(_00885_));
 sg13g2_mux2_1 _21185_ (.A0(\cpu.ex.r_15[9] ),
    .A1(net874),
    .S(_03650_),
    .X(_00886_));
 sg13g2_nor3_1 _21186_ (.A(net1142),
    .B(net1043),
    .C(_03607_),
    .Y(_03652_));
 sg13g2_buf_1 _21187_ (.A(_03652_),
    .X(_03653_));
 sg13g2_buf_1 _21188_ (.A(net611),
    .X(_03654_));
 sg13g2_mux2_1 _21189_ (.A0(\cpu.ex.r_8[0] ),
    .A1(net876),
    .S(net528),
    .X(_00887_));
 sg13g2_mux2_1 _21190_ (.A0(\cpu.ex.r_8[10] ),
    .A1(_03104_),
    .S(net528),
    .X(_00888_));
 sg13g2_mux2_1 _21191_ (.A0(\cpu.ex.r_8[11] ),
    .A1(_03105_),
    .S(net528),
    .X(_00889_));
 sg13g2_mux2_1 _21192_ (.A0(\cpu.ex.r_8[12] ),
    .A1(_03629_),
    .S(net528),
    .X(_00890_));
 sg13g2_buf_1 _21193_ (.A(net536),
    .X(_03655_));
 sg13g2_mux2_1 _21194_ (.A0(\cpu.ex.r_8[13] ),
    .A1(net466),
    .S(net528),
    .X(_00891_));
 sg13g2_inv_1 _21195_ (.Y(_03656_),
    .A(\cpu.ex.r_8[14] ));
 sg13g2_nand2_1 _21196_ (.Y(_03657_),
    .A(_03615_),
    .B(net611));
 sg13g2_o21ai_1 _21197_ (.B1(_03657_),
    .Y(_00892_),
    .A1(_03656_),
    .A2(net528));
 sg13g2_buf_1 _21198_ (.A(net617),
    .X(_03658_));
 sg13g2_mux2_1 _21199_ (.A0(\cpu.ex.r_8[15] ),
    .A1(net527),
    .S(_03654_),
    .X(_00893_));
 sg13g2_mux2_1 _21200_ (.A0(\cpu.ex.r_8[1] ),
    .A1(net470),
    .S(net528),
    .X(_00894_));
 sg13g2_mux2_1 _21201_ (.A0(\cpu.ex.r_8[2] ),
    .A1(net469),
    .S(net528),
    .X(_00895_));
 sg13g2_mux2_1 _21202_ (.A0(\cpu.ex.r_8[3] ),
    .A1(net378),
    .S(net611),
    .X(_00896_));
 sg13g2_mux2_1 _21203_ (.A0(\cpu.ex.r_8[4] ),
    .A1(net532),
    .S(net611),
    .X(_00897_));
 sg13g2_inv_1 _21204_ (.Y(_03659_),
    .A(\cpu.ex.r_8[5] ));
 sg13g2_nand2_1 _21205_ (.Y(_03660_),
    .A(net530),
    .B(net611));
 sg13g2_o21ai_1 _21206_ (.B1(_03660_),
    .Y(_00898_),
    .A1(_03659_),
    .A2(_03654_));
 sg13g2_mux2_1 _21207_ (.A0(\cpu.ex.r_8[6] ),
    .A1(net749),
    .S(net611),
    .X(_00899_));
 sg13g2_mux2_1 _21208_ (.A0(\cpu.ex.r_8[7] ),
    .A1(_03078_),
    .S(net611),
    .X(_00900_));
 sg13g2_mux2_1 _21209_ (.A0(\cpu.ex.r_8[8] ),
    .A1(net875),
    .S(net611),
    .X(_00901_));
 sg13g2_mux2_1 _21210_ (.A0(\cpu.ex.r_8[9] ),
    .A1(net874),
    .S(_03653_),
    .X(_00902_));
 sg13g2_nor2_1 _21211_ (.A(_03607_),
    .B(_03638_),
    .Y(_03661_));
 sg13g2_buf_2 _21212_ (.A(_03661_),
    .X(_03662_));
 sg13g2_buf_1 _21213_ (.A(_03662_),
    .X(_03663_));
 sg13g2_mux2_1 _21214_ (.A0(\cpu.ex.r_9[0] ),
    .A1(net876),
    .S(net526),
    .X(_00903_));
 sg13g2_mux2_1 _21215_ (.A0(\cpu.ex.r_9[10] ),
    .A1(_03104_),
    .S(net526),
    .X(_00904_));
 sg13g2_mux2_1 _21216_ (.A0(\cpu.ex.r_9[11] ),
    .A1(_03105_),
    .S(net526),
    .X(_00905_));
 sg13g2_buf_1 _21217_ (.A(net627),
    .X(_03664_));
 sg13g2_mux2_1 _21218_ (.A0(\cpu.ex.r_9[12] ),
    .A1(_03664_),
    .S(_03663_),
    .X(_00906_));
 sg13g2_mux2_1 _21219_ (.A0(\cpu.ex.r_9[13] ),
    .A1(net466),
    .S(_03663_),
    .X(_00907_));
 sg13g2_mux2_1 _21220_ (.A0(\cpu.ex.r_9[14] ),
    .A1(_03616_),
    .S(net526),
    .X(_00908_));
 sg13g2_mux2_1 _21221_ (.A0(\cpu.ex.r_9[15] ),
    .A1(net527),
    .S(net526),
    .X(_00909_));
 sg13g2_mux2_1 _21222_ (.A0(\cpu.ex.r_9[1] ),
    .A1(net470),
    .S(net526),
    .X(_00910_));
 sg13g2_mux2_1 _21223_ (.A0(\cpu.ex.r_9[2] ),
    .A1(net469),
    .S(net526),
    .X(_00911_));
 sg13g2_mux2_1 _21224_ (.A0(\cpu.ex.r_9[3] ),
    .A1(net378),
    .S(net526),
    .X(_00912_));
 sg13g2_mux2_1 _21225_ (.A0(\cpu.ex.r_9[4] ),
    .A1(net532),
    .S(_03662_),
    .X(_00913_));
 sg13g2_mux2_1 _21226_ (.A0(\cpu.ex.r_9[5] ),
    .A1(net467),
    .S(_03662_),
    .X(_00914_));
 sg13g2_mux2_1 _21227_ (.A0(\cpu.ex.r_9[6] ),
    .A1(_03102_),
    .S(_03662_),
    .X(_00915_));
 sg13g2_buf_1 _21228_ (.A(net997),
    .X(_03665_));
 sg13g2_mux2_1 _21229_ (.A0(\cpu.ex.r_9[7] ),
    .A1(net873),
    .S(_03662_),
    .X(_00916_));
 sg13g2_mux2_1 _21230_ (.A0(\cpu.ex.r_9[8] ),
    .A1(net875),
    .S(_03662_),
    .X(_00917_));
 sg13g2_mux2_1 _21231_ (.A0(\cpu.ex.r_9[9] ),
    .A1(net874),
    .S(_03662_),
    .X(_00918_));
 sg13g2_nand4_1 _21232_ (.B(net1043),
    .C(_10150_),
    .A(net1142),
    .Y(_03666_),
    .D(_10149_));
 sg13g2_nand2b_1 _21233_ (.Y(_03667_),
    .B(_08266_),
    .A_N(_03666_));
 sg13g2_buf_1 _21234_ (.A(_03667_),
    .X(_03668_));
 sg13g2_buf_1 _21235_ (.A(_03668_),
    .X(_03669_));
 sg13g2_buf_1 _21236_ (.A(_03668_),
    .X(_03670_));
 sg13g2_nand2_1 _21237_ (.Y(_03671_),
    .A(\cpu.ex.r_epc[1] ),
    .B(_03670_));
 sg13g2_o21ai_1 _21238_ (.B1(_03671_),
    .Y(_00920_),
    .A1(_10041_),
    .A2(net610));
 sg13g2_mux2_1 _21239_ (.A0(_03071_),
    .A1(\cpu.ex.r_epc[11] ),
    .S(net610),
    .X(_00921_));
 sg13g2_buf_1 _21240_ (.A(net537),
    .X(_03672_));
 sg13g2_mux2_1 _21241_ (.A0(_03672_),
    .A1(\cpu.ex.r_epc[12] ),
    .S(net610),
    .X(_00922_));
 sg13g2_buf_1 _21242_ (.A(net536),
    .X(_03673_));
 sg13g2_mux2_1 _21243_ (.A0(_03673_),
    .A1(\cpu.ex.r_epc[13] ),
    .S(net610),
    .X(_00923_));
 sg13g2_buf_1 _21244_ (.A(net618),
    .X(_03674_));
 sg13g2_mux2_1 _21245_ (.A0(_03674_),
    .A1(\cpu.ex.r_epc[14] ),
    .S(net609),
    .X(_00924_));
 sg13g2_buf_1 _21246_ (.A(net617),
    .X(_03675_));
 sg13g2_mux2_1 _21247_ (.A0(_03675_),
    .A1(\cpu.ex.r_epc[15] ),
    .S(net609),
    .X(_00925_));
 sg13g2_nand2_1 _21248_ (.Y(_03676_),
    .A(\cpu.ex.r_epc[2] ),
    .B(net609));
 sg13g2_o21ai_1 _21249_ (.B1(_03676_),
    .Y(_00926_),
    .A1(net767),
    .A2(net610));
 sg13g2_mux2_1 _21250_ (.A0(net378),
    .A1(\cpu.ex.r_epc[3] ),
    .S(net609),
    .X(_00927_));
 sg13g2_buf_1 _21251_ (.A(net679),
    .X(_03677_));
 sg13g2_buf_1 _21252_ (.A(net608),
    .X(_03678_));
 sg13g2_nand2_1 _21253_ (.Y(_03679_),
    .A(\cpu.ex.r_epc[4] ),
    .B(net609));
 sg13g2_o21ai_1 _21254_ (.B1(_03679_),
    .Y(_00928_),
    .A1(_03678_),
    .A2(net610));
 sg13g2_nand2_1 _21255_ (.Y(_03680_),
    .A(\cpu.ex.r_epc[5] ),
    .B(net609));
 sg13g2_o21ai_1 _21256_ (.B1(_03680_),
    .Y(_00929_),
    .A1(net674),
    .A2(_03669_));
 sg13g2_mux2_1 _21257_ (.A0(_03058_),
    .A1(\cpu.ex.r_epc[6] ),
    .S(_03670_),
    .X(_00930_));
 sg13g2_nand2_1 _21258_ (.Y(_03681_),
    .A(\cpu.ex.r_epc[7] ),
    .B(net609));
 sg13g2_o21ai_1 _21259_ (.B1(_03681_),
    .Y(_00931_),
    .A1(net753),
    .A2(net610));
 sg13g2_nand2_1 _21260_ (.Y(_03682_),
    .A(\cpu.ex.r_epc[8] ),
    .B(_03668_));
 sg13g2_o21ai_1 _21261_ (.B1(_03682_),
    .Y(_00932_),
    .A1(net752),
    .A2(net610));
 sg13g2_nand2_1 _21262_ (.Y(_03683_),
    .A(\cpu.ex.r_epc[9] ),
    .B(_03668_));
 sg13g2_o21ai_1 _21263_ (.B1(_03683_),
    .Y(_00933_),
    .A1(net751),
    .A2(_03669_));
 sg13g2_mux2_1 _21264_ (.A0(_03069_),
    .A1(\cpu.ex.r_epc[10] ),
    .S(net609),
    .X(_00934_));
 sg13g2_nand4_1 _21265_ (.B(net1043),
    .C(_10150_),
    .A(_03637_),
    .Y(_03684_),
    .D(_10149_));
 sg13g2_buf_1 _21266_ (.A(_03684_),
    .X(_03685_));
 sg13g2_buf_1 _21267_ (.A(_03685_),
    .X(_03686_));
 sg13g2_buf_1 _21268_ (.A(_03685_),
    .X(_03687_));
 sg13g2_nand2_1 _21269_ (.Y(_03688_),
    .A(\cpu.ex.r_lr[1] ),
    .B(net672));
 sg13g2_o21ai_1 _21270_ (.B1(_03688_),
    .Y(_00940_),
    .A1(_10041_),
    .A2(_03686_));
 sg13g2_mux2_1 _21271_ (.A0(_03071_),
    .A1(\cpu.ex.r_lr[11] ),
    .S(net673),
    .X(_00941_));
 sg13g2_mux2_1 _21272_ (.A0(_03672_),
    .A1(\cpu.ex.r_lr[12] ),
    .S(net673),
    .X(_00942_));
 sg13g2_mux2_1 _21273_ (.A0(net464),
    .A1(\cpu.ex.r_lr[13] ),
    .S(net673),
    .X(_00943_));
 sg13g2_mux2_1 _21274_ (.A0(_03674_),
    .A1(\cpu.ex.r_lr[14] ),
    .S(net672),
    .X(_00944_));
 sg13g2_mux2_1 _21275_ (.A0(_03675_),
    .A1(\cpu.ex.r_lr[15] ),
    .S(net672),
    .X(_00945_));
 sg13g2_nand2_1 _21276_ (.Y(_03689_),
    .A(\cpu.ex.r_lr[2] ),
    .B(net672));
 sg13g2_o21ai_1 _21277_ (.B1(_03689_),
    .Y(_00946_),
    .A1(net767),
    .A2(net673));
 sg13g2_mux2_1 _21278_ (.A0(net378),
    .A1(\cpu.ex.r_lr[3] ),
    .S(net672),
    .X(_00947_));
 sg13g2_nand2_1 _21279_ (.Y(_03690_),
    .A(\cpu.ex.r_lr[4] ),
    .B(net672));
 sg13g2_o21ai_1 _21280_ (.B1(_03690_),
    .Y(_00948_),
    .A1(_03678_),
    .A2(net673));
 sg13g2_nand2_1 _21281_ (.Y(_03691_),
    .A(\cpu.ex.r_lr[5] ),
    .B(_03687_));
 sg13g2_o21ai_1 _21282_ (.B1(_03691_),
    .Y(_00949_),
    .A1(net674),
    .A2(net673));
 sg13g2_mux2_1 _21283_ (.A0(_03058_),
    .A1(\cpu.ex.r_lr[6] ),
    .S(net672),
    .X(_00950_));
 sg13g2_nand2_1 _21284_ (.Y(_03692_),
    .A(\cpu.ex.r_lr[7] ),
    .B(net672));
 sg13g2_o21ai_1 _21285_ (.B1(_03692_),
    .Y(_00951_),
    .A1(net753),
    .A2(net673));
 sg13g2_nand2_1 _21286_ (.Y(_03693_),
    .A(\cpu.ex.r_lr[8] ),
    .B(_03685_));
 sg13g2_o21ai_1 _21287_ (.B1(_03693_),
    .Y(_00952_),
    .A1(net752),
    .A2(net673));
 sg13g2_nand2_1 _21288_ (.Y(_03694_),
    .A(\cpu.ex.r_lr[9] ),
    .B(_03685_));
 sg13g2_o21ai_1 _21289_ (.B1(_03694_),
    .Y(_00953_),
    .A1(net751),
    .A2(_03686_));
 sg13g2_mux2_1 _21290_ (.A0(_03069_),
    .A1(\cpu.ex.r_lr[10] ),
    .S(_03687_),
    .X(_00954_));
 sg13g2_nor2b_1 _21291_ (.A(net74),
    .B_N(net348),
    .Y(_03695_));
 sg13g2_buf_1 _21292_ (.A(_03695_),
    .X(_03696_));
 sg13g2_nor2_1 _21293_ (.A(_11397_),
    .B(_11411_),
    .Y(_03697_));
 sg13g2_buf_8 _21294_ (.A(_03697_),
    .X(_03698_));
 sg13g2_buf_8 _21295_ (.A(net29),
    .X(_03699_));
 sg13g2_nor2_1 _21296_ (.A(net258),
    .B(net27),
    .Y(_03700_));
 sg13g2_xnor2_1 _21297_ (.Y(_03701_),
    .A(net91),
    .B(_03700_));
 sg13g2_mux2_1 _21298_ (.A0(_11980_),
    .A1(_11951_),
    .S(_11360_),
    .X(_03702_));
 sg13g2_a22oi_1 _21299_ (.Y(_03703_),
    .B1(_03702_),
    .B2(_11996_),
    .A2(_11360_),
    .A1(net626));
 sg13g2_inv_1 _21300_ (.Y(_03704_),
    .A(_11951_));
 sg13g2_inv_1 _21301_ (.Y(_03705_),
    .A(_11360_));
 sg13g2_or4_1 _21302_ (.A(_03704_),
    .B(_03705_),
    .C(_11386_),
    .D(_11954_),
    .X(_03706_));
 sg13g2_o21ai_1 _21303_ (.B1(_03706_),
    .Y(_03707_),
    .A1(_11387_),
    .A2(_03703_));
 sg13g2_nand2_1 _21304_ (.Y(_03708_),
    .A(_03705_),
    .B(_11387_));
 sg13g2_nand3_1 _21305_ (.B(_03704_),
    .C(net554),
    .A(_11938_),
    .Y(_03709_));
 sg13g2_a21oi_1 _21306_ (.A1(_11643_),
    .A2(_03708_),
    .Y(_03710_),
    .B1(_03709_));
 sg13g2_a21o_1 _21307_ (.A2(_03707_),
    .A1(net90),
    .B1(_03710_),
    .X(_03711_));
 sg13g2_a22oi_1 _21308_ (.Y(_03712_),
    .B1(_11386_),
    .B2(_11938_),
    .A2(_11360_),
    .A1(_03704_));
 sg13g2_a21oi_1 _21309_ (.A1(_11951_),
    .A2(_03705_),
    .Y(_03713_),
    .B1(_03712_));
 sg13g2_nor2b_1 _21310_ (.A(_11879_),
    .B_N(_03713_),
    .Y(_03714_));
 sg13g2_a221oi_1 _21311_ (.B2(_03711_),
    .C1(_03714_),
    .B1(_11975_),
    .A1(\cpu.ex.r_mult[15] ),
    .Y(_03715_),
    .A2(_11660_));
 sg13g2_nand3_1 _21312_ (.B(net90),
    .C(_03713_),
    .A(net554),
    .Y(_03716_));
 sg13g2_and2_1 _21313_ (.A(_11974_),
    .B(_03716_),
    .X(_03717_));
 sg13g2_and2_1 _21314_ (.A(\cpu.ex.r_mult[15] ),
    .B(net554),
    .X(_03718_));
 sg13g2_o21ai_1 _21315_ (.B1(_03718_),
    .Y(_03719_),
    .A1(_03711_),
    .A2(_03714_));
 sg13g2_a21o_1 _21316_ (.A2(_03717_),
    .A1(_11969_),
    .B1(_03719_),
    .X(_03720_));
 sg13g2_buf_1 _21317_ (.A(_03720_),
    .X(_03721_));
 sg13g2_nand2_1 _21318_ (.Y(_03722_),
    .A(net492),
    .B(_03721_));
 sg13g2_nand2_1 _21319_ (.Y(_03723_),
    .A(_10561_),
    .B(net385));
 sg13g2_o21ai_1 _21320_ (.B1(_03723_),
    .Y(_03724_),
    .A1(_03715_),
    .A2(_03722_));
 sg13g2_a21oi_1 _21321_ (.A1(net32),
    .A2(_03701_),
    .Y(_03725_),
    .B1(_03724_));
 sg13g2_buf_1 _21322_ (.A(net486),
    .X(_03726_));
 sg13g2_nand2_1 _21323_ (.Y(_03727_),
    .A(_03603_),
    .B(net417));
 sg13g2_o21ai_1 _21324_ (.B1(_03727_),
    .Y(_00955_),
    .A1(net485),
    .A2(_03725_));
 sg13g2_inv_1 _21325_ (.Y(_03728_),
    .A(net1044));
 sg13g2_nand2_2 _21326_ (.Y(_03729_),
    .A(net646),
    .B(_11626_));
 sg13g2_nor2_1 _21327_ (.A(net485),
    .B(_03729_),
    .Y(_03730_));
 sg13g2_buf_1 _21328_ (.A(_03730_),
    .X(_03731_));
 sg13g2_buf_1 _21329_ (.A(_11475_),
    .X(_03732_));
 sg13g2_buf_1 _21330_ (.A(net193),
    .X(_03733_));
 sg13g2_buf_1 _21331_ (.A(_11413_),
    .X(_03734_));
 sg13g2_buf_1 _21332_ (.A(net248),
    .X(_03735_));
 sg13g2_nand2_1 _21333_ (.Y(_03736_),
    .A(_03735_),
    .B(net91));
 sg13g2_xnor2_1 _21334_ (.Y(_03737_),
    .A(net172),
    .B(_03736_));
 sg13g2_o21ai_1 _21335_ (.B1(_11167_),
    .Y(_03738_),
    .A1(_03699_),
    .A2(_03737_));
 sg13g2_or3_1 _21336_ (.A(_11167_),
    .B(net29),
    .C(_03737_),
    .X(_03739_));
 sg13g2_nand2_1 _21337_ (.Y(_03740_),
    .A(net348),
    .B(_11427_));
 sg13g2_a21oi_1 _21338_ (.A1(_03738_),
    .A2(_03739_),
    .Y(_03741_),
    .B1(_03740_));
 sg13g2_nand2_2 _21339_ (.Y(_03742_),
    .A(net1034),
    .B(net435));
 sg13g2_xnor2_1 _21340_ (.Y(_03743_),
    .A(_10562_),
    .B(_03721_));
 sg13g2_o21ai_1 _21341_ (.B1(_03729_),
    .Y(_03744_),
    .A1(_03742_),
    .A2(_03743_));
 sg13g2_o21ai_1 _21342_ (.B1(_11435_),
    .Y(_03745_),
    .A1(_03741_),
    .A2(_03744_));
 sg13g2_nand2_1 _21343_ (.Y(_03746_),
    .A(_03619_),
    .B(net417));
 sg13g2_a22oi_1 _21344_ (.Y(_00956_),
    .B1(_03745_),
    .B2(_03746_),
    .A2(net377),
    .A1(_03728_));
 sg13g2_buf_1 _21345_ (.A(_10540_),
    .X(_03747_));
 sg13g2_nor2_1 _21346_ (.A(net172),
    .B(_03736_),
    .Y(_03748_));
 sg13g2_a21oi_1 _21347_ (.A1(net172),
    .A2(_03736_),
    .Y(_03749_),
    .B1(_11167_));
 sg13g2_nor2_1 _21348_ (.A(_03748_),
    .B(_03749_),
    .Y(_03750_));
 sg13g2_xnor2_1 _21349_ (.Y(_03751_),
    .A(net259),
    .B(_03750_));
 sg13g2_nor2_1 _21350_ (.A(net29),
    .B(_03751_),
    .Y(_03752_));
 sg13g2_xnor2_1 _21351_ (.Y(_03753_),
    .A(_10558_),
    .B(_03752_));
 sg13g2_nor2_1 _21352_ (.A(_10562_),
    .B(_03721_),
    .Y(_03754_));
 sg13g2_nand3b_1 _21353_ (.B(net1044),
    .C(net435),
    .Y(_03755_),
    .A_N(_03754_));
 sg13g2_nand2_1 _21354_ (.Y(_03756_),
    .A(_03728_),
    .B(_03754_));
 sg13g2_a21oi_1 _21355_ (.A1(_03755_),
    .A2(_03756_),
    .Y(_03757_),
    .B1(_09294_));
 sg13g2_a221oi_1 _21356_ (.B2(_03753_),
    .C1(_03757_),
    .B1(net32),
    .A1(net991),
    .Y(_03758_),
    .A2(net385));
 sg13g2_nand2_1 _21357_ (.Y(_03759_),
    .A(net533),
    .B(net417));
 sg13g2_o21ai_1 _21358_ (.B1(_03759_),
    .Y(_00957_),
    .A1(net485),
    .A2(_03758_));
 sg13g2_a22oi_1 _21359_ (.Y(_03760_),
    .B1(net377),
    .B2(net1131),
    .A2(net417),
    .A1(net418));
 sg13g2_nor2_1 _21360_ (.A(net485),
    .B(_03742_),
    .Y(_03761_));
 sg13g2_buf_2 _21361_ (.A(_03761_),
    .X(_03762_));
 sg13g2_nand2_1 _21362_ (.Y(_03763_),
    .A(net1044),
    .B(_03754_));
 sg13g2_xnor2_1 _21363_ (.Y(_03764_),
    .A(net991),
    .B(_03763_));
 sg13g2_nor2_1 _21364_ (.A(net434),
    .B(net555),
    .Y(_03765_));
 sg13g2_and2_1 _21365_ (.A(_03695_),
    .B(_03765_),
    .X(_03766_));
 sg13g2_buf_1 _21366_ (.A(_03766_),
    .X(_03767_));
 sg13g2_or4_1 _21367_ (.A(_10841_),
    .B(_10958_),
    .C(_11164_),
    .D(_11188_),
    .X(_03768_));
 sg13g2_nand2_1 _21368_ (.Y(_03769_),
    .A(net231),
    .B(_10560_));
 sg13g2_a21oi_1 _21369_ (.A1(_10601_),
    .A2(_03768_),
    .Y(_03770_),
    .B1(_03769_));
 sg13g2_nand2_1 _21370_ (.Y(_03771_),
    .A(_10601_),
    .B(_03768_));
 sg13g2_a21oi_1 _21371_ (.A1(_10560_),
    .A2(_03771_),
    .Y(_03772_),
    .B1(net199));
 sg13g2_nor3_1 _21372_ (.A(net27),
    .B(_03770_),
    .C(_03772_),
    .Y(_03773_));
 sg13g2_xnor2_1 _21373_ (.Y(_03774_),
    .A(_10603_),
    .B(_03773_));
 sg13g2_a22oi_1 _21374_ (.Y(_03775_),
    .B1(_03767_),
    .B2(_03774_),
    .A2(_03764_),
    .A1(_03762_));
 sg13g2_nand2_1 _21375_ (.Y(_00958_),
    .A(_03760_),
    .B(_03775_));
 sg13g2_a22oi_1 _21376_ (.Y(_03776_),
    .B1(net377),
    .B2(net1130),
    .A2(net417),
    .A1(net616));
 sg13g2_and3_1 _21377_ (.X(_03777_),
    .A(net1044),
    .B(net991),
    .C(_03754_));
 sg13g2_xnor2_1 _21378_ (.Y(_03778_),
    .A(_11065_),
    .B(_03777_));
 sg13g2_buf_1 _21379_ (.A(net489),
    .X(_03779_));
 sg13g2_nand2_1 _21380_ (.Y(_03780_),
    .A(net1131),
    .B(net416));
 sg13g2_xnor2_1 _21381_ (.Y(_03781_),
    .A(net253),
    .B(_11230_));
 sg13g2_nor2_1 _21382_ (.A(_03699_),
    .B(_03781_),
    .Y(_03782_));
 sg13g2_xnor2_1 _21383_ (.Y(_03783_),
    .A(_03780_),
    .B(_03782_));
 sg13g2_a22oi_1 _21384_ (.Y(_03784_),
    .B1(_03783_),
    .B2(_03767_),
    .A2(_03778_),
    .A1(_03762_));
 sg13g2_nand2_1 _21385_ (.Y(_00959_),
    .A(_03776_),
    .B(_03784_));
 sg13g2_nand3_1 _21386_ (.B(net416),
    .C(net32),
    .A(net1130),
    .Y(_03785_));
 sg13g2_nand2_1 _21387_ (.Y(_03786_),
    .A(_10513_),
    .B(net32));
 sg13g2_buf_1 _21388_ (.A(_11694_),
    .X(_03787_));
 sg13g2_nand3_1 _21389_ (.B(net192),
    .C(net303),
    .A(net1131),
    .Y(_03788_));
 sg13g2_xnor2_1 _21390_ (.Y(_03789_),
    .A(_10450_),
    .B(net303));
 sg13g2_nand3_1 _21391_ (.B(net231),
    .C(_03789_),
    .A(net991),
    .Y(_03790_));
 sg13g2_o21ai_1 _21392_ (.B1(_03790_),
    .Y(_03791_),
    .A1(net991),
    .A2(_03788_));
 sg13g2_o21ai_1 _21393_ (.B1(net489),
    .Y(_03792_),
    .A1(net991),
    .A2(net1131));
 sg13g2_nor2_1 _21394_ (.A(net199),
    .B(net253),
    .Y(_03793_));
 sg13g2_a22oi_1 _21395_ (.Y(_03794_),
    .B1(_03792_),
    .B2(_03793_),
    .A2(_03791_),
    .A1(net489));
 sg13g2_nor2_2 _21396_ (.A(_11663_),
    .B(net200),
    .Y(_03795_));
 sg13g2_o21ai_1 _21397_ (.B1(_11442_),
    .Y(_03796_),
    .A1(_10561_),
    .A2(net1044));
 sg13g2_nand3_1 _21398_ (.B(_10557_),
    .C(net226),
    .A(_10562_),
    .Y(_03797_));
 sg13g2_xnor2_1 _21399_ (.Y(_03798_),
    .A(_03728_),
    .B(net259));
 sg13g2_nand3_1 _21400_ (.B(net200),
    .C(_03798_),
    .A(_10561_),
    .Y(_03799_));
 sg13g2_o21ai_1 _21401_ (.B1(_03799_),
    .Y(_03800_),
    .A1(net200),
    .A2(_03797_));
 sg13g2_a22oi_1 _21402_ (.Y(_03801_),
    .B1(_03800_),
    .B2(_11442_),
    .A2(_03796_),
    .A1(_03795_));
 sg13g2_nor2_1 _21403_ (.A(_03794_),
    .B(_03801_),
    .Y(_03802_));
 sg13g2_a22oi_1 _21404_ (.Y(_03803_),
    .B1(net193),
    .B2(_10561_),
    .A2(net259),
    .A1(_10557_));
 sg13g2_nand2_1 _21405_ (.Y(_03804_),
    .A(_03747_),
    .B(net225));
 sg13g2_o21ai_1 _21406_ (.B1(_03804_),
    .Y(_03805_),
    .A1(_10599_),
    .A2(_03803_));
 sg13g2_o21ai_1 _21407_ (.B1(_03805_),
    .Y(_03806_),
    .A1(_03747_),
    .A2(net192));
 sg13g2_a21o_1 _21408_ (.A2(_03806_),
    .A1(net253),
    .B1(_11065_),
    .X(_03807_));
 sg13g2_o21ai_1 _21409_ (.B1(_03807_),
    .Y(_03808_),
    .A1(net253),
    .A2(_03806_));
 sg13g2_a22oi_1 _21410_ (.Y(_03809_),
    .B1(_03808_),
    .B2(_03779_),
    .A2(_03802_),
    .A1(_03736_));
 sg13g2_xnor2_1 _21411_ (.Y(_03810_),
    .A(net232),
    .B(_03809_));
 sg13g2_nor2_1 _21412_ (.A(net29),
    .B(_03810_),
    .Y(_03811_));
 sg13g2_mux2_1 _21413_ (.A0(_03785_),
    .A1(_03786_),
    .S(_03811_),
    .X(_03812_));
 sg13g2_nor2_1 _21414_ (.A(_09294_),
    .B(net434),
    .Y(_03813_));
 sg13g2_nand4_1 _21415_ (.B(net1044),
    .C(net991),
    .A(_10561_),
    .Y(_03814_),
    .D(net1131));
 sg13g2_nor2_1 _21416_ (.A(_03721_),
    .B(_03814_),
    .Y(_03815_));
 sg13g2_buf_1 _21417_ (.A(_03815_),
    .X(_03816_));
 sg13g2_xnor2_1 _21418_ (.Y(_03817_),
    .A(_10513_),
    .B(net30));
 sg13g2_a22oi_1 _21419_ (.Y(_03818_),
    .B1(_03813_),
    .B2(_03817_),
    .A2(net385),
    .A1(net1133));
 sg13g2_a21oi_1 _21420_ (.A1(_03812_),
    .A2(_03818_),
    .Y(_03819_),
    .B1(net485));
 sg13g2_a21o_1 _21421_ (.A2(net417),
    .A1(net542),
    .B1(_03819_),
    .X(_00960_));
 sg13g2_o21ai_1 _21422_ (.B1(_11435_),
    .Y(_03820_),
    .A1(net1132),
    .A2(_03729_));
 sg13g2_nor2_1 _21423_ (.A(_11235_),
    .B(net434),
    .Y(_03821_));
 sg13g2_nand2_1 _21424_ (.Y(_03822_),
    .A(net1130),
    .B(net30));
 sg13g2_mux2_1 _21425_ (.A0(_11235_),
    .A1(_03821_),
    .S(_03822_),
    .X(_03823_));
 sg13g2_nand2b_1 _21426_ (.Y(_03824_),
    .B(net991),
    .A_N(_10523_));
 sg13g2_a21oi_1 _21427_ (.A1(_11231_),
    .A2(_11232_),
    .Y(_03825_),
    .B1(_11233_));
 sg13g2_o21ai_1 _21428_ (.B1(_03825_),
    .Y(_03826_),
    .A1(_03770_),
    .A2(_03824_));
 sg13g2_nor2_1 _21429_ (.A(net199),
    .B(_10523_),
    .Y(_03827_));
 sg13g2_nand2_1 _21430_ (.Y(_03828_),
    .A(_10560_),
    .B(_03771_));
 sg13g2_a22oi_1 _21431_ (.Y(_03829_),
    .B1(_03827_),
    .B2(_03828_),
    .A2(_03826_),
    .A1(net489));
 sg13g2_buf_1 _21432_ (.A(_03829_),
    .X(_03830_));
 sg13g2_xnor2_1 _21433_ (.Y(_03831_),
    .A(net252),
    .B(_03830_));
 sg13g2_nor2_1 _21434_ (.A(net29),
    .B(_03831_),
    .Y(_03832_));
 sg13g2_nand2_1 _21435_ (.Y(_03833_),
    .A(net1133),
    .B(net489));
 sg13g2_xnor2_1 _21436_ (.Y(_03834_),
    .A(_03832_),
    .B(_03833_));
 sg13g2_a221oi_1 _21437_ (.B2(net32),
    .C1(net385),
    .B1(_03834_),
    .A1(net1034),
    .Y(_03835_),
    .A2(_03823_));
 sg13g2_nand2_1 _21438_ (.Y(_03836_),
    .A(net890),
    .B(net417));
 sg13g2_o21ai_1 _21439_ (.B1(_03836_),
    .Y(_00961_),
    .A1(_03820_),
    .A2(_03835_));
 sg13g2_nand2_1 _21440_ (.Y(_03837_),
    .A(net252),
    .B(_03830_));
 sg13g2_o21ai_1 _21441_ (.B1(_03833_),
    .Y(_03838_),
    .A1(net252),
    .A2(_03830_));
 sg13g2_nand2_1 _21442_ (.Y(_03839_),
    .A(_03837_),
    .B(_03838_));
 sg13g2_xnor2_1 _21443_ (.Y(_03840_),
    .A(_11776_),
    .B(_03839_));
 sg13g2_nor2_1 _21444_ (.A(net27),
    .B(_03840_),
    .Y(_03841_));
 sg13g2_nor2_1 _21445_ (.A(_10377_),
    .B(net568),
    .Y(_03842_));
 sg13g2_xnor2_1 _21446_ (.Y(_03843_),
    .A(_03841_),
    .B(_03842_));
 sg13g2_a21oi_1 _21447_ (.A1(_09167_),
    .A2(net486),
    .Y(_03844_),
    .B1(_11458_));
 sg13g2_nand2_1 _21448_ (.Y(_03845_),
    .A(net32),
    .B(_03844_));
 sg13g2_nor2_1 _21449_ (.A(_10377_),
    .B(net434),
    .Y(_03846_));
 sg13g2_nor4_1 _21450_ (.A(_10513_),
    .B(_11235_),
    .C(_03721_),
    .D(_03814_),
    .Y(_03847_));
 sg13g2_mux2_1 _21451_ (.A0(_03846_),
    .A1(_10377_),
    .S(_03847_),
    .X(_03848_));
 sg13g2_a221oi_1 _21452_ (.B2(net1034),
    .C1(net486),
    .B1(_03848_),
    .A1(net1136),
    .Y(_03849_),
    .A2(net385));
 sg13g2_nand2b_1 _21453_ (.Y(_03850_),
    .B(_03844_),
    .A_N(_03849_));
 sg13g2_o21ai_1 _21454_ (.B1(_03850_),
    .Y(_00962_),
    .A1(_03843_),
    .A2(_03845_));
 sg13g2_nand2_1 _21455_ (.Y(_03851_),
    .A(_11435_),
    .B(net385));
 sg13g2_and4_1 _21456_ (.A(_10455_),
    .B(net1133),
    .C(net1132),
    .D(net30),
    .X(_03852_));
 sg13g2_xor2_1 _21457_ (.B(_03852_),
    .A(net1136),
    .X(_03853_));
 sg13g2_nor2_1 _21458_ (.A(net229),
    .B(_11243_),
    .Y(_03854_));
 sg13g2_and2_1 _21459_ (.A(net229),
    .B(_11243_),
    .X(_03855_));
 sg13g2_nor3_1 _21460_ (.A(net29),
    .B(_03854_),
    .C(_03855_),
    .Y(_03856_));
 sg13g2_nand2_1 _21461_ (.Y(_03857_),
    .A(net1136),
    .B(net489));
 sg13g2_xnor2_1 _21462_ (.Y(_03858_),
    .A(_03856_),
    .B(_03857_));
 sg13g2_nor2_1 _21463_ (.A(_10920_),
    .B(_11433_),
    .Y(_03859_));
 sg13g2_a221oi_1 _21464_ (.B2(_03767_),
    .C1(_03859_),
    .B1(_03858_),
    .A1(_03762_),
    .Y(_03860_),
    .A2(_03853_));
 sg13g2_nor2_1 _21465_ (.A(_10233_),
    .B(_03851_),
    .Y(_03861_));
 sg13g2_a21oi_1 _21466_ (.A1(_03851_),
    .A2(_03860_),
    .Y(_00963_),
    .B1(_03861_));
 sg13g2_nand3_1 _21467_ (.B(net1132),
    .C(net1136),
    .A(net1133),
    .Y(_03862_));
 sg13g2_nor2_1 _21468_ (.A(_03822_),
    .B(_03862_),
    .Y(_03863_));
 sg13g2_xnor2_1 _21469_ (.Y(_03864_),
    .A(_11259_),
    .B(_03863_));
 sg13g2_nand2_1 _21470_ (.Y(_03865_),
    .A(_03696_),
    .B(_03765_));
 sg13g2_nand2_1 _21471_ (.Y(_03866_),
    .A(net229),
    .B(_11243_));
 sg13g2_a21oi_1 _21472_ (.A1(_03866_),
    .A2(_03857_),
    .Y(_03867_),
    .B1(_03854_));
 sg13g2_xnor2_1 _21473_ (.Y(_03868_),
    .A(net208),
    .B(_03867_));
 sg13g2_nor2_1 _21474_ (.A(_03698_),
    .B(_03868_),
    .Y(_03869_));
 sg13g2_xor2_1 _21475_ (.B(_03869_),
    .A(_11251_),
    .X(_03870_));
 sg13g2_a22oi_1 _21476_ (.Y(_03871_),
    .B1(net377),
    .B2(net1052),
    .A2(net486),
    .A1(_10234_));
 sg13g2_o21ai_1 _21477_ (.B1(_03871_),
    .Y(_03872_),
    .A1(_03865_),
    .A2(_03870_));
 sg13g2_a21o_1 _21478_ (.A2(_03864_),
    .A1(_03762_),
    .B1(_03872_),
    .X(_00964_));
 sg13g2_nand2_1 _21479_ (.Y(_03873_),
    .A(_10366_),
    .B(_11243_));
 sg13g2_xnor2_1 _21480_ (.Y(_03874_),
    .A(net255),
    .B(_03873_));
 sg13g2_nand3_1 _21481_ (.B(_11250_),
    .C(_11265_),
    .A(_11249_),
    .Y(_03875_));
 sg13g2_buf_1 _21482_ (.A(_03875_),
    .X(_03876_));
 sg13g2_o21ai_1 _21483_ (.B1(_03873_),
    .Y(_03877_),
    .A1(net568),
    .A2(_03876_));
 sg13g2_nor2_1 _21484_ (.A(net1052),
    .B(net255),
    .Y(_03878_));
 sg13g2_nand2_1 _21485_ (.Y(_03879_),
    .A(_03876_),
    .B(_03873_));
 sg13g2_nor3_1 _21486_ (.A(net1052),
    .B(net230),
    .C(_03879_),
    .Y(_03880_));
 sg13g2_a221oi_1 _21487_ (.B2(_03878_),
    .C1(_03880_),
    .B1(_03877_),
    .A1(net568),
    .Y(_03881_),
    .A2(_03874_));
 sg13g2_xnor2_1 _21488_ (.Y(_03882_),
    .A(net255),
    .B(_03879_));
 sg13g2_and2_1 _21489_ (.A(net1052),
    .B(_03779_),
    .X(_03883_));
 sg13g2_o21ai_1 _21490_ (.B1(_03883_),
    .Y(_03884_),
    .A1(net29),
    .A2(_03882_));
 sg13g2_o21ai_1 _21491_ (.B1(_03884_),
    .Y(_03885_),
    .A1(net27),
    .A2(_03881_));
 sg13g2_nor2_1 _21492_ (.A(net1052),
    .B(_03742_),
    .Y(_03886_));
 sg13g2_and2_1 _21493_ (.A(net1052),
    .B(_03813_),
    .X(_03887_));
 sg13g2_nor3_1 _21494_ (.A(_10513_),
    .B(_11259_),
    .C(_03862_),
    .Y(_03888_));
 sg13g2_nand2_1 _21495_ (.Y(_03889_),
    .A(net30),
    .B(_03888_));
 sg13g2_mux2_1 _21496_ (.A0(_03886_),
    .A1(_03887_),
    .S(_03889_),
    .X(_03890_));
 sg13g2_a221oi_1 _21497_ (.B2(_03885_),
    .C1(_03890_),
    .B1(net32),
    .A1(net646),
    .Y(_03891_),
    .A2(_11626_));
 sg13g2_o21ai_1 _21498_ (.B1(_11435_),
    .Y(_03892_),
    .A1(net1045),
    .A2(_03729_));
 sg13g2_nand2_1 _21499_ (.Y(_03893_),
    .A(net999),
    .B(net417));
 sg13g2_o21ai_1 _21500_ (.B1(_03893_),
    .Y(_00965_),
    .A1(_03891_),
    .A2(_03892_));
 sg13g2_and2_1 _21501_ (.A(net1052),
    .B(_03888_),
    .X(_03894_));
 sg13g2_buf_1 _21502_ (.A(_03894_),
    .X(_03895_));
 sg13g2_nand2_1 _21503_ (.Y(_03896_),
    .A(net30),
    .B(_03895_));
 sg13g2_xnor2_1 _21504_ (.Y(_03897_),
    .A(net1045),
    .B(_03896_));
 sg13g2_nand2_1 _21505_ (.Y(_03898_),
    .A(net1045),
    .B(net416));
 sg13g2_nand3b_1 _21506_ (.B(_03876_),
    .C(_03873_),
    .Y(_03899_),
    .A_N(net1052));
 sg13g2_buf_1 _21507_ (.A(_03899_),
    .X(_03900_));
 sg13g2_a21oi_1 _21508_ (.A1(_10366_),
    .A2(_11243_),
    .Y(_03901_),
    .B1(net255));
 sg13g2_nand3_1 _21509_ (.B(net255),
    .C(_11243_),
    .A(_10366_),
    .Y(_03902_));
 sg13g2_a221oi_1 _21510_ (.B2(net568),
    .C1(_03878_),
    .B1(_03902_),
    .A1(_03876_),
    .Y(_03903_),
    .A2(_03901_));
 sg13g2_buf_2 _21511_ (.A(_03903_),
    .X(_03904_));
 sg13g2_a21o_1 _21512_ (.A2(_03904_),
    .A1(_03900_),
    .B1(net201),
    .X(_03905_));
 sg13g2_nand3_1 _21513_ (.B(_03900_),
    .C(_03904_),
    .A(net201),
    .Y(_03906_));
 sg13g2_a21oi_1 _21514_ (.A1(_03905_),
    .A2(_03906_),
    .Y(_03907_),
    .B1(net29));
 sg13g2_xor2_1 _21515_ (.B(_03907_),
    .A(_03898_),
    .X(_03908_));
 sg13g2_a22oi_1 _21516_ (.Y(_03909_),
    .B1(net377),
    .B2(net1134),
    .A2(net486),
    .A1(net1135));
 sg13g2_o21ai_1 _21517_ (.B1(_03909_),
    .Y(_03910_),
    .A1(_03865_),
    .A2(_03908_));
 sg13g2_a21o_1 _21518_ (.A2(_03897_),
    .A1(_03762_),
    .B1(_03910_),
    .X(_00966_));
 sg13g2_and2_1 _21519_ (.A(_11244_),
    .B(_11266_),
    .X(_03911_));
 sg13g2_buf_1 _21520_ (.A(_03911_),
    .X(_03912_));
 sg13g2_xnor2_1 _21521_ (.Y(_03913_),
    .A(net177),
    .B(_03912_));
 sg13g2_nor2_1 _21522_ (.A(_03698_),
    .B(_03913_),
    .Y(_03914_));
 sg13g2_nand2_1 _21523_ (.Y(_03915_),
    .A(net1134),
    .B(net489));
 sg13g2_xnor2_1 _21524_ (.Y(_03916_),
    .A(_03914_),
    .B(_03915_));
 sg13g2_nor2_1 _21525_ (.A(net1134),
    .B(_03742_),
    .Y(_03917_));
 sg13g2_nor2_1 _21526_ (.A(_11267_),
    .B(_03742_),
    .Y(_03918_));
 sg13g2_nand3_1 _21527_ (.B(net30),
    .C(_03895_),
    .A(net1045),
    .Y(_03919_));
 sg13g2_mux2_1 _21528_ (.A0(_03917_),
    .A1(_03918_),
    .S(_03919_),
    .X(_03920_));
 sg13g2_a221oi_1 _21529_ (.B2(_03916_),
    .C1(_03920_),
    .B1(_03696_),
    .A1(net1037),
    .Y(_03921_),
    .A2(net385));
 sg13g2_nand2_1 _21530_ (.Y(_03922_),
    .A(net537),
    .B(_03726_));
 sg13g2_o21ai_1 _21531_ (.B1(_03922_),
    .Y(_00967_),
    .A1(net485),
    .A2(_03921_));
 sg13g2_nand2_1 _21532_ (.Y(_03923_),
    .A(net1037),
    .B(net416));
 sg13g2_o21ai_1 _21533_ (.B1(_03923_),
    .Y(_03924_),
    .A1(_11397_),
    .A2(_11411_));
 sg13g2_nand3_1 _21534_ (.B(_03900_),
    .C(_03904_),
    .A(_11577_),
    .Y(_03925_));
 sg13g2_nor2_1 _21535_ (.A(net201),
    .B(_03915_),
    .Y(_03926_));
 sg13g2_nand3_1 _21536_ (.B(_03904_),
    .C(_03926_),
    .A(_03900_),
    .Y(_03927_));
 sg13g2_o21ai_1 _21537_ (.B1(_10316_),
    .Y(_03928_),
    .A1(_10338_),
    .A2(net150));
 sg13g2_nor2_1 _21538_ (.A(_09291_),
    .B(_03928_),
    .Y(_03929_));
 sg13g2_nand3_1 _21539_ (.B(_03904_),
    .C(_03929_),
    .A(_03900_),
    .Y(_03930_));
 sg13g2_nor2_1 _21540_ (.A(net177),
    .B(_03915_),
    .Y(_03931_));
 sg13g2_nor3_1 _21541_ (.A(net568),
    .B(net201),
    .C(_03928_),
    .Y(_03932_));
 sg13g2_nor2_1 _21542_ (.A(_03931_),
    .B(_03932_),
    .Y(_03933_));
 sg13g2_nand4_1 _21543_ (.B(_03927_),
    .C(_03930_),
    .A(_03925_),
    .Y(_03934_),
    .D(_03933_));
 sg13g2_xnor2_1 _21544_ (.Y(_03935_),
    .A(net206),
    .B(_03934_));
 sg13g2_mux2_1 _21545_ (.A0(_03923_),
    .A1(_03924_),
    .S(_03935_),
    .X(_03936_));
 sg13g2_and2_1 _21546_ (.A(net1045),
    .B(_10338_),
    .X(_03937_));
 sg13g2_nand3_1 _21547_ (.B(_03895_),
    .C(_03937_),
    .A(net30),
    .Y(_03938_));
 sg13g2_xnor2_1 _21548_ (.Y(_03939_),
    .A(net1037),
    .B(_03938_));
 sg13g2_a22oi_1 _21549_ (.Y(_03940_),
    .B1(net377),
    .B2(net1036),
    .A2(net486),
    .A1(net628));
 sg13g2_and2_1 _21550_ (.A(net1037),
    .B(net416),
    .X(_03941_));
 sg13g2_nand3_1 _21551_ (.B(_03767_),
    .C(_03941_),
    .A(net27),
    .Y(_03942_));
 sg13g2_nand2_1 _21552_ (.Y(_03943_),
    .A(_03940_),
    .B(_03942_));
 sg13g2_a21oi_1 _21553_ (.A1(_03762_),
    .A2(_03939_),
    .Y(_03944_),
    .B1(_03943_));
 sg13g2_o21ai_1 _21554_ (.B1(_03944_),
    .Y(_00968_),
    .A1(_03865_),
    .A2(_03936_));
 sg13g2_and3_1 _21555_ (.X(_03945_),
    .A(net1037),
    .B(net435),
    .C(_03937_));
 sg13g2_nand3_1 _21556_ (.B(_03895_),
    .C(_03945_),
    .A(net30),
    .Y(_03946_));
 sg13g2_xnor2_1 _21557_ (.Y(_03947_),
    .A(net1036),
    .B(_03946_));
 sg13g2_a22oi_1 _21558_ (.Y(_03948_),
    .B1(_03762_),
    .B2(_03947_),
    .A2(_03726_),
    .A1(net618));
 sg13g2_a21oi_1 _21559_ (.A1(net177),
    .A2(_03912_),
    .Y(_03949_),
    .B1(_11403_));
 sg13g2_o21ai_1 _21560_ (.B1(net206),
    .Y(_03950_),
    .A1(net177),
    .A2(_03912_));
 sg13g2_nor2_1 _21561_ (.A(_11422_),
    .B(_03912_),
    .Y(_03951_));
 sg13g2_a221oi_1 _21562_ (.B2(_03941_),
    .C1(_03951_),
    .B1(_03950_),
    .A1(net416),
    .Y(_03952_),
    .A2(_03949_));
 sg13g2_xnor2_1 _21563_ (.Y(_03953_),
    .A(net179),
    .B(_03952_));
 sg13g2_nand2_1 _21564_ (.Y(_03954_),
    .A(net1036),
    .B(net416));
 sg13g2_nand3_1 _21565_ (.B(_03767_),
    .C(_03954_),
    .A(_03851_),
    .Y(_03955_));
 sg13g2_or3_1 _21566_ (.A(net27),
    .B(_03953_),
    .C(_03955_),
    .X(_03956_));
 sg13g2_nor3_1 _21567_ (.A(net377),
    .B(_03865_),
    .C(_03954_),
    .Y(_03957_));
 sg13g2_o21ai_1 _21568_ (.B1(_03957_),
    .Y(_03958_),
    .A1(net27),
    .A2(_03953_));
 sg13g2_nand2_1 _21569_ (.Y(_03959_),
    .A(net1126),
    .B(_03731_));
 sg13g2_nand4_1 _21570_ (.B(_03956_),
    .C(_03958_),
    .A(_03948_),
    .Y(_00969_),
    .D(_03959_));
 sg13g2_inv_1 _21571_ (.Y(_03960_),
    .A(\cpu.ex.r_mult[31] ));
 sg13g2_nand2_1 _21572_ (.Y(_03961_),
    .A(net687),
    .B(net486));
 sg13g2_nand4_1 _21573_ (.B(_03816_),
    .C(_03895_),
    .A(net1036),
    .Y(_03962_),
    .D(_03945_));
 sg13g2_xnor2_1 _21574_ (.Y(_03963_),
    .A(net1126),
    .B(_03962_));
 sg13g2_o21ai_1 _21575_ (.B1(_03765_),
    .Y(_03964_),
    .A1(_09294_),
    .A2(_03963_));
 sg13g2_and3_1 _21576_ (.X(_03965_),
    .A(_10662_),
    .B(net416),
    .C(net32));
 sg13g2_nand2_1 _21577_ (.Y(_03966_),
    .A(_03705_),
    .B(_11398_));
 sg13g2_a21oi_1 _21578_ (.A1(net1036),
    .A2(_11394_),
    .Y(_03967_),
    .B1(net27));
 sg13g2_o21ai_1 _21579_ (.B1(_03967_),
    .Y(_03968_),
    .A1(_03952_),
    .A2(_03966_));
 sg13g2_nand3_1 _21580_ (.B(_03851_),
    .C(_03961_),
    .A(_11445_),
    .Y(_03969_));
 sg13g2_a21oi_1 _21581_ (.A1(_03965_),
    .A2(_03968_),
    .Y(_03970_),
    .B1(_03969_));
 sg13g2_a221oi_1 _21582_ (.B2(_03964_),
    .C1(_03970_),
    .B1(_03961_),
    .A1(_03960_),
    .Y(_00970_),
    .A2(net377));
 sg13g2_and2_1 _21583_ (.A(net358),
    .B(_11012_),
    .X(_03971_));
 sg13g2_buf_1 _21584_ (.A(_03971_),
    .X(_03972_));
 sg13g2_nor2b_1 _21585_ (.A(_11619_),
    .B_N(net1161),
    .Y(_03973_));
 sg13g2_mux2_1 _21586_ (.A0(_08353_),
    .A1(_03973_),
    .S(_12036_),
    .X(_03974_));
 sg13g2_nand3_1 _21587_ (.B(net247),
    .C(_03974_),
    .A(net814),
    .Y(_03975_));
 sg13g2_buf_1 _21588_ (.A(_03975_),
    .X(_03976_));
 sg13g2_buf_1 _21589_ (.A(_03976_),
    .X(_03977_));
 sg13g2_nand2b_1 _21590_ (.Y(_03978_),
    .B(_11627_),
    .A_N(_11626_));
 sg13g2_buf_1 _21591_ (.A(_03978_),
    .X(_03979_));
 sg13g2_and2_1 _21592_ (.A(net1156),
    .B(_11455_),
    .X(_03980_));
 sg13g2_buf_1 _21593_ (.A(_03980_),
    .X(_03981_));
 sg13g2_o21ai_1 _21594_ (.B1(net172),
    .Y(_03982_),
    .A1(net248),
    .A2(_03981_));
 sg13g2_or3_1 _21595_ (.A(_11495_),
    .B(_11497_),
    .C(_11500_),
    .X(_03983_));
 sg13g2_buf_2 _21596_ (.A(_03983_),
    .X(_03984_));
 sg13g2_buf_1 _21597_ (.A(_03984_),
    .X(_03985_));
 sg13g2_nand2_1 _21598_ (.Y(_03986_),
    .A(net215),
    .B(net214));
 sg13g2_a21oi_1 _21599_ (.A1(_03982_),
    .A2(_03986_),
    .Y(_03987_),
    .B1(net205));
 sg13g2_nand2_2 _21600_ (.Y(_03988_),
    .A(net231),
    .B(net254));
 sg13g2_nor3_1 _21601_ (.A(net248),
    .B(net228),
    .C(_03988_),
    .Y(_03989_));
 sg13g2_buf_2 _21602_ (.A(_03989_),
    .X(_03990_));
 sg13g2_nor2_1 _21603_ (.A(_11415_),
    .B(net254),
    .Y(_03991_));
 sg13g2_nand2_1 _21604_ (.Y(_03992_),
    .A(_11413_),
    .B(_03991_));
 sg13g2_nor2_1 _21605_ (.A(net227),
    .B(_03992_),
    .Y(_03993_));
 sg13g2_buf_1 _21606_ (.A(_03993_),
    .X(_03994_));
 sg13g2_buf_1 _21607_ (.A(net204),
    .X(_03995_));
 sg13g2_buf_8 _21608_ (.A(_11585_),
    .X(_03996_));
 sg13g2_nor3_1 _21609_ (.A(_03996_),
    .B(net200),
    .C(_03992_),
    .Y(_03997_));
 sg13g2_a221oi_1 _21610_ (.B2(net171),
    .C1(_03997_),
    .B1(net142),
    .A1(net109),
    .Y(_03998_),
    .A2(_03990_));
 sg13g2_nand3_1 _21611_ (.B(_10897_),
    .C(_10898_),
    .A(_10896_),
    .Y(_03999_));
 sg13g2_buf_1 _21612_ (.A(_03999_),
    .X(_04000_));
 sg13g2_buf_1 _21613_ (.A(_04000_),
    .X(_04001_));
 sg13g2_nor3_1 _21614_ (.A(net248),
    .B(net225),
    .C(_10598_),
    .Y(_04002_));
 sg13g2_buf_1 _21615_ (.A(_04002_),
    .X(_04003_));
 sg13g2_buf_1 _21616_ (.A(_04003_),
    .X(_04004_));
 sg13g2_nand2_1 _21617_ (.Y(_04005_),
    .A(net245),
    .B(net141));
 sg13g2_buf_1 _21618_ (.A(net300),
    .X(_04006_));
 sg13g2_nand2_1 _21619_ (.Y(_04007_),
    .A(net225),
    .B(_11662_));
 sg13g2_nor3_1 _21620_ (.A(_11413_),
    .B(net227),
    .C(_04007_),
    .Y(_04008_));
 sg13g2_buf_1 _21621_ (.A(_04008_),
    .X(_04009_));
 sg13g2_buf_1 _21622_ (.A(net140),
    .X(_04010_));
 sg13g2_nor3_1 _21623_ (.A(_11187_),
    .B(net228),
    .C(_04007_),
    .Y(_04011_));
 sg13g2_buf_1 _21624_ (.A(_04011_),
    .X(_04012_));
 sg13g2_buf_1 _21625_ (.A(net139),
    .X(_04013_));
 sg13g2_buf_1 _21626_ (.A(_11541_),
    .X(_04014_));
 sg13g2_a22oi_1 _21627_ (.Y(_04015_),
    .B1(net105),
    .B2(net169),
    .A2(net106),
    .A1(net244));
 sg13g2_nor3_2 _21628_ (.A(net258),
    .B(net228),
    .C(_03988_),
    .Y(_04016_));
 sg13g2_nor3_2 _21629_ (.A(_03734_),
    .B(net193),
    .C(_03988_),
    .Y(_04017_));
 sg13g2_o21ai_1 _21630_ (.B1(_11070_),
    .Y(_04018_),
    .A1(net778),
    .A2(_10726_));
 sg13g2_o21ai_1 _21631_ (.B1(_04018_),
    .Y(_04019_),
    .A1(_11073_),
    .A2(_10838_));
 sg13g2_buf_1 _21632_ (.A(_04019_),
    .X(_04020_));
 sg13g2_nor3_1 _21633_ (.A(_11413_),
    .B(_11417_),
    .C(net227),
    .Y(_04021_));
 sg13g2_buf_1 _21634_ (.A(_04021_),
    .X(_04022_));
 sg13g2_and2_1 _21635_ (.A(net191),
    .B(net168),
    .X(_04023_));
 sg13g2_a221oi_1 _21636_ (.B2(_11455_),
    .C1(_04023_),
    .B1(_04017_),
    .A1(net176),
    .Y(_04024_),
    .A2(_04016_));
 sg13g2_buf_1 _21637_ (.A(_10872_),
    .X(_04025_));
 sg13g2_nor2_1 _21638_ (.A(net248),
    .B(net227),
    .Y(_04026_));
 sg13g2_and2_1 _21639_ (.A(_03991_),
    .B(_04026_),
    .X(_04027_));
 sg13g2_buf_1 _21640_ (.A(_04027_),
    .X(_04028_));
 sg13g2_buf_1 _21641_ (.A(_04028_),
    .X(_04029_));
 sg13g2_nor3_1 _21642_ (.A(net258),
    .B(net193),
    .C(_03988_),
    .Y(_04030_));
 sg13g2_a22oi_1 _21643_ (.Y(_04031_),
    .B1(_04030_),
    .B2(_03981_),
    .A2(net104),
    .A1(net243));
 sg13g2_nor3_1 _21644_ (.A(_11413_),
    .B(_11419_),
    .C(_04007_),
    .Y(_04032_));
 sg13g2_buf_1 _21645_ (.A(_04032_),
    .X(_04033_));
 sg13g2_nand2b_1 _21646_ (.Y(_04034_),
    .B(net138),
    .A_N(net256));
 sg13g2_nor3_1 _21647_ (.A(_11187_),
    .B(_11475_),
    .C(_04007_),
    .Y(_04035_));
 sg13g2_buf_2 _21648_ (.A(_04035_),
    .X(_04036_));
 sg13g2_nand2_1 _21649_ (.Y(_04037_),
    .A(_11472_),
    .B(_04036_));
 sg13g2_and4_1 _21650_ (.A(_04024_),
    .B(_04031_),
    .C(_04034_),
    .D(_04037_),
    .X(_04038_));
 sg13g2_nand4_1 _21651_ (.B(_04005_),
    .C(_04015_),
    .A(_03998_),
    .Y(_04039_),
    .D(_04038_));
 sg13g2_nor3_1 _21652_ (.A(_11187_),
    .B(net205),
    .C(net228),
    .Y(_04040_));
 sg13g2_buf_1 _21653_ (.A(_04040_),
    .X(_04041_));
 sg13g2_buf_1 _21654_ (.A(_04041_),
    .X(_04042_));
 sg13g2_buf_1 _21655_ (.A(_04042_),
    .X(_04043_));
 sg13g2_nor2_1 _21656_ (.A(net1156),
    .B(net1146),
    .Y(_04044_));
 sg13g2_buf_1 _21657_ (.A(_04044_),
    .X(_04045_));
 sg13g2_a21oi_1 _21658_ (.A1(_11510_),
    .A2(net87),
    .Y(_04046_),
    .B1(net872));
 sg13g2_o21ai_1 _21659_ (.B1(_04046_),
    .Y(_04047_),
    .A1(_03987_),
    .A2(_04039_));
 sg13g2_nand4_1 _21660_ (.B(_10621_),
    .C(_10985_),
    .A(_08300_),
    .Y(_04048_),
    .D(_11006_));
 sg13g2_nor3_1 _21661_ (.A(_08359_),
    .B(_08415_),
    .C(_04048_),
    .Y(_04049_));
 sg13g2_a221oi_1 _21662_ (.B2(_11015_),
    .C1(_04049_),
    .B1(net347),
    .A1(net778),
    .Y(_04050_),
    .A2(_11486_));
 sg13g2_buf_2 _21663_ (.A(_04050_),
    .X(_04051_));
 sg13g2_nor2b_1 _21664_ (.A(_04051_),
    .B_N(_09844_),
    .Y(_04052_));
 sg13g2_buf_1 _21665_ (.A(_11629_),
    .X(_04053_));
 sg13g2_a221oi_1 _21666_ (.B2(_04052_),
    .C1(net213),
    .B1(net87),
    .A1(net1073),
    .Y(_04054_),
    .A2(_10360_));
 sg13g2_inv_1 _21667_ (.Y(_04055_),
    .A(net1155));
 sg13g2_buf_1 _21668_ (.A(_04055_),
    .X(_04056_));
 sg13g2_nor2_1 _21669_ (.A(net1072),
    .B(_11484_),
    .Y(_04057_));
 sg13g2_a21oi_1 _21670_ (.A1(net871),
    .A2(_11484_),
    .Y(_04058_),
    .B1(_04057_));
 sg13g2_nand2_1 _21671_ (.Y(_04059_),
    .A(net172),
    .B(_11482_));
 sg13g2_o21ai_1 _21672_ (.B1(_04059_),
    .Y(_04060_),
    .A1(net1063),
    .A2(_04058_));
 sg13g2_xnor2_1 _21673_ (.Y(_04061_),
    .A(net172),
    .B(_11482_));
 sg13g2_nor4_1 _21674_ (.A(net1157),
    .B(net1155),
    .C(net1145),
    .D(_09844_),
    .Y(_04062_));
 sg13g2_nand2_1 _21675_ (.Y(_04063_),
    .A(net872),
    .B(_04062_));
 sg13g2_nor4_2 _21676_ (.A(_08242_),
    .B(_09085_),
    .C(_09092_),
    .Y(_04064_),
    .D(_09813_));
 sg13g2_nor2b_1 _21677_ (.A(_04063_),
    .B_N(_04064_),
    .Y(_04065_));
 sg13g2_buf_1 _21678_ (.A(_04065_),
    .X(_04066_));
 sg13g2_nor3_1 _21679_ (.A(_09085_),
    .B(_09813_),
    .C(net607),
    .Y(_04067_));
 sg13g2_a21oi_1 _21680_ (.A1(_04051_),
    .A2(_04061_),
    .Y(_04068_),
    .B1(_04067_));
 sg13g2_nor2_1 _21681_ (.A(_08242_),
    .B(_04051_),
    .Y(_04069_));
 sg13g2_a21oi_1 _21682_ (.A1(_04051_),
    .A2(_04067_),
    .Y(_04070_),
    .B1(_04069_));
 sg13g2_nor2_1 _21683_ (.A(_04061_),
    .B(_04070_),
    .Y(_04071_));
 sg13g2_or3_1 _21684_ (.A(_09085_),
    .B(_09813_),
    .C(net607),
    .X(_04072_));
 sg13g2_buf_1 _21685_ (.A(_04072_),
    .X(_04073_));
 sg13g2_o21ai_1 _21686_ (.B1(net215),
    .Y(_04074_),
    .A1(_04051_),
    .A2(_04073_));
 sg13g2_a22oi_1 _21687_ (.Y(_04075_),
    .B1(_04074_),
    .B2(_04061_),
    .A2(_04071_),
    .A1(net215));
 sg13g2_o21ai_1 _21688_ (.B1(_04075_),
    .Y(_04076_),
    .A1(net1091),
    .A2(_04068_));
 sg13g2_nand4_1 _21689_ (.B(_04054_),
    .C(_04060_),
    .A(_04047_),
    .Y(_04077_),
    .D(_04076_));
 sg13g2_o21ai_1 _21690_ (.B1(_04077_),
    .Y(_04078_),
    .A1(net246),
    .A2(\cpu.ex.c_mult[1] ));
 sg13g2_and4_1 _21691_ (.A(net1161),
    .B(net814),
    .C(net247),
    .D(_12037_),
    .X(_04079_));
 sg13g2_buf_1 _21692_ (.A(_04079_),
    .X(_04080_));
 sg13g2_nand3_1 _21693_ (.B(net350),
    .C(_12024_),
    .A(_09110_),
    .Y(_04081_));
 sg13g2_o21ai_1 _21694_ (.B1(_04081_),
    .Y(_04082_),
    .A1(net350),
    .A2(_12024_));
 sg13g2_nor3_1 _21695_ (.A(_09110_),
    .B(_09160_),
    .C(_11624_),
    .Y(_04083_));
 sg13g2_a221oi_1 _21696_ (.B2(net350),
    .C1(_09258_),
    .B1(_04083_),
    .A1(_08353_),
    .Y(_04084_),
    .A2(_04082_));
 sg13g2_nand2_1 _21697_ (.Y(_04085_),
    .A(_03976_),
    .B(_04084_));
 sg13g2_nor2_1 _21698_ (.A(net81),
    .B(_04085_),
    .Y(_04086_));
 sg13g2_buf_1 _21699_ (.A(_04086_),
    .X(_04087_));
 sg13g2_buf_1 _21700_ (.A(_04087_),
    .X(_04088_));
 sg13g2_a22oi_1 _21701_ (.Y(_04089_),
    .B1(net31),
    .B2(net819),
    .A2(net81),
    .A1(_10563_));
 sg13g2_o21ai_1 _21702_ (.B1(_04089_),
    .Y(_00971_),
    .A1(net71),
    .A2(_04078_));
 sg13g2_buf_1 _21703_ (.A(net213),
    .X(_04090_));
 sg13g2_nand3_1 _21704_ (.B(_04062_),
    .C(_04064_),
    .A(net872),
    .Y(_04091_));
 sg13g2_buf_1 _21705_ (.A(_04091_),
    .X(_04092_));
 sg13g2_nand2_1 _21706_ (.Y(_04093_),
    .A(net223),
    .B(_11571_));
 sg13g2_nand2_1 _21707_ (.Y(_04094_),
    .A(net261),
    .B(net300));
 sg13g2_nand2_1 _21708_ (.Y(_04095_),
    .A(_04093_),
    .B(_04094_));
 sg13g2_nand2_1 _21709_ (.Y(_04096_),
    .A(net259),
    .B(net203));
 sg13g2_nor2_1 _21710_ (.A(net302),
    .B(net203),
    .Y(_04097_));
 sg13g2_or3_1 _21711_ (.A(_04097_),
    .B(_11484_),
    .C(_11490_),
    .X(_04098_));
 sg13g2_buf_1 _21712_ (.A(_04098_),
    .X(_04099_));
 sg13g2_nand3_1 _21713_ (.B(_04096_),
    .C(_04099_),
    .A(net191),
    .Y(_04100_));
 sg13g2_or2_1 _21714_ (.X(_04101_),
    .B(net256),
    .A(_11522_));
 sg13g2_nand2_1 _21715_ (.Y(_04102_),
    .A(_11493_),
    .B(net257));
 sg13g2_nand2_1 _21716_ (.Y(_04103_),
    .A(net232),
    .B(_04102_));
 sg13g2_a21oi_1 _21717_ (.A1(_04096_),
    .A2(_04099_),
    .Y(_04104_),
    .B1(net191));
 sg13g2_a221oi_1 _21718_ (.B2(_04103_),
    .C1(_04104_),
    .B1(_04101_),
    .A1(net225),
    .Y(_04105_),
    .A2(_04100_));
 sg13g2_nor2b_1 _21719_ (.A(_04105_),
    .B_N(_11553_),
    .Y(_04106_));
 sg13g2_nor2_1 _21720_ (.A(net252),
    .B(_04014_),
    .Y(_04107_));
 sg13g2_a21oi_1 _21721_ (.A1(_11542_),
    .A2(_04106_),
    .Y(_04108_),
    .B1(_04107_));
 sg13g2_xor2_1 _21722_ (.B(_04108_),
    .A(_04095_),
    .X(_04109_));
 sg13g2_nand2_1 _21723_ (.Y(_04110_),
    .A(_09813_),
    .B(_04109_));
 sg13g2_buf_1 _21724_ (.A(net138),
    .X(_04111_));
 sg13g2_nand2_1 _21725_ (.Y(_04112_),
    .A(net244),
    .B(_04111_));
 sg13g2_nor3_2 _21726_ (.A(_11187_),
    .B(net205),
    .C(net193),
    .Y(_04113_));
 sg13g2_a21oi_1 _21727_ (.A1(_11472_),
    .A2(_04113_),
    .Y(_04114_),
    .B1(_04041_));
 sg13g2_a22oi_1 _21728_ (.Y(_04115_),
    .B1(_04036_),
    .B2(_03984_),
    .A2(_04003_),
    .A1(net191));
 sg13g2_nand3_1 _21729_ (.B(_11478_),
    .C(_11480_),
    .A(_11477_),
    .Y(_04116_));
 sg13g2_buf_2 _21730_ (.A(_04116_),
    .X(_04117_));
 sg13g2_and2_1 _21731_ (.A(_04000_),
    .B(net168),
    .X(_04118_));
 sg13g2_a21oi_1 _21732_ (.A1(_04117_),
    .A2(_04028_),
    .Y(_04119_),
    .B1(_04118_));
 sg13g2_nand2_1 _21733_ (.Y(_04120_),
    .A(net301),
    .B(_11503_));
 sg13g2_o21ai_1 _21734_ (.B1(_04120_),
    .Y(_04121_),
    .A1(_11464_),
    .A2(_10983_));
 sg13g2_buf_1 _21735_ (.A(_04121_),
    .X(_04122_));
 sg13g2_nor2_1 _21736_ (.A(net228),
    .B(_03992_),
    .Y(_04123_));
 sg13g2_nor2b_1 _21737_ (.A(net256),
    .B_N(net140),
    .Y(_04124_));
 sg13g2_a21oi_1 _21738_ (.A1(_04122_),
    .A2(_04123_),
    .Y(_04125_),
    .B1(_04124_));
 sg13g2_and4_1 _21739_ (.A(_04114_),
    .B(_04115_),
    .C(_04119_),
    .D(_04125_),
    .X(_04126_));
 sg13g2_nand2_1 _21740_ (.Y(_04127_),
    .A(_11488_),
    .B(_11487_));
 sg13g2_buf_1 _21741_ (.A(_04127_),
    .X(_04128_));
 sg13g2_buf_1 _21742_ (.A(_04128_),
    .X(_04129_));
 sg13g2_a22oi_1 _21743_ (.Y(_04130_),
    .B1(_04013_),
    .B2(net169),
    .A2(net142),
    .A1(net189));
 sg13g2_nand3_1 _21744_ (.B(_04126_),
    .C(_04130_),
    .A(_04112_),
    .Y(_04131_));
 sg13g2_nand2_1 _21745_ (.Y(_04132_),
    .A(_03996_),
    .B(net103));
 sg13g2_nand3_1 _21746_ (.B(_04131_),
    .C(_04132_),
    .A(net1062),
    .Y(_04133_));
 sg13g2_buf_1 _21747_ (.A(net171),
    .X(_04134_));
 sg13g2_nor2_1 _21748_ (.A(_11226_),
    .B(_11662_),
    .Y(_04135_));
 sg13g2_buf_2 _21749_ (.A(_04135_),
    .X(_04136_));
 sg13g2_nand3_1 _21750_ (.B(_04136_),
    .C(net193),
    .A(net248),
    .Y(_04137_));
 sg13g2_buf_1 _21751_ (.A(_04137_),
    .X(_04138_));
 sg13g2_buf_1 _21752_ (.A(_04138_),
    .X(_04139_));
 sg13g2_nor2_2 _21753_ (.A(_11187_),
    .B(net227),
    .Y(_04140_));
 sg13g2_nand2_2 _21754_ (.Y(_04141_),
    .A(_04136_),
    .B(_04140_));
 sg13g2_nand2_1 _21755_ (.Y(_04142_),
    .A(net1156),
    .B(_11455_));
 sg13g2_buf_1 _21756_ (.A(_04142_),
    .X(_04143_));
 sg13g2_a21oi_1 _21757_ (.A1(net205),
    .A2(_04143_),
    .Y(_04144_),
    .B1(net872));
 sg13g2_o21ai_1 _21758_ (.B1(_04144_),
    .Y(_04145_),
    .A1(net148),
    .A2(_04141_));
 sg13g2_nor3_1 _21759_ (.A(net149),
    .B(net205),
    .C(net193),
    .Y(_04146_));
 sg13g2_a21oi_1 _21760_ (.A1(net172),
    .A2(_04143_),
    .Y(_04147_),
    .B1(_04146_));
 sg13g2_nor2_1 _21761_ (.A(net215),
    .B(_04147_),
    .Y(_04148_));
 sg13g2_nand3_1 _21762_ (.B(net178),
    .C(net102),
    .A(_09815_),
    .Y(_04149_));
 sg13g2_o21ai_1 _21763_ (.B1(_04149_),
    .Y(_04150_),
    .A1(_04145_),
    .A2(_04148_));
 sg13g2_o21ai_1 _21764_ (.B1(_04150_),
    .Y(_04151_),
    .A1(net137),
    .A2(net86));
 sg13g2_nand2_1 _21765_ (.Y(_04152_),
    .A(net1073),
    .B(net199));
 sg13g2_nand2_1 _21766_ (.Y(_04153_),
    .A(net243),
    .B(net201));
 sg13g2_nand2_1 _21767_ (.Y(_04154_),
    .A(net1072),
    .B(_04153_));
 sg13g2_o21ai_1 _21768_ (.B1(_04154_),
    .Y(_04155_),
    .A1(_04056_),
    .A2(_04153_));
 sg13g2_nand2_1 _21769_ (.Y(_04156_),
    .A(net299),
    .B(_10369_));
 sg13g2_o21ai_1 _21770_ (.B1(_04156_),
    .Y(_04157_),
    .A1(net1063),
    .A2(_04155_));
 sg13g2_and4_1 _21771_ (.A(_04133_),
    .B(_04151_),
    .C(_04152_),
    .D(_04157_),
    .X(_04158_));
 sg13g2_nor2_1 _21772_ (.A(net299),
    .B(_11594_),
    .Y(_04159_));
 sg13g2_nor2_2 _21773_ (.A(net243),
    .B(_10369_),
    .Y(_04160_));
 sg13g2_nor2_1 _21774_ (.A(_04159_),
    .B(_04160_),
    .Y(_04161_));
 sg13g2_nand2_1 _21775_ (.Y(_04162_),
    .A(net1091),
    .B(_04161_));
 sg13g2_o21ai_1 _21776_ (.B1(net1091),
    .Y(_04163_),
    .A1(_04159_),
    .A2(_04160_));
 sg13g2_nand4_1 _21777_ (.B(net303),
    .C(_11517_),
    .A(_11225_),
    .Y(_04164_),
    .D(net256));
 sg13g2_nand4_1 _21778_ (.B(net257),
    .C(_11516_),
    .A(_11225_),
    .Y(_04165_),
    .D(_11549_));
 sg13g2_nand3_1 _21779_ (.B(net257),
    .C(net256),
    .A(_10517_),
    .Y(_04166_));
 sg13g2_and2_1 _21780_ (.A(_10481_),
    .B(_10519_),
    .X(_04167_));
 sg13g2_a22oi_1 _21781_ (.Y(_04168_),
    .B1(_04167_),
    .B2(_11502_),
    .A2(_11549_),
    .A1(_10519_));
 sg13g2_nand4_1 _21782_ (.B(_04165_),
    .C(_04166_),
    .A(_04164_),
    .Y(_04169_),
    .D(_04168_));
 sg13g2_buf_1 _21783_ (.A(_04169_),
    .X(_04170_));
 sg13g2_nor2_1 _21784_ (.A(_11561_),
    .B(_04170_),
    .Y(_04171_));
 sg13g2_nor2_1 _21785_ (.A(net252),
    .B(_04170_),
    .Y(_04172_));
 sg13g2_a22oi_1 _21786_ (.Y(_04173_),
    .B1(_04051_),
    .B2(_11413_),
    .A2(_11482_),
    .A1(_10594_));
 sg13g2_buf_1 _21787_ (.A(_04173_),
    .X(_04174_));
 sg13g2_o21ai_1 _21788_ (.B1(net203),
    .Y(_04175_),
    .A1(_10594_),
    .A2(_11482_));
 sg13g2_nand2_1 _21789_ (.Y(_04176_),
    .A(net254),
    .B(net203));
 sg13g2_o21ai_1 _21790_ (.B1(_04176_),
    .Y(_04177_),
    .A1(_04174_),
    .A2(_04175_));
 sg13g2_nor2_1 _21791_ (.A(net231),
    .B(net202),
    .Y(_04178_));
 sg13g2_o21ai_1 _21792_ (.B1(net256),
    .Y(_04179_),
    .A1(_10517_),
    .A2(net257));
 sg13g2_nor2_1 _21793_ (.A(_04178_),
    .B(_04179_),
    .Y(_04180_));
 sg13g2_nor3_1 _21794_ (.A(net302),
    .B(_04178_),
    .C(_04179_),
    .Y(_04181_));
 sg13g2_a21oi_2 _21795_ (.B1(_04174_),
    .Y(_04182_),
    .A2(_04117_),
    .A1(net227));
 sg13g2_a21oi_1 _21796_ (.A1(_11493_),
    .A2(_03984_),
    .Y(_04183_),
    .B1(_11722_));
 sg13g2_a221oi_1 _21797_ (.B2(_04182_),
    .C1(_04183_),
    .B1(_04181_),
    .A1(_04177_),
    .Y(_04184_),
    .A2(_04180_));
 sg13g2_o21ai_1 _21798_ (.B1(_04184_),
    .Y(_04185_),
    .A1(_04171_),
    .A2(_04172_));
 sg13g2_buf_2 _21799_ (.A(_04185_),
    .X(_04186_));
 sg13g2_o21ai_1 _21800_ (.B1(_04174_),
    .Y(_04187_),
    .A1(net302),
    .A2(_04122_));
 sg13g2_nor2_1 _21801_ (.A(net254),
    .B(net203),
    .Y(_04188_));
 sg13g2_nor3_1 _21802_ (.A(net254),
    .B(net228),
    .C(_11482_),
    .Y(_04189_));
 sg13g2_nor3_1 _21803_ (.A(net228),
    .B(net203),
    .C(_11482_),
    .Y(_04190_));
 sg13g2_nor4_1 _21804_ (.A(_04188_),
    .B(_04178_),
    .C(_04189_),
    .D(_04190_),
    .Y(_04191_));
 sg13g2_o21ai_1 _21805_ (.B1(_11541_),
    .Y(_04192_),
    .A1(_11415_),
    .A2(net191));
 sg13g2_o21ai_1 _21806_ (.B1(net260),
    .Y(_04193_),
    .A1(_11415_),
    .A2(net191));
 sg13g2_a221oi_1 _21807_ (.B2(_04193_),
    .C1(_04170_),
    .B1(_04192_),
    .A1(_04187_),
    .Y(_04194_),
    .A2(_04191_));
 sg13g2_a21oi_2 _21808_ (.B1(_04194_),
    .Y(_04195_),
    .A2(_11541_),
    .A1(net260));
 sg13g2_nor2_2 _21809_ (.A(_10927_),
    .B(_10365_),
    .Y(_04196_));
 sg13g2_nor3_1 _21810_ (.A(net208),
    .B(net300),
    .C(_04196_),
    .Y(_04197_));
 sg13g2_nand3_1 _21811_ (.B(_04195_),
    .C(_04197_),
    .A(_04186_),
    .Y(_04198_));
 sg13g2_nor3_1 _21812_ (.A(net208),
    .B(net261),
    .C(_04196_),
    .Y(_04199_));
 sg13g2_nand3_1 _21813_ (.B(_04195_),
    .C(_04199_),
    .A(_04186_),
    .Y(_04200_));
 sg13g2_nand2_2 _21814_ (.Y(_04201_),
    .A(_10927_),
    .B(net233));
 sg13g2_inv_1 _21815_ (.Y(_04202_),
    .A(_04201_));
 sg13g2_a22oi_1 _21816_ (.Y(_04203_),
    .B1(_04197_),
    .B2(net223),
    .A2(_04202_),
    .A1(_10360_));
 sg13g2_nand4_1 _21817_ (.B(_04198_),
    .C(_04200_),
    .A(_04000_),
    .Y(_04204_),
    .D(_04203_));
 sg13g2_buf_1 _21818_ (.A(_04204_),
    .X(_04205_));
 sg13g2_nand3_1 _21819_ (.B(net300),
    .C(_04201_),
    .A(net208),
    .Y(_04206_));
 sg13g2_nand3_1 _21820_ (.B(_10444_),
    .C(_04201_),
    .A(net208),
    .Y(_04207_));
 sg13g2_a22oi_1 _21821_ (.Y(_04208_),
    .B1(_04206_),
    .B2(_04207_),
    .A2(_04195_),
    .A1(_04186_));
 sg13g2_nand2_1 _21822_ (.Y(_04209_),
    .A(net208),
    .B(_04196_));
 sg13g2_o21ai_1 _21823_ (.B1(_04209_),
    .Y(_04210_),
    .A1(_11776_),
    .A2(_04206_));
 sg13g2_nor2_1 _21824_ (.A(_11585_),
    .B(_10232_),
    .Y(_04211_));
 sg13g2_nor3_1 _21825_ (.A(_04208_),
    .B(_04210_),
    .C(_04211_),
    .Y(_04212_));
 sg13g2_and2_1 _21826_ (.A(_11585_),
    .B(_10232_),
    .X(_04213_));
 sg13g2_buf_1 _21827_ (.A(_04213_),
    .X(_04214_));
 sg13g2_a21oi_1 _21828_ (.A1(_04205_),
    .A2(_04212_),
    .Y(_04215_),
    .B1(_04214_));
 sg13g2_mux2_1 _21829_ (.A0(_04162_),
    .A1(_04163_),
    .S(_04215_),
    .X(_04216_));
 sg13g2_nand4_1 _21830_ (.B(_04110_),
    .C(_04158_),
    .A(net671),
    .Y(_04217_),
    .D(_04216_));
 sg13g2_a21oi_2 _21831_ (.B1(_11587_),
    .Y(_04218_),
    .A2(_11576_),
    .A1(net230));
 sg13g2_xnor2_1 _21832_ (.Y(_04219_),
    .A(_04218_),
    .B(_04161_));
 sg13g2_a21oi_1 _21833_ (.A1(net607),
    .A2(_04219_),
    .Y(_04220_),
    .B1(net190));
 sg13g2_a22oi_1 _21834_ (.Y(_04221_),
    .B1(_04217_),
    .B2(_04220_),
    .A2(\cpu.ex.c_mult[11] ),
    .A1(net190));
 sg13g2_buf_1 _21835_ (.A(_08795_),
    .X(_04222_));
 sg13g2_nor2_1 _21836_ (.A(net934),
    .B(_08522_),
    .Y(_04223_));
 sg13g2_and2_1 _21837_ (.A(net1159),
    .B(_04223_),
    .X(_04224_));
 sg13g2_buf_1 _21838_ (.A(_04224_),
    .X(_04225_));
 sg13g2_nand4_1 _21839_ (.B(_08819_),
    .C(_08785_),
    .A(_08804_),
    .Y(_04226_),
    .D(_04225_));
 sg13g2_nor2_1 _21840_ (.A(net990),
    .B(_04226_),
    .Y(_04227_));
 sg13g2_nand3_1 _21841_ (.B(_08829_),
    .C(_04227_),
    .A(_08845_),
    .Y(_04228_));
 sg13g2_xor2_1 _21842_ (.B(_04228_),
    .A(_10319_),
    .X(_04229_));
 sg13g2_buf_1 _21843_ (.A(net81),
    .X(_04230_));
 sg13g2_a22oi_1 _21844_ (.Y(_04231_),
    .B1(_04229_),
    .B2(net70),
    .A2(net31),
    .A1(_08837_));
 sg13g2_o21ai_1 _21845_ (.B1(_04231_),
    .Y(_00972_),
    .A1(net71),
    .A2(_04221_));
 sg13g2_nand2_1 _21846_ (.Y(_04232_),
    .A(net299),
    .B(_04218_));
 sg13g2_o21ai_1 _21847_ (.B1(_10369_),
    .Y(_04233_),
    .A1(net299),
    .A2(_04218_));
 sg13g2_nand2_1 _21848_ (.Y(_04234_),
    .A(_04232_),
    .B(_04233_));
 sg13g2_xnor2_1 _21849_ (.Y(_04235_),
    .A(net204),
    .B(_11296_));
 sg13g2_xor2_1 _21850_ (.B(_04235_),
    .A(_04234_),
    .X(_04236_));
 sg13g2_a21oi_1 _21851_ (.A1(net607),
    .A2(_04236_),
    .Y(_04237_),
    .B1(net190));
 sg13g2_nor2b_1 _21852_ (.A(_04160_),
    .B_N(_04235_),
    .Y(_04238_));
 sg13g2_nor3_1 _21853_ (.A(_04215_),
    .B(_04159_),
    .C(_04235_),
    .Y(_04239_));
 sg13g2_a21o_1 _21854_ (.A2(_04238_),
    .A1(_04215_),
    .B1(_04239_),
    .X(_04240_));
 sg13g2_nor2_1 _21855_ (.A(net1156),
    .B(net200),
    .Y(_04241_));
 sg13g2_nor3_1 _21856_ (.A(net148),
    .B(net205),
    .C(net172),
    .Y(_04242_));
 sg13g2_o21ai_1 _21857_ (.B1(net258),
    .Y(_04243_),
    .A1(_04241_),
    .A2(_04242_));
 sg13g2_buf_1 _21858_ (.A(net178),
    .X(_04244_));
 sg13g2_or3_1 _21859_ (.A(net258),
    .B(_11602_),
    .C(net205),
    .X(_04245_));
 sg13g2_o21ai_1 _21860_ (.B1(_04245_),
    .Y(_04246_),
    .A1(net215),
    .A2(net136));
 sg13g2_nand2_1 _21861_ (.Y(_04247_),
    .A(net1146),
    .B(_04136_));
 sg13g2_inv_1 _21862_ (.Y(_04248_),
    .A(net1156));
 sg13g2_a21oi_1 _21863_ (.A1(_04136_),
    .A2(_04141_),
    .Y(_04249_),
    .B1(net136));
 sg13g2_a221oi_1 _21864_ (.B2(_04248_),
    .C1(_04249_),
    .B1(_04247_),
    .A1(_03733_),
    .Y(_04250_),
    .A2(_04246_));
 sg13g2_nand3_1 _21865_ (.B(net137),
    .C(net177),
    .A(net871),
    .Y(_04251_));
 sg13g2_a21o_1 _21866_ (.A2(net177),
    .A1(net171),
    .B1(net1072),
    .X(_04252_));
 sg13g2_a21oi_1 _21867_ (.A1(_04251_),
    .A2(_04252_),
    .Y(_04253_),
    .B1(net1063));
 sg13g2_mux2_1 _21868_ (.A0(_04160_),
    .A1(_04159_),
    .S(_04235_),
    .X(_04254_));
 sg13g2_a22oi_1 _21869_ (.Y(_04255_),
    .B1(_04254_),
    .B2(_08242_),
    .A2(net253),
    .A1(net1157));
 sg13g2_o21ai_1 _21870_ (.B1(_04255_),
    .Y(_04256_),
    .A1(_11469_),
    .A2(_04253_));
 sg13g2_a21oi_1 _21871_ (.A1(_04243_),
    .A2(_04250_),
    .Y(_04257_),
    .B1(_04256_));
 sg13g2_nand2b_1 _21872_ (.Y(_04258_),
    .B(net168),
    .A_N(net170));
 sg13g2_nand2_1 _21873_ (.Y(_04259_),
    .A(_11537_),
    .B(net139));
 sg13g2_buf_1 _21874_ (.A(_04122_),
    .X(_04260_));
 sg13g2_buf_1 _21875_ (.A(_11551_),
    .X(_04261_));
 sg13g2_buf_1 _21876_ (.A(_04036_),
    .X(_04262_));
 sg13g2_nor2b_1 _21877_ (.A(net212),
    .B_N(_04262_),
    .Y(_04263_));
 sg13g2_a21oi_1 _21878_ (.A1(net167),
    .A2(net104),
    .Y(_04264_),
    .B1(_04263_));
 sg13g2_buf_1 _21879_ (.A(net191),
    .X(_04265_));
 sg13g2_buf_1 _21880_ (.A(_04123_),
    .X(_04266_));
 sg13g2_and2_1 _21881_ (.A(_11472_),
    .B(net138),
    .X(_04267_));
 sg13g2_a221oi_1 _21882_ (.B2(_04117_),
    .C1(_04267_),
    .B1(net142),
    .A1(net166),
    .Y(_04268_),
    .A2(net135));
 sg13g2_buf_1 _21883_ (.A(_04113_),
    .X(_04269_));
 sg13g2_a22oi_1 _21884_ (.Y(_04270_),
    .B1(net134),
    .B2(net245),
    .A2(_03990_),
    .A1(net189));
 sg13g2_nand2_1 _21885_ (.Y(_04271_),
    .A(net214),
    .B(net141));
 sg13g2_a21oi_1 _21886_ (.A1(_11541_),
    .A2(net140),
    .Y(_04272_),
    .B1(_04041_));
 sg13g2_and4_1 _21887_ (.A(_04268_),
    .B(_04270_),
    .C(_04271_),
    .D(_04272_),
    .X(_04273_));
 sg13g2_nand4_1 _21888_ (.B(_04259_),
    .C(_04264_),
    .A(_04258_),
    .Y(_04274_),
    .D(_04273_));
 sg13g2_nand2_1 _21889_ (.Y(_04275_),
    .A(_11590_),
    .B(net87));
 sg13g2_nand3_1 _21890_ (.B(_04274_),
    .C(_04275_),
    .A(net1062),
    .Y(_04276_));
 sg13g2_nand4_1 _21891_ (.B(_04110_),
    .C(_04257_),
    .A(net671),
    .Y(_04277_),
    .D(_04276_));
 sg13g2_a21o_1 _21892_ (.A2(_04240_),
    .A1(net951),
    .B1(_04277_),
    .X(_04278_));
 sg13g2_a22oi_1 _21893_ (.Y(_04279_),
    .B1(_04237_),
    .B2(_04278_),
    .A2(\cpu.ex.c_mult[12] ),
    .A1(net190));
 sg13g2_inv_1 _21894_ (.Y(_04280_),
    .A(_08837_));
 sg13g2_nor2_2 _21895_ (.A(net989),
    .B(_04228_),
    .Y(_04281_));
 sg13g2_xnor2_1 _21896_ (.Y(_04282_),
    .A(_10778_),
    .B(_04281_));
 sg13g2_a22oi_1 _21897_ (.Y(_04283_),
    .B1(_04282_),
    .B2(net70),
    .A2(net31),
    .A1(net733));
 sg13g2_o21ai_1 _21898_ (.B1(_04283_),
    .Y(_00973_),
    .A1(net71),
    .A2(_04279_));
 sg13g2_inv_1 _21899_ (.Y(_04284_),
    .A(_03976_));
 sg13g2_a21oi_2 _21900_ (.B1(net213),
    .Y(_04285_),
    .A2(_04109_),
    .A1(_09813_));
 sg13g2_buf_1 _21901_ (.A(_04117_),
    .X(_04286_));
 sg13g2_nand2_1 _21902_ (.Y(_04287_),
    .A(net242),
    .B(_03990_));
 sg13g2_a22oi_1 _21903_ (.Y(_04288_),
    .B1(_04262_),
    .B2(net169),
    .A2(_04016_),
    .A1(net189));
 sg13g2_and2_1 _21904_ (.A(net245),
    .B(net138),
    .X(_04289_));
 sg13g2_a21oi_1 _21905_ (.A1(_04006_),
    .A2(net106),
    .Y(_04290_),
    .B1(_04289_));
 sg13g2_buf_1 _21906_ (.A(_11472_),
    .X(_04291_));
 sg13g2_a22oi_1 _21907_ (.Y(_04292_),
    .B1(_04029_),
    .B2(net166),
    .A2(net105),
    .A1(net165));
 sg13g2_nand4_1 _21908_ (.B(_04288_),
    .C(_04290_),
    .A(_04287_),
    .Y(_04293_),
    .D(_04292_));
 sg13g2_o21ai_1 _21909_ (.B1(_04138_),
    .Y(_04294_),
    .A1(_11585_),
    .A2(_04141_));
 sg13g2_buf_1 _21910_ (.A(net168),
    .X(_04295_));
 sg13g2_nand2_1 _21911_ (.Y(_04296_),
    .A(net243),
    .B(net133));
 sg13g2_a22oi_1 _21912_ (.Y(_04297_),
    .B1(net142),
    .B2(_04260_),
    .A2(net135),
    .A1(net214));
 sg13g2_nand2b_1 _21913_ (.Y(_04298_),
    .B(_04004_),
    .A_N(_04261_));
 sg13g2_nand3_1 _21914_ (.B(_04297_),
    .C(_04298_),
    .A(_04296_),
    .Y(_04299_));
 sg13g2_nor3_1 _21915_ (.A(_04293_),
    .B(_04294_),
    .C(_04299_),
    .Y(_04300_));
 sg13g2_o21ai_1 _21916_ (.B1(net1062),
    .Y(_04301_),
    .A1(net137),
    .A2(net86));
 sg13g2_nor2_1 _21917_ (.A(_04300_),
    .B(_04301_),
    .Y(_04302_));
 sg13g2_nand2b_1 _21918_ (.Y(_04303_),
    .B(net150),
    .A_N(net137));
 sg13g2_nand2_1 _21919_ (.Y(_04304_),
    .A(net150),
    .B(_04153_));
 sg13g2_nor2_1 _21920_ (.A(net150),
    .B(_04153_),
    .Y(_04305_));
 sg13g2_a21oi_1 _21921_ (.A1(net137),
    .A2(_04304_),
    .Y(_04306_),
    .B1(_04305_));
 sg13g2_and2_1 _21922_ (.A(_11601_),
    .B(net207),
    .X(_04307_));
 sg13g2_buf_2 _21923_ (.A(_04307_),
    .X(_04308_));
 sg13g2_nor2_2 _21924_ (.A(net149),
    .B(_11321_),
    .Y(_04309_));
 sg13g2_nor2_2 _21925_ (.A(_04308_),
    .B(_04309_),
    .Y(_04310_));
 sg13g2_mux2_1 _21926_ (.A0(_04303_),
    .A1(_04306_),
    .S(_04310_),
    .X(_04311_));
 sg13g2_nor2_1 _21927_ (.A(net671),
    .B(_04311_),
    .Y(_04312_));
 sg13g2_a22oi_1 _21928_ (.Y(_04313_),
    .B1(_04043_),
    .B2(net148),
    .A2(net133),
    .A1(net136));
 sg13g2_nor2b_1 _21929_ (.A(_04313_),
    .B_N(net1146),
    .Y(_04314_));
 sg13g2_nand2_1 _21930_ (.Y(_04315_),
    .A(net1072),
    .B(_11603_));
 sg13g2_o21ai_1 _21931_ (.B1(_04315_),
    .Y(_04316_),
    .A1(net871),
    .A2(_11603_));
 sg13g2_nor2_1 _21932_ (.A(_09819_),
    .B(_04316_),
    .Y(_04317_));
 sg13g2_nand2_1 _21933_ (.Y(_04318_),
    .A(_10718_),
    .B(net103));
 sg13g2_o21ai_1 _21934_ (.B1(_04318_),
    .Y(_04319_),
    .A1(net136),
    .A2(net103));
 sg13g2_inv_1 _21935_ (.Y(_04320_),
    .A(_04319_));
 sg13g2_a22oi_1 _21936_ (.Y(_04321_),
    .B1(_04320_),
    .B2(net1156),
    .A2(net232),
    .A1(net1073));
 sg13g2_o21ai_1 _21937_ (.B1(_04321_),
    .Y(_04322_),
    .A1(_11605_),
    .A2(_04317_));
 sg13g2_nor4_1 _21938_ (.A(_04302_),
    .B(_04312_),
    .C(_04314_),
    .D(_04322_),
    .Y(_04323_));
 sg13g2_nand2_1 _21939_ (.Y(_04324_),
    .A(_04303_),
    .B(_04310_));
 sg13g2_nor3_1 _21940_ (.A(_04218_),
    .B(_04161_),
    .C(_04324_),
    .Y(_04325_));
 sg13g2_a21oi_1 _21941_ (.A1(_04232_),
    .A2(_04233_),
    .Y(_04326_),
    .B1(_04310_));
 sg13g2_a21oi_1 _21942_ (.A1(net137),
    .A2(_11468_),
    .Y(_04327_),
    .B1(net671));
 sg13g2_o21ai_1 _21943_ (.B1(_04327_),
    .Y(_04328_),
    .A1(_04325_),
    .A2(_04326_));
 sg13g2_o21ai_1 _21944_ (.B1(net951),
    .Y(_04329_),
    .A1(_04308_),
    .A2(_04309_));
 sg13g2_nand2_1 _21945_ (.Y(_04330_),
    .A(net951),
    .B(_04310_));
 sg13g2_a221oi_1 _21946_ (.B2(_04212_),
    .C1(net299),
    .B1(_04205_),
    .A1(net170),
    .Y(_04331_),
    .A2(_11245_));
 sg13g2_a21o_1 _21947_ (.A2(net150),
    .A1(net171),
    .B1(_10369_),
    .X(_04332_));
 sg13g2_nor3_1 _21948_ (.A(_04001_),
    .B(_04208_),
    .C(_04210_),
    .Y(_04333_));
 sg13g2_nor2_1 _21949_ (.A(net204),
    .B(_11331_),
    .Y(_04334_));
 sg13g2_nor2_1 _21950_ (.A(_04214_),
    .B(_04334_),
    .Y(_04335_));
 sg13g2_nand4_1 _21951_ (.B(_04200_),
    .C(_04203_),
    .A(_04198_),
    .Y(_04336_),
    .D(_04335_));
 sg13g2_nand2b_1 _21952_ (.Y(_04337_),
    .B(net299),
    .A_N(_04211_));
 sg13g2_a21o_1 _21953_ (.A2(_04337_),
    .A1(net171),
    .B1(_11331_),
    .X(_04338_));
 sg13g2_o21ai_1 _21954_ (.B1(_04338_),
    .Y(_04339_),
    .A1(net171),
    .A2(_04337_));
 sg13g2_o21ai_1 _21955_ (.B1(_04339_),
    .Y(_04340_),
    .A1(_04333_),
    .A2(_04336_));
 sg13g2_o21ai_1 _21956_ (.B1(_04340_),
    .Y(_04341_),
    .A1(_04331_),
    .A2(_04332_));
 sg13g2_buf_2 _21957_ (.A(_04341_),
    .X(_04342_));
 sg13g2_mux2_1 _21958_ (.A0(_04329_),
    .A1(_04330_),
    .S(_04342_),
    .X(_04343_));
 sg13g2_nand4_1 _21959_ (.B(_04323_),
    .C(_04328_),
    .A(_04285_),
    .Y(_04344_),
    .D(_04343_));
 sg13g2_o21ai_1 _21960_ (.B1(net190),
    .Y(_04345_),
    .A1(_11942_),
    .A2(_11949_));
 sg13g2_nand3_1 _21961_ (.B(_04344_),
    .C(_04345_),
    .A(_04284_),
    .Y(_04346_));
 sg13g2_nand2_1 _21962_ (.Y(_04347_),
    .A(net733),
    .B(_04281_));
 sg13g2_xnor2_1 _21963_ (.Y(_04348_),
    .A(_11324_),
    .B(_04347_));
 sg13g2_a22oi_1 _21964_ (.Y(_04349_),
    .B1(_04348_),
    .B2(net70),
    .A2(net31),
    .A1(net735));
 sg13g2_nand2_1 _21965_ (.Y(_00974_),
    .A(_04346_),
    .B(_04349_));
 sg13g2_nor2_1 _21966_ (.A(_11610_),
    .B(net147),
    .Y(_04350_));
 sg13g2_nand2_1 _21967_ (.Y(_04351_),
    .A(net176),
    .B(net147));
 sg13g2_nand2b_1 _21968_ (.Y(_04352_),
    .B(_04351_),
    .A_N(_04350_));
 sg13g2_buf_1 _21969_ (.A(_04352_),
    .X(_04353_));
 sg13g2_nor2b_1 _21970_ (.A(_04309_),
    .B_N(_04353_),
    .Y(_04354_));
 sg13g2_nor2_1 _21971_ (.A(_04308_),
    .B(_04353_),
    .Y(_04355_));
 sg13g2_mux2_1 _21972_ (.A0(_04354_),
    .A1(_04355_),
    .S(_04342_),
    .X(_04356_));
 sg13g2_and2_1 _21973_ (.A(net951),
    .B(_04356_),
    .X(_04357_));
 sg13g2_o21ai_1 _21974_ (.B1(_09845_),
    .Y(_04358_),
    .A1(net109),
    .A2(_04139_));
 sg13g2_a21oi_1 _21975_ (.A1(_10872_),
    .A2(_04113_),
    .Y(_04359_),
    .B1(_04041_));
 sg13g2_a22oi_1 _21976_ (.Y(_04360_),
    .B1(_04295_),
    .B2(net171),
    .A2(net142),
    .A1(net166));
 sg13g2_nor3_1 _21977_ (.A(net200),
    .B(net256),
    .C(_03992_),
    .Y(_04361_));
 sg13g2_a21oi_1 _21978_ (.A1(net169),
    .A2(net141),
    .Y(_04362_),
    .B1(_04361_));
 sg13g2_nor2b_1 _21979_ (.A(net170),
    .B_N(net138),
    .Y(_04363_));
 sg13g2_a21oi_1 _21980_ (.A1(net242),
    .A2(_04016_),
    .Y(_04364_),
    .B1(_04363_));
 sg13g2_a22oi_1 _21981_ (.Y(_04365_),
    .B1(_04017_),
    .B2(net189),
    .A2(_03990_),
    .A1(_04260_));
 sg13g2_and4_1 _21982_ (.A(_04360_),
    .B(_04362_),
    .C(_04364_),
    .D(_04365_),
    .X(_04366_));
 sg13g2_a22oi_1 _21983_ (.Y(_04367_),
    .B1(_04029_),
    .B2(net214),
    .A2(net106),
    .A1(net165));
 sg13g2_a22oi_1 _21984_ (.Y(_04368_),
    .B1(net101),
    .B2(net244),
    .A2(net105),
    .A1(net245));
 sg13g2_nand4_1 _21985_ (.B(_04366_),
    .C(_04367_),
    .A(_04359_),
    .Y(_04369_),
    .D(_04368_));
 sg13g2_nand2b_1 _21986_ (.Y(_04370_),
    .B(_04369_),
    .A_N(_04358_));
 sg13g2_mux2_1 _21987_ (.A0(_04309_),
    .A1(_04308_),
    .S(_04353_),
    .X(_04371_));
 sg13g2_nand2_1 _21988_ (.Y(_04372_),
    .A(net176),
    .B(net179));
 sg13g2_nand2_1 _21989_ (.Y(_04373_),
    .A(_09092_),
    .B(_04372_));
 sg13g2_o21ai_1 _21990_ (.B1(_04373_),
    .Y(_04374_),
    .A1(net871),
    .A2(_04372_));
 sg13g2_nand2_1 _21991_ (.Y(_04375_),
    .A(_10718_),
    .B(_11955_));
 sg13g2_o21ai_1 _21992_ (.B1(_04375_),
    .Y(_04376_),
    .A1(_09818_),
    .A2(_04374_));
 sg13g2_nand3_1 _21993_ (.B(net136),
    .C(net87),
    .A(net1146),
    .Y(_04377_));
 sg13g2_nand2_1 _21994_ (.Y(_04378_),
    .A(net1157),
    .B(_11749_));
 sg13g2_nand3_1 _21995_ (.B(_04377_),
    .C(_04378_),
    .A(_04376_),
    .Y(_04379_));
 sg13g2_a21oi_1 _21996_ (.A1(_08243_),
    .A2(_04371_),
    .Y(_04380_),
    .B1(_04379_));
 sg13g2_nand4_1 _21997_ (.B(_04285_),
    .C(_04370_),
    .A(_04143_),
    .Y(_04381_),
    .D(_04380_));
 sg13g2_and4_1 _21998_ (.A(_11597_),
    .B(_11603_),
    .C(net607),
    .D(_04353_),
    .X(_04382_));
 sg13g2_nor4_1 _21999_ (.A(_11597_),
    .B(_11605_),
    .C(_04092_),
    .D(_04353_),
    .Y(_04383_));
 sg13g2_or2_1 _22000_ (.X(_04384_),
    .B(_04353_),
    .A(_11603_));
 sg13g2_nand3_1 _22001_ (.B(net607),
    .C(_04353_),
    .A(_11605_),
    .Y(_04385_));
 sg13g2_o21ai_1 _22002_ (.B1(_04385_),
    .Y(_04386_),
    .A1(net671),
    .A2(_04384_));
 sg13g2_or4_1 _22003_ (.A(_04381_),
    .B(_04382_),
    .C(_04383_),
    .D(_04386_),
    .X(_04387_));
 sg13g2_nor2_1 _22004_ (.A(_04357_),
    .B(_04387_),
    .Y(_04388_));
 sg13g2_o21ai_1 _22005_ (.B1(_04284_),
    .Y(_04389_),
    .A1(net246),
    .A2(\cpu.ex.c_mult[14] ));
 sg13g2_nand3_1 _22006_ (.B(net735),
    .C(_04281_),
    .A(net733),
    .Y(_04390_));
 sg13g2_xnor2_1 _22007_ (.Y(_04391_),
    .A(_11362_),
    .B(_04390_));
 sg13g2_a22oi_1 _22008_ (.Y(_04392_),
    .B1(_04391_),
    .B2(_04230_),
    .A2(_04088_),
    .A1(net821));
 sg13g2_o21ai_1 _22009_ (.B1(_04392_),
    .Y(_00975_),
    .A1(_04388_),
    .A2(_04389_));
 sg13g2_xnor2_1 _22010_ (.Y(_04393_),
    .A(_11455_),
    .B(_11361_));
 sg13g2_buf_1 _22011_ (.A(_04393_),
    .X(_04394_));
 sg13g2_nand3_1 _22012_ (.B(_04351_),
    .C(_04394_),
    .A(net951),
    .Y(_04395_));
 sg13g2_or2_1 _22013_ (.X(_04396_),
    .B(_04342_),
    .A(_04309_));
 sg13g2_o21ai_1 _22014_ (.B1(_08242_),
    .Y(_04397_),
    .A1(net148),
    .A2(net147));
 sg13g2_or2_1 _22015_ (.X(_04398_),
    .B(_04397_),
    .A(_04394_));
 sg13g2_mux2_1 _22016_ (.A0(_04398_),
    .A1(net109),
    .S(_04342_),
    .X(_04399_));
 sg13g2_nand2_1 _22017_ (.Y(_04400_),
    .A(net109),
    .B(_04398_));
 sg13g2_nor2_1 _22018_ (.A(_04342_),
    .B(_04400_),
    .Y(_04401_));
 sg13g2_a221oi_1 _22019_ (.B2(_11321_),
    .C1(_04401_),
    .B1(_04399_),
    .A1(_04395_),
    .Y(_04402_),
    .A2(_04396_));
 sg13g2_a21oi_1 _22020_ (.A1(net148),
    .A2(_11389_),
    .Y(_04403_),
    .B1(_04394_));
 sg13g2_and2_1 _22021_ (.A(_04375_),
    .B(_04394_),
    .X(_04404_));
 sg13g2_mux2_1 _22022_ (.A0(_04403_),
    .A1(_04404_),
    .S(_11606_),
    .X(_04405_));
 sg13g2_o21ai_1 _22023_ (.B1(net148),
    .Y(_04406_),
    .A1(_11955_),
    .A2(_04308_));
 sg13g2_nand2_1 _22024_ (.Y(_04407_),
    .A(net147),
    .B(_04308_));
 sg13g2_nand2_1 _22025_ (.Y(_04408_),
    .A(_04406_),
    .B(_04407_));
 sg13g2_mux2_1 _22026_ (.A0(_04408_),
    .A1(_04350_),
    .S(_04394_),
    .X(_04409_));
 sg13g2_mux2_1 _22027_ (.A0(_04375_),
    .A1(_04372_),
    .S(_04394_),
    .X(_04410_));
 sg13g2_nor2_1 _22028_ (.A(_09092_),
    .B(_11457_),
    .Y(_04411_));
 sg13g2_a21oi_1 _22029_ (.A1(_04056_),
    .A2(_11457_),
    .Y(_04412_),
    .B1(_04411_));
 sg13g2_o21ai_1 _22030_ (.B1(_11462_),
    .Y(_04413_),
    .A1(_09819_),
    .A2(_04412_));
 sg13g2_o21ai_1 _22031_ (.B1(_04413_),
    .Y(_04414_),
    .A1(_04092_),
    .A2(_04410_));
 sg13g2_a221oi_1 _22032_ (.B2(_08243_),
    .C1(_04414_),
    .B1(_04409_),
    .A1(net1073),
    .Y(_04415_),
    .A2(net223));
 sg13g2_nor2_1 _22033_ (.A(net225),
    .B(net259),
    .Y(_04416_));
 sg13g2_nor2_1 _22034_ (.A(_03732_),
    .B(_04128_),
    .Y(_04417_));
 sg13g2_a21oi_1 _22035_ (.A1(_03732_),
    .A2(net203),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_a22oi_1 _22036_ (.Y(_04419_),
    .B1(_04416_),
    .B2(_04418_),
    .A2(_03795_),
    .A1(net192));
 sg13g2_a22oi_1 _22037_ (.Y(_04420_),
    .B1(net102),
    .B2(net243),
    .A2(net135),
    .A1(net169));
 sg13g2_a22oi_1 _22038_ (.Y(_04421_),
    .B1(net141),
    .B2(net244),
    .A2(net142),
    .A1(net214));
 sg13g2_nand2_1 _22039_ (.Y(_04422_),
    .A(_04420_),
    .B(_04421_));
 sg13g2_nand2b_1 _22040_ (.Y(_04423_),
    .B(net104),
    .A_N(net212));
 sg13g2_nand2_1 _22041_ (.Y(_04424_),
    .A(_03995_),
    .B(net134));
 sg13g2_a22oi_1 _22042_ (.Y(_04425_),
    .B1(_04017_),
    .B2(_04117_),
    .A2(net133),
    .A1(net149));
 sg13g2_nand3_1 _22043_ (.B(_04424_),
    .C(_04425_),
    .A(_04423_),
    .Y(_04426_));
 sg13g2_nand2b_1 _22044_ (.Y(_04427_),
    .B(net139),
    .A_N(_11585_));
 sg13g2_and2_1 _22045_ (.A(_04001_),
    .B(net140),
    .X(_04428_));
 sg13g2_a21oi_1 _22046_ (.A1(net166),
    .A2(_03990_),
    .Y(_04429_),
    .B1(_04428_));
 sg13g2_nand3_1 _22047_ (.B(_04427_),
    .C(_04429_),
    .A(_04037_),
    .Y(_04430_));
 sg13g2_nor3_1 _22048_ (.A(_04422_),
    .B(_04426_),
    .C(_04430_),
    .Y(_04431_));
 sg13g2_o21ai_1 _22049_ (.B1(_04431_),
    .Y(_04432_),
    .A1(net258),
    .A2(_04419_));
 sg13g2_nand3_1 _22050_ (.B(_04318_),
    .C(_04432_),
    .A(net1062),
    .Y(_04433_));
 sg13g2_nand4_1 _22051_ (.B(_04285_),
    .C(_04415_),
    .A(_04143_),
    .Y(_04434_),
    .D(_04433_));
 sg13g2_a21o_1 _22052_ (.A2(_04405_),
    .A1(_04066_),
    .B1(_04434_),
    .X(_04435_));
 sg13g2_o21ai_1 _22053_ (.B1(net190),
    .Y(_04436_),
    .A1(_12010_),
    .A2(_12012_));
 sg13g2_o21ai_1 _22054_ (.B1(_04436_),
    .Y(_04437_),
    .A1(_04402_),
    .A2(_04435_));
 sg13g2_nand4_1 _22055_ (.B(net735),
    .C(net821),
    .A(net733),
    .Y(_04438_),
    .D(_04281_));
 sg13g2_xor2_1 _22056_ (.B(_04438_),
    .A(_00192_),
    .X(_04439_));
 sg13g2_a22oi_1 _22057_ (.Y(_04440_),
    .B1(_04439_),
    .B2(net70),
    .A2(net31),
    .A1(_08637_));
 sg13g2_o21ai_1 _22058_ (.B1(_04440_),
    .Y(_00976_),
    .A1(_03977_),
    .A2(_04437_));
 sg13g2_nand2_1 _22059_ (.Y(_04441_),
    .A(_04244_),
    .B(_04016_));
 sg13g2_a22oi_1 _22060_ (.Y(_04442_),
    .B1(net142),
    .B2(net109),
    .A2(net135),
    .A1(net243));
 sg13g2_nand2b_1 _22061_ (.Y(_04443_),
    .B(net141),
    .A_N(net170));
 sg13g2_o21ai_1 _22062_ (.B1(_04259_),
    .Y(_04444_),
    .A1(net212),
    .A2(_04141_));
 sg13g2_a221oi_1 _22063_ (.B2(net214),
    .C1(_04444_),
    .B1(net133),
    .A1(net165),
    .Y(_04445_),
    .A2(net106));
 sg13g2_nand4_1 _22064_ (.B(_04442_),
    .C(_04443_),
    .A(_04441_),
    .Y(_04446_),
    .D(_04445_));
 sg13g2_nor2_1 _22065_ (.A(_03734_),
    .B(net200),
    .Y(_04447_));
 sg13g2_nand3_1 _22066_ (.B(_04447_),
    .C(net169),
    .A(net192),
    .Y(_04448_));
 sg13g2_nor2_1 _22067_ (.A(net192),
    .B(_04143_),
    .Y(_04449_));
 sg13g2_nand2_1 _22068_ (.Y(_04450_),
    .A(_11645_),
    .B(_04449_));
 sg13g2_a21oi_1 _22069_ (.A1(_04448_),
    .A2(_04450_),
    .Y(_04451_),
    .B1(_11416_));
 sg13g2_and2_1 _22070_ (.A(net148),
    .B(_03990_),
    .X(_04452_));
 sg13g2_a221oi_1 _22071_ (.B2(net245),
    .C1(_04452_),
    .B1(net101),
    .A1(net137),
    .Y(_04453_),
    .A2(net104));
 sg13g2_o21ai_1 _22072_ (.B1(_04453_),
    .Y(_04454_),
    .A1(_11418_),
    .A2(_03982_));
 sg13g2_nor3_1 _22073_ (.A(_04446_),
    .B(_04451_),
    .C(_04454_),
    .Y(_04455_));
 sg13g2_inv_1 _22074_ (.Y(_04456_),
    .A(_04045_));
 sg13g2_o21ai_1 _22075_ (.B1(_04456_),
    .Y(_04457_),
    .A1(net166),
    .A2(net86));
 sg13g2_nor2_1 _22076_ (.A(_11484_),
    .B(_11490_),
    .Y(_04458_));
 sg13g2_xnor2_1 _22077_ (.Y(_04459_),
    .A(net226),
    .B(_11510_));
 sg13g2_xnor2_1 _22078_ (.Y(_04460_),
    .A(_04458_),
    .B(_04459_));
 sg13g2_xor2_1 _22079_ (.B(_04459_),
    .A(_04182_),
    .X(_04461_));
 sg13g2_a221oi_1 _22080_ (.B2(net1155),
    .C1(_11629_),
    .B1(_04097_),
    .A1(net1157),
    .Y(_04462_),
    .A2(net230));
 sg13g2_nor2b_1 _22081_ (.A(_04097_),
    .B_N(net1072),
    .Y(_04463_));
 sg13g2_o21ai_1 _22082_ (.B1(_04096_),
    .Y(_04464_),
    .A1(net1145),
    .A2(_04463_));
 sg13g2_a22oi_1 _22083_ (.Y(_04465_),
    .B1(net103),
    .B2(net242),
    .A2(net133),
    .A1(net189));
 sg13g2_nand2b_1 _22084_ (.Y(_04466_),
    .B(_09844_),
    .A_N(_04465_));
 sg13g2_nand3_1 _22085_ (.B(_04464_),
    .C(_04466_),
    .A(_04462_),
    .Y(_04467_));
 sg13g2_a221oi_1 _22086_ (.B2(net1091),
    .C1(_04467_),
    .B1(_04461_),
    .A1(_04073_),
    .Y(_04468_),
    .A2(_04460_));
 sg13g2_o21ai_1 _22087_ (.B1(_04468_),
    .Y(_04469_),
    .A1(_04455_),
    .A2(_04457_));
 sg13g2_o21ai_1 _22088_ (.B1(_04469_),
    .Y(_04470_),
    .A1(net246),
    .A2(\cpu.ex.c_mult[2] ));
 sg13g2_a21o_1 _22089_ (.A2(net81),
    .A1(net934),
    .B1(_04087_),
    .X(_04471_));
 sg13g2_nor2_1 _22090_ (.A(net718),
    .B(net934),
    .Y(_04472_));
 sg13g2_nor4_1 _22091_ (.A(net1081),
    .B(_11011_),
    .C(_08419_),
    .D(_12025_),
    .Y(_04473_));
 sg13g2_a221oi_1 _22092_ (.B2(_04080_),
    .C1(_04473_),
    .B1(_04472_),
    .A1(net718),
    .Y(_04474_),
    .A2(_04471_));
 sg13g2_o21ai_1 _22093_ (.B1(_04474_),
    .Y(_00977_),
    .A1(_03977_),
    .A2(_04470_));
 sg13g2_nor4_1 _22094_ (.A(net1081),
    .B(_11011_),
    .C(_00267_),
    .D(_12025_),
    .Y(_04475_));
 sg13g2_buf_1 _22095_ (.A(net350),
    .X(_04476_));
 sg13g2_o21ai_1 _22096_ (.B1(net292),
    .Y(_04477_),
    .A1(_04083_),
    .A2(_04475_));
 sg13g2_nand2_1 _22097_ (.Y(_04478_),
    .A(net718),
    .B(net819));
 sg13g2_a21o_1 _22098_ (.A2(_04478_),
    .A1(net81),
    .B1(_04087_),
    .X(_04479_));
 sg13g2_nor2_1 _22099_ (.A(net649),
    .B(_04478_),
    .Y(_04480_));
 sg13g2_a22oi_1 _22100_ (.Y(_04481_),
    .B1(_04480_),
    .B2(_04080_),
    .A2(_04479_),
    .A1(net649));
 sg13g2_nor2b_1 _22101_ (.A(net212),
    .B_N(_04022_),
    .Y(_04482_));
 sg13g2_a221oi_1 _22102_ (.B2(_11612_),
    .C1(_04482_),
    .B1(_03994_),
    .A1(net137),
    .Y(_04483_),
    .A2(_04266_));
 sg13g2_a21oi_1 _22103_ (.A1(net165),
    .A2(net139),
    .Y(_04484_),
    .B1(_04428_));
 sg13g2_a21oi_1 _22104_ (.A1(_04014_),
    .A2(net134),
    .Y(_04485_),
    .B1(_04041_));
 sg13g2_nand2_1 _22105_ (.Y(_04486_),
    .A(_04484_),
    .B(_04485_));
 sg13g2_a21oi_1 _22106_ (.A1(_04025_),
    .A2(_04004_),
    .Y(_04487_),
    .B1(_04486_));
 sg13g2_nor2b_1 _22107_ (.A(net170),
    .B_N(net101),
    .Y(_04488_));
 sg13g2_a221oi_1 _22108_ (.B2(net244),
    .C1(_04488_),
    .B1(net102),
    .A1(net109),
    .Y(_04489_),
    .A2(net104));
 sg13g2_nor2_1 _22109_ (.A(_11420_),
    .B(_04416_),
    .Y(_04490_));
 sg13g2_nor2_1 _22110_ (.A(_04248_),
    .B(_04490_),
    .Y(_04491_));
 sg13g2_o21ai_1 _22111_ (.B1(net136),
    .Y(_04492_),
    .A1(_03990_),
    .A2(_04491_));
 sg13g2_nand4_1 _22112_ (.B(_04487_),
    .C(_04489_),
    .A(_04483_),
    .Y(_04493_),
    .D(_04492_));
 sg13g2_nor2_1 _22113_ (.A(net214),
    .B(net86),
    .Y(_04494_));
 sg13g2_nor2_1 _22114_ (.A(net872),
    .B(_04494_),
    .Y(_04495_));
 sg13g2_nor2_1 _22115_ (.A(net192),
    .B(net202),
    .Y(_04496_));
 sg13g2_nor2_1 _22116_ (.A(_09092_),
    .B(_04496_),
    .Y(_04497_));
 sg13g2_a21oi_1 _22117_ (.A1(net871),
    .A2(_04496_),
    .Y(_04498_),
    .B1(_04497_));
 sg13g2_nand2_1 _22118_ (.Y(_04499_),
    .A(net225),
    .B(net202));
 sg13g2_o21ai_1 _22119_ (.B1(_04499_),
    .Y(_04500_),
    .A1(net1145),
    .A2(_04498_));
 sg13g2_a21oi_1 _22120_ (.A1(net1157),
    .A2(_11594_),
    .Y(_04501_),
    .B1(net213));
 sg13g2_mux2_1 _22121_ (.A0(_11484_),
    .A1(_04418_),
    .S(net215),
    .X(_04502_));
 sg13g2_nand3_1 _22122_ (.B(_04136_),
    .C(_04502_),
    .A(_09844_),
    .Y(_04503_));
 sg13g2_nand3_1 _22123_ (.B(_04501_),
    .C(_04503_),
    .A(_04500_),
    .Y(_04504_));
 sg13g2_a21oi_1 _22124_ (.A1(_04493_),
    .A2(_04495_),
    .Y(_04505_),
    .B1(_04504_));
 sg13g2_and2_1 _22125_ (.A(_04096_),
    .B(_04099_),
    .X(_04506_));
 sg13g2_xnor2_1 _22126_ (.Y(_04507_),
    .A(net199),
    .B(_11517_));
 sg13g2_xor2_1 _22127_ (.B(_04507_),
    .A(_04506_),
    .X(_04508_));
 sg13g2_a21oi_1 _22128_ (.A1(net226),
    .A2(_04182_),
    .Y(_04509_),
    .B1(_04177_));
 sg13g2_xnor2_1 _22129_ (.Y(_04510_),
    .A(_04509_),
    .B(_04507_));
 sg13g2_a22oi_1 _22130_ (.Y(_04511_),
    .B1(_04510_),
    .B2(net1091),
    .A2(_04508_),
    .A1(_04073_));
 sg13g2_a22oi_1 _22131_ (.Y(_04512_),
    .B1(_04505_),
    .B2(_04511_),
    .A2(_11703_),
    .A1(net213));
 sg13g2_nand2_1 _22132_ (.Y(_04513_),
    .A(_04284_),
    .B(_04512_));
 sg13g2_nand3_1 _22133_ (.B(_04481_),
    .C(_04513_),
    .A(_04477_),
    .Y(_00978_));
 sg13g2_a21oi_1 _22134_ (.A1(_04506_),
    .A2(_04499_),
    .Y(_04514_),
    .B1(_04496_));
 sg13g2_nand2_1 _22135_ (.Y(_04515_),
    .A(_11704_),
    .B(net257));
 sg13g2_nand2_1 _22136_ (.Y(_04516_),
    .A(_11493_),
    .B(_03984_));
 sg13g2_nand2_1 _22137_ (.Y(_04517_),
    .A(_04515_),
    .B(_04516_));
 sg13g2_xor2_1 _22138_ (.B(_04517_),
    .A(_04514_),
    .X(_04518_));
 sg13g2_a22oi_1 _22139_ (.Y(_04519_),
    .B1(_04187_),
    .B2(_04191_),
    .A2(net202),
    .A1(net231));
 sg13g2_buf_1 _22140_ (.A(_04519_),
    .X(_04520_));
 sg13g2_xnor2_1 _22141_ (.Y(_04521_),
    .A(_04520_),
    .B(_04517_));
 sg13g2_a21oi_1 _22142_ (.A1(_11541_),
    .A2(net168),
    .Y(_04522_),
    .B1(_04041_));
 sg13g2_nor2b_1 _22143_ (.A(net170),
    .B_N(_04009_),
    .Y(_04523_));
 sg13g2_a21oi_1 _22144_ (.A1(net149),
    .A2(net135),
    .Y(_04524_),
    .B1(_04523_));
 sg13g2_nand2_1 _22145_ (.Y(_04525_),
    .A(_04522_),
    .B(_04524_));
 sg13g2_a221oi_1 _22146_ (.B2(_04025_),
    .C1(_04525_),
    .B1(net101),
    .A1(_11612_),
    .Y(_04526_),
    .A2(net104));
 sg13g2_a22oi_1 _22147_ (.Y(_04527_),
    .B1(_04269_),
    .B2(_04006_),
    .A2(net141),
    .A1(_04134_));
 sg13g2_a22oi_1 _22148_ (.Y(_04528_),
    .B1(net102),
    .B2(net165),
    .A2(net105),
    .A1(net245));
 sg13g2_o21ai_1 _22149_ (.B1(_04244_),
    .Y(_04529_),
    .A1(_03994_),
    .A2(_04491_));
 sg13g2_nand4_1 _22150_ (.B(_04527_),
    .C(_04528_),
    .A(_04526_),
    .Y(_04530_),
    .D(_04529_));
 sg13g2_a21oi_1 _22151_ (.A1(net212),
    .A2(net87),
    .Y(_04531_),
    .B1(net872));
 sg13g2_mux2_1 _22152_ (.A0(_09092_),
    .A1(net1155),
    .S(_11543_),
    .X(_04532_));
 sg13g2_o21ai_1 _22153_ (.B1(_04102_),
    .Y(_04533_),
    .A1(net1145),
    .A2(_04532_));
 sg13g2_a21oi_1 _22154_ (.A1(net1157),
    .A2(_11468_),
    .Y(_04534_),
    .B1(net213));
 sg13g2_a22oi_1 _22155_ (.Y(_04535_),
    .B1(net134),
    .B2(net242),
    .A2(net133),
    .A1(net167));
 sg13g2_a21oi_1 _22156_ (.A1(_04128_),
    .A2(net102),
    .Y(_04536_),
    .B1(net103));
 sg13g2_o21ai_1 _22157_ (.B1(_09844_),
    .Y(_04537_),
    .A1(net166),
    .A2(_04138_));
 sg13g2_a21o_1 _22158_ (.A2(_04536_),
    .A1(_04535_),
    .B1(_04537_),
    .X(_04538_));
 sg13g2_nand3_1 _22159_ (.B(_04534_),
    .C(_04538_),
    .A(_04533_),
    .Y(_04539_));
 sg13g2_a221oi_1 _22160_ (.B2(_04531_),
    .C1(_04539_),
    .B1(_04530_),
    .A1(net1091),
    .Y(_04540_),
    .A2(_04521_));
 sg13g2_o21ai_1 _22161_ (.B1(_04540_),
    .Y(_04541_),
    .A1(_04067_),
    .A2(_04518_));
 sg13g2_o21ai_1 _22162_ (.B1(_04541_),
    .Y(_04542_),
    .A1(net246),
    .A2(\cpu.ex.c_mult[4] ));
 sg13g2_nand2b_1 _22163_ (.Y(_04543_),
    .B(net81),
    .A_N(_04223_));
 sg13g2_nand2b_1 _22164_ (.Y(_04544_),
    .B(_04543_),
    .A_N(_04087_));
 sg13g2_nor3_1 _22165_ (.A(net1159),
    .B(net934),
    .C(_08522_),
    .Y(_04545_));
 sg13g2_nor4_1 _22166_ (.A(_08378_),
    .B(net350),
    .C(net815),
    .D(_12024_),
    .Y(_04546_));
 sg13g2_a221oi_1 _22167_ (.B2(net81),
    .C1(_04546_),
    .B1(_04545_),
    .A1(net1159),
    .Y(_04547_),
    .A2(_04544_));
 sg13g2_o21ai_1 _22168_ (.B1(_04547_),
    .Y(_00979_),
    .A1(net71),
    .A2(_04542_));
 sg13g2_xnor2_1 _22169_ (.Y(_04548_),
    .A(net232),
    .B(net212));
 sg13g2_inv_1 _22170_ (.Y(_04549_),
    .A(_04516_));
 sg13g2_o21ai_1 _22171_ (.B1(_04515_),
    .Y(_04550_),
    .A1(_04549_),
    .A2(_04520_));
 sg13g2_xor2_1 _22172_ (.B(_04550_),
    .A(_04548_),
    .X(_04551_));
 sg13g2_nand2_1 _22173_ (.Y(_04552_),
    .A(_11704_),
    .B(net214));
 sg13g2_a21oi_1 _22174_ (.A1(_04514_),
    .A2(_04552_),
    .Y(_04553_),
    .B1(_11522_));
 sg13g2_xor2_1 _22175_ (.B(_04548_),
    .A(_04553_),
    .X(_04554_));
 sg13g2_a221oi_1 _22176_ (.B2(net167),
    .C1(_04023_),
    .B1(net134),
    .A1(net242),
    .Y(_04555_),
    .A2(net102));
 sg13g2_a21oi_1 _22177_ (.A1(_04129_),
    .A2(net105),
    .Y(_04556_),
    .B1(net103));
 sg13g2_nand2_1 _22178_ (.Y(_04557_),
    .A(_04555_),
    .B(_04556_));
 sg13g2_nand3b_1 _22179_ (.B(_04557_),
    .C(net1062),
    .Y(_04558_),
    .A_N(_04494_));
 sg13g2_mux2_1 _22180_ (.A0(net1072),
    .A1(net1155),
    .S(_11550_),
    .X(_04559_));
 sg13g2_o21ai_1 _22181_ (.B1(_11552_),
    .Y(_04560_),
    .A1(net1063),
    .A2(_04559_));
 sg13g2_a21oi_1 _22182_ (.A1(net1073),
    .A2(net206),
    .Y(_04561_),
    .B1(net213));
 sg13g2_nor2_1 _22183_ (.A(net248),
    .B(net192),
    .Y(_04562_));
 sg13g2_a22oi_1 _22184_ (.Y(_04563_),
    .B1(_04562_),
    .B2(net149),
    .A2(_03981_),
    .A1(net192));
 sg13g2_a221oi_1 _22185_ (.B2(_03995_),
    .C1(_04289_),
    .B1(net101),
    .A1(_11460_),
    .Y(_04564_),
    .A2(net104));
 sg13g2_o21ai_1 _22186_ (.B1(_04564_),
    .Y(_04565_),
    .A1(_10598_),
    .A2(_04563_));
 sg13g2_o21ai_1 _22187_ (.B1(_04449_),
    .Y(_04566_),
    .A1(net226),
    .A2(_04140_));
 sg13g2_nand2_1 _22188_ (.Y(_04567_),
    .A(_11537_),
    .B(net168));
 sg13g2_nand2_1 _22189_ (.Y(_04568_),
    .A(_04427_),
    .B(_04567_));
 sg13g2_a221oi_1 _22190_ (.B2(net243),
    .C1(_04568_),
    .B1(net140),
    .A1(net176),
    .Y(_04569_),
    .A2(net135));
 sg13g2_nand3_1 _22191_ (.B(_04566_),
    .C(_04569_),
    .A(_04114_),
    .Y(_04570_));
 sg13g2_a21oi_1 _22192_ (.A1(_11561_),
    .A2(net103),
    .Y(_04571_),
    .B1(net872));
 sg13g2_o21ai_1 _22193_ (.B1(_04571_),
    .Y(_04572_),
    .A1(_04565_),
    .A2(_04570_));
 sg13g2_nand4_1 _22194_ (.B(_04560_),
    .C(_04561_),
    .A(_04558_),
    .Y(_04573_),
    .D(_04572_));
 sg13g2_a221oi_1 _22195_ (.B2(_04073_),
    .C1(_04573_),
    .B1(_04554_),
    .A1(net1091),
    .Y(_04574_),
    .A2(_04551_));
 sg13g2_a21oi_1 _22196_ (.A1(net190),
    .A2(_11743_),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_inv_1 _22197_ (.Y(_04576_),
    .A(_04575_));
 sg13g2_buf_1 _22198_ (.A(_08804_),
    .X(_04577_));
 sg13g2_xnor2_1 _22199_ (.Y(_04578_),
    .A(_10507_),
    .B(_04225_));
 sg13g2_a22oi_1 _22200_ (.Y(_04579_),
    .B1(_04578_),
    .B2(net70),
    .A2(net31),
    .A1(net988));
 sg13g2_o21ai_1 _22201_ (.B1(_04579_),
    .Y(_00980_),
    .A1(net71),
    .A2(_04576_));
 sg13g2_nor2_1 _22202_ (.A(_04549_),
    .B(_04520_),
    .Y(_04580_));
 sg13g2_o21ai_1 _22203_ (.B1(net212),
    .Y(_04581_),
    .A1(net199),
    .A2(net202));
 sg13g2_o21ai_1 _22204_ (.B1(_11722_),
    .Y(_04582_),
    .A1(_04509_),
    .A2(_04581_));
 sg13g2_a21oi_1 _22205_ (.A1(_04580_),
    .A2(_04582_),
    .Y(_04583_),
    .B1(_04170_));
 sg13g2_xnor2_1 _22206_ (.Y(_04584_),
    .A(net252),
    .B(_11561_));
 sg13g2_xnor2_1 _22207_ (.Y(_04585_),
    .A(_04583_),
    .B(_04584_));
 sg13g2_xnor2_1 _22208_ (.Y(_04586_),
    .A(_04106_),
    .B(_04584_));
 sg13g2_nand2_1 _22209_ (.Y(_04587_),
    .A(net212),
    .B(_04043_));
 sg13g2_a22oi_1 _22210_ (.Y(_04588_),
    .B1(_04269_),
    .B2(net166),
    .A2(net133),
    .A1(_03985_));
 sg13g2_a22oi_1 _22211_ (.Y(_04589_),
    .B1(_04111_),
    .B2(net167),
    .A2(_04010_),
    .A1(net189));
 sg13g2_a21oi_1 _22212_ (.A1(net242),
    .A2(_04013_),
    .Y(_04590_),
    .B1(net103));
 sg13g2_nand3_1 _22213_ (.B(_04589_),
    .C(_04590_),
    .A(_04588_),
    .Y(_04591_));
 sg13g2_nand3_1 _22214_ (.B(_04587_),
    .C(_04591_),
    .A(net1062),
    .Y(_04592_));
 sg13g2_nand2_1 _22215_ (.Y(_04593_),
    .A(net1072),
    .B(_11542_));
 sg13g2_o21ai_1 _22216_ (.B1(_04593_),
    .Y(_04594_),
    .A1(net871),
    .A2(_11542_));
 sg13g2_o21ai_1 _22217_ (.B1(_11562_),
    .Y(_04595_),
    .A1(net1063),
    .A2(_04594_));
 sg13g2_a21oi_1 _22218_ (.A1(net1073),
    .A2(_11389_),
    .Y(_04596_),
    .B1(_04053_));
 sg13g2_nand2_1 _22219_ (.Y(_04597_),
    .A(_03735_),
    .B(net245));
 sg13g2_a21oi_1 _22220_ (.A1(_03982_),
    .A2(_04597_),
    .Y(_04598_),
    .B1(_11418_));
 sg13g2_nand3_1 _22221_ (.B(net176),
    .C(_03795_),
    .A(net258),
    .Y(_04599_));
 sg13g2_o21ai_1 _22222_ (.B1(_04599_),
    .Y(_04600_),
    .A1(_03795_),
    .A2(_04143_));
 sg13g2_nand2_1 _22223_ (.Y(_04601_),
    .A(_11684_),
    .B(_04600_));
 sg13g2_a21oi_1 _22224_ (.A1(net165),
    .A2(_04295_),
    .Y(_04602_),
    .B1(_04363_));
 sg13g2_a22oi_1 _22225_ (.Y(_04603_),
    .B1(net101),
    .B2(net109),
    .A2(net105),
    .A1(net243));
 sg13g2_a22oi_1 _22226_ (.Y(_04604_),
    .B1(_04010_),
    .B2(_04134_),
    .A2(_04266_),
    .A1(net178));
 sg13g2_nand4_1 _22227_ (.B(_04602_),
    .C(_04603_),
    .A(_04601_),
    .Y(_04605_),
    .D(_04604_));
 sg13g2_a21oi_1 _22228_ (.A1(_11571_),
    .A2(net87),
    .Y(_04606_),
    .B1(net872));
 sg13g2_o21ai_1 _22229_ (.B1(_04606_),
    .Y(_04607_),
    .A1(_04598_),
    .A2(_04605_));
 sg13g2_nand4_1 _22230_ (.B(_04595_),
    .C(_04596_),
    .A(_04592_),
    .Y(_04608_),
    .D(_04607_));
 sg13g2_a221oi_1 _22231_ (.B2(_04073_),
    .C1(_04608_),
    .B1(_04586_),
    .A1(_08244_),
    .Y(_04609_),
    .A2(_04585_));
 sg13g2_a21o_1 _22232_ (.A2(_11764_),
    .A1(_04090_),
    .B1(_04609_),
    .X(_04610_));
 sg13g2_buf_1 _22233_ (.A(_08819_),
    .X(_04611_));
 sg13g2_nand2_1 _22234_ (.Y(_04612_),
    .A(_08804_),
    .B(_04225_));
 sg13g2_xnor2_1 _22235_ (.Y(_04613_),
    .A(_10434_),
    .B(_04612_));
 sg13g2_a22oi_1 _22236_ (.Y(_04614_),
    .B1(_04613_),
    .B2(net70),
    .A2(net31),
    .A1(net987));
 sg13g2_o21ai_1 _22237_ (.B1(_04614_),
    .Y(_00981_),
    .A1(net71),
    .A2(_04610_));
 sg13g2_nand2_1 _22238_ (.Y(_04615_),
    .A(_04186_),
    .B(_04195_));
 sg13g2_xnor2_1 _22239_ (.Y(_04616_),
    .A(_04095_),
    .B(_04615_));
 sg13g2_nor2_1 _22240_ (.A(_04291_),
    .B(net86),
    .Y(_04617_));
 sg13g2_a22oi_1 _22241_ (.Y(_04618_),
    .B1(_04012_),
    .B2(net204),
    .A2(net140),
    .A1(net149));
 sg13g2_a221oi_1 _22242_ (.B2(_11610_),
    .C1(_04118_),
    .B1(_04036_),
    .A1(_10872_),
    .Y(_04619_),
    .A2(net138));
 sg13g2_nand3b_1 _22243_ (.B(_04618_),
    .C(_04619_),
    .Y(_04620_),
    .A_N(_04294_));
 sg13g2_a21o_1 _22244_ (.A2(net141),
    .A1(net178),
    .B1(_04620_),
    .X(_04621_));
 sg13g2_o21ai_1 _22245_ (.B1(_03787_),
    .Y(_04622_),
    .A1(net248),
    .A2(_10598_));
 sg13g2_nand2_1 _22246_ (.Y(_04623_),
    .A(net178),
    .B(_04622_));
 sg13g2_nand2b_1 _22247_ (.Y(_04624_),
    .B(_04623_),
    .A_N(_04620_));
 sg13g2_a22oi_1 _22248_ (.Y(_04625_),
    .B1(_04624_),
    .B2(_09082_),
    .A2(_04621_),
    .A1(net1146));
 sg13g2_mux2_1 _22249_ (.A0(_09092_),
    .A1(net1155),
    .S(_11539_),
    .X(_04626_));
 sg13g2_nor2_1 _22250_ (.A(net1145),
    .B(_04626_),
    .Y(_04627_));
 sg13g2_a21oi_1 _22251_ (.A1(net1157),
    .A2(_11361_),
    .Y(_04628_),
    .B1(_11629_));
 sg13g2_o21ai_1 _22252_ (.B1(_04628_),
    .Y(_04629_),
    .A1(_11569_),
    .A2(_04627_));
 sg13g2_a221oi_1 _22253_ (.B2(net166),
    .C1(_04482_),
    .B1(net102),
    .A1(net167),
    .Y(_04630_),
    .A2(net105));
 sg13g2_a21o_1 _22254_ (.A2(_04036_),
    .A1(_04128_),
    .B1(_04041_),
    .X(_04631_));
 sg13g2_a221oi_1 _22255_ (.B2(_03985_),
    .C1(_04631_),
    .B1(net134),
    .A1(net242),
    .Y(_04632_),
    .A2(net106));
 sg13g2_o21ai_1 _22256_ (.B1(_09844_),
    .Y(_04633_),
    .A1(net169),
    .A2(net86));
 sg13g2_a21oi_1 _22257_ (.A1(_04630_),
    .A2(_04632_),
    .Y(_04634_),
    .B1(_04633_));
 sg13g2_nor2_1 _22258_ (.A(_04629_),
    .B(_04634_),
    .Y(_04635_));
 sg13g2_o21ai_1 _22259_ (.B1(_04635_),
    .Y(_04636_),
    .A1(_04617_),
    .A2(_04625_));
 sg13g2_a221oi_1 _22260_ (.B2(net951),
    .C1(_04636_),
    .B1(_04616_),
    .A1(_04073_),
    .Y(_04637_),
    .A2(_04109_));
 sg13g2_a21o_1 _22261_ (.A2(_11783_),
    .A1(_04090_),
    .B1(_04637_),
    .X(_04638_));
 sg13g2_buf_1 _22262_ (.A(_08785_),
    .X(_04639_));
 sg13g2_nand3_1 _22263_ (.B(_08819_),
    .C(_04225_),
    .A(_08804_),
    .Y(_04640_));
 sg13g2_xor2_1 _22264_ (.B(_04640_),
    .A(_10411_),
    .X(_04641_));
 sg13g2_a22oi_1 _22265_ (.Y(_04642_),
    .B1(_04641_),
    .B2(net70),
    .A2(net31),
    .A1(net986));
 sg13g2_o21ai_1 _22266_ (.B1(_04642_),
    .Y(_00982_),
    .A1(net71),
    .A2(_04638_));
 sg13g2_or2_1 _22267_ (.X(_04643_),
    .B(_04196_),
    .A(_04202_));
 sg13g2_buf_1 _22268_ (.A(_04643_),
    .X(_04644_));
 sg13g2_nor2_1 _22269_ (.A(_11569_),
    .B(_11568_),
    .Y(_04645_));
 sg13g2_xor2_1 _22270_ (.B(_04645_),
    .A(_04644_),
    .X(_04646_));
 sg13g2_inv_1 _22271_ (.Y(_04647_),
    .A(_04094_));
 sg13g2_o21ai_1 _22272_ (.B1(_04093_),
    .Y(_04648_),
    .A1(_04647_),
    .A2(_04615_));
 sg13g2_xor2_1 _22273_ (.B(_04644_),
    .A(_04648_),
    .X(_04649_));
 sg13g2_nand2_1 _22274_ (.Y(_04650_),
    .A(net951),
    .B(_04649_));
 sg13g2_nor2_1 _22275_ (.A(_04261_),
    .B(_04141_),
    .Y(_04651_));
 sg13g2_a221oi_1 _22276_ (.B2(_04286_),
    .C1(_04651_),
    .B1(net101),
    .A1(_04129_),
    .Y(_04652_),
    .A2(net141));
 sg13g2_and2_1 _22277_ (.A(_03984_),
    .B(net138),
    .X(_04653_));
 sg13g2_a221oi_1 _22278_ (.B2(_04265_),
    .C1(_04653_),
    .B1(net105),
    .A1(net167),
    .Y(_04654_),
    .A2(net106));
 sg13g2_and3_1 _22279_ (.X(_04655_),
    .A(_04522_),
    .B(_04652_),
    .C(_04654_));
 sg13g2_o21ai_1 _22280_ (.B1(_09845_),
    .Y(_04656_),
    .A1(net244),
    .A2(_04139_));
 sg13g2_nand2_1 _22281_ (.Y(_04657_),
    .A(_10927_),
    .B(net229));
 sg13g2_o21ai_1 _22282_ (.B1(_09093_),
    .Y(_04658_),
    .A1(_10927_),
    .A2(net229));
 sg13g2_nand3_1 _22283_ (.B(net165),
    .C(_10365_),
    .A(net1155),
    .Y(_04659_));
 sg13g2_nand3b_1 _22284_ (.B(_04658_),
    .C(_04659_),
    .Y(_04660_),
    .A_N(_09818_));
 sg13g2_a22oi_1 _22285_ (.Y(_04661_),
    .B1(_04657_),
    .B2(_04660_),
    .A2(net215),
    .A1(net1073));
 sg13g2_o21ai_1 _22286_ (.B1(_04661_),
    .Y(_04662_),
    .A1(_04655_),
    .A2(_04656_));
 sg13g2_a22oi_1 _22287_ (.Y(_04663_),
    .B1(_04033_),
    .B2(net204),
    .A2(_04012_),
    .A1(_11601_));
 sg13g2_a22oi_1 _22288_ (.Y(_04664_),
    .B1(_04036_),
    .B2(_11455_),
    .A2(net140),
    .A1(net176));
 sg13g2_nand4_1 _22289_ (.B(_04359_),
    .C(_04663_),
    .A(_04258_),
    .Y(_04665_),
    .D(_04664_));
 sg13g2_nand2b_1 _22290_ (.Y(_04666_),
    .B(_04623_),
    .A_N(_04665_));
 sg13g2_a22oi_1 _22291_ (.Y(_04667_),
    .B1(_04666_),
    .B2(net1156),
    .A2(_04665_),
    .A1(net1146));
 sg13g2_a21oi_1 _22292_ (.A1(_10900_),
    .A2(net87),
    .Y(_04668_),
    .B1(_04667_));
 sg13g2_nor2_1 _22293_ (.A(_04662_),
    .B(_04668_),
    .Y(_04669_));
 sg13g2_nand4_1 _22294_ (.B(_04110_),
    .C(_04650_),
    .A(net671),
    .Y(_04670_),
    .D(_04669_));
 sg13g2_o21ai_1 _22295_ (.B1(_04670_),
    .Y(_04671_),
    .A1(net671),
    .A2(_04646_));
 sg13g2_mux2_1 _22296_ (.A0(_11810_),
    .A1(_04671_),
    .S(net246),
    .X(_04672_));
 sg13g2_inv_1 _22297_ (.Y(_04673_),
    .A(_00282_));
 sg13g2_xnor2_1 _22298_ (.Y(_04674_),
    .A(_04673_),
    .B(_04226_));
 sg13g2_a22oi_1 _22299_ (.Y(_04675_),
    .B1(_04674_),
    .B2(_04230_),
    .A2(_04088_),
    .A1(\cpu.ex.pc[8] ));
 sg13g2_o21ai_1 _22300_ (.B1(_04675_),
    .Y(_00983_),
    .A1(net71),
    .A2(_04672_));
 sg13g2_or2_1 _22301_ (.X(_04676_),
    .B(\cpu.ex.c_mult[9] ),
    .A(_03979_));
 sg13g2_xnor2_1 _22302_ (.Y(_04677_),
    .A(_10900_),
    .B(net208));
 sg13g2_nor3_1 _22303_ (.A(net229),
    .B(_11569_),
    .C(_11568_),
    .Y(_04678_));
 sg13g2_o21ai_1 _22304_ (.B1(net229),
    .Y(_04679_),
    .A1(_11569_),
    .A2(_11568_));
 sg13g2_o21ai_1 _22305_ (.B1(_04679_),
    .Y(_04680_),
    .A1(net165),
    .A2(_04678_));
 sg13g2_xor2_1 _22306_ (.B(_04680_),
    .A(_04677_),
    .X(_04681_));
 sg13g2_nor2_1 _22307_ (.A(net1072),
    .B(_11473_),
    .Y(_04682_));
 sg13g2_a21oi_1 _22308_ (.A1(net871),
    .A2(_11473_),
    .Y(_04683_),
    .B1(_04682_));
 sg13g2_o21ai_1 _22309_ (.B1(_11574_),
    .Y(_04684_),
    .A1(net1063),
    .A2(_04683_));
 sg13g2_nand2_1 _22310_ (.Y(_04685_),
    .A(_09055_),
    .B(_11645_));
 sg13g2_nand2_1 _22311_ (.Y(_04686_),
    .A(_04034_),
    .B(_04567_));
 sg13g2_a221oi_1 _22312_ (.B2(net167),
    .C1(_04686_),
    .B1(net101),
    .A1(_03984_),
    .Y(_04687_),
    .A2(net139));
 sg13g2_nand2_1 _22313_ (.Y(_04688_),
    .A(_04286_),
    .B(_04003_));
 sg13g2_a22oi_1 _22314_ (.Y(_04689_),
    .B1(net106),
    .B2(_04265_),
    .A2(net135),
    .A1(_04128_));
 sg13g2_nand4_1 _22315_ (.B(_04687_),
    .C(_04688_),
    .A(_04485_),
    .Y(_04690_),
    .D(_04689_));
 sg13g2_nand3b_1 _22316_ (.B(_04690_),
    .C(net1062),
    .Y(_04691_),
    .A_N(_04617_));
 sg13g2_a21oi_1 _22317_ (.A1(_11611_),
    .A2(net139),
    .Y(_04692_),
    .B1(_04449_));
 sg13g2_a22oi_1 _22318_ (.Y(_04693_),
    .B1(_03981_),
    .B2(net226),
    .A2(_04136_),
    .A1(_11467_));
 sg13g2_nand2b_1 _22319_ (.Y(_04694_),
    .B(_04140_),
    .A_N(_04693_));
 sg13g2_a22oi_1 _22320_ (.Y(_04695_),
    .B1(_04033_),
    .B2(_11604_),
    .A2(net106),
    .A1(net178));
 sg13g2_nor2_1 _22321_ (.A(_11436_),
    .B(_11226_),
    .Y(_04696_));
 sg13g2_o21ai_1 _22322_ (.B1(net193),
    .Y(_04697_),
    .A1(_03981_),
    .A2(_04696_));
 sg13g2_nand3_1 _22323_ (.B(_11694_),
    .C(_04026_),
    .A(_10872_),
    .Y(_04698_));
 sg13g2_a21o_1 _22324_ (.A2(_04698_),
    .A1(_04697_),
    .B1(_11663_),
    .X(_04699_));
 sg13g2_nand4_1 _22325_ (.B(_04694_),
    .C(_04695_),
    .A(_04692_),
    .Y(_04700_),
    .D(_04699_));
 sg13g2_nand3_1 _22326_ (.B(_04132_),
    .C(_04700_),
    .A(_04456_),
    .Y(_04701_));
 sg13g2_nand4_1 _22327_ (.B(_04685_),
    .C(_04691_),
    .A(_04684_),
    .Y(_04702_),
    .D(_04701_));
 sg13g2_a21oi_1 _22328_ (.A1(net607),
    .A2(_04681_),
    .Y(_04703_),
    .B1(_04702_));
 sg13g2_nand2_1 _22329_ (.Y(_04704_),
    .A(net300),
    .B(_04201_));
 sg13g2_nand2_1 _22330_ (.Y(_04705_),
    .A(net261),
    .B(_04201_));
 sg13g2_a22oi_1 _22331_ (.Y(_04706_),
    .B1(_04704_),
    .B2(_04705_),
    .A2(_04195_),
    .A1(_04186_));
 sg13g2_nor2_1 _22332_ (.A(_04094_),
    .B(_04202_),
    .Y(_04707_));
 sg13g2_nor3_1 _22333_ (.A(_04196_),
    .B(_04706_),
    .C(_04707_),
    .Y(_04708_));
 sg13g2_xnor2_1 _22334_ (.Y(_04709_),
    .A(_04708_),
    .B(_04677_));
 sg13g2_nand2_1 _22335_ (.Y(_04710_),
    .A(net951),
    .B(_04709_));
 sg13g2_nand3_1 _22336_ (.B(_04703_),
    .C(_04710_),
    .A(_04285_),
    .Y(_04711_));
 sg13g2_nand2_1 _22337_ (.Y(_04712_),
    .A(_04676_),
    .B(_04711_));
 sg13g2_buf_1 _22338_ (.A(_08845_),
    .X(_04713_));
 sg13g2_xnor2_1 _22339_ (.Y(_04714_),
    .A(_00287_),
    .B(_04227_));
 sg13g2_a22oi_1 _22340_ (.Y(_04715_),
    .B1(_04714_),
    .B2(net70),
    .A2(_04087_),
    .A1(net985));
 sg13g2_o21ai_1 _22341_ (.B1(_04715_),
    .Y(_00984_),
    .A1(_03976_),
    .A2(_04712_));
 sg13g2_nor2_1 _22342_ (.A(_04211_),
    .B(_04214_),
    .Y(_04716_));
 sg13g2_nand2_1 _22343_ (.Y(_04717_),
    .A(_08242_),
    .B(_04716_));
 sg13g2_o21ai_1 _22344_ (.B1(_08242_),
    .Y(_04718_),
    .A1(_04211_),
    .A2(_04214_));
 sg13g2_o21ai_1 _22345_ (.B1(_04205_),
    .Y(_04719_),
    .A1(_10360_),
    .A2(_04708_));
 sg13g2_mux2_1 _22346_ (.A0(_04717_),
    .A1(_04718_),
    .S(_04719_),
    .X(_04720_));
 sg13g2_or2_1 _22347_ (.X(_04721_),
    .B(_04696_),
    .A(net178));
 sg13g2_o21ai_1 _22348_ (.B1(_03787_),
    .Y(_04722_),
    .A1(_11416_),
    .A2(_03733_));
 sg13g2_a22oi_1 _22349_ (.Y(_04723_),
    .B1(_04722_),
    .B2(net136),
    .A2(_04721_),
    .A1(_03795_));
 sg13g2_nand2_1 _22350_ (.Y(_04724_),
    .A(net171),
    .B(net133));
 sg13g2_a22oi_1 _22351_ (.Y(_04725_),
    .B1(net102),
    .B2(net176),
    .A2(net139),
    .A1(net178));
 sg13g2_a22oi_1 _22352_ (.Y(_04726_),
    .B1(net134),
    .B2(_11604_),
    .A2(_04042_),
    .A1(net1146));
 sg13g2_nand3_1 _22353_ (.B(_04725_),
    .C(_04726_),
    .A(_04724_),
    .Y(_04727_));
 sg13g2_nand2_1 _22354_ (.Y(_04728_),
    .A(_04456_),
    .B(_04727_));
 sg13g2_o21ai_1 _22355_ (.B1(_04728_),
    .Y(_04729_),
    .A1(_04248_),
    .A2(_04723_));
 sg13g2_nand2b_1 _22356_ (.Y(_04730_),
    .B(net139),
    .A_N(_11551_));
 sg13g2_inv_1 _22357_ (.Y(_04731_),
    .A(_04730_));
 sg13g2_a22oi_1 _22358_ (.Y(_04732_),
    .B1(net134),
    .B2(net244),
    .A2(net168),
    .A1(_11472_));
 sg13g2_a22oi_1 _22359_ (.Y(_04733_),
    .B1(net104),
    .B2(_04128_),
    .A2(net135),
    .A1(_04117_));
 sg13g2_a22oi_1 _22360_ (.Y(_04734_),
    .B1(_04036_),
    .B2(net191),
    .A2(_04003_),
    .A1(_04122_));
 sg13g2_a22oi_1 _22361_ (.Y(_04735_),
    .B1(net138),
    .B2(net169),
    .A2(net140),
    .A1(_03984_));
 sg13g2_nand4_1 _22362_ (.B(_04733_),
    .C(_04734_),
    .A(_04732_),
    .Y(_04736_),
    .D(_04735_));
 sg13g2_nor3_1 _22363_ (.A(net87),
    .B(_04731_),
    .C(_04736_),
    .Y(_04737_));
 sg13g2_o21ai_1 _22364_ (.B1(_09844_),
    .Y(_04738_),
    .A1(net245),
    .A2(net86));
 sg13g2_nor2_1 _22365_ (.A(_11585_),
    .B(net255),
    .Y(_04739_));
 sg13g2_mux2_1 _22366_ (.A0(_09092_),
    .A1(net1155),
    .S(_04739_),
    .X(_04740_));
 sg13g2_nor2_1 _22367_ (.A(net1145),
    .B(_04740_),
    .Y(_04741_));
 sg13g2_a21oi_1 _22368_ (.A1(net170),
    .A2(net255),
    .Y(_04742_),
    .B1(_04741_));
 sg13g2_a21oi_1 _22369_ (.A1(net1157),
    .A2(net226),
    .Y(_04743_),
    .B1(_04742_));
 sg13g2_o21ai_1 _22370_ (.B1(_04743_),
    .Y(_04744_),
    .A1(_04737_),
    .A2(_04738_));
 sg13g2_a21oi_1 _22371_ (.A1(_04275_),
    .A2(_04729_),
    .Y(_04745_),
    .B1(_04744_));
 sg13g2_nand4_1 _22372_ (.B(_04110_),
    .C(_04720_),
    .A(net671),
    .Y(_04746_),
    .D(_04745_));
 sg13g2_xor2_1 _22373_ (.B(_04716_),
    .A(_11576_),
    .X(_04747_));
 sg13g2_a21oi_1 _22374_ (.A1(net607),
    .A2(_04747_),
    .Y(_04748_),
    .B1(net213));
 sg13g2_a22oi_1 _22375_ (.Y(_04749_),
    .B1(_04746_),
    .B2(_04748_),
    .A2(\cpu.ex.c_mult[10] ),
    .A1(net190));
 sg13g2_buf_1 _22376_ (.A(_08829_),
    .X(_04750_));
 sg13g2_nand2_1 _22377_ (.Y(_04751_),
    .A(_08845_),
    .B(_04227_));
 sg13g2_xor2_1 _22378_ (.B(_04751_),
    .A(_10136_),
    .X(_04752_));
 sg13g2_a22oi_1 _22379_ (.Y(_04753_),
    .B1(_04752_),
    .B2(net81),
    .A2(_04087_),
    .A1(net984));
 sg13g2_o21ai_1 _22380_ (.B1(_04753_),
    .Y(_00985_),
    .A1(_03976_),
    .A2(_04749_));
 sg13g2_buf_1 _22381_ (.A(_00248_),
    .X(_04754_));
 sg13g2_nor4_1 _22382_ (.A(net1141),
    .B(_10148_),
    .C(_04754_),
    .D(_03605_),
    .Y(_04755_));
 sg13g2_buf_1 _22383_ (.A(_04755_),
    .X(_04756_));
 sg13g2_buf_1 _22384_ (.A(net606),
    .X(_04757_));
 sg13g2_mux2_1 _22385_ (.A0(_10570_),
    .A1(_03619_),
    .S(net521),
    .X(_00988_));
 sg13g2_buf_1 _22386_ (.A(net998),
    .X(_04758_));
 sg13g2_mux2_1 _22387_ (.A0(_10347_),
    .A1(_04758_),
    .S(net521),
    .X(_00989_));
 sg13g2_nand2_1 _22388_ (.Y(_04759_),
    .A(net537),
    .B(net606));
 sg13g2_o21ai_1 _22389_ (.B1(_04759_),
    .Y(_00990_),
    .A1(_11272_),
    .A2(net521));
 sg13g2_mux2_1 _22390_ (.A0(_10791_),
    .A1(net466),
    .S(net521),
    .X(_00991_));
 sg13g2_buf_1 _22391_ (.A(net698),
    .X(_04760_));
 sg13g2_mux2_1 _22392_ (.A0(_10697_),
    .A1(_04760_),
    .S(net521),
    .X(_00992_));
 sg13g2_mux2_1 _22393_ (.A0(_10734_),
    .A1(net527),
    .S(_04757_),
    .X(_00993_));
 sg13g2_mux2_1 _22394_ (.A0(_10529_),
    .A1(net469),
    .S(net521),
    .X(_00994_));
 sg13g2_nand2_1 _22395_ (.Y(_04761_),
    .A(net418),
    .B(net606));
 sg13g2_o21ai_1 _22396_ (.B1(_04761_),
    .Y(_00995_),
    .A1(_11197_),
    .A2(net521));
 sg13g2_mux2_1 _22397_ (.A0(_10457_),
    .A1(net532),
    .S(net606),
    .X(_00996_));
 sg13g2_inv_1 _22398_ (.Y(_04762_),
    .A(_10484_));
 sg13g2_nand2_1 _22399_ (.Y(_04763_),
    .A(net530),
    .B(net606));
 sg13g2_o21ai_1 _22400_ (.B1(_04763_),
    .Y(_00997_),
    .A1(_04762_),
    .A2(net521));
 sg13g2_nand2_1 _22401_ (.Y(_04764_),
    .A(net890),
    .B(_04756_));
 sg13g2_o21ai_1 _22402_ (.B1(_04764_),
    .Y(_00998_),
    .A1(_11149_),
    .A2(_04757_));
 sg13g2_mux2_1 _22403_ (.A0(_10391_),
    .A1(net873),
    .S(net606),
    .X(_00999_));
 sg13g2_mux2_1 _22404_ (.A0(_10301_),
    .A1(net875),
    .S(net606),
    .X(_01000_));
 sg13g2_mux2_1 _22405_ (.A0(_10265_),
    .A1(net874),
    .S(_04756_),
    .X(_01001_));
 sg13g2_buf_1 _22406_ (.A(net1143),
    .X(_04765_));
 sg13g2_mux2_1 _22407_ (.A0(_10211_),
    .A1(_04765_),
    .S(net606),
    .X(_01002_));
 sg13g2_or2_1 _22408_ (.X(_04766_),
    .B(_03605_),
    .A(_11450_));
 sg13g2_buf_1 _22409_ (.A(_04766_),
    .X(_04767_));
 sg13g2_buf_1 _22410_ (.A(_04767_),
    .X(_04768_));
 sg13g2_nor2_1 _22411_ (.A(_08560_),
    .B(_04754_),
    .Y(_04769_));
 sg13g2_nand2_1 _22412_ (.Y(_04770_),
    .A(_03603_),
    .B(_04769_));
 sg13g2_nor2_1 _22413_ (.A(net825),
    .B(_11430_),
    .Y(_04771_));
 sg13g2_a21oi_1 _22414_ (.A1(_11430_),
    .A2(\cpu.ex.r_wb_swapsp ),
    .Y(_04772_),
    .B1(_04771_));
 sg13g2_or4_1 _22415_ (.A(net1141),
    .B(_04754_),
    .C(_03605_),
    .D(_04772_),
    .X(_04773_));
 sg13g2_buf_2 _22416_ (.A(_04773_),
    .X(_04774_));
 sg13g2_buf_1 _22417_ (.A(_04774_),
    .X(_04775_));
 sg13g2_nand2_1 _22418_ (.Y(_04776_),
    .A(\cpu.ex.r_stmp[0] ),
    .B(net415));
 sg13g2_o21ai_1 _22419_ (.B1(_04776_),
    .Y(_01003_),
    .A1(net520),
    .A2(_04770_));
 sg13g2_mux2_1 _22420_ (.A0(net1143),
    .A1(_10211_),
    .S(net520),
    .X(_04777_));
 sg13g2_buf_1 _22421_ (.A(_04774_),
    .X(_04778_));
 sg13g2_mux2_1 _22422_ (.A0(_04777_),
    .A1(\cpu.ex.r_stmp[10] ),
    .S(net414),
    .X(_01004_));
 sg13g2_mux2_1 _22423_ (.A0(net1135),
    .A1(_10347_),
    .S(net520),
    .X(_04779_));
 sg13g2_mux2_1 _22424_ (.A0(_04779_),
    .A1(\cpu.ex.r_stmp[11] ),
    .S(net415),
    .X(_01005_));
 sg13g2_buf_1 _22425_ (.A(_04767_),
    .X(_04780_));
 sg13g2_mux2_1 _22426_ (.A0(net627),
    .A1(\cpu.ex.r_sp[12] ),
    .S(net519),
    .X(_04781_));
 sg13g2_mux2_1 _22427_ (.A0(_04781_),
    .A1(\cpu.ex.r_stmp[12] ),
    .S(net415),
    .X(_01006_));
 sg13g2_mux2_1 _22428_ (.A0(net628),
    .A1(_10791_),
    .S(_04767_),
    .X(_04782_));
 sg13g2_nor2_1 _22429_ (.A(_04774_),
    .B(_04782_),
    .Y(_04783_));
 sg13g2_a21oi_1 _22430_ (.A1(_11304_),
    .A2(net414),
    .Y(_01007_),
    .B1(_04783_));
 sg13g2_mux2_1 _22431_ (.A0(net698),
    .A1(_10697_),
    .S(_04780_),
    .X(_04784_));
 sg13g2_mux2_1 _22432_ (.A0(_04784_),
    .A1(\cpu.ex.r_stmp[14] ),
    .S(_04775_),
    .X(_01008_));
 sg13g2_mux2_1 _22433_ (.A0(net687),
    .A1(_10734_),
    .S(net519),
    .X(_04785_));
 sg13g2_mux2_1 _22434_ (.A0(_04785_),
    .A1(\cpu.ex.r_stmp[15] ),
    .S(net415),
    .X(_01009_));
 sg13g2_nor2_1 _22435_ (.A(_10040_),
    .B(net519),
    .Y(_04786_));
 sg13g2_a21oi_1 _22436_ (.A1(_10570_),
    .A2(net520),
    .Y(_04787_),
    .B1(_04786_));
 sg13g2_nand2_1 _22437_ (.Y(_04788_),
    .A(\cpu.ex.r_stmp[1] ),
    .B(net415));
 sg13g2_o21ai_1 _22438_ (.B1(_04788_),
    .Y(_01010_),
    .A1(net414),
    .A2(_04787_));
 sg13g2_nor2_1 _22439_ (.A(_12122_),
    .B(net519),
    .Y(_04789_));
 sg13g2_a21oi_1 _22440_ (.A1(_10529_),
    .A2(net520),
    .Y(_04790_),
    .B1(_04789_));
 sg13g2_nand2_1 _22441_ (.Y(_04791_),
    .A(\cpu.ex.r_stmp[2] ),
    .B(net415));
 sg13g2_o21ai_1 _22442_ (.B1(_04791_),
    .Y(_01011_),
    .A1(net414),
    .A2(_04790_));
 sg13g2_mux2_1 _22443_ (.A0(net418),
    .A1(\cpu.ex.r_sp[3] ),
    .S(net519),
    .X(_04792_));
 sg13g2_mux2_1 _22444_ (.A0(_04792_),
    .A1(\cpu.ex.r_stmp[3] ),
    .S(net415),
    .X(_01012_));
 sg13g2_nor2_1 _22445_ (.A(net608),
    .B(net519),
    .Y(_04793_));
 sg13g2_a21oi_1 _22446_ (.A1(_10457_),
    .A2(_04768_),
    .Y(_04794_),
    .B1(_04793_));
 sg13g2_nand2_1 _22447_ (.Y(_04795_),
    .A(\cpu.ex.r_stmp[4] ),
    .B(_04775_));
 sg13g2_o21ai_1 _22448_ (.B1(_04795_),
    .Y(_01013_),
    .A1(net414),
    .A2(_04794_));
 sg13g2_nor2_1 _22449_ (.A(_12074_),
    .B(net519),
    .Y(_04796_));
 sg13g2_a21oi_1 _22450_ (.A1(_10484_),
    .A2(_04768_),
    .Y(_04797_),
    .B1(_04796_));
 sg13g2_nand2_1 _22451_ (.Y(_04798_),
    .A(\cpu.ex.r_stmp[5] ),
    .B(net415));
 sg13g2_o21ai_1 _22452_ (.B1(_04798_),
    .Y(_01014_),
    .A1(net414),
    .A2(_04797_));
 sg13g2_inv_1 _22453_ (.Y(_04799_),
    .A(\cpu.ex.r_stmp[6] ));
 sg13g2_mux2_1 _22454_ (.A0(net1000),
    .A1(\cpu.ex.r_sp[6] ),
    .S(_04767_),
    .X(_04800_));
 sg13g2_nor2_1 _22455_ (.A(_04774_),
    .B(_04800_),
    .Y(_04801_));
 sg13g2_a21oi_1 _22456_ (.A1(_04799_),
    .A2(net414),
    .Y(_01015_),
    .B1(_04801_));
 sg13g2_nor2_1 _22457_ (.A(_09167_),
    .B(net519),
    .Y(_04802_));
 sg13g2_a21oi_1 _22458_ (.A1(_10391_),
    .A2(net520),
    .Y(_04803_),
    .B1(_04802_));
 sg13g2_nand2_1 _22459_ (.Y(_04804_),
    .A(\cpu.ex.r_stmp[7] ),
    .B(_04774_));
 sg13g2_o21ai_1 _22460_ (.B1(_04804_),
    .Y(_01016_),
    .A1(net414),
    .A2(_04803_));
 sg13g2_nor2_1 _22461_ (.A(_10920_),
    .B(_04780_),
    .Y(_04805_));
 sg13g2_a21oi_1 _22462_ (.A1(_10301_),
    .A2(net520),
    .Y(_04806_),
    .B1(_04805_));
 sg13g2_nand2_1 _22463_ (.Y(_04807_),
    .A(\cpu.ex.r_stmp[8] ),
    .B(_04774_));
 sg13g2_o21ai_1 _22464_ (.B1(_04807_),
    .Y(_01017_),
    .A1(_04778_),
    .A2(_04806_));
 sg13g2_nor2_1 _22465_ (.A(_10876_),
    .B(_04767_),
    .Y(_04808_));
 sg13g2_a21oi_1 _22466_ (.A1(_10265_),
    .A2(net520),
    .Y(_04809_),
    .B1(_04808_));
 sg13g2_nand2_1 _22467_ (.Y(_04810_),
    .A(\cpu.ex.r_stmp[9] ),
    .B(_04774_));
 sg13g2_o21ai_1 _22468_ (.B1(_04810_),
    .Y(_01018_),
    .A1(_04778_),
    .A2(_04809_));
 sg13g2_nor2_1 _22469_ (.A(\cpu.ex.c_mult[0] ),
    .B(net246),
    .Y(_04811_));
 sg13g2_nor2_1 _22470_ (.A(net242),
    .B(net86),
    .Y(_04812_));
 sg13g2_a22oi_1 _22471_ (.Y(_04813_),
    .B1(_04140_),
    .B2(_11455_),
    .A2(_04447_),
    .A1(_11467_));
 sg13g2_nand2b_1 _22472_ (.Y(_04814_),
    .B(_04416_),
    .A_N(_04813_));
 sg13g2_nor2b_1 _22473_ (.A(net170),
    .B_N(_04028_),
    .Y(_04815_));
 sg13g2_a221oi_1 _22474_ (.B2(_11611_),
    .C1(_04815_),
    .B1(_04017_),
    .A1(_11602_),
    .Y(_04816_),
    .A2(_04016_));
 sg13g2_a21o_1 _22475_ (.A2(_04113_),
    .A1(_04020_),
    .B1(_04653_),
    .X(_04817_));
 sg13g2_a221oi_1 _22476_ (.B2(net244),
    .C1(_04817_),
    .B1(_04036_),
    .A1(net167),
    .Y(_04818_),
    .A2(net168));
 sg13g2_a22oi_1 _22477_ (.Y(_04819_),
    .B1(net142),
    .B2(_10872_),
    .A2(_04123_),
    .A1(_04000_));
 sg13g2_nand3_1 _22478_ (.B(_04730_),
    .C(_04819_),
    .A(_04272_),
    .Y(_04820_));
 sg13g2_a21oi_1 _22479_ (.A1(_04291_),
    .A2(_04003_),
    .Y(_04821_),
    .B1(_04820_));
 sg13g2_nand4_1 _22480_ (.B(_04816_),
    .C(_04818_),
    .A(_04814_),
    .Y(_04822_),
    .D(_04821_));
 sg13g2_a21o_1 _22481_ (.A2(_11420_),
    .A1(net136),
    .B1(_04822_),
    .X(_04823_));
 sg13g2_a22oi_1 _22482_ (.Y(_04824_),
    .B1(_04823_),
    .B2(net1156),
    .A2(_04822_),
    .A1(net1146));
 sg13g2_nand2_1 _22483_ (.Y(_04825_),
    .A(_04063_),
    .B(_04064_));
 sg13g2_nand3_1 _22484_ (.B(net215),
    .C(net189),
    .A(net871),
    .Y(_04826_));
 sg13g2_o21ai_1 _22485_ (.B1(_04826_),
    .Y(_04827_),
    .A1(net189),
    .A2(_04825_));
 sg13g2_nand2b_1 _22486_ (.Y(_04828_),
    .B(_04827_),
    .A_N(net1063));
 sg13g2_nor2_1 _22487_ (.A(net1145),
    .B(_04825_),
    .Y(_04829_));
 sg13g2_o21ai_1 _22488_ (.B1(_11436_),
    .Y(_04830_),
    .A1(_04051_),
    .A2(_04829_));
 sg13g2_a221oi_1 _22489_ (.B2(_04830_),
    .C1(_04053_),
    .B1(_04828_),
    .A1(net1073),
    .Y(_04831_),
    .A2(net233));
 sg13g2_o21ai_1 _22490_ (.B1(_04831_),
    .Y(_04832_),
    .A1(_04812_),
    .A2(_04824_));
 sg13g2_a21o_1 _22491_ (.A2(_11630_),
    .A1(_11617_),
    .B1(_09258_),
    .X(_04833_));
 sg13g2_buf_1 _22492_ (.A(_04833_),
    .X(_04834_));
 sg13g2_nand2_1 _22493_ (.Y(_04835_),
    .A(net247),
    .B(_11622_));
 sg13g2_nor2_2 _22494_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 sg13g2_nand2_1 _22495_ (.Y(_04837_),
    .A(_04832_),
    .B(_04836_));
 sg13g2_buf_1 _22496_ (.A(net175),
    .X(_04838_));
 sg13g2_nand2_1 _22497_ (.Y(_04839_),
    .A(_08378_),
    .B(_11636_));
 sg13g2_buf_2 _22498_ (.A(_04839_),
    .X(_04840_));
 sg13g2_buf_2 _22499_ (.A(\cpu.gpio.r_uart_rx_src[0] ),
    .X(_04841_));
 sg13g2_nor3_1 _22500_ (.A(net1061),
    .B(net1069),
    .C(_09556_),
    .Y(_04842_));
 sg13g2_buf_1 _22501_ (.A(_04842_),
    .X(_04843_));
 sg13g2_buf_1 _22502_ (.A(_09563_),
    .X(_04844_));
 sg13g2_buf_1 _22503_ (.A(net982),
    .X(_04845_));
 sg13g2_nor2_1 _22504_ (.A(net923),
    .B(net924),
    .Y(_04846_));
 sg13g2_buf_1 _22505_ (.A(_04846_),
    .X(_04847_));
 sg13g2_nand2_1 _22506_ (.Y(_04848_),
    .A(_04845_),
    .B(_04847_));
 sg13g2_inv_1 _22507_ (.Y(_04849_),
    .A(_04848_));
 sg13g2_buf_2 _22508_ (.A(\cpu.gpio.r_spi_miso_src[0][0] ),
    .X(_04850_));
 sg13g2_a22oi_1 _22509_ (.Y(_04851_),
    .B1(_04849_),
    .B2(_04850_),
    .A2(net670),
    .A1(_04841_));
 sg13g2_buf_1 _22510_ (.A(_09443_),
    .X(_04852_));
 sg13g2_buf_2 _22511_ (.A(\cpu.gpio.r_src_o[6][0] ),
    .X(_04853_));
 sg13g2_nand3_1 _22512_ (.B(net676),
    .C(_04853_),
    .A(net899),
    .Y(_04854_));
 sg13g2_nand3_1 _22513_ (.B(net900),
    .C(net923),
    .A(_09149_),
    .Y(_04855_));
 sg13g2_nand2_1 _22514_ (.Y(_04856_),
    .A(_04854_),
    .B(_04855_));
 sg13g2_nand3_1 _22515_ (.B(net669),
    .C(_04856_),
    .A(net533),
    .Y(_04857_));
 sg13g2_buf_2 _22516_ (.A(\cpu.gpio.r_src_o[4][0] ),
    .X(_04858_));
 sg13g2_buf_1 _22517_ (.A(_09335_),
    .X(_04859_));
 sg13g2_nand2_1 _22518_ (.Y(_04860_),
    .A(net817),
    .B(_09888_));
 sg13g2_buf_1 _22519_ (.A(_04860_),
    .X(_04861_));
 sg13g2_nor3_1 _22520_ (.A(net982),
    .B(net747),
    .C(net604),
    .Y(_04862_));
 sg13g2_buf_1 _22521_ (.A(_04862_),
    .X(_04863_));
 sg13g2_nand2_1 _22522_ (.Y(_04864_),
    .A(_04858_),
    .B(_04863_));
 sg13g2_buf_2 _22523_ (.A(\cpu.gpio.r_src_io[6][0] ),
    .X(_04865_));
 sg13g2_nand2_2 _22524_ (.Y(_04866_),
    .A(net817),
    .B(_09177_));
 sg13g2_nand2_1 _22525_ (.Y(_04867_),
    .A(_09454_),
    .B(net715));
 sg13g2_buf_1 _22526_ (.A(_04867_),
    .X(_04868_));
 sg13g2_nor3_2 _22527_ (.A(_04845_),
    .B(_04866_),
    .C(net518),
    .Y(_04869_));
 sg13g2_nor3_1 _22528_ (.A(net982),
    .B(net604),
    .C(net518),
    .Y(_04870_));
 sg13g2_buf_1 _22529_ (.A(_04870_),
    .X(_04871_));
 sg13g2_buf_2 _22530_ (.A(\cpu.gpio.r_src_io[4][0] ),
    .X(_04872_));
 sg13g2_a22oi_1 _22531_ (.Y(_04873_),
    .B1(net413),
    .B2(_04872_),
    .A2(_04869_),
    .A1(_04865_));
 sg13g2_nand4_1 _22532_ (.B(_04857_),
    .C(_04864_),
    .A(_04851_),
    .Y(_04874_),
    .D(_04873_));
 sg13g2_nand2_1 _22533_ (.Y(_04875_),
    .A(net925),
    .B(_09564_));
 sg13g2_nand2_1 _22534_ (.Y(_04876_),
    .A(net648),
    .B(_04844_));
 sg13g2_a21oi_1 _22535_ (.A1(_04875_),
    .A2(_04876_),
    .Y(_04877_),
    .B1(net926));
 sg13g2_o21ai_1 _22536_ (.B1(_09563_),
    .Y(_04878_),
    .A1(_09177_),
    .A2(net925));
 sg13g2_nor2_1 _22537_ (.A(_09893_),
    .B(net715),
    .Y(_04879_));
 sg13g2_and2_1 _22538_ (.A(_09893_),
    .B(net648),
    .X(_04880_));
 sg13g2_a21oi_1 _22539_ (.A1(_04878_),
    .A2(_04879_),
    .Y(_04881_),
    .B1(_04880_));
 sg13g2_a21o_1 _22540_ (.A2(_04879_),
    .A1(_09564_),
    .B1(_09568_),
    .X(_04882_));
 sg13g2_nand2_1 _22541_ (.Y(_04883_),
    .A(net771),
    .B(_09563_));
 sg13g2_o21ai_1 _22542_ (.B1(_04875_),
    .Y(_04884_),
    .A1(_04860_),
    .A2(_04883_));
 sg13g2_a22oi_1 _22543_ (.Y(_04885_),
    .B1(_04884_),
    .B2(net1061),
    .A2(_04882_),
    .A1(net1069));
 sg13g2_o21ai_1 _22544_ (.B1(_04885_),
    .Y(_04886_),
    .A1(net716),
    .A2(_04881_));
 sg13g2_or2_1 _22545_ (.X(_04887_),
    .B(_04886_),
    .A(_04877_));
 sg13g2_buf_2 _22546_ (.A(_04887_),
    .X(_04888_));
 sg13g2_nor3_1 _22547_ (.A(net817),
    .B(net1069),
    .C(net518),
    .Y(_04889_));
 sg13g2_and2_1 _22548_ (.A(_11080_),
    .B(_04889_),
    .X(_04890_));
 sg13g2_buf_1 _22549_ (.A(_04890_),
    .X(_04891_));
 sg13g2_a21oi_1 _22550_ (.A1(_09149_),
    .A2(_04888_),
    .Y(_04892_),
    .B1(_04891_));
 sg13g2_nor2b_1 _22551_ (.A(_04892_),
    .B_N(\cpu.gpio.r_enable_in[0] ),
    .Y(_04893_));
 sg13g2_nand2_1 _22552_ (.Y(_04894_),
    .A(_10920_),
    .B(net1154));
 sg13g2_nor2_1 _22553_ (.A(_09164_),
    .B(_04894_),
    .Y(_04895_));
 sg13g2_buf_1 _22554_ (.A(_04895_),
    .X(_04896_));
 sg13g2_o21ai_1 _22555_ (.B1(_04896_),
    .Y(_04897_),
    .A1(_04874_),
    .A2(_04893_));
 sg13g2_nor2_1 _22556_ (.A(_09114_),
    .B(_09115_),
    .Y(_04898_));
 sg13g2_nand2_1 _22557_ (.Y(_04899_),
    .A(net926),
    .B(_09177_));
 sg13g2_buf_1 _22558_ (.A(_04899_),
    .X(_04900_));
 sg13g2_a21oi_1 _22559_ (.A1(net604),
    .A2(_04900_),
    .Y(_04901_),
    .B1(net648));
 sg13g2_nor2_1 _22560_ (.A(net925),
    .B(_04901_),
    .Y(_04902_));
 sg13g2_buf_2 _22561_ (.A(_04902_),
    .X(_04903_));
 sg13g2_nor2_1 _22562_ (.A(net747),
    .B(net668),
    .Y(_04904_));
 sg13g2_buf_1 _22563_ (.A(_04904_),
    .X(_04905_));
 sg13g2_a21oi_1 _22564_ (.A1(_09116_),
    .A2(_04903_),
    .Y(_04906_),
    .B1(net517));
 sg13g2_a22oi_1 _22565_ (.Y(_04907_),
    .B1(net420),
    .B2(\cpu.intr.r_timer_reload[16] ),
    .A2(net422),
    .A1(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_inv_1 _22566_ (.Y(_04908_),
    .A(_00278_));
 sg13g2_a221oi_1 _22567_ (.B2(_04908_),
    .C1(net796),
    .B1(net380),
    .A1(\cpu.intr.r_clock_cmp[0] ),
    .Y(_04909_),
    .A2(net422));
 sg13g2_a21oi_1 _22568_ (.A1(net695),
    .A2(_04907_),
    .Y(_04910_),
    .B1(_04909_));
 sg13g2_nand3_1 _22569_ (.B(_09904_),
    .C(net380),
    .A(net676),
    .Y(_04911_));
 sg13g2_nor2_1 _22570_ (.A(net747),
    .B(net604),
    .Y(_04912_));
 sg13g2_buf_2 _22571_ (.A(_04912_),
    .X(_04913_));
 sg13g2_nor2_1 _22572_ (.A(net771),
    .B(net648),
    .Y(_04914_));
 sg13g2_nor2_2 _22573_ (.A(net817),
    .B(_09888_),
    .Y(_04915_));
 sg13g2_and2_1 _22574_ (.A(_04914_),
    .B(_04915_),
    .X(_04916_));
 sg13g2_buf_1 _22575_ (.A(_04916_),
    .X(_04917_));
 sg13g2_buf_2 _22576_ (.A(_04917_),
    .X(_04918_));
 sg13g2_buf_1 _22577_ (.A(\cpu.intr.r_clock_count[16] ),
    .X(_04919_));
 sg13g2_a22oi_1 _22578_ (.Y(_04920_),
    .B1(net376),
    .B2(_04919_),
    .A2(_04913_),
    .A1(_09116_));
 sg13g2_nor2_1 _22579_ (.A(net796),
    .B(_09892_),
    .Y(_04921_));
 sg13g2_nor2_1 _22580_ (.A(_09178_),
    .B(_10031_),
    .Y(_04922_));
 sg13g2_buf_1 _22581_ (.A(_04922_),
    .X(_04923_));
 sg13g2_a22oi_1 _22582_ (.Y(_04924_),
    .B1(net412),
    .B2(_10036_),
    .A2(_04921_),
    .A1(\cpu.intr.r_timer_reload[0] ));
 sg13g2_nand3_1 _22583_ (.B(_04920_),
    .C(_04924_),
    .A(_04911_),
    .Y(_04925_));
 sg13g2_nor2_1 _22584_ (.A(_04910_),
    .B(_04925_),
    .Y(_04926_));
 sg13g2_o21ai_1 _22585_ (.B1(_04926_),
    .Y(_04927_),
    .A1(_04898_),
    .A2(_04906_));
 sg13g2_nor2_1 _22586_ (.A(net931),
    .B(_09556_),
    .Y(_04928_));
 sg13g2_buf_1 _22587_ (.A(_04928_),
    .X(_04929_));
 sg13g2_buf_1 _22588_ (.A(_04889_),
    .X(_04930_));
 sg13g2_buf_1 _22589_ (.A(net411),
    .X(_04931_));
 sg13g2_nor3_1 _22590_ (.A(_00295_),
    .B(net518),
    .C(net668),
    .Y(_04932_));
 sg13g2_a221oi_1 _22591_ (.B2(_12105_),
    .C1(_04932_),
    .B1(_04931_),
    .A1(\cpu.spi.r_mode[1][0] ),
    .Y(_04933_),
    .A2(net667));
 sg13g2_nand2_1 _22592_ (.Y(_04934_),
    .A(net648),
    .B(_04875_));
 sg13g2_or2_1 _22593_ (.X(_04935_),
    .B(_09171_),
    .A(net648));
 sg13g2_o21ai_1 _22594_ (.B1(_04935_),
    .Y(_04936_),
    .A1(net817),
    .A2(_04883_));
 sg13g2_a21oi_1 _22595_ (.A1(net817),
    .A2(_09191_),
    .Y(_04937_),
    .B1(_09346_));
 sg13g2_nor2_1 _22596_ (.A(net1069),
    .B(_04937_),
    .Y(_04938_));
 sg13g2_a221oi_1 _22597_ (.B2(_09178_),
    .C1(_04938_),
    .B1(_04936_),
    .A1(net926),
    .Y(_04939_),
    .A2(_04934_));
 sg13g2_nor3_1 _22598_ (.A(_09894_),
    .B(net518),
    .C(_04899_),
    .Y(_04940_));
 sg13g2_buf_1 _22599_ (.A(_04940_),
    .X(_04941_));
 sg13g2_nor3_1 _22600_ (.A(net670),
    .B(_04939_),
    .C(net410),
    .Y(_04942_));
 sg13g2_buf_2 _22601_ (.A(_04942_),
    .X(_04943_));
 sg13g2_a22oi_1 _22602_ (.Y(_04944_),
    .B1(\cpu.spi.r_timeout[0] ),
    .B2(net493),
    .A2(_09171_),
    .A1(_09119_));
 sg13g2_inv_1 _22603_ (.Y(_04945_),
    .A(\cpu.spi.r_ready ));
 sg13g2_or3_1 _22604_ (.A(net796),
    .B(net493),
    .C(_04945_),
    .X(_04946_));
 sg13g2_o21ai_1 _22605_ (.B1(_04946_),
    .Y(_04947_),
    .A1(net923),
    .A2(_04944_));
 sg13g2_nand3_1 _22606_ (.B(net982),
    .C(net544),
    .A(net1069),
    .Y(_04948_));
 sg13g2_buf_2 _22607_ (.A(_04948_),
    .X(_04949_));
 sg13g2_buf_1 _22608_ (.A(\cpu.spi.r_clk_count[2][0] ),
    .X(_04950_));
 sg13g2_nor3_1 _22609_ (.A(net982),
    .B(net518),
    .C(net668),
    .Y(_04951_));
 sg13g2_buf_2 _22610_ (.A(_04951_),
    .X(_04952_));
 sg13g2_and2_1 _22611_ (.A(net1061),
    .B(\cpu.spi.r_mode[2][0] ),
    .X(_04953_));
 sg13g2_a22oi_1 _22612_ (.Y(_04954_),
    .B1(_04953_),
    .B2(net411),
    .A2(_04952_),
    .A1(_04950_));
 sg13g2_o21ai_1 _22613_ (.B1(_04954_),
    .Y(_04955_),
    .A1(_00294_),
    .A2(_04949_));
 sg13g2_a221oi_1 _22614_ (.B2(net622),
    .C1(_04955_),
    .B1(_04947_),
    .A1(_09217_),
    .Y(_04956_),
    .A2(_04943_));
 sg13g2_o21ai_1 _22615_ (.B1(_04956_),
    .Y(_04957_),
    .A1(net769),
    .A2(_04933_));
 sg13g2_nand2_1 _22616_ (.Y(_04958_),
    .A(_09164_),
    .B(_09895_));
 sg13g2_buf_1 _22617_ (.A(_04958_),
    .X(_04959_));
 sg13g2_nand2_1 _22618_ (.Y(_04960_),
    .A(_04894_),
    .B(_04959_));
 sg13g2_buf_1 _22619_ (.A(_04960_),
    .X(_04961_));
 sg13g2_buf_1 _22620_ (.A(_09513_),
    .X(_04962_));
 sg13g2_o21ai_1 _22621_ (.B1(_12075_),
    .Y(_04963_),
    .A1(_04962_),
    .A2(_09517_));
 sg13g2_buf_2 _22622_ (.A(_04963_),
    .X(_04964_));
 sg13g2_nor2_1 _22623_ (.A(_04868_),
    .B(_04899_),
    .Y(_04965_));
 sg13g2_buf_1 _22624_ (.A(_04965_),
    .X(_04966_));
 sg13g2_nor2_1 _22625_ (.A(net747),
    .B(_04866_),
    .Y(_04967_));
 sg13g2_buf_1 _22626_ (.A(_04967_),
    .X(_04968_));
 sg13g2_buf_2 _22627_ (.A(\cpu.uart.r_x_invert ),
    .X(_04969_));
 sg13g2_a22oi_1 _22628_ (.Y(_04970_),
    .B1(net515),
    .B2(_04969_),
    .A2(net409),
    .A1(\cpu.uart.r_div_value[8] ));
 sg13g2_a22oi_1 _22629_ (.Y(_04971_),
    .B1(_04930_),
    .B2(\cpu.uart.r_div_value[0] ),
    .A2(_04913_),
    .A1(_09114_));
 sg13g2_nand2_1 _22630_ (.Y(_04972_),
    .A(_04970_),
    .B(_04971_));
 sg13g2_a21oi_1 _22631_ (.A1(\cpu.uart.r_in[0] ),
    .A2(_04964_),
    .Y(_04973_),
    .B1(_04972_));
 sg13g2_o21ai_1 _22632_ (.B1(net1166),
    .Y(_04974_),
    .A1(net516),
    .A2(_04973_));
 sg13g2_a221oi_1 _22633_ (.B2(_09170_),
    .C1(_04974_),
    .B1(_04957_),
    .A1(_09897_),
    .Y(_04975_),
    .A2(_04927_));
 sg13g2_nand2_1 _22634_ (.Y(_04976_),
    .A(net1081),
    .B(net1067));
 sg13g2_nor3_1 _22635_ (.A(net994),
    .B(net1161),
    .C(_04976_),
    .Y(_04977_));
 sg13g2_buf_2 _22636_ (.A(_04977_),
    .X(_04978_));
 sg13g2_a22oi_1 _22637_ (.Y(_04979_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][16] ),
    .A2(net638),
    .A1(\cpu.dcache.r_data[0][16] ));
 sg13g2_a22oi_1 _22638_ (.Y(_04980_),
    .B1(net567),
    .B2(\cpu.dcache.r_data[4][16] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[1][16] ));
 sg13g2_a22oi_1 _22639_ (.Y(_04981_),
    .B1(net546),
    .B2(\cpu.dcache.r_data[3][16] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[6][16] ));
 sg13g2_a22oi_1 _22640_ (.Y(_04982_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][16] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[5][16] ));
 sg13g2_and4_1 _22641_ (.A(_04979_),
    .B(_04980_),
    .C(_04981_),
    .D(_04982_),
    .X(_04983_));
 sg13g2_nor2_1 _22642_ (.A(net923),
    .B(_04983_),
    .Y(_04984_));
 sg13g2_a21o_1 _22643_ (.A2(net994),
    .A1(_10984_),
    .B1(_04976_),
    .X(_04985_));
 sg13g2_buf_1 _22644_ (.A(_04985_),
    .X(_04986_));
 sg13g2_mux2_1 _22645_ (.A0(\cpu.dcache.r_data[1][24] ),
    .A1(\cpu.dcache.r_data[3][24] ),
    .S(net569),
    .X(_04987_));
 sg13g2_a22oi_1 _22646_ (.Y(_04988_),
    .B1(_04987_),
    .B2(net716),
    .A2(net666),
    .A1(\cpu.dcache.r_data[2][24] ));
 sg13g2_inv_1 _22647_ (.Y(_04989_),
    .A(_00292_));
 sg13g2_mux2_1 _22648_ (.A0(\cpu.dcache.r_data[4][24] ),
    .A1(\cpu.dcache.r_data[6][24] ),
    .S(_09191_),
    .X(_04990_));
 sg13g2_a22oi_1 _22649_ (.Y(_04991_),
    .B1(_04990_),
    .B2(net767),
    .A2(_09517_),
    .A1(\cpu.dcache.r_data[5][24] ));
 sg13g2_nor2_1 _22650_ (.A(net771),
    .B(_04991_),
    .Y(_04992_));
 sg13g2_a221oi_1 _22651_ (.B2(\cpu.dcache.r_data[7][24] ),
    .C1(_04992_),
    .B1(_03045_),
    .A1(_04989_),
    .Y(_04993_),
    .A2(_09641_));
 sg13g2_o21ai_1 _22652_ (.B1(_04993_),
    .Y(_04994_),
    .A1(_09511_),
    .A2(_04988_));
 sg13g2_nor2b_1 _22653_ (.A(net665),
    .B_N(_04994_),
    .Y(_04995_));
 sg13g2_a21oi_1 _22654_ (.A1(_04984_),
    .A2(net665),
    .Y(_04996_),
    .B1(_04995_));
 sg13g2_inv_1 _22655_ (.Y(_04997_),
    .A(_00293_));
 sg13g2_a22oi_1 _22656_ (.Y(_04998_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][8] ),
    .A2(net638),
    .A1(_04997_));
 sg13g2_a22oi_1 _22657_ (.Y(_04999_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][8] ),
    .A2(net543),
    .A1(\cpu.dcache.r_data[7][8] ));
 sg13g2_a22oi_1 _22658_ (.Y(_05000_),
    .B1(net567),
    .B2(\cpu.dcache.r_data[4][8] ),
    .A2(net548),
    .A1(\cpu.dcache.r_data[1][8] ));
 sg13g2_a22oi_1 _22659_ (.Y(_05001_),
    .B1(net481),
    .B2(\cpu.dcache.r_data[3][8] ),
    .A2(net479),
    .A1(\cpu.dcache.r_data[6][8] ));
 sg13g2_nand4_1 _22660_ (.B(_04999_),
    .C(_05000_),
    .A(_04998_),
    .Y(_05002_),
    .D(_05001_));
 sg13g2_nor2_1 _22661_ (.A(_12224_),
    .B(net665),
    .Y(_05003_));
 sg13g2_and2_1 _22662_ (.A(_12139_),
    .B(net665),
    .X(_05004_));
 sg13g2_buf_1 _22663_ (.A(_05004_),
    .X(_05005_));
 sg13g2_nand2_1 _22664_ (.Y(_05006_),
    .A(\cpu.dcache.r_data[4][0] ),
    .B(net640));
 sg13g2_a22oi_1 _22665_ (.Y(_05007_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][0] ),
    .A2(net644),
    .A1(\cpu.dcache.r_data[6][0] ));
 sg13g2_a22oi_1 _22666_ (.Y(_05008_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][0] ),
    .A2(net639),
    .A1(\cpu.dcache.r_data[5][0] ));
 sg13g2_a22oi_1 _22667_ (.Y(_05009_),
    .B1(_03031_),
    .B2(\cpu.dcache.r_data[3][0] ),
    .A2(net643),
    .A1(\cpu.dcache.r_data[1][0] ));
 sg13g2_nand4_1 _22668_ (.B(_05007_),
    .C(_05008_),
    .A(_05006_),
    .Y(_05010_),
    .D(_05009_));
 sg13g2_mux2_1 _22669_ (.A0(\cpu.dcache.r_data[0][0] ),
    .A1(_05010_),
    .S(_09460_),
    .X(_05011_));
 sg13g2_buf_1 _22670_ (.A(_05011_),
    .X(_05012_));
 sg13g2_a22oi_1 _22671_ (.Y(_05013_),
    .B1(_05005_),
    .B2(_05012_),
    .A2(_05003_),
    .A1(_05002_));
 sg13g2_o21ai_1 _22672_ (.B1(_05013_),
    .Y(_05014_),
    .A1(net1030),
    .A2(_04996_));
 sg13g2_a21oi_1 _22673_ (.A1(net798),
    .A2(_05012_),
    .Y(_05015_),
    .B1(_04984_));
 sg13g2_nand2_1 _22674_ (.Y(_05016_),
    .A(_05015_),
    .B(_04978_));
 sg13g2_o21ai_1 _22675_ (.B1(_05016_),
    .Y(_05017_),
    .A1(_04978_),
    .A2(_05014_));
 sg13g2_a221oi_1 _22676_ (.B2(net1067),
    .C1(_04840_),
    .B1(_05017_),
    .A1(_04897_),
    .Y(_05018_),
    .A2(_04975_));
 sg13g2_a21oi_1 _22677_ (.A1(net992),
    .A2(_04840_),
    .Y(_05019_),
    .B1(_05018_));
 sg13g2_nand3_1 _22678_ (.B(net175),
    .C(_04835_),
    .A(net993),
    .Y(_05020_));
 sg13g2_o21ai_1 _22679_ (.B1(_05020_),
    .Y(_05021_),
    .A1(net132),
    .A2(_05019_));
 sg13g2_inv_1 _22680_ (.Y(_05022_),
    .A(_05021_));
 sg13g2_o21ai_1 _22681_ (.B1(_05022_),
    .Y(_01019_),
    .A1(_04811_),
    .A2(_04837_));
 sg13g2_buf_1 _22682_ (.A(net164),
    .X(_05023_));
 sg13g2_buf_1 _22683_ (.A(_04840_),
    .X(_05024_));
 sg13g2_buf_2 _22684_ (.A(_04840_),
    .X(_05025_));
 sg13g2_or3_1 _22685_ (.A(net994),
    .B(net1161),
    .C(_04976_),
    .X(_05026_));
 sg13g2_buf_1 _22686_ (.A(_05026_),
    .X(_05027_));
 sg13g2_inv_1 _22687_ (.Y(_05028_),
    .A(_00145_));
 sg13g2_a22oi_1 _22688_ (.Y(_05029_),
    .B1(net639),
    .B2(\cpu.dcache.r_data[5][7] ),
    .A2(net638),
    .A1(_05028_));
 sg13g2_a22oi_1 _22689_ (.Y(_05030_),
    .B1(net643),
    .B2(\cpu.dcache.r_data[1][7] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[6][7] ));
 sg13g2_a22oi_1 _22690_ (.Y(_05031_),
    .B1(net640),
    .B2(\cpu.dcache.r_data[4][7] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][7] ));
 sg13g2_a22oi_1 _22691_ (.Y(_05032_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][7] ),
    .A2(net621),
    .A1(\cpu.dcache.r_data[7][7] ));
 sg13g2_nand4_1 _22692_ (.B(_05030_),
    .C(_05031_),
    .A(_05029_),
    .Y(_05033_),
    .D(_05032_));
 sg13g2_buf_1 _22693_ (.A(_05033_),
    .X(_05034_));
 sg13g2_inv_1 _22694_ (.Y(_05035_),
    .A(_00146_));
 sg13g2_a22oi_1 _22695_ (.Y(_05036_),
    .B1(net639),
    .B2(\cpu.dcache.r_data[5][23] ),
    .A2(net638),
    .A1(_05035_));
 sg13g2_a22oi_1 _22696_ (.Y(_05037_),
    .B1(net643),
    .B2(\cpu.dcache.r_data[1][23] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[6][23] ));
 sg13g2_a22oi_1 _22697_ (.Y(_05038_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][23] ),
    .A2(net640),
    .A1(\cpu.dcache.r_data[4][23] ));
 sg13g2_a22oi_1 _22698_ (.Y(_05039_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][23] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][23] ));
 sg13g2_nand4_1 _22699_ (.B(_05037_),
    .C(_05038_),
    .A(_05036_),
    .Y(_05040_),
    .D(_05039_));
 sg13g2_buf_1 _22700_ (.A(_05040_),
    .X(_05041_));
 sg13g2_nor2_2 _22701_ (.A(_09888_),
    .B(_12139_),
    .Y(_05042_));
 sg13g2_a22oi_1 _22702_ (.Y(_05043_),
    .B1(_05041_),
    .B2(_05042_),
    .A2(_05034_),
    .A1(_12139_));
 sg13g2_a22oi_1 _22703_ (.Y(_05044_),
    .B1(net546),
    .B2(\cpu.dcache.r_data[3][15] ),
    .A2(net644),
    .A1(\cpu.dcache.r_data[6][15] ));
 sg13g2_a22oi_1 _22704_ (.Y(_05045_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][15] ),
    .A2(net640),
    .A1(\cpu.dcache.r_data[4][15] ));
 sg13g2_a22oi_1 _22705_ (.Y(_05046_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][15] ),
    .A2(net639),
    .A1(\cpu.dcache.r_data[5][15] ));
 sg13g2_nand3_1 _22706_ (.B(_05045_),
    .C(_05046_),
    .A(_05044_),
    .Y(_05047_));
 sg13g2_nand2_1 _22707_ (.Y(_05048_),
    .A(_00148_),
    .B(net669));
 sg13g2_o21ai_1 _22708_ (.B1(_05048_),
    .Y(_05049_),
    .A1(net669),
    .A2(_05047_));
 sg13g2_o21ai_1 _22709_ (.B1(net548),
    .Y(_05050_),
    .A1(\cpu.dcache.r_data[1][15] ),
    .A2(_05047_));
 sg13g2_o21ai_1 _22710_ (.B1(_05050_),
    .Y(_05051_),
    .A1(net548),
    .A2(_05049_));
 sg13g2_inv_1 _22711_ (.Y(_05052_),
    .A(_00147_));
 sg13g2_a22oi_1 _22712_ (.Y(_05053_),
    .B1(_03027_),
    .B2(\cpu.dcache.r_data[2][31] ),
    .A2(net638),
    .A1(_05052_));
 sg13g2_a22oi_1 _22713_ (.Y(_05054_),
    .B1(net548),
    .B2(\cpu.dcache.r_data[1][31] ),
    .A2(_03040_),
    .A1(\cpu.dcache.r_data[6][31] ));
 sg13g2_a22oi_1 _22714_ (.Y(_05055_),
    .B1(_03045_),
    .B2(\cpu.dcache.r_data[7][31] ),
    .A2(net639),
    .A1(\cpu.dcache.r_data[5][31] ));
 sg13g2_a22oi_1 _22715_ (.Y(_05056_),
    .B1(net640),
    .B2(\cpu.dcache.r_data[4][31] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][31] ));
 sg13g2_nand4_1 _22716_ (.B(_05054_),
    .C(_05055_),
    .A(_05053_),
    .Y(_05057_),
    .D(_05056_));
 sg13g2_a221oi_1 _22717_ (.B2(net898),
    .C1(net665),
    .B1(_05057_),
    .A1(net923),
    .Y(_05058_),
    .A2(_05051_));
 sg13g2_a21oi_1 _22718_ (.A1(net665),
    .A2(_05043_),
    .Y(_05059_),
    .B1(_05058_));
 sg13g2_nor2_1 _22719_ (.A(_10025_),
    .B(_05034_),
    .Y(_05060_));
 sg13g2_nor2_1 _22720_ (.A(_09889_),
    .B(_05041_),
    .Y(_05061_));
 sg13g2_nor3_1 _22721_ (.A(_05027_),
    .B(_05060_),
    .C(_05061_),
    .Y(_05062_));
 sg13g2_a21oi_1 _22722_ (.A1(_05027_),
    .A2(_05059_),
    .Y(_05063_),
    .B1(_05062_));
 sg13g2_a22oi_1 _22723_ (.Y(_05064_),
    .B1(_04964_),
    .B2(\cpu.uart.r_in[7] ),
    .A2(_04930_),
    .A1(\cpu.uart.r_div_value[7] ));
 sg13g2_and2_1 _22724_ (.A(net931),
    .B(\cpu.intr.r_clock_cmp[23] ),
    .X(_05065_));
 sg13g2_a21oi_1 _22725_ (.A1(_09888_),
    .A2(\cpu.intr.r_clock_cmp[7] ),
    .Y(_05066_),
    .B1(_05065_));
 sg13g2_buf_1 _22726_ (.A(\cpu.intr.r_clock_count[23] ),
    .X(_05067_));
 sg13g2_mux2_1 _22727_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(\cpu.intr.r_timer_reload[23] ),
    .S(net931),
    .X(_05068_));
 sg13g2_a22oi_1 _22728_ (.Y(_05069_),
    .B1(_05068_),
    .B2(net543),
    .A2(net376),
    .A1(_05067_));
 sg13g2_o21ai_1 _22729_ (.B1(_05069_),
    .Y(_05070_),
    .A1(net924),
    .A2(_05066_));
 sg13g2_a22oi_1 _22730_ (.Y(_05071_),
    .B1(net567),
    .B2(_10072_),
    .A2(net544),
    .A1(_09906_));
 sg13g2_nand3_1 _22731_ (.B(_09926_),
    .C(net479),
    .A(net931),
    .Y(_05072_));
 sg13g2_o21ai_1 _22732_ (.B1(_05072_),
    .Y(_05073_),
    .A1(net931),
    .A2(_05071_));
 sg13g2_nor2_1 _22733_ (.A(_04959_),
    .B(_04903_),
    .Y(_05074_));
 sg13g2_o21ai_1 _22734_ (.B1(_05074_),
    .Y(_05075_),
    .A1(_05070_),
    .A2(_05073_));
 sg13g2_o21ai_1 _22735_ (.B1(_05075_),
    .Y(_05076_),
    .A1(net516),
    .A2(_05064_));
 sg13g2_inv_1 _22736_ (.Y(_05077_),
    .A(_04896_));
 sg13g2_buf_1 _22737_ (.A(\cpu.gpio.r_src_io[5][3] ),
    .X(_05078_));
 sg13g2_or3_1 _22738_ (.A(net982),
    .B(_04866_),
    .C(net518),
    .X(_05079_));
 sg13g2_buf_1 _22739_ (.A(_05079_),
    .X(_05080_));
 sg13g2_nand2_1 _22740_ (.Y(_05081_),
    .A(_09139_),
    .B(_11080_));
 sg13g2_o21ai_1 _22741_ (.B1(_05081_),
    .Y(_05082_),
    .A1(net982),
    .A2(_00153_));
 sg13g2_and2_1 _22742_ (.A(_09132_),
    .B(net982),
    .X(_05083_));
 sg13g2_a22oi_1 _22743_ (.Y(_05084_),
    .B1(_05083_),
    .B2(net515),
    .A2(_05082_),
    .A1(_04913_));
 sg13g2_o21ai_1 _22744_ (.B1(_05084_),
    .Y(_05085_),
    .A1(_00151_),
    .A2(_05080_));
 sg13g2_a221oi_1 _22745_ (.B2(_09138_),
    .C1(_05085_),
    .B1(_04891_),
    .A1(_05078_),
    .Y(_05086_),
    .A2(net413));
 sg13g2_or2_1 _22746_ (.X(_05087_),
    .B(_04866_),
    .A(net747));
 sg13g2_buf_1 _22747_ (.A(_05087_),
    .X(_05088_));
 sg13g2_nor2_1 _22748_ (.A(_00152_),
    .B(_05088_),
    .Y(_05089_));
 sg13g2_nor3_1 _22749_ (.A(_00154_),
    .B(net747),
    .C(net668),
    .Y(_05090_));
 sg13g2_o21ai_1 _22750_ (.B1(net1061),
    .Y(_05091_),
    .A1(_05089_),
    .A2(_05090_));
 sg13g2_nand2b_1 _22751_ (.Y(_05092_),
    .B(net1069),
    .A_N(_00155_));
 sg13g2_nand2_1 _22752_ (.Y(_05093_),
    .A(_09888_),
    .B(net10));
 sg13g2_a21oi_1 _22753_ (.A1(_05092_),
    .A2(_05093_),
    .Y(_05094_),
    .B1(net924));
 sg13g2_a221oi_1 _22754_ (.B2(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .C1(_05094_),
    .B1(net412),
    .A1(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .Y(_05095_),
    .A2(_04917_));
 sg13g2_inv_1 _22755_ (.Y(_05096_),
    .A(_05095_));
 sg13g2_nor3_1 _22756_ (.A(_09564_),
    .B(net747),
    .C(net668),
    .Y(_05097_));
 sg13g2_a21o_1 _22757_ (.A2(_05097_),
    .A1(_09132_),
    .B1(net410),
    .X(_05098_));
 sg13g2_a22oi_1 _22758_ (.Y(_05099_),
    .B1(_05098_),
    .B2(\cpu.gpio.r_enable_io[7] ),
    .A2(_05096_),
    .A1(_04844_));
 sg13g2_nand3_1 _22759_ (.B(_09139_),
    .C(_04888_),
    .A(_09138_),
    .Y(_05100_));
 sg13g2_and4_1 _22760_ (.A(_05086_),
    .B(_05091_),
    .C(_05099_),
    .D(_05100_),
    .X(_05101_));
 sg13g2_nor2b_1 _22761_ (.A(_00214_),
    .B_N(_04943_),
    .Y(_05102_));
 sg13g2_buf_1 _22762_ (.A(\cpu.spi.r_clk_count[2][7] ),
    .X(_05103_));
 sg13g2_and3_1 _22763_ (.X(_05104_),
    .A(net716),
    .B(net1069),
    .C(net648));
 sg13g2_buf_2 _22764_ (.A(_05104_),
    .X(_05105_));
 sg13g2_nand2_1 _22765_ (.Y(_05106_),
    .A(_11080_),
    .B(_04965_));
 sg13g2_buf_2 _22766_ (.A(_05106_),
    .X(_05107_));
 sg13g2_nor2_1 _22767_ (.A(_00150_),
    .B(_05107_),
    .Y(_05108_));
 sg13g2_a221oi_1 _22768_ (.B2(\cpu.spi.r_timeout[7] ),
    .C1(_05108_),
    .B1(_05105_),
    .A1(_05103_),
    .Y(_05109_),
    .A2(_04952_));
 sg13g2_o21ai_1 _22769_ (.B1(_05109_),
    .Y(_05110_),
    .A1(_00149_),
    .A2(_04949_));
 sg13g2_o21ai_1 _22770_ (.B1(_09170_),
    .Y(_05111_),
    .A1(_05102_),
    .A2(_05110_));
 sg13g2_o21ai_1 _22771_ (.B1(_05111_),
    .Y(_05112_),
    .A1(_05077_),
    .A2(_05101_));
 sg13g2_nor3_1 _22772_ (.A(net1067),
    .B(_05076_),
    .C(_05112_),
    .Y(_05113_));
 sg13g2_a21oi_2 _22773_ (.B1(_05113_),
    .Y(_05114_),
    .A2(_05063_),
    .A1(_09194_));
 sg13g2_nand2b_1 _22774_ (.Y(_05115_),
    .B(net994),
    .A_N(_05114_));
 sg13g2_inv_1 _22775_ (.Y(_05116_),
    .A(_05115_));
 sg13g2_buf_1 _22776_ (.A(_04978_),
    .X(_05117_));
 sg13g2_inv_1 _22777_ (.Y(_05118_),
    .A(_00094_));
 sg13g2_buf_1 _22778_ (.A(net638),
    .X(_05119_));
 sg13g2_a22oi_1 _22779_ (.Y(_05120_),
    .B1(_03028_),
    .B2(\cpu.dcache.r_data[2][26] ),
    .A2(_05119_),
    .A1(_05118_));
 sg13g2_a22oi_1 _22780_ (.Y(_05121_),
    .B1(net483),
    .B2(\cpu.dcache.r_data[1][26] ),
    .A2(net479),
    .A1(\cpu.dcache.r_data[6][26] ));
 sg13g2_a22oi_1 _22781_ (.Y(_05122_),
    .B1(net478),
    .B2(\cpu.dcache.r_data[7][26] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[5][26] ));
 sg13g2_a22oi_1 _22782_ (.Y(_05123_),
    .B1(net491),
    .B2(\cpu.dcache.r_data[4][26] ),
    .A2(_03032_),
    .A1(\cpu.dcache.r_data[3][26] ));
 sg13g2_nand4_1 _22783_ (.B(_05121_),
    .C(_05122_),
    .A(_05120_),
    .Y(_05124_),
    .D(_05123_));
 sg13g2_buf_1 _22784_ (.A(net514),
    .X(_05125_));
 sg13g2_a22oi_1 _22785_ (.Y(_05126_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][10] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][10] ));
 sg13g2_a22oi_1 _22786_ (.Y(_05127_),
    .B1(net483),
    .B2(\cpu.dcache.r_data[1][10] ),
    .A2(net480),
    .A1(\cpu.dcache.r_data[5][10] ));
 sg13g2_nor2b_1 _22787_ (.A(net569),
    .B_N(\cpu.dcache.r_data[4][10] ),
    .Y(_05128_));
 sg13g2_a21oi_1 _22788_ (.A1(net569),
    .A2(\cpu.dcache.r_data[6][10] ),
    .Y(_05129_),
    .B1(_05128_));
 sg13g2_nand3_1 _22789_ (.B(_09192_),
    .C(\cpu.dcache.r_data[7][10] ),
    .A(net716),
    .Y(_05130_));
 sg13g2_o21ai_1 _22790_ (.B1(_05130_),
    .Y(_05131_),
    .A1(_09176_),
    .A2(_05129_));
 sg13g2_nand2_1 _22791_ (.Y(_05132_),
    .A(net925),
    .B(_05131_));
 sg13g2_and4_1 _22792_ (.A(_09460_),
    .B(_05126_),
    .C(_05127_),
    .D(_05132_),
    .X(_05133_));
 sg13g2_a21oi_1 _22793_ (.A1(_00095_),
    .A2(net463),
    .Y(_05134_),
    .B1(_05133_));
 sg13g2_mux2_1 _22794_ (.A0(_05124_),
    .A1(_05134_),
    .S(net694),
    .X(_05135_));
 sg13g2_nor3_1 _22795_ (.A(net1067),
    .B(_04959_),
    .C(_04903_),
    .Y(_05136_));
 sg13g2_buf_2 _22796_ (.A(_05136_),
    .X(_05137_));
 sg13g2_buf_1 _22797_ (.A(_04847_),
    .X(_05138_));
 sg13g2_buf_1 _22798_ (.A(_04921_),
    .X(_05139_));
 sg13g2_a22oi_1 _22799_ (.Y(_05140_),
    .B1(net341),
    .B2(\cpu.intr.r_timer_reload[10] ),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_buf_1 _22800_ (.A(net376),
    .X(_05141_));
 sg13g2_buf_2 _22801_ (.A(\cpu.intr.r_clock_count[26] ),
    .X(_05142_));
 sg13g2_a22oi_1 _22802_ (.Y(_05143_),
    .B1(net340),
    .B2(_05142_),
    .A2(net667),
    .A1(_09905_));
 sg13g2_buf_1 _22803_ (.A(net412),
    .X(_05144_));
 sg13g2_nor2_1 _22804_ (.A(net796),
    .B(net924),
    .Y(_05145_));
 sg13g2_buf_1 _22805_ (.A(_05145_),
    .X(_05146_));
 sg13g2_a22oi_1 _22806_ (.Y(_05147_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[10] ),
    .A2(net374),
    .A1(_10088_));
 sg13g2_nand3_1 _22807_ (.B(_05143_),
    .C(_05147_),
    .A(_05140_),
    .Y(_05148_));
 sg13g2_a221oi_1 _22808_ (.B2(_05148_),
    .C1(net994),
    .B1(_05137_),
    .A1(net603),
    .Y(_05149_),
    .A2(_05135_));
 sg13g2_nor3_1 _22809_ (.A(net68),
    .B(_05116_),
    .C(_05149_),
    .Y(_05150_));
 sg13g2_a21oi_1 _22810_ (.A1(net1143),
    .A2(_05024_),
    .Y(_05151_),
    .B1(_05150_));
 sg13g2_buf_1 _22811_ (.A(_11622_),
    .X(_05152_));
 sg13g2_nor2_1 _22812_ (.A(_05152_),
    .B(_04752_),
    .Y(_05153_));
 sg13g2_a21o_1 _22813_ (.A2(_04749_),
    .A1(_05152_),
    .B1(_05153_),
    .X(_05154_));
 sg13g2_buf_1 _22814_ (.A(net347),
    .X(_05155_));
 sg13g2_nor2_1 _22815_ (.A(net291),
    .B(net164),
    .Y(_05156_));
 sg13g2_buf_1 _22816_ (.A(net247),
    .X(_05157_));
 sg13g2_nor3_1 _22817_ (.A(net984),
    .B(net211),
    .C(net164),
    .Y(_05158_));
 sg13g2_a221oi_1 _22818_ (.B2(_05156_),
    .C1(_05158_),
    .B1(_05154_),
    .A1(_05023_),
    .Y(_01020_),
    .A2(_05151_));
 sg13g2_a21oi_1 _22819_ (.A1(_11619_),
    .A2(_11620_),
    .Y(_05159_),
    .B1(_08375_));
 sg13g2_buf_1 _22820_ (.A(_05159_),
    .X(_05160_));
 sg13g2_buf_1 _22821_ (.A(net664),
    .X(_05161_));
 sg13g2_nand2_1 _22822_ (.Y(_05162_),
    .A(net599),
    .B(_04229_));
 sg13g2_o21ai_1 _22823_ (.B1(_05162_),
    .Y(_05163_),
    .A1(net599),
    .A2(_04221_));
 sg13g2_a22oi_1 _22824_ (.Y(_05164_),
    .B1(net374),
    .B2(_10093_),
    .A2(net341),
    .A1(\cpu.intr.r_timer_reload[11] ));
 sg13g2_buf_2 _22825_ (.A(\cpu.intr.r_clock_count[27] ),
    .X(_05165_));
 sg13g2_a22oi_1 _22826_ (.Y(_05166_),
    .B1(net340),
    .B2(_05165_),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_a22oi_1 _22827_ (.Y(_05167_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[11] ),
    .A2(net667),
    .A1(\cpu.intr.r_timer_count[11] ));
 sg13g2_nand3_1 _22828_ (.B(_05166_),
    .C(_05167_),
    .A(_05164_),
    .Y(_05168_));
 sg13g2_inv_1 _22829_ (.Y(_05169_),
    .A(_00106_));
 sg13g2_a22oi_1 _22830_ (.Y(_05170_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][11] ),
    .A2(net463),
    .A1(_05169_));
 sg13g2_a22oi_1 _22831_ (.Y(_05171_),
    .B1(net425),
    .B2(\cpu.dcache.r_data[1][11] ),
    .A2(_03043_),
    .A1(\cpu.dcache.r_data[6][11] ));
 sg13g2_a22oi_1 _22832_ (.Y(_05172_),
    .B1(_03048_),
    .B2(\cpu.dcache.r_data[7][11] ),
    .A2(net480),
    .A1(\cpu.dcache.r_data[5][11] ));
 sg13g2_a22oi_1 _22833_ (.Y(_05173_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][11] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][11] ));
 sg13g2_nand4_1 _22834_ (.B(_05171_),
    .C(_05172_),
    .A(_05170_),
    .Y(_05174_),
    .D(_05173_));
 sg13g2_a22oi_1 _22835_ (.Y(_05175_),
    .B1(net543),
    .B2(\cpu.dcache.r_data[7][27] ),
    .A2(_03032_),
    .A1(\cpu.dcache.r_data[3][27] ));
 sg13g2_a22oi_1 _22836_ (.Y(_05176_),
    .B1(net479),
    .B2(\cpu.dcache.r_data[6][27] ),
    .A2(_03036_),
    .A1(\cpu.dcache.r_data[5][27] ));
 sg13g2_a22oi_1 _22837_ (.Y(_05177_),
    .B1(_03028_),
    .B2(\cpu.dcache.r_data[2][27] ),
    .A2(net567),
    .A1(\cpu.dcache.r_data[4][27] ));
 sg13g2_nand3_1 _22838_ (.B(_05176_),
    .C(_05177_),
    .A(_05175_),
    .Y(_05178_));
 sg13g2_nand2_1 _22839_ (.Y(_05179_),
    .A(_00105_),
    .B(net669));
 sg13g2_o21ai_1 _22840_ (.B1(_05179_),
    .Y(_05180_),
    .A1(net669),
    .A2(_05178_));
 sg13g2_o21ai_1 _22841_ (.B1(net425),
    .Y(_05181_),
    .A1(\cpu.dcache.r_data[1][27] ),
    .A2(_05178_));
 sg13g2_o21ai_1 _22842_ (.B1(_05181_),
    .Y(_05182_),
    .A1(net425),
    .A2(_05180_));
 sg13g2_mux2_1 _22843_ (.A0(_05174_),
    .A1(_05182_),
    .S(net695),
    .X(_05183_));
 sg13g2_a22oi_1 _22844_ (.Y(_05184_),
    .B1(_05183_),
    .B2(_04978_),
    .A2(_05168_),
    .A1(_05137_));
 sg13g2_a21oi_2 _22845_ (.B1(net175),
    .Y(_05185_),
    .A2(_05114_),
    .A1(_03140_));
 sg13g2_o21ai_1 _22846_ (.B1(_05185_),
    .Y(_05186_),
    .A1(_03140_),
    .A2(_05184_));
 sg13g2_nor2b_1 _22847_ (.A(_04840_),
    .B_N(_05186_),
    .Y(_05187_));
 sg13g2_a21oi_1 _22848_ (.A1(net1135),
    .A2(net68),
    .Y(_05188_),
    .B1(_05187_));
 sg13g2_nand3_1 _22849_ (.B(net291),
    .C(net175),
    .A(_08837_),
    .Y(_05189_));
 sg13g2_o21ai_1 _22850_ (.B1(_05189_),
    .Y(_05190_),
    .A1(net132),
    .A2(_05188_));
 sg13g2_a21o_1 _22851_ (.A2(_05163_),
    .A1(_05156_),
    .B1(_05190_),
    .X(_01021_));
 sg13g2_inv_1 _22852_ (.Y(_05191_),
    .A(_00116_));
 sg13g2_a22oi_1 _22853_ (.Y(_05192_),
    .B1(_03027_),
    .B2(\cpu.dcache.r_data[2][28] ),
    .A2(net638),
    .A1(_05191_));
 sg13g2_a22oi_1 _22854_ (.Y(_05193_),
    .B1(net548),
    .B2(\cpu.dcache.r_data[1][28] ),
    .A2(_03040_),
    .A1(\cpu.dcache.r_data[6][28] ));
 sg13g2_a22oi_1 _22855_ (.Y(_05194_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][28] ),
    .A2(_09414_),
    .A1(\cpu.dcache.r_data[5][28] ));
 sg13g2_a22oi_1 _22856_ (.Y(_05195_),
    .B1(net640),
    .B2(\cpu.dcache.r_data[4][28] ),
    .A2(_03031_),
    .A1(\cpu.dcache.r_data[3][28] ));
 sg13g2_and4_1 _22857_ (.A(_05192_),
    .B(_05193_),
    .C(_05194_),
    .D(_05195_),
    .X(_05196_));
 sg13g2_buf_1 _22858_ (.A(_05196_),
    .X(_05197_));
 sg13g2_nor2_1 _22859_ (.A(net694),
    .B(_05197_),
    .Y(_05198_));
 sg13g2_inv_1 _22860_ (.Y(_05199_),
    .A(_00117_));
 sg13g2_a22oi_1 _22861_ (.Y(_05200_),
    .B1(net482),
    .B2(\cpu.dcache.r_data[2][12] ),
    .A2(net514),
    .A1(_05199_));
 sg13g2_a22oi_1 _22862_ (.Y(_05201_),
    .B1(_03023_),
    .B2(\cpu.dcache.r_data[1][12] ),
    .A2(_03041_),
    .A1(\cpu.dcache.r_data[6][12] ));
 sg13g2_a22oi_1 _22863_ (.Y(_05202_),
    .B1(_03046_),
    .B2(\cpu.dcache.r_data[7][12] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[5][12] ));
 sg13g2_a22oi_1 _22864_ (.Y(_05203_),
    .B1(net567),
    .B2(\cpu.dcache.r_data[4][12] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[3][12] ));
 sg13g2_nand4_1 _22865_ (.B(_05201_),
    .C(_05202_),
    .A(_05200_),
    .Y(_05204_),
    .D(_05203_));
 sg13g2_and2_1 _22866_ (.A(_09889_),
    .B(_05204_),
    .X(_05205_));
 sg13g2_or2_1 _22867_ (.X(_05206_),
    .B(_05205_),
    .A(_05198_));
 sg13g2_a22oi_1 _22868_ (.Y(_05207_),
    .B1(net374),
    .B2(_10100_),
    .A2(net341),
    .A1(\cpu.intr.r_timer_reload[12] ));
 sg13g2_buf_1 _22869_ (.A(\cpu.intr.r_clock_count[28] ),
    .X(_05208_));
 sg13g2_a22oi_1 _22870_ (.Y(_05209_),
    .B1(net340),
    .B2(_05208_),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_a22oi_1 _22871_ (.Y(_05210_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[12] ),
    .A2(net667),
    .A1(\cpu.intr.r_timer_count[12] ));
 sg13g2_nand3_1 _22872_ (.B(_05209_),
    .C(_05210_),
    .A(_05207_),
    .Y(_05211_));
 sg13g2_a221oi_1 _22873_ (.B2(_05137_),
    .C1(net877),
    .B1(_05211_),
    .A1(net603),
    .Y(_05212_),
    .A2(_05206_));
 sg13g2_nor3_1 _22874_ (.A(net68),
    .B(_05116_),
    .C(_05212_),
    .Y(_05213_));
 sg13g2_a21oi_1 _22875_ (.A1(net627),
    .A2(net69),
    .Y(_05214_),
    .B1(_05213_));
 sg13g2_nor4_1 _22876_ (.A(net347),
    .B(net600),
    .C(net164),
    .D(_04282_),
    .Y(_05215_));
 sg13g2_nor3_1 _22877_ (.A(_08494_),
    .B(_03972_),
    .C(net164),
    .Y(_05216_));
 sg13g2_or2_1 _22878_ (.X(_05217_),
    .B(_05216_),
    .A(_05215_));
 sg13g2_a221oi_1 _22879_ (.B2(net131),
    .C1(_05217_),
    .B1(_05214_),
    .A1(_04279_),
    .Y(_01022_),
    .A2(_04836_));
 sg13g2_nand3_1 _22880_ (.B(_05155_),
    .C(_04838_),
    .A(_08423_),
    .Y(_05218_));
 sg13g2_buf_1 _22881_ (.A(net164),
    .X(_05219_));
 sg13g2_a22oi_1 _22882_ (.Y(_05220_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[13] ),
    .A2(net341),
    .A1(\cpu.intr.r_timer_reload[13] ));
 sg13g2_a22oi_1 _22883_ (.Y(_05221_),
    .B1(net412),
    .B2(_10105_),
    .A2(_05138_),
    .A1(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_buf_1 _22884_ (.A(\cpu.intr.r_clock_count[29] ),
    .X(_05222_));
 sg13g2_a22oi_1 _22885_ (.Y(_05223_),
    .B1(_04918_),
    .B2(_05222_),
    .A2(net667),
    .A1(\cpu.intr.r_timer_count[13] ));
 sg13g2_nand3_1 _22886_ (.B(_05221_),
    .C(_05223_),
    .A(_05220_),
    .Y(_05224_));
 sg13g2_inv_1 _22887_ (.Y(_05225_),
    .A(_00123_));
 sg13g2_a22oi_1 _22888_ (.Y(_05226_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][29] ),
    .A2(net514),
    .A1(_05225_));
 sg13g2_a22oi_1 _22889_ (.Y(_05227_),
    .B1(net483),
    .B2(\cpu.dcache.r_data[1][29] ),
    .A2(_03042_),
    .A1(\cpu.dcache.r_data[6][29] ));
 sg13g2_a22oi_1 _22890_ (.Y(_05228_),
    .B1(net478),
    .B2(\cpu.dcache.r_data[7][29] ),
    .A2(net480),
    .A1(\cpu.dcache.r_data[5][29] ));
 sg13g2_a22oi_1 _22891_ (.Y(_05229_),
    .B1(_10018_),
    .B2(\cpu.dcache.r_data[4][29] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][29] ));
 sg13g2_nand4_1 _22892_ (.B(_05227_),
    .C(_05228_),
    .A(_05226_),
    .Y(_05230_),
    .D(_05229_));
 sg13g2_mux2_1 _22893_ (.A0(\cpu.dcache.r_data[1][13] ),
    .A1(\cpu.dcache.r_data[3][13] ),
    .S(net493),
    .X(_05231_));
 sg13g2_a22oi_1 _22894_ (.Y(_05232_),
    .B1(_05231_),
    .B2(_12563_),
    .A2(net666),
    .A1(\cpu.dcache.r_data[2][13] ));
 sg13g2_inv_1 _22895_ (.Y(_05233_),
    .A(_00124_));
 sg13g2_mux2_1 _22896_ (.A0(\cpu.dcache.r_data[4][13] ),
    .A1(\cpu.dcache.r_data[6][13] ),
    .S(net569),
    .X(_05234_));
 sg13g2_a22oi_1 _22897_ (.Y(_05235_),
    .B1(_05234_),
    .B2(net767),
    .A2(_09517_),
    .A1(\cpu.dcache.r_data[5][13] ));
 sg13g2_nor2_1 _22898_ (.A(_12075_),
    .B(_05235_),
    .Y(_05236_));
 sg13g2_a221oi_1 _22899_ (.B2(\cpu.dcache.r_data[7][13] ),
    .C1(_05236_),
    .B1(net478),
    .A1(_05233_),
    .Y(_05237_),
    .A2(_05119_));
 sg13g2_o21ai_1 _22900_ (.B1(_05237_),
    .Y(_05238_),
    .A1(_09511_),
    .A2(_05232_));
 sg13g2_mux2_1 _22901_ (.A0(_05230_),
    .A1(_05238_),
    .S(net798),
    .X(_05239_));
 sg13g2_a22oi_1 _22902_ (.Y(_05240_),
    .B1(_05239_),
    .B2(_04978_),
    .A2(_05224_),
    .A1(_05137_));
 sg13g2_nor2_1 _22903_ (.A(net994),
    .B(_05240_),
    .Y(_05241_));
 sg13g2_nor2b_1 _22904_ (.A(_05241_),
    .B_N(_05185_),
    .Y(_05242_));
 sg13g2_nand2_1 _22905_ (.Y(_05243_),
    .A(net628),
    .B(_04840_));
 sg13g2_o21ai_1 _22906_ (.B1(_05243_),
    .Y(_05244_),
    .A1(net68),
    .A2(_05242_));
 sg13g2_nand2_1 _22907_ (.Y(_05245_),
    .A(net130),
    .B(_05244_));
 sg13g2_a21oi_2 _22908_ (.B1(_11632_),
    .Y(_05246_),
    .A2(_11636_),
    .A1(net1081));
 sg13g2_nor3_1 _22909_ (.A(net347),
    .B(_05242_),
    .C(_05246_),
    .Y(_05247_));
 sg13g2_nand4_1 _22910_ (.B(_04344_),
    .C(_04345_),
    .A(net600),
    .Y(_05248_),
    .D(_05247_));
 sg13g2_nand3_1 _22911_ (.B(_04348_),
    .C(_05247_),
    .A(net599),
    .Y(_05249_));
 sg13g2_nand4_1 _22912_ (.B(_05245_),
    .C(_05248_),
    .A(_05218_),
    .Y(_01023_),
    .D(_05249_));
 sg13g2_nor4_1 _22913_ (.A(net246),
    .B(net664),
    .C(_11976_),
    .D(_11978_),
    .Y(_05250_));
 sg13g2_o21ai_1 _22914_ (.B1(_03972_),
    .Y(_05251_),
    .A1(_11622_),
    .A2(_04391_));
 sg13g2_nand2_1 _22915_ (.Y(_05252_),
    .A(_08636_),
    .B(net347));
 sg13g2_o21ai_1 _22916_ (.B1(_05252_),
    .Y(_05253_),
    .A1(_05250_),
    .A2(_05251_));
 sg13g2_nand2_1 _22917_ (.Y(_05254_),
    .A(net132),
    .B(_05253_));
 sg13g2_nor3_1 _22918_ (.A(_04357_),
    .B(_04387_),
    .C(_04835_),
    .Y(_05255_));
 sg13g2_inv_1 _22919_ (.Y(_05256_),
    .A(_00135_));
 sg13g2_a22oi_1 _22920_ (.Y(_05257_),
    .B1(_03036_),
    .B2(\cpu.dcache.r_data[5][30] ),
    .A2(net514),
    .A1(_05256_));
 sg13g2_a22oi_1 _22921_ (.Y(_05258_),
    .B1(net567),
    .B2(\cpu.dcache.r_data[4][30] ),
    .A2(_03023_),
    .A1(\cpu.dcache.r_data[1][30] ));
 sg13g2_a22oi_1 _22922_ (.Y(_05259_),
    .B1(net481),
    .B2(\cpu.dcache.r_data[3][30] ),
    .A2(_03041_),
    .A1(\cpu.dcache.r_data[6][30] ));
 sg13g2_a22oi_1 _22923_ (.Y(_05260_),
    .B1(net482),
    .B2(\cpu.dcache.r_data[2][30] ),
    .A2(_03046_),
    .A1(\cpu.dcache.r_data[7][30] ));
 sg13g2_nand4_1 _22924_ (.B(_05258_),
    .C(_05259_),
    .A(_05257_),
    .Y(_05261_),
    .D(_05260_));
 sg13g2_a22oi_1 _22925_ (.Y(_05262_),
    .B1(net547),
    .B2(\cpu.dcache.r_data[2][14] ),
    .A2(net544),
    .A1(\cpu.dcache.r_data[6][14] ));
 sg13g2_a22oi_1 _22926_ (.Y(_05263_),
    .B1(_10017_),
    .B2(\cpu.dcache.r_data[4][14] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][14] ));
 sg13g2_a22oi_1 _22927_ (.Y(_05264_),
    .B1(net621),
    .B2(\cpu.dcache.r_data[7][14] ),
    .A2(net639),
    .A1(\cpu.dcache.r_data[5][14] ));
 sg13g2_nand3_1 _22928_ (.B(_05263_),
    .C(_05264_),
    .A(_05262_),
    .Y(_05265_));
 sg13g2_nand2_1 _22929_ (.Y(_05266_),
    .A(_00136_),
    .B(net669));
 sg13g2_o21ai_1 _22930_ (.B1(_05266_),
    .Y(_05267_),
    .A1(net669),
    .A2(_05265_));
 sg13g2_o21ai_1 _22931_ (.B1(_03024_),
    .Y(_05268_),
    .A1(\cpu.dcache.r_data[1][14] ),
    .A2(_05265_));
 sg13g2_o21ai_1 _22932_ (.B1(_05268_),
    .Y(_05269_),
    .A1(_03025_),
    .A2(_05267_));
 sg13g2_mux2_1 _22933_ (.A0(_05261_),
    .A1(_05269_),
    .S(net798),
    .X(_05270_));
 sg13g2_a22oi_1 _22934_ (.Y(_05271_),
    .B1(net380),
    .B2(\cpu.intr.r_timer_count[14] ),
    .A2(_03038_),
    .A1(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_buf_1 _22935_ (.A(\cpu.intr.r_clock_count[30] ),
    .X(_05272_));
 sg13g2_a22oi_1 _22936_ (.Y(_05273_),
    .B1(net374),
    .B2(_10110_),
    .A2(net340),
    .A1(_05272_));
 sg13g2_a22oi_1 _22937_ (.Y(_05274_),
    .B1(net341),
    .B2(\cpu.intr.r_timer_reload[14] ),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_and2_1 _22938_ (.A(_05273_),
    .B(_05274_),
    .X(_05275_));
 sg13g2_o21ai_1 _22939_ (.B1(_05275_),
    .Y(_05276_),
    .A1(net636),
    .A2(_05271_));
 sg13g2_a221oi_1 _22940_ (.B2(_05137_),
    .C1(net994),
    .B1(_05276_),
    .A1(net603),
    .Y(_05277_),
    .A2(_05270_));
 sg13g2_nor3_1 _22941_ (.A(_04840_),
    .B(_05116_),
    .C(_05277_),
    .Y(_05278_));
 sg13g2_a21oi_1 _22942_ (.A1(net698),
    .A2(net68),
    .Y(_05279_),
    .B1(_05278_));
 sg13g2_or2_1 _22943_ (.X(_05280_),
    .B(_05279_),
    .A(net132));
 sg13g2_o21ai_1 _22944_ (.B1(_05280_),
    .Y(_01024_),
    .A1(_05254_),
    .A2(_05255_));
 sg13g2_a22oi_1 _22945_ (.Y(_05281_),
    .B1(net374),
    .B2(_10116_),
    .A2(net341),
    .A1(\cpu.intr.r_timer_reload[15] ));
 sg13g2_buf_1 _22946_ (.A(\cpu.intr.r_clock_count[31] ),
    .X(_05282_));
 sg13g2_a22oi_1 _22947_ (.Y(_05283_),
    .B1(net340),
    .B2(_05282_),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_a22oi_1 _22948_ (.Y(_05284_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[15] ),
    .A2(net667),
    .A1(\cpu.intr.r_timer_count[15] ));
 sg13g2_nand3_1 _22949_ (.B(_05283_),
    .C(_05284_),
    .A(_05281_),
    .Y(_05285_));
 sg13g2_mux2_1 _22950_ (.A0(_05051_),
    .A1(_05057_),
    .S(net636),
    .X(_05286_));
 sg13g2_a22oi_1 _22951_ (.Y(_05287_),
    .B1(_05286_),
    .B2(net603),
    .A2(_05285_),
    .A1(_05137_));
 sg13g2_o21ai_1 _22952_ (.B1(_05185_),
    .Y(_05288_),
    .A1(net877),
    .A2(_05287_));
 sg13g2_mux2_1 _22953_ (.A0(_05288_),
    .A1(net687),
    .S(_05025_),
    .X(_05289_));
 sg13g2_nor2_1 _22954_ (.A(_08637_),
    .B(net247),
    .Y(_05290_));
 sg13g2_nor3_1 _22955_ (.A(net347),
    .B(net600),
    .C(_04439_),
    .Y(_05291_));
 sg13g2_nor3_1 _22956_ (.A(net164),
    .B(_05290_),
    .C(_05291_),
    .Y(_05292_));
 sg13g2_a21oi_1 _22957_ (.A1(net130),
    .A2(_05289_),
    .Y(_05293_),
    .B1(_05292_));
 sg13g2_a21oi_1 _22958_ (.A1(_04437_),
    .A2(_04836_),
    .Y(_01025_),
    .B1(_05293_));
 sg13g2_nand2_1 _22959_ (.Y(_05294_),
    .A(_10563_),
    .B(net664));
 sg13g2_o21ai_1 _22960_ (.B1(_05294_),
    .Y(_05295_),
    .A1(net664),
    .A2(_04078_));
 sg13g2_nor2_1 _22961_ (.A(net934),
    .B(_05157_),
    .Y(_05296_));
 sg13g2_a21oi_1 _22962_ (.A1(net211),
    .A2(_05295_),
    .Y(_05297_),
    .B1(_05296_));
 sg13g2_mux2_1 _22963_ (.A0(\cpu.dcache.r_data[1][1] ),
    .A1(\cpu.dcache.r_data[3][1] ),
    .S(net493),
    .X(_05298_));
 sg13g2_a22oi_1 _22964_ (.Y(_05299_),
    .B1(_05298_),
    .B2(net622),
    .A2(_04962_),
    .A1(\cpu.dcache.r_data[2][1] ));
 sg13g2_mux2_1 _22965_ (.A0(\cpu.dcache.r_data[5][1] ),
    .A1(\cpu.dcache.r_data[7][1] ),
    .S(net569),
    .X(_05300_));
 sg13g2_a22oi_1 _22966_ (.Y(_05301_),
    .B1(_05300_),
    .B2(net716),
    .A2(net666),
    .A1(\cpu.dcache.r_data[6][1] ));
 sg13g2_nor2_1 _22967_ (.A(net771),
    .B(_05301_),
    .Y(_05302_));
 sg13g2_a221oi_1 _22968_ (.B2(\cpu.dcache.r_data[4][1] ),
    .C1(_05302_),
    .B1(net491),
    .A1(\cpu.dcache.r_data[0][1] ),
    .Y(_05303_),
    .A2(net463));
 sg13g2_o21ai_1 _22969_ (.B1(_05303_),
    .Y(_05304_),
    .A1(_09511_),
    .A2(_05299_));
 sg13g2_inv_1 _22970_ (.Y(_05305_),
    .A(_00296_));
 sg13g2_a22oi_1 _22971_ (.Y(_05306_),
    .B1(net480),
    .B2(\cpu.dcache.r_data[5][17] ),
    .A2(net514),
    .A1(_05305_));
 sg13g2_a22oi_1 _22972_ (.Y(_05307_),
    .B1(net491),
    .B2(\cpu.dcache.r_data[4][17] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[1][17] ));
 sg13g2_a22oi_1 _22973_ (.Y(_05308_),
    .B1(net423),
    .B2(\cpu.dcache.r_data[3][17] ),
    .A2(net421),
    .A1(\cpu.dcache.r_data[6][17] ));
 sg13g2_a22oi_1 _22974_ (.Y(_05309_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][17] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[7][17] ));
 sg13g2_and4_1 _22975_ (.A(_05306_),
    .B(_05307_),
    .C(_05308_),
    .D(_05309_),
    .X(_05310_));
 sg13g2_nand2_1 _22976_ (.Y(_05311_),
    .A(net636),
    .B(_05310_));
 sg13g2_o21ai_1 _22977_ (.B1(_05311_),
    .Y(_05312_),
    .A1(net566),
    .A2(_05304_));
 sg13g2_buf_1 _22978_ (.A(net665),
    .X(_05313_));
 sg13g2_inv_1 _22979_ (.Y(_05314_),
    .A(_05310_));
 sg13g2_a22oi_1 _22980_ (.Y(_05315_),
    .B1(_05314_),
    .B2(_05042_),
    .A2(_05304_),
    .A1(net1030));
 sg13g2_inv_1 _22981_ (.Y(_05316_),
    .A(_00298_));
 sg13g2_a22oi_1 _22982_ (.Y(_05317_),
    .B1(_03037_),
    .B2(\cpu.dcache.r_data[5][9] ),
    .A2(_05125_),
    .A1(_05316_));
 sg13g2_a22oi_1 _22983_ (.Y(_05318_),
    .B1(_03024_),
    .B2(\cpu.dcache.r_data[1][9] ),
    .A2(net421),
    .A1(\cpu.dcache.r_data[6][9] ));
 sg13g2_a22oi_1 _22984_ (.Y(_05319_),
    .B1(_10018_),
    .B2(\cpu.dcache.r_data[4][9] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][9] ));
 sg13g2_a22oi_1 _22985_ (.Y(_05320_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][9] ),
    .A2(_03047_),
    .A1(\cpu.dcache.r_data[7][9] ));
 sg13g2_nand4_1 _22986_ (.B(_05318_),
    .C(_05319_),
    .A(_05317_),
    .Y(_05321_),
    .D(_05320_));
 sg13g2_inv_1 _22987_ (.Y(_05322_),
    .A(_00297_));
 sg13g2_a22oi_1 _22988_ (.Y(_05323_),
    .B1(_03037_),
    .B2(\cpu.dcache.r_data[5][25] ),
    .A2(_05125_),
    .A1(_05322_));
 sg13g2_a22oi_1 _22989_ (.Y(_05324_),
    .B1(net491),
    .B2(\cpu.dcache.r_data[4][25] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[1][25] ));
 sg13g2_a22oi_1 _22990_ (.Y(_05325_),
    .B1(_03033_),
    .B2(\cpu.dcache.r_data[3][25] ),
    .A2(_03042_),
    .A1(\cpu.dcache.r_data[6][25] ));
 sg13g2_a22oi_1 _22991_ (.Y(_05326_),
    .B1(_03029_),
    .B2(\cpu.dcache.r_data[2][25] ),
    .A2(_03047_),
    .A1(\cpu.dcache.r_data[7][25] ));
 sg13g2_nand4_1 _22992_ (.B(_05324_),
    .C(_05325_),
    .A(_05323_),
    .Y(_05327_),
    .D(_05326_));
 sg13g2_a221oi_1 _22993_ (.B2(net898),
    .C1(_05313_),
    .B1(_05327_),
    .A1(net798),
    .Y(_05328_),
    .A2(_05321_));
 sg13g2_a21oi_1 _22994_ (.A1(_05313_),
    .A2(_05315_),
    .Y(_05329_),
    .B1(_05328_));
 sg13g2_nor2_1 _22995_ (.A(_04978_),
    .B(_05329_),
    .Y(_05330_));
 sg13g2_a21oi_1 _22996_ (.A1(net603),
    .A2(_05312_),
    .Y(_05331_),
    .B1(_05330_));
 sg13g2_nor2_1 _22997_ (.A(net1001),
    .B(_05331_),
    .Y(_05332_));
 sg13g2_nor2b_1 _22998_ (.A(_00304_),
    .B_N(net670),
    .Y(_05333_));
 sg13g2_buf_1 _22999_ (.A(_04913_),
    .X(_05334_));
 sg13g2_a22oi_1 _23000_ (.Y(_05335_),
    .B1(net411),
    .B2(_09125_),
    .A2(_05334_),
    .A1(_09126_));
 sg13g2_or2_1 _23001_ (.X(_05336_),
    .B(_04848_),
    .A(_00305_));
 sg13g2_o21ai_1 _23002_ (.B1(_05336_),
    .Y(_05337_),
    .A1(net769),
    .A2(_05335_));
 sg13g2_nand2b_1 _23003_ (.Y(_05338_),
    .B(_04863_),
    .A_N(_00303_));
 sg13g2_o21ai_1 _23004_ (.B1(_05338_),
    .Y(_05339_),
    .A1(_00301_),
    .A2(_05080_));
 sg13g2_nand2_2 _23005_ (.Y(_05340_),
    .A(net1061),
    .B(_04968_));
 sg13g2_buf_2 _23006_ (.A(\cpu.gpio.r_src_io[4][1] ),
    .X(_05341_));
 sg13g2_nand2_1 _23007_ (.Y(_05342_),
    .A(_05341_),
    .B(net413));
 sg13g2_o21ai_1 _23008_ (.B1(_05342_),
    .Y(_05343_),
    .A1(_00302_),
    .A2(_05340_));
 sg13g2_nor4_1 _23009_ (.A(_05333_),
    .B(_05337_),
    .C(_05339_),
    .D(_05343_),
    .Y(_05344_));
 sg13g2_nand3_1 _23010_ (.B(_09126_),
    .C(_04888_),
    .A(_09125_),
    .Y(_05345_));
 sg13g2_a21oi_1 _23011_ (.A1(_05344_),
    .A2(_05345_),
    .Y(_05346_),
    .B1(_05077_));
 sg13g2_nand3_1 _23012_ (.B(\cpu.intr.r_clock_cmp[1] ),
    .C(_04914_),
    .A(net798),
    .Y(_05347_));
 sg13g2_o21ai_1 _23013_ (.B1(_12076_),
    .Y(_05348_),
    .A1(\cpu.intr.r_enable[1] ),
    .A2(net695));
 sg13g2_a21oi_1 _23014_ (.A1(_05347_),
    .A2(_05348_),
    .Y(_05349_),
    .B1(net767));
 sg13g2_a221oi_1 _23015_ (.B2(\cpu.intr.r_clock ),
    .C1(_05349_),
    .B1(net517),
    .A1(_09907_),
    .Y(_05350_),
    .A2(net667));
 sg13g2_nand3_1 _23016_ (.B(\cpu.intr.r_clock_cmp[17] ),
    .C(_04914_),
    .A(net622),
    .Y(_05351_));
 sg13g2_nand2_1 _23017_ (.Y(_05352_),
    .A(_09903_),
    .B(net666));
 sg13g2_nand2_1 _23018_ (.Y(_05353_),
    .A(_05351_),
    .B(_05352_));
 sg13g2_and2_1 _23019_ (.A(net796),
    .B(\cpu.intr.r_timer_reload[17] ),
    .X(_05354_));
 sg13g2_a21oi_1 _23020_ (.A1(net923),
    .A2(\cpu.intr.r_timer_reload[1] ),
    .Y(_05355_),
    .B1(_05354_));
 sg13g2_o21ai_1 _23021_ (.B1(_12077_),
    .Y(_05356_),
    .A1(net767),
    .A2(_05355_));
 sg13g2_nor2b_1 _23022_ (.A(net493),
    .B_N(_10037_),
    .Y(_05357_));
 sg13g2_nor3_1 _23023_ (.A(net695),
    .B(net771),
    .C(_05357_),
    .Y(_05358_));
 sg13g2_buf_1 _23024_ (.A(\cpu.intr.r_clock_count[17] ),
    .X(_05359_));
 sg13g2_a21oi_1 _23025_ (.A1(_05359_),
    .A2(_04914_),
    .Y(_05360_),
    .B1(net798));
 sg13g2_nor3_1 _23026_ (.A(net533),
    .B(_05358_),
    .C(_05360_),
    .Y(_05361_));
 sg13g2_a221oi_1 _23027_ (.B2(net418),
    .C1(_05361_),
    .B1(_05356_),
    .A1(net636),
    .Y(_05362_),
    .A2(_05353_));
 sg13g2_a221oi_1 _23028_ (.B2(_05362_),
    .C1(_04959_),
    .B1(_05350_),
    .A1(_09111_),
    .Y(_05363_),
    .A2(_04903_));
 sg13g2_a22oi_1 _23029_ (.Y(_05364_),
    .B1(net515),
    .B2(\cpu.uart.r_r_invert ),
    .A2(net409),
    .A1(\cpu.uart.r_div_value[9] ));
 sg13g2_a22oi_1 _23030_ (.Y(_05365_),
    .B1(net375),
    .B2(\cpu.uart.r_div_value[1] ),
    .A2(net408),
    .A1(_09115_));
 sg13g2_nand2_1 _23031_ (.Y(_05366_),
    .A(_05364_),
    .B(_05365_));
 sg13g2_a21oi_1 _23032_ (.A1(\cpu.uart.r_in[1] ),
    .A2(_04964_),
    .Y(_05367_),
    .B1(_05366_));
 sg13g2_o21ai_1 _23033_ (.B1(net1001),
    .Y(_05368_),
    .A1(_04961_),
    .A2(_05367_));
 sg13g2_nand2_1 _23034_ (.Y(_05369_),
    .A(net1000),
    .B(_09168_));
 sg13g2_buf_1 _23035_ (.A(\cpu.spi.r_clk_count[2][1] ),
    .X(_05370_));
 sg13g2_mux2_1 _23036_ (.A0(_12066_),
    .A1(_12067_),
    .S(net1061),
    .X(_05371_));
 sg13g2_a22oi_1 _23037_ (.Y(_05372_),
    .B1(_05371_),
    .B2(net411),
    .A2(_05105_),
    .A1(\cpu.spi.r_timeout[1] ));
 sg13g2_o21ai_1 _23038_ (.B1(_05372_),
    .Y(_05373_),
    .A1(_00300_),
    .A2(_05107_));
 sg13g2_a21oi_1 _23039_ (.A1(_05370_),
    .A2(_04952_),
    .Y(_05374_),
    .B1(_05373_));
 sg13g2_nor2_1 _23040_ (.A(_00299_),
    .B(_04949_),
    .Y(_05375_));
 sg13g2_a21oi_1 _23041_ (.A1(_12071_),
    .A2(net670),
    .Y(_05376_),
    .B1(_05375_));
 sg13g2_nand2_1 _23042_ (.Y(_05377_),
    .A(_05374_),
    .B(_05376_));
 sg13g2_a21oi_1 _23043_ (.A1(_09216_),
    .A2(_04943_),
    .Y(_05378_),
    .B1(_05377_));
 sg13g2_nor2_1 _23044_ (.A(_05369_),
    .B(_05378_),
    .Y(_05379_));
 sg13g2_nor4_1 _23045_ (.A(_05346_),
    .B(_05363_),
    .C(_05368_),
    .D(_05379_),
    .Y(_05380_));
 sg13g2_nor3_1 _23046_ (.A(net68),
    .B(_05332_),
    .C(_05380_),
    .Y(_05381_));
 sg13g2_a21oi_1 _23047_ (.A1(net1081),
    .A2(_11636_),
    .Y(_05382_),
    .B1(net635));
 sg13g2_o21ai_1 _23048_ (.B1(net130),
    .Y(_05383_),
    .A1(_05381_),
    .A2(_05382_));
 sg13g2_o21ai_1 _23049_ (.B1(_05383_),
    .Y(_01026_),
    .A1(net131),
    .A2(_05297_));
 sg13g2_mux2_1 _23050_ (.A0(\cpu.dcache.r_data[1][2] ),
    .A1(\cpu.dcache.r_data[3][2] ),
    .S(net493),
    .X(_05384_));
 sg13g2_a22oi_1 _23051_ (.Y(_05385_),
    .B1(_05384_),
    .B2(net622),
    .A2(net666),
    .A1(\cpu.dcache.r_data[2][2] ));
 sg13g2_inv_1 _23052_ (.Y(_05386_),
    .A(_05385_));
 sg13g2_mux2_1 _23053_ (.A0(\cpu.dcache.r_data[5][2] ),
    .A1(\cpu.dcache.r_data[7][2] ),
    .S(_09193_),
    .X(_05387_));
 sg13g2_a22oi_1 _23054_ (.Y(_05388_),
    .B1(_05387_),
    .B2(net622),
    .A2(net666),
    .A1(\cpu.dcache.r_data[6][2] ));
 sg13g2_a22oi_1 _23055_ (.Y(_05389_),
    .B1(net491),
    .B2(\cpu.dcache.r_data[4][2] ),
    .A2(net514),
    .A1(\cpu.dcache.r_data[0][2] ));
 sg13g2_o21ai_1 _23056_ (.B1(_05389_),
    .Y(_05390_),
    .A1(net771),
    .A2(_05388_));
 sg13g2_a21oi_1 _23057_ (.A1(net1065),
    .A2(_05386_),
    .Y(_05391_),
    .B1(_05390_));
 sg13g2_nand2_1 _23058_ (.Y(_05392_),
    .A(\cpu.dcache.r_data[2][18] ),
    .B(net482));
 sg13g2_a22oi_1 _23059_ (.Y(_05393_),
    .B1(net491),
    .B2(\cpu.dcache.r_data[4][18] ),
    .A2(net483),
    .A1(\cpu.dcache.r_data[1][18] ));
 sg13g2_a22oi_1 _23060_ (.Y(_05394_),
    .B1(net543),
    .B2(\cpu.dcache.r_data[7][18] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[5][18] ));
 sg13g2_a22oi_1 _23061_ (.Y(_05395_),
    .B1(net481),
    .B2(\cpu.dcache.r_data[3][18] ),
    .A2(net479),
    .A1(\cpu.dcache.r_data[6][18] ));
 sg13g2_nand4_1 _23062_ (.B(_05393_),
    .C(_05394_),
    .A(_05392_),
    .Y(_05396_),
    .D(_05395_));
 sg13g2_nor2_1 _23063_ (.A(net463),
    .B(_05396_),
    .Y(_05397_));
 sg13g2_a21oi_1 _23064_ (.A1(_00093_),
    .A2(net463),
    .Y(_05398_),
    .B1(_05397_));
 sg13g2_nand2_1 _23065_ (.Y(_05399_),
    .A(net695),
    .B(_05398_));
 sg13g2_mux2_1 _23066_ (.A0(_05391_),
    .A1(_05399_),
    .S(net898),
    .X(_05400_));
 sg13g2_a221oi_1 _23067_ (.B2(net694),
    .C1(net598),
    .B1(_05134_),
    .A1(net898),
    .Y(_05401_),
    .A2(_05124_));
 sg13g2_a21oi_1 _23068_ (.A1(net598),
    .A2(_05400_),
    .Y(_05402_),
    .B1(_05401_));
 sg13g2_o21ai_1 _23069_ (.B1(_05399_),
    .Y(_05403_),
    .A1(net566),
    .A2(_05391_));
 sg13g2_mux2_1 _23070_ (.A0(_05402_),
    .A1(_05403_),
    .S(net603),
    .X(_05404_));
 sg13g2_a22oi_1 _23071_ (.Y(_05405_),
    .B1(net420),
    .B2(\cpu.intr.r_timer_reload[18] ),
    .A2(net380),
    .A1(_09902_));
 sg13g2_a221oi_1 _23072_ (.B2(\cpu.intr.r_timer_reload[2] ),
    .C1(net636),
    .B1(net420),
    .A1(\cpu.intr.r_clock_cmp[2] ),
    .Y(_05406_),
    .A2(net422));
 sg13g2_a21oi_1 _23073_ (.A1(net636),
    .A2(_05405_),
    .Y(_05407_),
    .B1(_05406_));
 sg13g2_buf_1 _23074_ (.A(\cpu.intr.r_clock_count[18] ),
    .X(_05408_));
 sg13g2_a22oi_1 _23075_ (.Y(_05409_),
    .B1(net517),
    .B2(_09112_),
    .A2(net340),
    .A1(_05408_));
 sg13g2_nand2_1 _23076_ (.Y(_05410_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(net602));
 sg13g2_a22oi_1 _23077_ (.Y(_05411_),
    .B1(net374),
    .B2(_10045_),
    .A2(net667),
    .A1(\cpu.intr.r_timer_count[2] ));
 sg13g2_nand3_1 _23078_ (.B(_05410_),
    .C(_05411_),
    .A(_05409_),
    .Y(_05412_));
 sg13g2_a21oi_1 _23079_ (.A1(_09112_),
    .A2(_04903_),
    .Y(_05413_),
    .B1(net408));
 sg13g2_nor2b_1 _23080_ (.A(_05413_),
    .B_N(\cpu.intr.r_enable[2] ),
    .Y(_05414_));
 sg13g2_nor3_1 _23081_ (.A(_05407_),
    .B(_05412_),
    .C(_05414_),
    .Y(_05415_));
 sg13g2_nor2_1 _23082_ (.A(_00099_),
    .B(_05088_),
    .Y(_05416_));
 sg13g2_nor2b_1 _23083_ (.A(net769),
    .B_N(_09137_),
    .Y(_05417_));
 sg13g2_nand2b_1 _23084_ (.Y(_05418_),
    .B(net670),
    .A_N(_00101_));
 sg13g2_o21ai_1 _23085_ (.B1(_05418_),
    .Y(_05419_),
    .A1(_00102_),
    .A2(_04848_));
 sg13g2_a221oi_1 _23086_ (.B2(_05334_),
    .C1(_05419_),
    .B1(_05417_),
    .A1(_12084_),
    .Y(_05420_),
    .A2(_05416_));
 sg13g2_buf_1 _23087_ (.A(\cpu.gpio.r_src_io[4][2] ),
    .X(_05421_));
 sg13g2_nand2b_1 _23088_ (.Y(_05422_),
    .B(_04863_),
    .A_N(_00100_));
 sg13g2_o21ai_1 _23089_ (.B1(_05422_),
    .Y(_05423_),
    .A1(_00098_),
    .A2(_05080_));
 sg13g2_a221oi_1 _23090_ (.B2(_09136_),
    .C1(_05423_),
    .B1(_04891_),
    .A1(_05421_),
    .Y(_05424_),
    .A2(net413));
 sg13g2_nand3_1 _23091_ (.B(_09137_),
    .C(_04888_),
    .A(_09136_),
    .Y(_05425_));
 sg13g2_nand3_1 _23092_ (.B(_05424_),
    .C(_05425_),
    .A(_05420_),
    .Y(_05426_));
 sg13g2_buf_1 _23093_ (.A(\cpu.spi.r_clk_count[2][2] ),
    .X(_05427_));
 sg13g2_nand2_1 _23094_ (.Y(_05428_),
    .A(net899),
    .B(_12056_));
 sg13g2_o21ai_1 _23095_ (.B1(_05428_),
    .Y(_05429_),
    .A1(net899),
    .A2(_12052_));
 sg13g2_a22oi_1 _23096_ (.Y(_05430_),
    .B1(_05429_),
    .B2(net411),
    .A2(_05105_),
    .A1(\cpu.spi.r_timeout[2] ));
 sg13g2_o21ai_1 _23097_ (.B1(_05430_),
    .Y(_05431_),
    .A1(_00097_),
    .A2(_05107_));
 sg13g2_a21oi_1 _23098_ (.A1(_05427_),
    .A2(_04952_),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_nand2b_1 _23099_ (.Y(_05433_),
    .B(net670),
    .A_N(_00276_));
 sg13g2_or2_1 _23100_ (.X(_05434_),
    .B(_04949_),
    .A(_00096_));
 sg13g2_nand2_1 _23101_ (.Y(_05435_),
    .A(_09220_),
    .B(_04943_));
 sg13g2_nand4_1 _23102_ (.B(_05433_),
    .C(_05434_),
    .A(_05432_),
    .Y(_05436_),
    .D(_05435_));
 sg13g2_nor3_1 _23103_ (.A(_09880_),
    .B(net518),
    .C(net668),
    .Y(_05437_));
 sg13g2_a221oi_1 _23104_ (.B2(\cpu.uart.r_in[2] ),
    .C1(_05437_),
    .B1(_04964_),
    .A1(\cpu.uart.r_div_value[2] ),
    .Y(_05438_),
    .A2(net375));
 sg13g2_o21ai_1 _23105_ (.B1(net1166),
    .Y(_05439_),
    .A1(net516),
    .A2(_05438_));
 sg13g2_a221oi_1 _23106_ (.B2(_09170_),
    .C1(_05439_),
    .B1(_05436_),
    .A1(_04896_),
    .Y(_05440_),
    .A2(_05426_));
 sg13g2_o21ai_1 _23107_ (.B1(_05440_),
    .Y(_05441_),
    .A1(_04959_),
    .A2(_05415_));
 sg13g2_o21ai_1 _23108_ (.B1(_05441_),
    .Y(_05442_),
    .A1(net1001),
    .A2(_05404_));
 sg13g2_mux2_1 _23109_ (.A0(_05442_),
    .A1(net767),
    .S(net69),
    .X(_05443_));
 sg13g2_o21ai_1 _23110_ (.B1(net247),
    .Y(_05444_),
    .A1(net819),
    .A2(net600));
 sg13g2_nand2_1 _23111_ (.Y(_05445_),
    .A(net664),
    .B(_04472_));
 sg13g2_o21ai_1 _23112_ (.B1(_05445_),
    .Y(_05446_),
    .A1(_05161_),
    .A2(_04470_));
 sg13g2_a221oi_1 _23113_ (.B2(net211),
    .C1(net130),
    .B1(_05446_),
    .A1(net718),
    .Y(_05447_),
    .A2(_05444_));
 sg13g2_a21oi_1 _23114_ (.A1(net131),
    .A2(_05443_),
    .Y(_01027_),
    .B1(_05447_));
 sg13g2_buf_1 _23115_ (.A(net132),
    .X(_05448_));
 sg13g2_a21oi_1 _23116_ (.A1(_05161_),
    .A2(_04478_),
    .Y(_05449_),
    .B1(net291));
 sg13g2_nand2_1 _23117_ (.Y(_05450_),
    .A(_05160_),
    .B(_04223_));
 sg13g2_o21ai_1 _23118_ (.B1(_05450_),
    .Y(_05451_),
    .A1(_05160_),
    .A2(_04512_));
 sg13g2_nand2_1 _23119_ (.Y(_05452_),
    .A(_05157_),
    .B(_05451_));
 sg13g2_o21ai_1 _23120_ (.B1(_05452_),
    .Y(_05453_),
    .A1(net649),
    .A2(_05449_));
 sg13g2_buf_1 _23121_ (.A(net175),
    .X(_05454_));
 sg13g2_a22oi_1 _23122_ (.Y(_05455_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][3] ),
    .A2(net463),
    .A1(\cpu.dcache.r_data[0][3] ));
 sg13g2_a22oi_1 _23123_ (.Y(_05456_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][3] ),
    .A2(net425),
    .A1(\cpu.dcache.r_data[1][3] ));
 sg13g2_a22oi_1 _23124_ (.Y(_05457_),
    .B1(net420),
    .B2(\cpu.dcache.r_data[7][3] ),
    .A2(net422),
    .A1(\cpu.dcache.r_data[5][3] ));
 sg13g2_a22oi_1 _23125_ (.Y(_05458_),
    .B1(net423),
    .B2(\cpu.dcache.r_data[3][3] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[6][3] ));
 sg13g2_nand4_1 _23126_ (.B(_05456_),
    .C(_05457_),
    .A(_05455_),
    .Y(_05459_),
    .D(_05458_));
 sg13g2_inv_1 _23127_ (.Y(_05460_),
    .A(_00104_));
 sg13g2_a22oi_1 _23128_ (.Y(_05461_),
    .B1(net480),
    .B2(\cpu.dcache.r_data[5][19] ),
    .A2(net463),
    .A1(_05460_));
 sg13g2_a22oi_1 _23129_ (.Y(_05462_),
    .B1(net425),
    .B2(\cpu.dcache.r_data[1][19] ),
    .A2(net421),
    .A1(\cpu.dcache.r_data[6][19] ));
 sg13g2_a22oi_1 _23130_ (.Y(_05463_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][19] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][19] ));
 sg13g2_a22oi_1 _23131_ (.Y(_05464_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][19] ),
    .A2(net478),
    .A1(\cpu.dcache.r_data[7][19] ));
 sg13g2_nand4_1 _23132_ (.B(_05462_),
    .C(_05463_),
    .A(_05461_),
    .Y(_05465_),
    .D(_05464_));
 sg13g2_buf_1 _23133_ (.A(_05465_),
    .X(_05466_));
 sg13g2_a22oi_1 _23134_ (.Y(_05467_),
    .B1(_05466_),
    .B2(_05042_),
    .A2(_05459_),
    .A1(net1030));
 sg13g2_a221oi_1 _23135_ (.B2(net898),
    .C1(net598),
    .B1(_05182_),
    .A1(_09890_),
    .Y(_05468_),
    .A2(_05174_));
 sg13g2_a21oi_1 _23136_ (.A1(net598),
    .A2(_05467_),
    .Y(_05469_),
    .B1(_05468_));
 sg13g2_mux2_1 _23137_ (.A0(_05459_),
    .A1(_05466_),
    .S(_10027_),
    .X(_05470_));
 sg13g2_mux2_1 _23138_ (.A0(_05469_),
    .A1(_05470_),
    .S(net603),
    .X(_05471_));
 sg13g2_buf_1 _23139_ (.A(\cpu.spi.r_clk_count[2][3] ),
    .X(_05472_));
 sg13g2_nor2_1 _23140_ (.A(_00108_),
    .B(_05107_),
    .Y(_05473_));
 sg13g2_a221oi_1 _23141_ (.B2(\cpu.spi.r_timeout[3] ),
    .C1(_05473_),
    .B1(_05105_),
    .A1(_05472_),
    .Y(_05474_),
    .A2(_04952_));
 sg13g2_o21ai_1 _23142_ (.B1(_05474_),
    .Y(_05475_),
    .A1(_00107_),
    .A2(_04949_));
 sg13g2_a21oi_1 _23143_ (.A1(_09215_),
    .A2(_04943_),
    .Y(_05476_),
    .B1(_05475_));
 sg13g2_nand2_1 _23144_ (.Y(_05477_),
    .A(net796),
    .B(net422));
 sg13g2_nand2_1 _23145_ (.Y(_05478_),
    .A(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .B(net412));
 sg13g2_o21ai_1 _23146_ (.B1(_05478_),
    .Y(_05479_),
    .A1(_00112_),
    .A2(_05477_));
 sg13g2_a22oi_1 _23147_ (.Y(_05480_),
    .B1(net411),
    .B2(_09144_),
    .A2(_04913_),
    .A1(_09145_));
 sg13g2_inv_1 _23148_ (.Y(_05481_),
    .A(_00109_));
 sg13g2_buf_1 _23149_ (.A(\cpu.gpio.r_src_io[4][3] ),
    .X(_05482_));
 sg13g2_nand2b_1 _23150_ (.Y(_05483_),
    .B(_04863_),
    .A_N(_00111_));
 sg13g2_o21ai_1 _23151_ (.B1(_05483_),
    .Y(_05484_),
    .A1(_00110_),
    .A2(_05340_));
 sg13g2_a221oi_1 _23152_ (.B2(_05482_),
    .C1(_05484_),
    .B1(net413),
    .A1(_05481_),
    .Y(_05485_),
    .A2(_04869_));
 sg13g2_o21ai_1 _23153_ (.B1(_05485_),
    .Y(_05486_),
    .A1(net899),
    .A2(_05480_));
 sg13g2_a21oi_1 _23154_ (.A1(net869),
    .A2(_05479_),
    .Y(_05487_),
    .B1(_05486_));
 sg13g2_nand3_1 _23155_ (.B(_09145_),
    .C(_04888_),
    .A(_09144_),
    .Y(_05488_));
 sg13g2_nand2_1 _23156_ (.Y(_05489_),
    .A(_05487_),
    .B(_05488_));
 sg13g2_mux2_1 _23157_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(\cpu.intr.r_clock_cmp[19] ),
    .S(net676),
    .X(_05490_));
 sg13g2_mux2_1 _23158_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(\cpu.intr.r_timer_reload[19] ),
    .S(net676),
    .X(_05491_));
 sg13g2_a22oi_1 _23159_ (.Y(_05492_),
    .B1(_05491_),
    .B2(net420),
    .A2(_05490_),
    .A1(net422));
 sg13g2_mux2_1 _23160_ (.A0(\cpu.intr.r_timer_count[3] ),
    .A1(_09901_),
    .S(net676),
    .X(_05493_));
 sg13g2_a22oi_1 _23161_ (.Y(_05494_),
    .B1(_05493_),
    .B2(net380),
    .A2(net517),
    .A1(_09118_));
 sg13g2_buf_1 _23162_ (.A(\cpu.intr.r_clock_count[19] ),
    .X(_05495_));
 sg13g2_a22oi_1 _23163_ (.Y(_05496_),
    .B1(net374),
    .B2(_10049_),
    .A2(net340),
    .A1(_05495_));
 sg13g2_a21oi_1 _23164_ (.A1(_09118_),
    .A2(_04903_),
    .Y(_05497_),
    .B1(net408));
 sg13g2_nand2b_1 _23165_ (.Y(_05498_),
    .B(\cpu.intr.r_enable[3] ),
    .A_N(_05497_));
 sg13g2_nand4_1 _23166_ (.B(_05494_),
    .C(_05496_),
    .A(_05492_),
    .Y(_05499_),
    .D(_05498_));
 sg13g2_and2_1 _23167_ (.A(\cpu.uart.r_div_value[11] ),
    .B(net409),
    .X(_05500_));
 sg13g2_a221oi_1 _23168_ (.B2(\cpu.uart.r_in[3] ),
    .C1(_05500_),
    .B1(_04964_),
    .A1(\cpu.uart.r_div_value[3] ),
    .Y(_05501_),
    .A2(net375));
 sg13g2_o21ai_1 _23169_ (.B1(net1166),
    .Y(_05502_),
    .A1(net516),
    .A2(_05501_));
 sg13g2_a221oi_1 _23170_ (.B2(_09897_),
    .C1(_05502_),
    .B1(_05499_),
    .A1(_04896_),
    .Y(_05503_),
    .A2(_05489_));
 sg13g2_o21ai_1 _23171_ (.B1(_05503_),
    .Y(_05504_),
    .A1(_05369_),
    .A2(_05476_));
 sg13g2_o21ai_1 _23172_ (.B1(_05504_),
    .Y(_05505_),
    .A1(net1001),
    .A2(_05471_));
 sg13g2_nand2_1 _23173_ (.Y(_05506_),
    .A(net418),
    .B(net68));
 sg13g2_o21ai_1 _23174_ (.B1(_05506_),
    .Y(_05507_),
    .A1(net69),
    .A2(_05505_));
 sg13g2_nor2_1 _23175_ (.A(net129),
    .B(_05507_),
    .Y(_05508_));
 sg13g2_a21oi_1 _23176_ (.A1(net100),
    .A2(_05453_),
    .Y(_01028_),
    .B1(_05508_));
 sg13g2_a22oi_1 _23177_ (.Y(_05509_),
    .B1(net640),
    .B2(\cpu.dcache.r_data[4][4] ),
    .A2(net546),
    .A1(\cpu.dcache.r_data[3][4] ));
 sg13g2_a22oi_1 _23178_ (.Y(_05510_),
    .B1(net544),
    .B2(\cpu.dcache.r_data[6][4] ),
    .A2(net639),
    .A1(\cpu.dcache.r_data[5][4] ));
 sg13g2_nand2_1 _23179_ (.Y(_05511_),
    .A(_05509_),
    .B(_05510_));
 sg13g2_a221oi_1 _23180_ (.B2(\cpu.dcache.r_data[2][4] ),
    .C1(_05511_),
    .B1(net482),
    .A1(\cpu.dcache.r_data[7][4] ),
    .Y(_05512_),
    .A2(net543));
 sg13g2_mux2_1 _23181_ (.A0(_00114_),
    .A1(_05512_),
    .S(_04859_),
    .X(_05513_));
 sg13g2_nor2_1 _23182_ (.A(\cpu.dcache.r_data[1][4] ),
    .B(net699),
    .Y(_05514_));
 sg13g2_a22oi_1 _23183_ (.Y(_05515_),
    .B1(_05514_),
    .B2(_05512_),
    .A2(_05513_),
    .A1(net699));
 sg13g2_inv_1 _23184_ (.Y(_05516_),
    .A(_00115_));
 sg13g2_a22oi_1 _23185_ (.Y(_05517_),
    .B1(net482),
    .B2(\cpu.dcache.r_data[2][20] ),
    .A2(net514),
    .A1(_05516_));
 sg13g2_a22oi_1 _23186_ (.Y(_05518_),
    .B1(net483),
    .B2(\cpu.dcache.r_data[1][20] ),
    .A2(net479),
    .A1(\cpu.dcache.r_data[6][20] ));
 sg13g2_a22oi_1 _23187_ (.Y(_05519_),
    .B1(net543),
    .B2(\cpu.dcache.r_data[7][20] ),
    .A2(net545),
    .A1(\cpu.dcache.r_data[5][20] ));
 sg13g2_a22oi_1 _23188_ (.Y(_05520_),
    .B1(net567),
    .B2(\cpu.dcache.r_data[4][20] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[3][20] ));
 sg13g2_nand4_1 _23189_ (.B(_05518_),
    .C(_05519_),
    .A(_05517_),
    .Y(_05521_),
    .D(_05520_));
 sg13g2_buf_1 _23190_ (.A(_05521_),
    .X(_05522_));
 sg13g2_and2_1 _23191_ (.A(_10027_),
    .B(_05522_),
    .X(_05523_));
 sg13g2_a21oi_1 _23192_ (.A1(net694),
    .A2(_05515_),
    .Y(_05524_),
    .B1(_05523_));
 sg13g2_a22oi_1 _23193_ (.Y(_05525_),
    .B1(_05522_),
    .B2(_05042_),
    .A2(_05515_),
    .A1(net1030));
 sg13g2_nor2_1 _23194_ (.A(net1030),
    .B(_05197_),
    .Y(_05526_));
 sg13g2_nor3_1 _23195_ (.A(net598),
    .B(_05205_),
    .C(_05526_),
    .Y(_05527_));
 sg13g2_a21oi_1 _23196_ (.A1(net598),
    .A2(_05525_),
    .Y(_05528_),
    .B1(_05527_));
 sg13g2_nor2_1 _23197_ (.A(_04978_),
    .B(_05528_),
    .Y(_05529_));
 sg13g2_a21oi_1 _23198_ (.A1(net603),
    .A2(_05524_),
    .Y(_05530_),
    .B1(_05529_));
 sg13g2_a22oi_1 _23199_ (.Y(_05531_),
    .B1(_04964_),
    .B2(\cpu.uart.r_in[4] ),
    .A2(net375),
    .A1(\cpu.uart.r_div_value[4] ));
 sg13g2_nor2_1 _23200_ (.A(net516),
    .B(_05531_),
    .Y(_05532_));
 sg13g2_buf_1 _23201_ (.A(\cpu.spi.r_clk_count[2][4] ),
    .X(_05533_));
 sg13g2_nor2_1 _23202_ (.A(_00119_),
    .B(_05107_),
    .Y(_05534_));
 sg13g2_a221oi_1 _23203_ (.B2(\cpu.spi.r_timeout[4] ),
    .C1(_05534_),
    .B1(_05105_),
    .A1(_05533_),
    .Y(_05535_),
    .A2(_04952_));
 sg13g2_o21ai_1 _23204_ (.B1(_05535_),
    .Y(_05536_),
    .A1(_00118_),
    .A2(_04949_));
 sg13g2_a21oi_1 _23205_ (.A1(_09222_),
    .A2(_04943_),
    .Y(_05537_),
    .B1(_05536_));
 sg13g2_a22oi_1 _23206_ (.Y(_05538_),
    .B1(net441),
    .B2(_10053_),
    .A2(net422),
    .A1(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_mux2_1 _23207_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(\cpu.intr.r_timer_reload[20] ),
    .S(net931),
    .X(_05539_));
 sg13g2_mux2_1 _23208_ (.A0(\cpu.intr.r_timer_count[4] ),
    .A1(_09925_),
    .S(net931),
    .X(_05540_));
 sg13g2_a22oi_1 _23209_ (.Y(_05541_),
    .B1(_05540_),
    .B2(net421),
    .A2(_05539_),
    .A1(net478));
 sg13g2_buf_2 _23210_ (.A(\cpu.intr.r_clock_count[20] ),
    .X(_05542_));
 sg13g2_a22oi_1 _23211_ (.Y(_05543_),
    .B1(net376),
    .B2(_05542_),
    .A2(_04913_),
    .A1(_09155_));
 sg13g2_nand2_1 _23212_ (.Y(_05544_),
    .A(_05541_),
    .B(_05543_));
 sg13g2_a21oi_1 _23213_ (.A1(\cpu.intr.r_clock_cmp[20] ),
    .A2(net602),
    .Y(_05545_),
    .B1(_05544_));
 sg13g2_o21ai_1 _23214_ (.B1(_05545_),
    .Y(_05546_),
    .A1(net695),
    .A2(_05538_));
 sg13g2_o21ai_1 _23215_ (.B1(net771),
    .Y(_05547_),
    .A1(net418),
    .A2(net604));
 sg13g2_a21oi_1 _23216_ (.A1(_09135_),
    .A2(_09154_),
    .Y(_05548_),
    .B1(_05547_));
 sg13g2_a21oi_1 _23217_ (.A1(_09156_),
    .A2(_04903_),
    .Y(_05549_),
    .B1(_04959_));
 sg13g2_o21ai_1 _23218_ (.B1(_05549_),
    .Y(_05550_),
    .A1(_05546_),
    .A2(_05548_));
 sg13g2_o21ai_1 _23219_ (.B1(_05550_),
    .Y(_05551_),
    .A1(_05369_),
    .A2(_05537_));
 sg13g2_a21o_1 _23220_ (.A2(_05097_),
    .A1(_09141_),
    .B1(net410),
    .X(_05552_));
 sg13g2_a22oi_1 _23221_ (.Y(_05553_),
    .B1(_05145_),
    .B2(net7),
    .A2(net412),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_buf_2 _23222_ (.A(\cpu.gpio.r_spi_miso_src[1][0] ),
    .X(_05554_));
 sg13g2_a22oi_1 _23223_ (.Y(_05555_),
    .B1(net376),
    .B2(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A2(_04847_),
    .A1(_05554_));
 sg13g2_nand2_1 _23224_ (.Y(_05556_),
    .A(_05553_),
    .B(_05555_));
 sg13g2_buf_2 _23225_ (.A(\cpu.gpio.r_src_io[7][0] ),
    .X(_05557_));
 sg13g2_buf_2 _23226_ (.A(\cpu.gpio.r_src_io[5][0] ),
    .X(_05558_));
 sg13g2_buf_2 _23227_ (.A(\cpu.gpio.r_src_o[7][0] ),
    .X(_05559_));
 sg13g2_a22oi_1 _23228_ (.Y(_05560_),
    .B1(_05559_),
    .B2(net1061),
    .A2(net869),
    .A1(_09141_));
 sg13g2_buf_2 _23229_ (.A(\cpu.gpio.r_src_o[5][0] ),
    .X(_05561_));
 sg13g2_a22oi_1 _23230_ (.Y(_05562_),
    .B1(_09564_),
    .B2(_05561_),
    .A2(net900),
    .A1(_09147_));
 sg13g2_nand2b_1 _23231_ (.Y(_05563_),
    .B(_04913_),
    .A_N(_05562_));
 sg13g2_o21ai_1 _23232_ (.B1(_05563_),
    .Y(_05564_),
    .A1(_05088_),
    .A2(_05560_));
 sg13g2_a221oi_1 _23233_ (.B2(_05558_),
    .C1(_05564_),
    .B1(_04871_),
    .A1(_05557_),
    .Y(_05565_),
    .A2(_04869_));
 sg13g2_nand3_1 _23234_ (.B(net900),
    .C(net411),
    .A(_09146_),
    .Y(_05566_));
 sg13g2_buf_2 _23235_ (.A(\cpu.gpio.r_src_o[3][0] ),
    .X(_05567_));
 sg13g2_nand3_1 _23236_ (.B(_05567_),
    .C(_04905_),
    .A(net899),
    .Y(_05568_));
 sg13g2_nand3_1 _23237_ (.B(_05566_),
    .C(_05568_),
    .A(_05565_),
    .Y(_05569_));
 sg13g2_a221oi_1 _23238_ (.B2(net869),
    .C1(_05569_),
    .B1(_05556_),
    .A1(\cpu.gpio.r_enable_io[4] ),
    .Y(_05570_),
    .A2(_05552_));
 sg13g2_nand3_1 _23239_ (.B(_09147_),
    .C(_04888_),
    .A(_09146_),
    .Y(_05571_));
 sg13g2_a21oi_1 _23240_ (.A1(_05570_),
    .A2(_05571_),
    .Y(_05572_),
    .B1(_05077_));
 sg13g2_or4_1 _23241_ (.A(net1067),
    .B(_05532_),
    .C(_05551_),
    .D(_05572_),
    .X(_05573_));
 sg13g2_o21ai_1 _23242_ (.B1(_05573_),
    .Y(_05574_),
    .A1(net1001),
    .A2(_05530_));
 sg13g2_nor2_1 _23243_ (.A(net69),
    .B(_05574_),
    .Y(_05575_));
 sg13g2_a21oi_1 _23244_ (.A1(net616),
    .A2(net69),
    .Y(_05576_),
    .B1(_05575_));
 sg13g2_o21ai_1 _23245_ (.B1(net247),
    .Y(_05577_),
    .A1(net600),
    .A2(_04223_));
 sg13g2_nand2_1 _23246_ (.Y(_05578_),
    .A(net664),
    .B(_04545_));
 sg13g2_o21ai_1 _23247_ (.B1(_05578_),
    .Y(_05579_),
    .A1(net599),
    .A2(_04542_));
 sg13g2_a221oi_1 _23248_ (.B2(net211),
    .C1(net130),
    .B1(_05579_),
    .A1(net1159),
    .Y(_05580_),
    .A2(_05577_));
 sg13g2_a21oi_1 _23249_ (.A1(net131),
    .A2(_05576_),
    .Y(_01029_),
    .B1(_05580_));
 sg13g2_and2_1 _23250_ (.A(net664),
    .B(_04578_),
    .X(_05581_));
 sg13g2_a21oi_1 _23251_ (.A1(net600),
    .A2(_04575_),
    .Y(_05582_),
    .B1(_05581_));
 sg13g2_nand2_1 _23252_ (.Y(_05583_),
    .A(net988),
    .B(net291));
 sg13g2_o21ai_1 _23253_ (.B1(_05583_),
    .Y(_05584_),
    .A1(net291),
    .A2(_05582_));
 sg13g2_inv_1 _23254_ (.Y(_05585_),
    .A(_00121_));
 sg13g2_a22oi_1 _23255_ (.Y(_05586_),
    .B1(net424),
    .B2(\cpu.dcache.r_data[2][5] ),
    .A2(net463),
    .A1(_05585_));
 sg13g2_a22oi_1 _23256_ (.Y(_05587_),
    .B1(net425),
    .B2(\cpu.dcache.r_data[1][5] ),
    .A2(net380),
    .A1(\cpu.dcache.r_data[6][5] ));
 sg13g2_a22oi_1 _23257_ (.Y(_05588_),
    .B1(net420),
    .B2(\cpu.dcache.r_data[7][5] ),
    .A2(net422),
    .A1(\cpu.dcache.r_data[5][5] ));
 sg13g2_a22oi_1 _23258_ (.Y(_05589_),
    .B1(net441),
    .B2(\cpu.dcache.r_data[4][5] ),
    .A2(net423),
    .A1(\cpu.dcache.r_data[3][5] ));
 sg13g2_and4_1 _23259_ (.A(_05586_),
    .B(_05587_),
    .C(_05588_),
    .D(_05589_),
    .X(_05590_));
 sg13g2_buf_1 _23260_ (.A(_05590_),
    .X(_05591_));
 sg13g2_a221oi_1 _23261_ (.B2(net694),
    .C1(net598),
    .B1(_05238_),
    .A1(net898),
    .Y(_05592_),
    .A2(_05230_));
 sg13g2_a21o_1 _23262_ (.A2(_05591_),
    .A1(_05005_),
    .B1(_05592_),
    .X(_05593_));
 sg13g2_a22oi_1 _23263_ (.Y(_05594_),
    .B1(net478),
    .B2(\cpu.dcache.r_data[7][21] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[3][21] ));
 sg13g2_a22oi_1 _23264_ (.Y(_05595_),
    .B1(net421),
    .B2(\cpu.dcache.r_data[6][21] ),
    .A2(net480),
    .A1(\cpu.dcache.r_data[5][21] ));
 sg13g2_a22oi_1 _23265_ (.Y(_05596_),
    .B1(net482),
    .B2(\cpu.dcache.r_data[2][21] ),
    .A2(net491),
    .A1(\cpu.dcache.r_data[4][21] ));
 sg13g2_nand3_1 _23266_ (.B(_05595_),
    .C(_05596_),
    .A(_05594_),
    .Y(_05597_));
 sg13g2_nand2_1 _23267_ (.Y(_05598_),
    .A(_00122_),
    .B(_04852_));
 sg13g2_o21ai_1 _23268_ (.B1(_05598_),
    .Y(_05599_),
    .A1(_04852_),
    .A2(_05597_));
 sg13g2_o21ai_1 _23269_ (.B1(net425),
    .Y(_05600_),
    .A1(\cpu.dcache.r_data[1][21] ),
    .A2(_05597_));
 sg13g2_o21ai_1 _23270_ (.B1(_05600_),
    .Y(_05601_),
    .A1(net425),
    .A2(_05599_));
 sg13g2_nand2_1 _23271_ (.Y(_05602_),
    .A(net898),
    .B(net598));
 sg13g2_o21ai_1 _23272_ (.B1(_04978_),
    .Y(_05603_),
    .A1(net566),
    .A2(_05591_));
 sg13g2_a22oi_1 _23273_ (.Y(_05604_),
    .B1(_05602_),
    .B2(_05603_),
    .A2(_05601_),
    .A1(net566));
 sg13g2_a21oi_1 _23274_ (.A1(_05027_),
    .A2(_05593_),
    .Y(_05605_),
    .B1(_05604_));
 sg13g2_buf_1 _23275_ (.A(\cpu.spi.r_clk_count[2][5] ),
    .X(_05606_));
 sg13g2_nor2_1 _23276_ (.A(_00126_),
    .B(_05107_),
    .Y(_05607_));
 sg13g2_a221oi_1 _23277_ (.B2(\cpu.spi.r_timeout[5] ),
    .C1(_05607_),
    .B1(_05105_),
    .A1(_05606_),
    .Y(_05608_),
    .A2(_04952_));
 sg13g2_o21ai_1 _23278_ (.B1(_05608_),
    .Y(_05609_),
    .A1(_00125_),
    .A2(_04949_));
 sg13g2_a21o_1 _23279_ (.A2(_04943_),
    .A1(_09221_),
    .B1(_05609_),
    .X(_05610_));
 sg13g2_nand3_1 _23280_ (.B(_09128_),
    .C(_04888_),
    .A(_09127_),
    .Y(_05611_));
 sg13g2_a21oi_1 _23281_ (.A1(_09142_),
    .A2(_05097_),
    .Y(_05612_),
    .B1(_04941_));
 sg13g2_nand2b_1 _23282_ (.Y(_05613_),
    .B(\cpu.gpio.r_enable_io[5] ),
    .A_N(_05612_));
 sg13g2_a22oi_1 _23283_ (.Y(_05614_),
    .B1(net515),
    .B2(_09142_),
    .A2(net376),
    .A1(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_nand2_1 _23284_ (.Y(_05615_),
    .A(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .B(net412));
 sg13g2_inv_1 _23285_ (.Y(_05616_),
    .A(_00131_));
 sg13g2_a22oi_1 _23286_ (.Y(_05617_),
    .B1(_05145_),
    .B2(net8),
    .A2(_04847_),
    .A1(_05616_));
 sg13g2_nand3_1 _23287_ (.B(_05615_),
    .C(_05617_),
    .A(_05614_),
    .Y(_05618_));
 sg13g2_nand2_1 _23288_ (.Y(_05619_),
    .A(net869),
    .B(_05618_));
 sg13g2_nand2_1 _23289_ (.Y(_05620_),
    .A(_12083_),
    .B(net517));
 sg13g2_inv_1 _23290_ (.Y(_05621_),
    .A(_00129_));
 sg13g2_buf_2 _23291_ (.A(\cpu.gpio.r_src_io[5][1] ),
    .X(_05622_));
 sg13g2_a22oi_1 _23292_ (.Y(_05623_),
    .B1(net413),
    .B2(_05622_),
    .A2(_04863_),
    .A1(_05621_));
 sg13g2_o21ai_1 _23293_ (.B1(_05623_),
    .Y(_05624_),
    .A1(_00130_),
    .A2(_05620_));
 sg13g2_a22oi_1 _23294_ (.Y(_05625_),
    .B1(net411),
    .B2(_09127_),
    .A2(_04913_),
    .A1(_09128_));
 sg13g2_nor2_1 _23295_ (.A(_12084_),
    .B(_05625_),
    .Y(_05626_));
 sg13g2_nor2_1 _23296_ (.A(_00128_),
    .B(_05340_),
    .Y(_05627_));
 sg13g2_nor2_1 _23297_ (.A(_00127_),
    .B(_05080_),
    .Y(_05628_));
 sg13g2_nor4_1 _23298_ (.A(_05624_),
    .B(_05626_),
    .C(_05627_),
    .D(_05628_),
    .Y(_05629_));
 sg13g2_nand4_1 _23299_ (.B(_05613_),
    .C(_05619_),
    .A(_05611_),
    .Y(_05630_),
    .D(_05629_));
 sg13g2_a22oi_1 _23300_ (.Y(_05631_),
    .B1(_04964_),
    .B2(\cpu.uart.r_in[5] ),
    .A2(net375),
    .A1(\cpu.uart.r_div_value[5] ));
 sg13g2_a22oi_1 _23301_ (.Y(_05632_),
    .B1(net420),
    .B2(\cpu.intr.r_timer_reload[21] ),
    .A2(net380),
    .A1(_09924_));
 sg13g2_a221oi_1 _23302_ (.B2(_10059_),
    .C1(net796),
    .B1(net441),
    .A1(\cpu.intr.r_timer_count[5] ),
    .Y(_05633_),
    .A2(net421));
 sg13g2_a21o_1 _23303_ (.A2(_05632_),
    .A1(net695),
    .B1(_05633_),
    .X(_05634_));
 sg13g2_nand2_1 _23304_ (.Y(_05635_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(net601));
 sg13g2_buf_1 _23305_ (.A(\cpu.intr.r_clock_count[21] ),
    .X(_05636_));
 sg13g2_a22oi_1 _23306_ (.Y(_05637_),
    .B1(net376),
    .B2(_05636_),
    .A2(net408),
    .A1(_09120_));
 sg13g2_a22oi_1 _23307_ (.Y(_05638_),
    .B1(net341),
    .B2(\cpu.intr.r_timer_reload[5] ),
    .A2(_04847_),
    .A1(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_nand4_1 _23308_ (.B(_05635_),
    .C(_05637_),
    .A(_05634_),
    .Y(_05639_),
    .D(_05638_));
 sg13g2_a21oi_1 _23309_ (.A1(_09120_),
    .A2(_04903_),
    .Y(_05640_),
    .B1(_04905_));
 sg13g2_nor2b_1 _23310_ (.A(_05640_),
    .B_N(_09119_),
    .Y(_05641_));
 sg13g2_o21ai_1 _23311_ (.B1(_09897_),
    .Y(_05642_),
    .A1(_05639_),
    .A2(_05641_));
 sg13g2_o21ai_1 _23312_ (.B1(_05642_),
    .Y(_05643_),
    .A1(net516),
    .A2(_05631_));
 sg13g2_a221oi_1 _23313_ (.B2(_04896_),
    .C1(_05643_),
    .B1(_05630_),
    .A1(_09170_),
    .Y(_05644_),
    .A2(_05610_));
 sg13g2_nand2_1 _23314_ (.Y(_05645_),
    .A(net1001),
    .B(_05644_));
 sg13g2_o21ai_1 _23315_ (.B1(_05645_),
    .Y(_05646_),
    .A1(_03011_),
    .A2(_05605_));
 sg13g2_nand2_1 _23316_ (.Y(_05647_),
    .A(net620),
    .B(net69));
 sg13g2_o21ai_1 _23317_ (.B1(_05647_),
    .Y(_05648_),
    .A1(net69),
    .A2(_05646_));
 sg13g2_mux2_1 _23318_ (.A0(_05584_),
    .A1(_05648_),
    .S(net131),
    .X(_01030_));
 sg13g2_a21oi_1 _23319_ (.A1(net599),
    .A2(_04613_),
    .Y(_05649_),
    .B1(net291));
 sg13g2_o21ai_1 _23320_ (.B1(_05649_),
    .Y(_05650_),
    .A1(net599),
    .A2(_04610_));
 sg13g2_o21ai_1 _23321_ (.B1(net175),
    .Y(_05651_),
    .A1(net987),
    .A2(net211));
 sg13g2_inv_1 _23322_ (.Y(_05652_),
    .A(_05651_));
 sg13g2_mux2_1 _23323_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(\cpu.intr.r_timer_reload[22] ),
    .S(net493),
    .X(_05653_));
 sg13g2_a22oi_1 _23324_ (.Y(_05654_),
    .B1(_05653_),
    .B2(net622),
    .A2(net666),
    .A1(_09927_));
 sg13g2_nand3b_1 _23325_ (.B(_12077_),
    .C(net695),
    .Y(_05655_),
    .A_N(_05654_));
 sg13g2_a22oi_1 _23326_ (.Y(_05656_),
    .B1(net420),
    .B2(\cpu.intr.r_timer_reload[6] ),
    .A2(net480),
    .A1(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_or2_1 _23327_ (.X(_05657_),
    .B(_05656_),
    .A(net676));
 sg13g2_nand2_1 _23328_ (.Y(_05658_),
    .A(_10065_),
    .B(_04923_));
 sg13g2_buf_1 _23329_ (.A(\cpu.intr.r_clock_count[22] ),
    .X(_05659_));
 sg13g2_a22oi_1 _23330_ (.Y(_05660_),
    .B1(_04918_),
    .B2(_05659_),
    .A2(_04928_),
    .A1(\cpu.intr.r_timer_count[6] ));
 sg13g2_nand4_1 _23331_ (.B(_05657_),
    .C(_05658_),
    .A(_05655_),
    .Y(_05661_),
    .D(_05660_));
 sg13g2_nor2_1 _23332_ (.A(_00139_),
    .B(_05080_),
    .Y(_05662_));
 sg13g2_a221oi_1 _23333_ (.B2(_09130_),
    .C1(_05662_),
    .B1(_04941_),
    .A1(_09150_),
    .Y(_05663_),
    .A2(_04891_));
 sg13g2_buf_1 _23334_ (.A(\cpu.gpio.r_src_io[5][2] ),
    .X(_05664_));
 sg13g2_nand2b_1 _23335_ (.Y(_05665_),
    .B(_04904_),
    .A_N(_00142_));
 sg13g2_o21ai_1 _23336_ (.B1(_05665_),
    .Y(_05666_),
    .A1(_00140_),
    .A2(_05088_));
 sg13g2_inv_1 _23337_ (.Y(_05667_),
    .A(_00141_));
 sg13g2_a22oi_1 _23338_ (.Y(_05668_),
    .B1(_09564_),
    .B2(_05667_),
    .A2(net900),
    .A1(_09151_));
 sg13g2_nor3_1 _23339_ (.A(net747),
    .B(net604),
    .C(_05668_),
    .Y(_05669_));
 sg13g2_a221oi_1 _23340_ (.B2(_12083_),
    .C1(_05669_),
    .B1(_05666_),
    .A1(_05664_),
    .Y(_05670_),
    .A2(net413));
 sg13g2_inv_1 _23341_ (.Y(_05671_),
    .A(_09131_));
 sg13g2_a21oi_1 _23342_ (.A1(_09130_),
    .A2(_04904_),
    .Y(_05672_),
    .B1(net515));
 sg13g2_nand2b_1 _23343_ (.Y(_05673_),
    .B(_09179_),
    .A_N(_00143_));
 sg13g2_nand2_1 _23344_ (.Y(_05674_),
    .A(net923),
    .B(net9));
 sg13g2_a21oi_1 _23345_ (.A1(_05673_),
    .A2(_05674_),
    .Y(_05675_),
    .B1(net924));
 sg13g2_a221oi_1 _23346_ (.B2(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .C1(_05675_),
    .B1(net412),
    .A1(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .Y(_05676_),
    .A2(net376));
 sg13g2_o21ai_1 _23347_ (.B1(_05676_),
    .Y(_05677_),
    .A1(_05671_),
    .A2(_05672_));
 sg13g2_nand2_1 _23348_ (.Y(_05678_),
    .A(net869),
    .B(_05677_));
 sg13g2_nand3_1 _23349_ (.B(_09151_),
    .C(_04888_),
    .A(_09150_),
    .Y(_05679_));
 sg13g2_nand4_1 _23350_ (.B(_05670_),
    .C(_05678_),
    .A(_05663_),
    .Y(_05680_),
    .D(_05679_));
 sg13g2_buf_1 _23351_ (.A(\cpu.spi.r_clk_count[2][6] ),
    .X(_05681_));
 sg13g2_nor2_1 _23352_ (.A(_00138_),
    .B(_05107_),
    .Y(_05682_));
 sg13g2_a221oi_1 _23353_ (.B2(\cpu.spi.r_timeout[6] ),
    .C1(_05682_),
    .B1(_05105_),
    .A1(_05681_),
    .Y(_05683_),
    .A2(_04952_));
 sg13g2_o21ai_1 _23354_ (.B1(_05683_),
    .Y(_05684_),
    .A1(_00137_),
    .A2(_04949_));
 sg13g2_a21oi_1 _23355_ (.A1(_09223_),
    .A2(_04943_),
    .Y(_05685_),
    .B1(_05684_));
 sg13g2_nor2_1 _23356_ (.A(_05369_),
    .B(_05685_),
    .Y(_05686_));
 sg13g2_a221oi_1 _23357_ (.B2(_04896_),
    .C1(_05686_),
    .B1(_05680_),
    .A1(_05074_),
    .Y(_05687_),
    .A2(_05661_));
 sg13g2_a221oi_1 _23358_ (.B2(\cpu.uart.r_in[6] ),
    .C1(net516),
    .B1(_04964_),
    .A1(\cpu.uart.r_div_value[6] ),
    .Y(_05688_),
    .A2(net375));
 sg13g2_a21oi_1 _23359_ (.A1(net516),
    .A2(_05687_),
    .Y(_05689_),
    .B1(_05688_));
 sg13g2_inv_1 _23360_ (.Y(_05690_),
    .A(_00134_));
 sg13g2_a22oi_1 _23361_ (.Y(_05691_),
    .B1(net545),
    .B2(\cpu.dcache.r_data[5][22] ),
    .A2(net638),
    .A1(_05690_));
 sg13g2_a22oi_1 _23362_ (.Y(_05692_),
    .B1(net548),
    .B2(\cpu.dcache.r_data[1][22] ),
    .A2(net479),
    .A1(\cpu.dcache.r_data[6][22] ));
 sg13g2_a22oi_1 _23363_ (.Y(_05693_),
    .B1(net482),
    .B2(\cpu.dcache.r_data[2][22] ),
    .A2(net567),
    .A1(\cpu.dcache.r_data[4][22] ));
 sg13g2_a22oi_1 _23364_ (.Y(_05694_),
    .B1(net543),
    .B2(\cpu.dcache.r_data[7][22] ),
    .A2(net481),
    .A1(\cpu.dcache.r_data[3][22] ));
 sg13g2_nand4_1 _23365_ (.B(_05692_),
    .C(_05693_),
    .A(_05691_),
    .Y(_05695_),
    .D(_05694_));
 sg13g2_mux2_1 _23366_ (.A0(\cpu.dcache.r_data[5][6] ),
    .A1(\cpu.dcache.r_data[7][6] ),
    .S(net569),
    .X(_05696_));
 sg13g2_a22oi_1 _23367_ (.Y(_05697_),
    .B1(_05696_),
    .B2(_12563_),
    .A2(_09592_),
    .A1(\cpu.dcache.r_data[4][6] ));
 sg13g2_nand2b_1 _23368_ (.Y(_05698_),
    .B(net925),
    .A_N(_05697_));
 sg13g2_mux2_1 _23369_ (.A0(\cpu.dcache.r_data[1][6] ),
    .A1(\cpu.dcache.r_data[3][6] ),
    .S(net569),
    .X(_05699_));
 sg13g2_a22oi_1 _23370_ (.Y(_05700_),
    .B1(_05699_),
    .B2(net716),
    .A2(net666),
    .A1(\cpu.dcache.r_data[2][6] ));
 sg13g2_nand2b_1 _23371_ (.Y(_05701_),
    .B(net1065),
    .A_N(_05700_));
 sg13g2_inv_1 _23372_ (.Y(_05702_),
    .A(_00133_));
 sg13g2_a22oi_1 _23373_ (.Y(_05703_),
    .B1(net421),
    .B2(\cpu.dcache.r_data[6][6] ),
    .A2(net514),
    .A1(_05702_));
 sg13g2_nand3_1 _23374_ (.B(_05701_),
    .C(_05703_),
    .A(_05698_),
    .Y(_05704_));
 sg13g2_mux2_1 _23375_ (.A0(_05695_),
    .A1(_05704_),
    .S(_09890_),
    .X(_05705_));
 sg13g2_nand2b_1 _23376_ (.Y(_05706_),
    .B(_05261_),
    .A_N(_04986_));
 sg13g2_nand3_1 _23377_ (.B(net665),
    .C(_05695_),
    .A(_12224_),
    .Y(_05707_));
 sg13g2_a21oi_1 _23378_ (.A1(_05706_),
    .A2(_05707_),
    .Y(_05708_),
    .B1(net1030));
 sg13g2_a221oi_1 _23379_ (.B2(_05005_),
    .C1(_05708_),
    .B1(_05704_),
    .A1(_05003_),
    .Y(_05709_),
    .A2(_05269_));
 sg13g2_nand2_1 _23380_ (.Y(_05710_),
    .A(_05027_),
    .B(_05709_));
 sg13g2_o21ai_1 _23381_ (.B1(_05710_),
    .Y(_05711_),
    .A1(_05027_),
    .A2(_05705_));
 sg13g2_nor2_1 _23382_ (.A(net1166),
    .B(_05711_),
    .Y(_05712_));
 sg13g2_a21oi_1 _23383_ (.A1(net1001),
    .A2(_05689_),
    .Y(_05713_),
    .B1(_05712_));
 sg13g2_nor2_1 _23384_ (.A(net68),
    .B(_05713_),
    .Y(_05714_));
 sg13g2_a21oi_1 _23385_ (.A1(net1000),
    .A2(net69),
    .Y(_05715_),
    .B1(_05714_));
 sg13g2_nor2_1 _23386_ (.A(net132),
    .B(_05715_),
    .Y(_05716_));
 sg13g2_a21o_1 _23387_ (.A2(_05652_),
    .A1(_05650_),
    .B1(_05716_),
    .X(_01031_));
 sg13g2_nand2_1 _23388_ (.Y(_05717_),
    .A(net664),
    .B(_04641_));
 sg13g2_o21ai_1 _23389_ (.B1(_05717_),
    .Y(_05718_),
    .A1(net599),
    .A2(_04638_));
 sg13g2_nor2_1 _23390_ (.A(net291),
    .B(_05718_),
    .Y(_05719_));
 sg13g2_o21ai_1 _23391_ (.B1(net132),
    .Y(_05720_),
    .A1(net986),
    .A2(net211));
 sg13g2_mux2_1 _23392_ (.A0(_05114_),
    .A1(net1154),
    .S(_05025_),
    .X(_05721_));
 sg13g2_nand2_1 _23393_ (.Y(_05722_),
    .A(_05219_),
    .B(_05721_));
 sg13g2_o21ai_1 _23394_ (.B1(_05722_),
    .Y(_01032_),
    .A1(_05719_),
    .A2(_05720_));
 sg13g2_nor3_1 _23395_ (.A(net347),
    .B(net600),
    .C(_04674_),
    .Y(_05723_));
 sg13g2_a21o_1 _23396_ (.A2(net291),
    .A1(net990),
    .B1(_05723_),
    .X(_05724_));
 sg13g2_buf_1 _23397_ (.A(net132),
    .X(_05725_));
 sg13g2_a22oi_1 _23398_ (.Y(_05726_),
    .B1(_05146_),
    .B2(\cpu.intr.r_clock_cmp[8] ),
    .A2(_05139_),
    .A1(\cpu.intr.r_timer_reload[8] ));
 sg13g2_buf_2 _23399_ (.A(\cpu.intr.r_clock_count[24] ),
    .X(_05727_));
 sg13g2_a22oi_1 _23400_ (.Y(_05728_),
    .B1(_05141_),
    .B2(_05727_),
    .A2(_05138_),
    .A1(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_a22oi_1 _23401_ (.Y(_05729_),
    .B1(_05144_),
    .B2(_10076_),
    .A2(_04929_),
    .A1(\cpu.intr.r_timer_count[8] ));
 sg13g2_nand3_1 _23402_ (.B(_05728_),
    .C(_05729_),
    .A(_05726_),
    .Y(_05730_));
 sg13g2_mux2_1 _23403_ (.A0(_05002_),
    .A1(_04994_),
    .S(net566),
    .X(_05731_));
 sg13g2_a22oi_1 _23404_ (.Y(_05732_),
    .B1(_05731_),
    .B2(_05117_),
    .A2(_05730_),
    .A1(_05137_));
 sg13g2_o21ai_1 _23405_ (.B1(_05185_),
    .Y(_05733_),
    .A1(_03141_),
    .A2(_05732_));
 sg13g2_nand2_1 _23406_ (.Y(_05734_),
    .A(net888),
    .B(_05246_));
 sg13g2_o21ai_1 _23407_ (.B1(_05734_),
    .Y(_05735_),
    .A1(_05246_),
    .A2(_05733_));
 sg13g2_a221oi_1 _23408_ (.B2(net99),
    .C1(_05735_),
    .B1(_05724_),
    .A1(_04672_),
    .Y(_01033_),
    .A2(_04836_));
 sg13g2_nor2_1 _23409_ (.A(net985),
    .B(net211),
    .Y(_05736_));
 sg13g2_and2_1 _23410_ (.A(net600),
    .B(_04711_),
    .X(_05737_));
 sg13g2_a22oi_1 _23411_ (.Y(_05738_),
    .B1(_05737_),
    .B2(_04676_),
    .A2(_04714_),
    .A1(net599));
 sg13g2_a22oi_1 _23412_ (.Y(_05739_),
    .B1(net601),
    .B2(\cpu.intr.r_clock_cmp[9] ),
    .A2(_05139_),
    .A1(\cpu.intr.r_timer_reload[9] ));
 sg13g2_buf_2 _23413_ (.A(\cpu.intr.r_clock_count[25] ),
    .X(_05740_));
 sg13g2_a22oi_1 _23414_ (.Y(_05741_),
    .B1(_05141_),
    .B2(_05740_),
    .A2(net602),
    .A1(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_a22oi_1 _23415_ (.Y(_05742_),
    .B1(_05144_),
    .B2(_10083_),
    .A2(_04929_),
    .A1(\cpu.intr.r_timer_count[9] ));
 sg13g2_nand3_1 _23416_ (.B(_05741_),
    .C(_05742_),
    .A(_05739_),
    .Y(_05743_));
 sg13g2_mux2_1 _23417_ (.A0(_05321_),
    .A1(_05327_),
    .S(net566),
    .X(_05744_));
 sg13g2_a22oi_1 _23418_ (.Y(_05745_),
    .B1(_05744_),
    .B2(_05117_),
    .A2(_05743_),
    .A1(_05137_));
 sg13g2_o21ai_1 _23419_ (.B1(_05185_),
    .Y(_05746_),
    .A1(_03141_),
    .A2(_05745_));
 sg13g2_nand2_1 _23420_ (.Y(_05747_),
    .A(_03065_),
    .B(_05246_));
 sg13g2_o21ai_1 _23421_ (.B1(_05747_),
    .Y(_05748_),
    .A1(_05246_),
    .A2(_05746_));
 sg13g2_a221oi_1 _23422_ (.B2(_05156_),
    .C1(_05748_),
    .B1(_05738_),
    .A1(net99),
    .Y(_01034_),
    .A2(_05736_));
 sg13g2_nand2b_1 _23423_ (.Y(_05749_),
    .B(\cpu.dec.r_rd[0] ),
    .A_N(_03558_));
 sg13g2_a21oi_1 _23424_ (.A1(net211),
    .A2(_05749_),
    .Y(_05750_),
    .B1(net164));
 sg13g2_a21o_1 _23425_ (.A2(_05023_),
    .A1(_10633_),
    .B1(_05750_),
    .X(_01035_));
 sg13g2_nor2b_1 _23426_ (.A(_03558_),
    .B_N(\cpu.dec.r_rd[1] ),
    .Y(_05751_));
 sg13g2_o21ai_1 _23427_ (.B1(_05454_),
    .Y(_05752_),
    .A1(_05155_),
    .A2(_05751_));
 sg13g2_o21ai_1 _23428_ (.B1(_05752_),
    .Y(_01036_),
    .A1(_03637_),
    .A2(_05448_));
 sg13g2_nor3_1 _23429_ (.A(_03558_),
    .B(net815),
    .C(_11014_),
    .Y(_05753_));
 sg13g2_nand3_1 _23430_ (.B(net129),
    .C(_05753_),
    .A(\cpu.dec.r_rd[2] ),
    .Y(_05754_));
 sg13g2_o21ai_1 _23431_ (.B1(_05754_),
    .Y(_01037_),
    .A1(_11430_),
    .A2(_05448_));
 sg13g2_inv_1 _23432_ (.Y(_05755_),
    .A(_10147_));
 sg13g2_nand3_1 _23433_ (.B(_04838_),
    .C(_05753_),
    .A(\cpu.dec.r_rd[3] ),
    .Y(_05756_));
 sg13g2_o21ai_1 _23434_ (.B1(_05756_),
    .Y(_01038_),
    .A1(_05755_),
    .A2(net100));
 sg13g2_mux2_1 _23435_ (.A0(\cpu.dec.r_swapsp ),
    .A1(\cpu.ex.r_wb_swapsp ),
    .S(_05219_),
    .X(_01039_));
 sg13g2_nand2_1 _23436_ (.Y(_05757_),
    .A(_11184_),
    .B(net129));
 sg13g2_o21ai_1 _23437_ (.B1(_05757_),
    .Y(_01040_),
    .A1(_12703_),
    .A2(net100));
 sg13g2_a22oi_1 _23438_ (.Y(_05758_),
    .B1(net440),
    .B2(_10226_),
    .A2(net490),
    .A1(net1143));
 sg13g2_nand2_1 _23439_ (.Y(_05759_),
    .A(net748),
    .B(_10550_));
 sg13g2_o21ai_1 _23440_ (.B1(_05759_),
    .Y(_05760_),
    .A1(net748),
    .A2(_05758_));
 sg13g2_mux2_1 _23441_ (.A0(_10091_),
    .A1(_05760_),
    .S(_05725_),
    .X(_01041_));
 sg13g2_inv_1 _23442_ (.Y(_05761_),
    .A(_10098_));
 sg13g2_a22oi_1 _23443_ (.Y(_05762_),
    .B1(net440),
    .B2(_10351_),
    .A2(net490),
    .A1(net1135));
 sg13g2_nand2_1 _23444_ (.Y(_05763_),
    .A(net877),
    .B(_11220_));
 sg13g2_o21ai_1 _23445_ (.B1(_05763_),
    .Y(_05764_),
    .A1(net748),
    .A2(_05762_));
 sg13g2_nand2_1 _23446_ (.Y(_05765_),
    .A(net99),
    .B(_05764_));
 sg13g2_o21ai_1 _23447_ (.B1(_05765_),
    .Y(_01042_),
    .A1(_05761_),
    .A2(net100));
 sg13g2_nand2b_1 _23448_ (.Y(_05766_),
    .B(_08375_),
    .A_N(_11290_));
 sg13g2_a22oi_1 _23449_ (.Y(_05767_),
    .B1(net440),
    .B2(_10476_),
    .A2(net490),
    .A1(_03624_));
 sg13g2_nand2_1 _23450_ (.Y(_05768_),
    .A(net748),
    .B(_05767_));
 sg13g2_nand3_1 _23451_ (.B(_05766_),
    .C(_05768_),
    .A(_05454_),
    .Y(_05769_));
 sg13g2_o21ai_1 _23452_ (.B1(_05769_),
    .Y(_01043_),
    .A1(_12192_),
    .A2(net100));
 sg13g2_nand2_1 _23453_ (.Y(_05770_),
    .A(net877),
    .B(_10506_));
 sg13g2_o21ai_1 _23454_ (.B1(_05770_),
    .Y(_05771_),
    .A1(net748),
    .A2(_11317_));
 sg13g2_nand2_1 _23455_ (.Y(_05772_),
    .A(net129),
    .B(_05771_));
 sg13g2_o21ai_1 _23456_ (.B1(_05772_),
    .Y(_01044_),
    .A1(_12203_),
    .A2(net100));
 sg13g2_a22oi_1 _23457_ (.Y(_05773_),
    .B1(net440),
    .B2(_10431_),
    .A2(net490),
    .A1(_03056_));
 sg13g2_mux2_1 _23458_ (.A0(_11382_),
    .A1(_05773_),
    .S(net748),
    .X(_05774_));
 sg13g2_nand2_1 _23459_ (.Y(_05775_),
    .A(_10114_),
    .B(net130));
 sg13g2_o21ai_1 _23460_ (.B1(_05775_),
    .Y(_01045_),
    .A1(net131),
    .A2(_05774_));
 sg13g2_nand2_1 _23461_ (.Y(_05776_),
    .A(_10378_),
    .B(_10409_));
 sg13g2_nand2_1 _23462_ (.Y(_05777_),
    .A(net748),
    .B(_05776_));
 sg13g2_o21ai_1 _23463_ (.B1(_05777_),
    .Y(_05778_),
    .A1(_03142_),
    .A2(_11356_));
 sg13g2_mux2_1 _23464_ (.A0(_10122_),
    .A1(_05778_),
    .S(net99),
    .X(_01046_));
 sg13g2_nand2_1 _23465_ (.Y(_05779_),
    .A(_10588_),
    .B(net129));
 sg13g2_o21ai_1 _23466_ (.B1(_05779_),
    .Y(_01047_),
    .A1(net759),
    .A2(net100));
 sg13g2_nand2_1 _23467_ (.Y(_05780_),
    .A(_10550_),
    .B(net129));
 sg13g2_o21ai_1 _23468_ (.B1(_05780_),
    .Y(_01048_),
    .A1(net758),
    .A2(net100));
 sg13g2_buf_1 _23469_ (.A(net1144),
    .X(_05781_));
 sg13g2_mux2_1 _23470_ (.A0(_05781_),
    .A1(_11220_),
    .S(net99),
    .X(_01049_));
 sg13g2_nand2_1 _23471_ (.Y(_05782_),
    .A(net1057),
    .B(net130));
 sg13g2_o21ai_1 _23472_ (.B1(_05782_),
    .Y(_01050_),
    .A1(_05767_),
    .A2(net131));
 sg13g2_nand2_1 _23473_ (.Y(_05783_),
    .A(_10506_),
    .B(net129));
 sg13g2_o21ai_1 _23474_ (.B1(_05783_),
    .Y(_01051_),
    .A1(net892),
    .A2(net99));
 sg13g2_nand2_1 _23475_ (.Y(_05784_),
    .A(net1053),
    .B(net130));
 sg13g2_o21ai_1 _23476_ (.B1(_05784_),
    .Y(_01052_),
    .A1(_05773_),
    .A2(net131));
 sg13g2_nand2_1 _23477_ (.Y(_05785_),
    .A(_05776_),
    .B(net129));
 sg13g2_o21ai_1 _23478_ (.B1(_05785_),
    .Y(_01053_),
    .A1(_02749_),
    .A2(net99));
 sg13g2_nand2_1 _23479_ (.Y(_05786_),
    .A(net877),
    .B(_11184_));
 sg13g2_o21ai_1 _23480_ (.B1(_05786_),
    .Y(_05787_),
    .A1(net748),
    .A2(_10361_));
 sg13g2_mux2_1 _23481_ (.A0(_10081_),
    .A1(_05787_),
    .S(net99),
    .X(_01054_));
 sg13g2_nand2_1 _23482_ (.Y(_05788_),
    .A(_10236_),
    .B(_10274_));
 sg13g2_mux2_1 _23483_ (.A0(_10588_),
    .A1(_05788_),
    .S(_08375_),
    .X(_05789_));
 sg13g2_mux2_1 _23484_ (.A0(_10086_),
    .A1(_05789_),
    .S(_05725_),
    .X(_01055_));
 sg13g2_mux2_1 _23485_ (.A0(_08494_),
    .A1(net627),
    .S(_08351_),
    .X(_05790_));
 sg13g2_or3_1 _23486_ (.A(_11168_),
    .B(_10551_),
    .C(_11221_),
    .X(_05791_));
 sg13g2_o21ai_1 _23487_ (.B1(_03447_),
    .Y(_05792_),
    .A1(_10589_),
    .A2(_05791_));
 sg13g2_buf_2 _23488_ (.A(_05792_),
    .X(_05793_));
 sg13g2_nor4_2 _23489_ (.A(_08265_),
    .B(_04754_),
    .C(_11450_),
    .Y(_05794_),
    .D(_03638_));
 sg13g2_and2_1 _23490_ (.A(_05793_),
    .B(_05794_),
    .X(_05795_));
 sg13g2_buf_1 _23491_ (.A(_05795_),
    .X(_05796_));
 sg13g2_buf_1 _23492_ (.A(_00281_),
    .X(_05797_));
 sg13g2_nand2b_1 _23493_ (.Y(_05798_),
    .B(net1162),
    .A_N(_05797_));
 sg13g2_o21ai_1 _23494_ (.B1(_05798_),
    .Y(_05799_),
    .A1(net992),
    .A2(net627));
 sg13g2_nand3_1 _23495_ (.B(_05796_),
    .C(_05799_),
    .A(net350),
    .Y(_05800_));
 sg13g2_o21ai_1 _23496_ (.B1(_05800_),
    .Y(_05801_),
    .A1(net292),
    .A2(_05790_));
 sg13g2_o21ai_1 _23497_ (.B1(net933),
    .Y(_05802_),
    .A1(_08419_),
    .A2(_05796_));
 sg13g2_buf_1 _23498_ (.A(_05802_),
    .X(_05803_));
 sg13g2_a22oi_1 _23499_ (.Y(_01058_),
    .B1(_05803_),
    .B2(_11268_),
    .A2(_05801_),
    .A1(net717));
 sg13g2_mux2_1 _23500_ (.A0(_08423_),
    .A1(_10807_),
    .S(_08351_),
    .X(_05804_));
 sg13g2_nor2_1 _23501_ (.A(_11268_),
    .B(_10799_),
    .Y(_05805_));
 sg13g2_buf_2 _23502_ (.A(_05805_),
    .X(_05806_));
 sg13g2_buf_1 _23503_ (.A(_10831_),
    .X(_05807_));
 sg13g2_nor2_2 _23504_ (.A(_05807_),
    .B(net1124),
    .Y(_05808_));
 sg13g2_o21ai_1 _23505_ (.B1(net992),
    .Y(_05809_),
    .A1(_05806_),
    .A2(_05808_));
 sg13g2_o21ai_1 _23506_ (.B1(_05809_),
    .Y(_05810_),
    .A1(net992),
    .A2(_10807_));
 sg13g2_nand3_1 _23507_ (.B(_05796_),
    .C(_05810_),
    .A(net292),
    .Y(_05811_));
 sg13g2_o21ai_1 _23508_ (.B1(_05811_),
    .Y(_05812_),
    .A1(net292),
    .A2(_05804_));
 sg13g2_buf_2 _23509_ (.A(net818),
    .X(_05813_));
 sg13g2_a22oi_1 _23510_ (.Y(_01059_),
    .B1(_05812_),
    .B2(net663),
    .A2(_05803_),
    .A1(_10799_));
 sg13g2_inv_1 _23511_ (.Y(_05814_),
    .A(net1123));
 sg13g2_buf_1 _23512_ (.A(_05814_),
    .X(_05815_));
 sg13g2_mux2_1 _23513_ (.A0(_08636_),
    .A1(net698),
    .S(_08351_),
    .X(_05816_));
 sg13g2_nand2_1 _23514_ (.Y(_05817_),
    .A(_10831_),
    .B(net1124));
 sg13g2_buf_1 _23515_ (.A(_05817_),
    .X(_05818_));
 sg13g2_nor2_2 _23516_ (.A(net868),
    .B(net867),
    .Y(_05819_));
 sg13g2_buf_1 _23517_ (.A(net1123),
    .X(_05820_));
 sg13g2_nor2_1 _23518_ (.A(net979),
    .B(_05806_),
    .Y(_05821_));
 sg13g2_o21ai_1 _23519_ (.B1(net992),
    .Y(_05822_),
    .A1(_05819_),
    .A2(_05821_));
 sg13g2_o21ai_1 _23520_ (.B1(_05822_),
    .Y(_05823_),
    .A1(net992),
    .A2(net698));
 sg13g2_nand3_1 _23521_ (.B(_05796_),
    .C(_05823_),
    .A(_09745_),
    .Y(_05824_));
 sg13g2_o21ai_1 _23522_ (.B1(_05824_),
    .Y(_05825_),
    .A1(_04476_),
    .A2(_05816_));
 sg13g2_a22oi_1 _23523_ (.Y(_01060_),
    .B1(_05825_),
    .B2(_05813_),
    .A2(_05803_),
    .A1(net868));
 sg13g2_mux2_1 _23524_ (.A0(net937),
    .A1(net687),
    .S(_08351_),
    .X(_05826_));
 sg13g2_xnor2_1 _23525_ (.Y(_05827_),
    .A(net1125),
    .B(_05819_));
 sg13g2_nand2_1 _23526_ (.Y(_05828_),
    .A(_03602_),
    .B(_05827_));
 sg13g2_o21ai_1 _23527_ (.B1(_05828_),
    .Y(_05829_),
    .A1(_03602_),
    .A2(net687));
 sg13g2_nand3_1 _23528_ (.B(_05796_),
    .C(_05829_),
    .A(_09745_),
    .Y(_05830_));
 sg13g2_o21ai_1 _23529_ (.B1(_05830_),
    .Y(_05831_),
    .A1(_04476_),
    .A2(_05826_));
 sg13g2_a22oi_1 _23530_ (.Y(_01061_),
    .B1(_05831_),
    .B2(_05813_),
    .A2(_05803_),
    .A1(net1035));
 sg13g2_buf_2 _23531_ (.A(_00186_),
    .X(_05832_));
 sg13g2_buf_1 _23532_ (.A(_10533_),
    .X(_05833_));
 sg13g2_nor2_1 _23533_ (.A(net978),
    .B(net1125),
    .Y(_05834_));
 sg13g2_buf_2 _23534_ (.A(_05834_),
    .X(_05835_));
 sg13g2_nand2_1 _23535_ (.Y(_05836_),
    .A(_05832_),
    .B(_05835_));
 sg13g2_nand4_1 _23536_ (.B(_11058_),
    .C(_05794_),
    .A(net1162),
    .Y(_05837_),
    .D(_05808_));
 sg13g2_buf_1 _23537_ (.A(_05837_),
    .X(_05838_));
 sg13g2_nor2_1 _23538_ (.A(_05836_),
    .B(_05838_),
    .Y(_05839_));
 sg13g2_buf_1 _23539_ (.A(_05839_),
    .X(_05840_));
 sg13g2_buf_1 _23540_ (.A(_05840_),
    .X(_05841_));
 sg13g2_mux2_1 _23541_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][0] ),
    .A1(_03625_),
    .S(net373),
    .X(_01129_));
 sg13g2_mux2_1 _23542_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][10] ),
    .A1(net605),
    .S(net373),
    .X(_01130_));
 sg13g2_mux2_1 _23543_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][11] ),
    .A1(net527),
    .S(net373),
    .X(_01131_));
 sg13g2_mux2_1 _23544_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][1] ),
    .A1(net467),
    .S(net373),
    .X(_01132_));
 sg13g2_mux2_1 _23545_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][2] ),
    .A1(_03102_),
    .S(net373),
    .X(_01133_));
 sg13g2_mux2_1 _23546_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][3] ),
    .A1(net873),
    .S(net373),
    .X(_01134_));
 sg13g2_mux2_1 _23547_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][4] ),
    .A1(net875),
    .S(net373),
    .X(_01135_));
 sg13g2_mux2_1 _23548_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][5] ),
    .A1(net874),
    .S(_05841_),
    .X(_01136_));
 sg13g2_mux2_1 _23549_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][6] ),
    .A1(net983),
    .S(net373),
    .X(_01137_));
 sg13g2_mux2_1 _23550_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][7] ),
    .A1(net870),
    .S(_05841_),
    .X(_01138_));
 sg13g2_mux2_1 _23551_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][8] ),
    .A1(_03664_),
    .S(_05840_),
    .X(_01139_));
 sg13g2_mux2_1 _23552_ (.A0(\cpu.genblk1.mmu.r_vtop_d[0][9] ),
    .A1(net466),
    .S(_05840_),
    .X(_01140_));
 sg13g2_buf_1 _23553_ (.A(net616),
    .X(_05842_));
 sg13g2_nand3_1 _23554_ (.B(_11058_),
    .C(_05794_),
    .A(_08376_),
    .Y(_05843_));
 sg13g2_buf_1 _23555_ (.A(_05843_),
    .X(_05844_));
 sg13g2_buf_1 _23556_ (.A(_05844_),
    .X(_05845_));
 sg13g2_nand2_1 _23557_ (.Y(_05846_),
    .A(_11268_),
    .B(net1124));
 sg13g2_buf_1 _23558_ (.A(_05846_),
    .X(_05847_));
 sg13g2_inv_1 _23559_ (.Y(_05848_),
    .A(net978));
 sg13g2_nand2_1 _23560_ (.Y(_05849_),
    .A(_05848_),
    .B(net1125));
 sg13g2_buf_2 _23561_ (.A(_05849_),
    .X(_05850_));
 sg13g2_nor3_2 _23562_ (.A(_05820_),
    .B(_05847_),
    .C(_05850_),
    .Y(_05851_));
 sg13g2_nor2b_1 _23563_ (.A(net462),
    .B_N(_05851_),
    .Y(_05852_));
 sg13g2_buf_1 _23564_ (.A(_05852_),
    .X(_05853_));
 sg13g2_buf_1 _23565_ (.A(_05853_),
    .X(_05854_));
 sg13g2_mux2_1 _23566_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][0] ),
    .A1(net513),
    .S(net339),
    .X(_01141_));
 sg13g2_mux2_1 _23567_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][10] ),
    .A1(net605),
    .S(net339),
    .X(_01142_));
 sg13g2_mux2_1 _23568_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][11] ),
    .A1(net527),
    .S(net339),
    .X(_01143_));
 sg13g2_mux2_1 _23569_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][1] ),
    .A1(net467),
    .S(net339),
    .X(_01144_));
 sg13g2_buf_1 _23570_ (.A(net1000),
    .X(_05855_));
 sg13g2_mux2_1 _23571_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][2] ),
    .A1(net866),
    .S(net339),
    .X(_01145_));
 sg13g2_mux2_1 _23572_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][3] ),
    .A1(net873),
    .S(net339),
    .X(_01146_));
 sg13g2_mux2_1 _23573_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][4] ),
    .A1(net875),
    .S(net339),
    .X(_01147_));
 sg13g2_mux2_1 _23574_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][5] ),
    .A1(net874),
    .S(_05854_),
    .X(_01148_));
 sg13g2_mux2_1 _23575_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][6] ),
    .A1(net983),
    .S(net339),
    .X(_01149_));
 sg13g2_mux2_1 _23576_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][7] ),
    .A1(net870),
    .S(_05854_),
    .X(_01150_));
 sg13g2_mux2_1 _23577_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][8] ),
    .A1(net525),
    .S(_05853_),
    .X(_01151_));
 sg13g2_mux2_1 _23578_ (.A0(\cpu.genblk1.mmu.r_vtop_d[10][9] ),
    .A1(net466),
    .S(_05853_),
    .X(_01152_));
 sg13g2_nor3_1 _23579_ (.A(net1123),
    .B(net867),
    .C(_05850_),
    .Y(_05856_));
 sg13g2_buf_2 _23580_ (.A(_05856_),
    .X(_05857_));
 sg13g2_nor2b_1 _23581_ (.A(net462),
    .B_N(_05857_),
    .Y(_05858_));
 sg13g2_buf_1 _23582_ (.A(_05858_),
    .X(_05859_));
 sg13g2_buf_1 _23583_ (.A(_05859_),
    .X(_05860_));
 sg13g2_mux2_1 _23584_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][0] ),
    .A1(net513),
    .S(net338),
    .X(_01153_));
 sg13g2_mux2_1 _23585_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][10] ),
    .A1(_04760_),
    .S(net338),
    .X(_01154_));
 sg13g2_mux2_1 _23586_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][11] ),
    .A1(net527),
    .S(net338),
    .X(_01155_));
 sg13g2_mux2_1 _23587_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][1] ),
    .A1(net467),
    .S(net338),
    .X(_01156_));
 sg13g2_mux2_1 _23588_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][2] ),
    .A1(net866),
    .S(net338),
    .X(_01157_));
 sg13g2_mux2_1 _23589_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][3] ),
    .A1(net873),
    .S(net338),
    .X(_01158_));
 sg13g2_mux2_1 _23590_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][4] ),
    .A1(net875),
    .S(net338),
    .X(_01159_));
 sg13g2_mux2_1 _23591_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][5] ),
    .A1(net874),
    .S(_05860_),
    .X(_01160_));
 sg13g2_mux2_1 _23592_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][6] ),
    .A1(_04765_),
    .S(net338),
    .X(_01161_));
 sg13g2_mux2_1 _23593_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][7] ),
    .A1(net870),
    .S(_05860_),
    .X(_01162_));
 sg13g2_mux2_1 _23594_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][8] ),
    .A1(net525),
    .S(_05859_),
    .X(_01163_));
 sg13g2_mux2_1 _23595_ (.A0(\cpu.genblk1.mmu.r_vtop_d[11][9] ),
    .A1(net466),
    .S(_05859_),
    .X(_01164_));
 sg13g2_nor2_2 _23596_ (.A(net978),
    .B(net1035),
    .Y(_05861_));
 sg13g2_nand2b_1 _23597_ (.Y(_05862_),
    .B(_05861_),
    .A_N(_05832_));
 sg13g2_buf_1 _23598_ (.A(_05862_),
    .X(_05863_));
 sg13g2_nor2_1 _23599_ (.A(_05838_),
    .B(_05863_),
    .Y(_05864_));
 sg13g2_buf_1 _23600_ (.A(_05864_),
    .X(_05865_));
 sg13g2_buf_1 _23601_ (.A(_05865_),
    .X(_05866_));
 sg13g2_mux2_1 _23602_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][0] ),
    .A1(net513),
    .S(net372),
    .X(_01165_));
 sg13g2_mux2_1 _23603_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][10] ),
    .A1(net605),
    .S(net372),
    .X(_01166_));
 sg13g2_mux2_1 _23604_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][11] ),
    .A1(net527),
    .S(net372),
    .X(_01167_));
 sg13g2_mux2_1 _23605_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][1] ),
    .A1(net467),
    .S(net372),
    .X(_01168_));
 sg13g2_mux2_1 _23606_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][2] ),
    .A1(net866),
    .S(net372),
    .X(_01169_));
 sg13g2_mux2_1 _23607_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][3] ),
    .A1(net873),
    .S(_05866_),
    .X(_01170_));
 sg13g2_mux2_1 _23608_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][4] ),
    .A1(_03647_),
    .S(_05866_),
    .X(_01171_));
 sg13g2_mux2_1 _23609_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][5] ),
    .A1(_03648_),
    .S(net372),
    .X(_01172_));
 sg13g2_mux2_1 _23610_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][6] ),
    .A1(net983),
    .S(net372),
    .X(_01173_));
 sg13g2_mux2_1 _23611_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][7] ),
    .A1(net870),
    .S(net372),
    .X(_01174_));
 sg13g2_mux2_1 _23612_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][8] ),
    .A1(net525),
    .S(_05865_),
    .X(_01175_));
 sg13g2_mux2_1 _23613_ (.A0(\cpu.genblk1.mmu.r_vtop_d[12][9] ),
    .A1(net466),
    .S(_05865_),
    .X(_01176_));
 sg13g2_nand2_2 _23614_ (.Y(_05867_),
    .A(net980),
    .B(_10799_));
 sg13g2_or2_1 _23615_ (.X(_05868_),
    .B(_05844_),
    .A(_05867_));
 sg13g2_buf_2 _23616_ (.A(_05868_),
    .X(_05869_));
 sg13g2_nor2_1 _23617_ (.A(_05863_),
    .B(_05869_),
    .Y(_05870_));
 sg13g2_buf_1 _23618_ (.A(_05870_),
    .X(_05871_));
 sg13g2_buf_1 _23619_ (.A(_05871_),
    .X(_05872_));
 sg13g2_mux2_1 _23620_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][0] ),
    .A1(net513),
    .S(net290),
    .X(_01177_));
 sg13g2_mux2_1 _23621_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][10] ),
    .A1(net605),
    .S(net290),
    .X(_01178_));
 sg13g2_mux2_1 _23622_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][11] ),
    .A1(net527),
    .S(net290),
    .X(_01179_));
 sg13g2_mux2_1 _23623_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][1] ),
    .A1(_03643_),
    .S(net290),
    .X(_01180_));
 sg13g2_mux2_1 _23624_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][2] ),
    .A1(net866),
    .S(net290),
    .X(_01181_));
 sg13g2_mux2_1 _23625_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][3] ),
    .A1(net873),
    .S(net290),
    .X(_01182_));
 sg13g2_mux2_1 _23626_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][4] ),
    .A1(_03647_),
    .S(_05872_),
    .X(_01183_));
 sg13g2_mux2_1 _23627_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][5] ),
    .A1(_03648_),
    .S(_05872_),
    .X(_01184_));
 sg13g2_mux2_1 _23628_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][6] ),
    .A1(net983),
    .S(net290),
    .X(_01185_));
 sg13g2_mux2_1 _23629_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][7] ),
    .A1(net870),
    .S(net290),
    .X(_01186_));
 sg13g2_mux2_1 _23630_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][8] ),
    .A1(net525),
    .S(_05871_),
    .X(_01187_));
 sg13g2_mux2_1 _23631_ (.A0(\cpu.genblk1.mmu.r_vtop_d[13][9] ),
    .A1(net466),
    .S(_05871_),
    .X(_01188_));
 sg13g2_buf_1 _23632_ (.A(_05844_),
    .X(_05873_));
 sg13g2_nor3_1 _23633_ (.A(net746),
    .B(_05873_),
    .C(_05863_),
    .Y(_05874_));
 sg13g2_buf_1 _23634_ (.A(_05874_),
    .X(_05875_));
 sg13g2_buf_1 _23635_ (.A(_05875_),
    .X(_05876_));
 sg13g2_mux2_1 _23636_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][0] ),
    .A1(_05842_),
    .S(net337),
    .X(_01189_));
 sg13g2_mux2_1 _23637_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][10] ),
    .A1(net605),
    .S(net337),
    .X(_01190_));
 sg13g2_mux2_1 _23638_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][11] ),
    .A1(_03658_),
    .S(net337),
    .X(_01191_));
 sg13g2_mux2_1 _23639_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][1] ),
    .A1(_03643_),
    .S(net337),
    .X(_01192_));
 sg13g2_mux2_1 _23640_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][2] ),
    .A1(net866),
    .S(net337),
    .X(_01193_));
 sg13g2_mux2_1 _23641_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][3] ),
    .A1(net873),
    .S(net337),
    .X(_01194_));
 sg13g2_buf_1 _23642_ (.A(net996),
    .X(_05877_));
 sg13g2_mux2_1 _23643_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][4] ),
    .A1(_05877_),
    .S(net337),
    .X(_01195_));
 sg13g2_buf_1 _23644_ (.A(net995),
    .X(_05878_));
 sg13g2_mux2_1 _23645_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][5] ),
    .A1(net864),
    .S(_05876_),
    .X(_01196_));
 sg13g2_mux2_1 _23646_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][6] ),
    .A1(net983),
    .S(net337),
    .X(_01197_));
 sg13g2_mux2_1 _23647_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][7] ),
    .A1(net870),
    .S(_05876_),
    .X(_01198_));
 sg13g2_mux2_1 _23648_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][8] ),
    .A1(net525),
    .S(_05875_),
    .X(_01199_));
 sg13g2_mux2_1 _23649_ (.A0(\cpu.genblk1.mmu.r_vtop_d[14][9] ),
    .A1(_03655_),
    .S(_05875_),
    .X(_01200_));
 sg13g2_nor3_1 _23650_ (.A(net867),
    .B(net461),
    .C(_05863_),
    .Y(_05879_));
 sg13g2_buf_1 _23651_ (.A(_05879_),
    .X(_05880_));
 sg13g2_buf_1 _23652_ (.A(_05880_),
    .X(_05881_));
 sg13g2_mux2_1 _23653_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][0] ),
    .A1(_05842_),
    .S(net336),
    .X(_01201_));
 sg13g2_mux2_1 _23654_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][10] ),
    .A1(net605),
    .S(net336),
    .X(_01202_));
 sg13g2_mux2_1 _23655_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][11] ),
    .A1(_03658_),
    .S(net336),
    .X(_01203_));
 sg13g2_buf_1 _23656_ (.A(net530),
    .X(_05882_));
 sg13g2_mux2_1 _23657_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][1] ),
    .A1(_05882_),
    .S(net336),
    .X(_01204_));
 sg13g2_mux2_1 _23658_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][2] ),
    .A1(net866),
    .S(net336),
    .X(_01205_));
 sg13g2_mux2_1 _23659_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][3] ),
    .A1(_03665_),
    .S(net336),
    .X(_01206_));
 sg13g2_mux2_1 _23660_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][4] ),
    .A1(_05877_),
    .S(net336),
    .X(_01207_));
 sg13g2_mux2_1 _23661_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][5] ),
    .A1(net864),
    .S(_05881_),
    .X(_01208_));
 sg13g2_mux2_1 _23662_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][6] ),
    .A1(net983),
    .S(net336),
    .X(_01209_));
 sg13g2_mux2_1 _23663_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][7] ),
    .A1(net870),
    .S(_05881_),
    .X(_01210_));
 sg13g2_mux2_1 _23664_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][8] ),
    .A1(net525),
    .S(_05880_),
    .X(_01211_));
 sg13g2_mux2_1 _23665_ (.A0(\cpu.genblk1.mmu.r_vtop_d[15][9] ),
    .A1(_03655_),
    .S(_05880_),
    .X(_01212_));
 sg13g2_nand2_1 _23666_ (.Y(_05883_),
    .A(net978),
    .B(net1035));
 sg13g2_buf_2 _23667_ (.A(_05883_),
    .X(_05884_));
 sg13g2_nand2_2 _23668_ (.Y(_05885_),
    .A(net868),
    .B(_05808_));
 sg13g2_nor3_1 _23669_ (.A(net461),
    .B(_05884_),
    .C(_05885_),
    .Y(_05886_));
 sg13g2_buf_1 _23670_ (.A(_05886_),
    .X(_05887_));
 sg13g2_buf_1 _23671_ (.A(_05887_),
    .X(_05888_));
 sg13g2_mux2_1 _23672_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][0] ),
    .A1(net513),
    .S(net335),
    .X(_01213_));
 sg13g2_mux2_1 _23673_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][10] ),
    .A1(net605),
    .S(net335),
    .X(_01214_));
 sg13g2_buf_1 _23674_ (.A(_10730_),
    .X(_05889_));
 sg13g2_mux2_1 _23675_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][11] ),
    .A1(net597),
    .S(net335),
    .X(_01215_));
 sg13g2_mux2_1 _23676_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][1] ),
    .A1(net460),
    .S(_05888_),
    .X(_01216_));
 sg13g2_mux2_1 _23677_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][2] ),
    .A1(net866),
    .S(net335),
    .X(_01217_));
 sg13g2_mux2_1 _23678_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][3] ),
    .A1(_03665_),
    .S(net335),
    .X(_01218_));
 sg13g2_mux2_1 _23679_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][4] ),
    .A1(net865),
    .S(_05888_),
    .X(_01219_));
 sg13g2_mux2_1 _23680_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][5] ),
    .A1(net864),
    .S(net335),
    .X(_01220_));
 sg13g2_mux2_1 _23681_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][6] ),
    .A1(net983),
    .S(net335),
    .X(_01221_));
 sg13g2_mux2_1 _23682_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][7] ),
    .A1(net870),
    .S(net335),
    .X(_01222_));
 sg13g2_mux2_1 _23683_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][8] ),
    .A1(net525),
    .S(_05887_),
    .X(_01223_));
 sg13g2_buf_1 _23684_ (.A(net628),
    .X(_05890_));
 sg13g2_mux2_1 _23685_ (.A0(\cpu.genblk1.mmu.r_vtop_d[16][9] ),
    .A1(net512),
    .S(_05887_),
    .X(_01224_));
 sg13g2_nor3_1 _23686_ (.A(net979),
    .B(_05869_),
    .C(_05884_),
    .Y(_05891_));
 sg13g2_buf_1 _23687_ (.A(_05891_),
    .X(_05892_));
 sg13g2_buf_1 _23688_ (.A(_05892_),
    .X(_05893_));
 sg13g2_mux2_1 _23689_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][0] ),
    .A1(net513),
    .S(net289),
    .X(_01225_));
 sg13g2_mux2_1 _23690_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][10] ),
    .A1(net605),
    .S(net289),
    .X(_01226_));
 sg13g2_mux2_1 _23691_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][11] ),
    .A1(net597),
    .S(net289),
    .X(_01227_));
 sg13g2_mux2_1 _23692_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][1] ),
    .A1(net460),
    .S(_05893_),
    .X(_01228_));
 sg13g2_mux2_1 _23693_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][2] ),
    .A1(net866),
    .S(net289),
    .X(_01229_));
 sg13g2_buf_1 _23694_ (.A(net997),
    .X(_05894_));
 sg13g2_mux2_1 _23695_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][3] ),
    .A1(net863),
    .S(net289),
    .X(_01230_));
 sg13g2_mux2_1 _23696_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][4] ),
    .A1(net865),
    .S(_05893_),
    .X(_01231_));
 sg13g2_mux2_1 _23697_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][5] ),
    .A1(net864),
    .S(net289),
    .X(_01232_));
 sg13g2_mux2_1 _23698_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][6] ),
    .A1(net983),
    .S(net289),
    .X(_01233_));
 sg13g2_mux2_1 _23699_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][7] ),
    .A1(_04758_),
    .S(net289),
    .X(_01234_));
 sg13g2_mux2_1 _23700_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][8] ),
    .A1(net525),
    .S(_05892_),
    .X(_01235_));
 sg13g2_mux2_1 _23701_ (.A0(\cpu.genblk1.mmu.r_vtop_d[17][9] ),
    .A1(net512),
    .S(_05892_),
    .X(_01236_));
 sg13g2_nor2_1 _23702_ (.A(_05848_),
    .B(net980),
    .Y(_05895_));
 sg13g2_nand3_1 _23703_ (.B(net868),
    .C(_05895_),
    .A(net1124),
    .Y(_05896_));
 sg13g2_nor2_2 _23704_ (.A(net1125),
    .B(_05896_),
    .Y(_05897_));
 sg13g2_nor2b_1 _23705_ (.A(net462),
    .B_N(_05897_),
    .Y(_05898_));
 sg13g2_buf_1 _23706_ (.A(_05898_),
    .X(_05899_));
 sg13g2_buf_1 _23707_ (.A(_05899_),
    .X(_05900_));
 sg13g2_mux2_1 _23708_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][0] ),
    .A1(net513),
    .S(net334),
    .X(_01237_));
 sg13g2_buf_1 _23709_ (.A(_09523_),
    .X(_05901_));
 sg13g2_mux2_1 _23710_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][10] ),
    .A1(net596),
    .S(net334),
    .X(_01238_));
 sg13g2_mux2_1 _23711_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][11] ),
    .A1(_05889_),
    .S(net334),
    .X(_01239_));
 sg13g2_mux2_1 _23712_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][1] ),
    .A1(net460),
    .S(_05900_),
    .X(_01240_));
 sg13g2_mux2_1 _23713_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][2] ),
    .A1(_05855_),
    .S(net334),
    .X(_01241_));
 sg13g2_mux2_1 _23714_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][3] ),
    .A1(_05894_),
    .S(net334),
    .X(_01242_));
 sg13g2_mux2_1 _23715_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][4] ),
    .A1(net865),
    .S(net334),
    .X(_01243_));
 sg13g2_mux2_1 _23716_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][5] ),
    .A1(_05878_),
    .S(_05900_),
    .X(_01244_));
 sg13g2_buf_1 _23717_ (.A(net1143),
    .X(_05902_));
 sg13g2_mux2_1 _23718_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][6] ),
    .A1(net977),
    .S(net334),
    .X(_01245_));
 sg13g2_buf_1 _23719_ (.A(net1135),
    .X(_05903_));
 sg13g2_mux2_1 _23720_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][7] ),
    .A1(net976),
    .S(net334),
    .X(_01246_));
 sg13g2_buf_1 _23721_ (.A(_10810_),
    .X(_05904_));
 sg13g2_mux2_1 _23722_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][8] ),
    .A1(net511),
    .S(_05899_),
    .X(_01247_));
 sg13g2_mux2_1 _23723_ (.A0(\cpu.genblk1.mmu.r_vtop_d[18][9] ),
    .A1(net512),
    .S(_05899_),
    .X(_01248_));
 sg13g2_nor3_1 _23724_ (.A(_11375_),
    .B(net867),
    .C(_05884_),
    .Y(_05905_));
 sg13g2_buf_2 _23725_ (.A(_05905_),
    .X(_05906_));
 sg13g2_nor2b_1 _23726_ (.A(net462),
    .B_N(_05906_),
    .Y(_05907_));
 sg13g2_buf_1 _23727_ (.A(_05907_),
    .X(_05908_));
 sg13g2_buf_1 _23728_ (.A(_05908_),
    .X(_05909_));
 sg13g2_mux2_1 _23729_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][0] ),
    .A1(net513),
    .S(net333),
    .X(_01249_));
 sg13g2_mux2_1 _23730_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][10] ),
    .A1(net596),
    .S(net333),
    .X(_01250_));
 sg13g2_mux2_1 _23731_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][11] ),
    .A1(net597),
    .S(net333),
    .X(_01251_));
 sg13g2_mux2_1 _23732_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][1] ),
    .A1(net460),
    .S(_05909_),
    .X(_01252_));
 sg13g2_mux2_1 _23733_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][2] ),
    .A1(_05855_),
    .S(net333),
    .X(_01253_));
 sg13g2_mux2_1 _23734_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][3] ),
    .A1(_05894_),
    .S(net333),
    .X(_01254_));
 sg13g2_mux2_1 _23735_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][4] ),
    .A1(net865),
    .S(net333),
    .X(_01255_));
 sg13g2_mux2_1 _23736_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][5] ),
    .A1(net864),
    .S(_05909_),
    .X(_01256_));
 sg13g2_mux2_1 _23737_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][6] ),
    .A1(_05902_),
    .S(net333),
    .X(_01257_));
 sg13g2_mux2_1 _23738_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][7] ),
    .A1(net976),
    .S(net333),
    .X(_01258_));
 sg13g2_mux2_1 _23739_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][8] ),
    .A1(net511),
    .S(_05908_),
    .X(_01259_));
 sg13g2_mux2_1 _23740_ (.A0(\cpu.genblk1.mmu.r_vtop_d[19][9] ),
    .A1(net512),
    .S(_05908_),
    .X(_01260_));
 sg13g2_buf_1 _23741_ (.A(net616),
    .X(_05910_));
 sg13g2_nor2_1 _23742_ (.A(_05836_),
    .B(_05869_),
    .Y(_05911_));
 sg13g2_buf_1 _23743_ (.A(_05911_),
    .X(_05912_));
 sg13g2_buf_1 _23744_ (.A(_05912_),
    .X(_05913_));
 sg13g2_mux2_1 _23745_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][0] ),
    .A1(net510),
    .S(net288),
    .X(_01261_));
 sg13g2_mux2_1 _23746_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][10] ),
    .A1(_05901_),
    .S(net288),
    .X(_01262_));
 sg13g2_mux2_1 _23747_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][11] ),
    .A1(_05889_),
    .S(net288),
    .X(_01263_));
 sg13g2_mux2_1 _23748_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][1] ),
    .A1(_05882_),
    .S(net288),
    .X(_01264_));
 sg13g2_buf_1 _23749_ (.A(_03056_),
    .X(_05914_));
 sg13g2_mux2_1 _23750_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][2] ),
    .A1(net862),
    .S(net288),
    .X(_01265_));
 sg13g2_mux2_1 _23751_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][3] ),
    .A1(net863),
    .S(net288),
    .X(_01266_));
 sg13g2_mux2_1 _23752_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][4] ),
    .A1(net865),
    .S(net288),
    .X(_01267_));
 sg13g2_mux2_1 _23753_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][5] ),
    .A1(_05878_),
    .S(_05913_),
    .X(_01268_));
 sg13g2_mux2_1 _23754_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][6] ),
    .A1(_05902_),
    .S(net288),
    .X(_01269_));
 sg13g2_mux2_1 _23755_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][7] ),
    .A1(net976),
    .S(_05913_),
    .X(_01270_));
 sg13g2_mux2_1 _23756_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][8] ),
    .A1(net511),
    .S(_05912_),
    .X(_01271_));
 sg13g2_mux2_1 _23757_ (.A0(\cpu.genblk1.mmu.r_vtop_d[1][9] ),
    .A1(_05890_),
    .S(_05912_),
    .X(_01272_));
 sg13g2_or2_1 _23758_ (.X(_05915_),
    .B(_05884_),
    .A(_05832_));
 sg13g2_buf_1 _23759_ (.A(_05915_),
    .X(_05916_));
 sg13g2_nor2_1 _23760_ (.A(_05838_),
    .B(_05916_),
    .Y(_05917_));
 sg13g2_buf_1 _23761_ (.A(_05917_),
    .X(_05918_));
 sg13g2_buf_1 _23762_ (.A(_05918_),
    .X(_05919_));
 sg13g2_mux2_1 _23763_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][0] ),
    .A1(net510),
    .S(_05919_),
    .X(_01273_));
 sg13g2_mux2_1 _23764_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][10] ),
    .A1(net596),
    .S(net371),
    .X(_01274_));
 sg13g2_mux2_1 _23765_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][11] ),
    .A1(net597),
    .S(net371),
    .X(_01275_));
 sg13g2_mux2_1 _23766_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][1] ),
    .A1(net460),
    .S(_05919_),
    .X(_01276_));
 sg13g2_mux2_1 _23767_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][2] ),
    .A1(net862),
    .S(net371),
    .X(_01277_));
 sg13g2_mux2_1 _23768_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][3] ),
    .A1(net863),
    .S(net371),
    .X(_01278_));
 sg13g2_mux2_1 _23769_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][4] ),
    .A1(net865),
    .S(net371),
    .X(_01279_));
 sg13g2_mux2_1 _23770_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][5] ),
    .A1(net864),
    .S(net371),
    .X(_01280_));
 sg13g2_mux2_1 _23771_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][6] ),
    .A1(net977),
    .S(net371),
    .X(_01281_));
 sg13g2_mux2_1 _23772_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][7] ),
    .A1(net976),
    .S(net371),
    .X(_01282_));
 sg13g2_mux2_1 _23773_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][8] ),
    .A1(net511),
    .S(_05918_),
    .X(_01283_));
 sg13g2_mux2_1 _23774_ (.A0(\cpu.genblk1.mmu.r_vtop_d[20][9] ),
    .A1(net512),
    .S(_05918_),
    .X(_01284_));
 sg13g2_nor2_1 _23775_ (.A(_05869_),
    .B(_05916_),
    .Y(_05920_));
 sg13g2_buf_1 _23776_ (.A(_05920_),
    .X(_05921_));
 sg13g2_buf_1 _23777_ (.A(_05921_),
    .X(_05922_));
 sg13g2_mux2_1 _23778_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][0] ),
    .A1(net510),
    .S(_05922_),
    .X(_01285_));
 sg13g2_mux2_1 _23779_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][10] ),
    .A1(net596),
    .S(net287),
    .X(_01286_));
 sg13g2_mux2_1 _23780_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][11] ),
    .A1(net597),
    .S(net287),
    .X(_01287_));
 sg13g2_mux2_1 _23781_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][1] ),
    .A1(net460),
    .S(_05922_),
    .X(_01288_));
 sg13g2_mux2_1 _23782_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][2] ),
    .A1(net862),
    .S(net287),
    .X(_01289_));
 sg13g2_mux2_1 _23783_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][3] ),
    .A1(net863),
    .S(net287),
    .X(_01290_));
 sg13g2_mux2_1 _23784_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][4] ),
    .A1(net865),
    .S(net287),
    .X(_01291_));
 sg13g2_mux2_1 _23785_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][5] ),
    .A1(net864),
    .S(net287),
    .X(_01292_));
 sg13g2_mux2_1 _23786_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][6] ),
    .A1(net977),
    .S(net287),
    .X(_01293_));
 sg13g2_mux2_1 _23787_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][7] ),
    .A1(net976),
    .S(net287),
    .X(_01294_));
 sg13g2_mux2_1 _23788_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][8] ),
    .A1(net511),
    .S(_05921_),
    .X(_01295_));
 sg13g2_mux2_1 _23789_ (.A0(\cpu.genblk1.mmu.r_vtop_d[21][9] ),
    .A1(net512),
    .S(_05921_),
    .X(_01296_));
 sg13g2_nor3_1 _23790_ (.A(net746),
    .B(net461),
    .C(_05916_),
    .Y(_05923_));
 sg13g2_buf_1 _23791_ (.A(_05923_),
    .X(_05924_));
 sg13g2_buf_1 _23792_ (.A(_05924_),
    .X(_05925_));
 sg13g2_mux2_1 _23793_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][0] ),
    .A1(net510),
    .S(_05925_),
    .X(_01297_));
 sg13g2_mux2_1 _23794_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][10] ),
    .A1(net596),
    .S(net332),
    .X(_01298_));
 sg13g2_mux2_1 _23795_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][11] ),
    .A1(net597),
    .S(net332),
    .X(_01299_));
 sg13g2_mux2_1 _23796_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][1] ),
    .A1(net460),
    .S(_05925_),
    .X(_01300_));
 sg13g2_mux2_1 _23797_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][2] ),
    .A1(net862),
    .S(net332),
    .X(_01301_));
 sg13g2_mux2_1 _23798_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][3] ),
    .A1(net863),
    .S(net332),
    .X(_01302_));
 sg13g2_mux2_1 _23799_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][4] ),
    .A1(net865),
    .S(net332),
    .X(_01303_));
 sg13g2_mux2_1 _23800_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][5] ),
    .A1(net864),
    .S(net332),
    .X(_01304_));
 sg13g2_mux2_1 _23801_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][6] ),
    .A1(net977),
    .S(net332),
    .X(_01305_));
 sg13g2_mux2_1 _23802_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][7] ),
    .A1(net976),
    .S(net332),
    .X(_01306_));
 sg13g2_mux2_1 _23803_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][8] ),
    .A1(net511),
    .S(_05924_),
    .X(_01307_));
 sg13g2_mux2_1 _23804_ (.A0(\cpu.genblk1.mmu.r_vtop_d[22][9] ),
    .A1(net512),
    .S(_05924_),
    .X(_01308_));
 sg13g2_nor3_1 _23805_ (.A(net867),
    .B(net461),
    .C(_05916_),
    .Y(_05926_));
 sg13g2_buf_1 _23806_ (.A(_05926_),
    .X(_05927_));
 sg13g2_buf_1 _23807_ (.A(_05927_),
    .X(_05928_));
 sg13g2_mux2_1 _23808_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][0] ),
    .A1(net510),
    .S(_05928_),
    .X(_01309_));
 sg13g2_mux2_1 _23809_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][10] ),
    .A1(net596),
    .S(net331),
    .X(_01310_));
 sg13g2_mux2_1 _23810_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][11] ),
    .A1(net597),
    .S(net331),
    .X(_01311_));
 sg13g2_mux2_1 _23811_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][1] ),
    .A1(net460),
    .S(_05928_),
    .X(_01312_));
 sg13g2_mux2_1 _23812_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][2] ),
    .A1(net862),
    .S(net331),
    .X(_01313_));
 sg13g2_mux2_1 _23813_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][3] ),
    .A1(net863),
    .S(net331),
    .X(_01314_));
 sg13g2_buf_1 _23814_ (.A(_09165_),
    .X(_05929_));
 sg13g2_mux2_1 _23815_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][4] ),
    .A1(net975),
    .S(net331),
    .X(_01315_));
 sg13g2_buf_1 _23816_ (.A(_10234_),
    .X(_05930_));
 sg13g2_mux2_1 _23817_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][5] ),
    .A1(net974),
    .S(net331),
    .X(_01316_));
 sg13g2_mux2_1 _23818_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][6] ),
    .A1(net977),
    .S(net331),
    .X(_01317_));
 sg13g2_mux2_1 _23819_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][7] ),
    .A1(net976),
    .S(net331),
    .X(_01318_));
 sg13g2_mux2_1 _23820_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][8] ),
    .A1(net511),
    .S(_05927_),
    .X(_01319_));
 sg13g2_mux2_1 _23821_ (.A0(\cpu.genblk1.mmu.r_vtop_d[23][9] ),
    .A1(net512),
    .S(_05927_),
    .X(_01320_));
 sg13g2_nand2_1 _23822_ (.Y(_05931_),
    .A(net978),
    .B(net1125));
 sg13g2_buf_2 _23823_ (.A(_05931_),
    .X(_05932_));
 sg13g2_nor3_1 _23824_ (.A(net461),
    .B(_05885_),
    .C(_05932_),
    .Y(_05933_));
 sg13g2_buf_1 _23825_ (.A(_05933_),
    .X(_05934_));
 sg13g2_buf_1 _23826_ (.A(_05934_),
    .X(_05935_));
 sg13g2_mux2_1 _23827_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][0] ),
    .A1(net510),
    .S(_05935_),
    .X(_01321_));
 sg13g2_mux2_1 _23828_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][10] ),
    .A1(net596),
    .S(net330),
    .X(_01322_));
 sg13g2_mux2_1 _23829_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][11] ),
    .A1(net597),
    .S(net330),
    .X(_01323_));
 sg13g2_buf_1 _23830_ (.A(_03072_),
    .X(_05936_));
 sg13g2_mux2_1 _23831_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][1] ),
    .A1(net509),
    .S(net330),
    .X(_01324_));
 sg13g2_mux2_1 _23832_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][2] ),
    .A1(_05914_),
    .S(_05935_),
    .X(_01325_));
 sg13g2_mux2_1 _23833_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][3] ),
    .A1(net863),
    .S(net330),
    .X(_01326_));
 sg13g2_mux2_1 _23834_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][4] ),
    .A1(net975),
    .S(net330),
    .X(_01327_));
 sg13g2_mux2_1 _23835_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][5] ),
    .A1(net974),
    .S(net330),
    .X(_01328_));
 sg13g2_mux2_1 _23836_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][6] ),
    .A1(net977),
    .S(net330),
    .X(_01329_));
 sg13g2_mux2_1 _23837_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][7] ),
    .A1(net976),
    .S(net330),
    .X(_01330_));
 sg13g2_mux2_1 _23838_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][8] ),
    .A1(_05904_),
    .S(_05934_),
    .X(_01331_));
 sg13g2_mux2_1 _23839_ (.A0(\cpu.genblk1.mmu.r_vtop_d[24][9] ),
    .A1(_05890_),
    .S(_05934_),
    .X(_01332_));
 sg13g2_nor3_1 _23840_ (.A(net979),
    .B(_05869_),
    .C(_05932_),
    .Y(_05937_));
 sg13g2_buf_1 _23841_ (.A(_05937_),
    .X(_05938_));
 sg13g2_buf_1 _23842_ (.A(_05938_),
    .X(_05939_));
 sg13g2_mux2_1 _23843_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][0] ),
    .A1(net510),
    .S(net286),
    .X(_01333_));
 sg13g2_mux2_1 _23844_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][10] ),
    .A1(_05901_),
    .S(net286),
    .X(_01334_));
 sg13g2_buf_1 _23845_ (.A(net687),
    .X(_05940_));
 sg13g2_mux2_1 _23846_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][11] ),
    .A1(net595),
    .S(net286),
    .X(_01335_));
 sg13g2_mux2_1 _23847_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][1] ),
    .A1(net509),
    .S(_05939_),
    .X(_01336_));
 sg13g2_mux2_1 _23848_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][2] ),
    .A1(_05914_),
    .S(_05939_),
    .X(_01337_));
 sg13g2_mux2_1 _23849_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][3] ),
    .A1(net863),
    .S(net286),
    .X(_01338_));
 sg13g2_mux2_1 _23850_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][4] ),
    .A1(net975),
    .S(net286),
    .X(_01339_));
 sg13g2_mux2_1 _23851_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][5] ),
    .A1(net974),
    .S(net286),
    .X(_01340_));
 sg13g2_mux2_1 _23852_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][6] ),
    .A1(net977),
    .S(net286),
    .X(_01341_));
 sg13g2_mux2_1 _23853_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][7] ),
    .A1(_05903_),
    .S(net286),
    .X(_01342_));
 sg13g2_mux2_1 _23854_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][8] ),
    .A1(_05904_),
    .S(_05938_),
    .X(_01343_));
 sg13g2_buf_1 _23855_ (.A(net628),
    .X(_05941_));
 sg13g2_mux2_1 _23856_ (.A0(\cpu.genblk1.mmu.r_vtop_d[25][9] ),
    .A1(net508),
    .S(_05938_),
    .X(_01344_));
 sg13g2_nor2_2 _23857_ (.A(net1035),
    .B(_05896_),
    .Y(_05942_));
 sg13g2_nor2b_1 _23858_ (.A(net462),
    .B_N(_05942_),
    .Y(_05943_));
 sg13g2_buf_1 _23859_ (.A(_05943_),
    .X(_05944_));
 sg13g2_buf_1 _23860_ (.A(_05944_),
    .X(_05945_));
 sg13g2_mux2_1 _23861_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][0] ),
    .A1(_05910_),
    .S(_05945_),
    .X(_01345_));
 sg13g2_mux2_1 _23862_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][10] ),
    .A1(net596),
    .S(net329),
    .X(_01346_));
 sg13g2_mux2_1 _23863_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][11] ),
    .A1(net595),
    .S(net329),
    .X(_01347_));
 sg13g2_mux2_1 _23864_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][1] ),
    .A1(net509),
    .S(_05945_),
    .X(_01348_));
 sg13g2_mux2_1 _23865_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][2] ),
    .A1(net862),
    .S(net329),
    .X(_01349_));
 sg13g2_buf_1 _23866_ (.A(net1154),
    .X(_05946_));
 sg13g2_mux2_1 _23867_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][3] ),
    .A1(net973),
    .S(net329),
    .X(_01350_));
 sg13g2_mux2_1 _23868_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][4] ),
    .A1(net975),
    .S(net329),
    .X(_01351_));
 sg13g2_mux2_1 _23869_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][5] ),
    .A1(net974),
    .S(net329),
    .X(_01352_));
 sg13g2_mux2_1 _23870_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][6] ),
    .A1(net977),
    .S(net329),
    .X(_01353_));
 sg13g2_mux2_1 _23871_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][7] ),
    .A1(_05903_),
    .S(net329),
    .X(_01354_));
 sg13g2_mux2_1 _23872_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][8] ),
    .A1(net511),
    .S(_05944_),
    .X(_01355_));
 sg13g2_mux2_1 _23873_ (.A0(\cpu.genblk1.mmu.r_vtop_d[26][9] ),
    .A1(net508),
    .S(_05944_),
    .X(_01356_));
 sg13g2_nor3_1 _23874_ (.A(_11375_),
    .B(_05818_),
    .C(_05932_),
    .Y(_05947_));
 sg13g2_buf_2 _23875_ (.A(_05947_),
    .X(_05948_));
 sg13g2_nor2b_1 _23876_ (.A(net462),
    .B_N(_05948_),
    .Y(_05949_));
 sg13g2_buf_1 _23877_ (.A(_05949_),
    .X(_05950_));
 sg13g2_buf_1 _23878_ (.A(_05950_),
    .X(_05951_));
 sg13g2_mux2_1 _23879_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][0] ),
    .A1(_05910_),
    .S(_05951_),
    .X(_01357_));
 sg13g2_buf_1 _23880_ (.A(_09523_),
    .X(_05952_));
 sg13g2_mux2_1 _23881_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][10] ),
    .A1(net594),
    .S(net328),
    .X(_01358_));
 sg13g2_mux2_1 _23882_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][11] ),
    .A1(net595),
    .S(net328),
    .X(_01359_));
 sg13g2_mux2_1 _23883_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][1] ),
    .A1(net509),
    .S(_05951_),
    .X(_01360_));
 sg13g2_mux2_1 _23884_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][2] ),
    .A1(net862),
    .S(net328),
    .X(_01361_));
 sg13g2_mux2_1 _23885_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][3] ),
    .A1(net973),
    .S(net328),
    .X(_01362_));
 sg13g2_mux2_1 _23886_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][4] ),
    .A1(net975),
    .S(net328),
    .X(_01363_));
 sg13g2_mux2_1 _23887_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][5] ),
    .A1(net974),
    .S(net328),
    .X(_01364_));
 sg13g2_buf_1 _23888_ (.A(_10143_),
    .X(_05953_));
 sg13g2_mux2_1 _23889_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][6] ),
    .A1(net972),
    .S(net328),
    .X(_01365_));
 sg13g2_buf_1 _23890_ (.A(_10322_),
    .X(_05954_));
 sg13g2_mux2_1 _23891_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][7] ),
    .A1(net971),
    .S(net328),
    .X(_01366_));
 sg13g2_buf_1 _23892_ (.A(_10810_),
    .X(_05955_));
 sg13g2_mux2_1 _23893_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][8] ),
    .A1(net507),
    .S(_05950_),
    .X(_01367_));
 sg13g2_mux2_1 _23894_ (.A0(\cpu.genblk1.mmu.r_vtop_d[27][9] ),
    .A1(net508),
    .S(_05950_),
    .X(_01368_));
 sg13g2_or2_1 _23895_ (.X(_05956_),
    .B(_05932_),
    .A(_05832_));
 sg13g2_buf_1 _23896_ (.A(_05956_),
    .X(_05957_));
 sg13g2_nor2_1 _23897_ (.A(_05838_),
    .B(_05957_),
    .Y(_05958_));
 sg13g2_buf_1 _23898_ (.A(_05958_),
    .X(_05959_));
 sg13g2_buf_1 _23899_ (.A(_05959_),
    .X(_05960_));
 sg13g2_mux2_1 _23900_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][0] ),
    .A1(net510),
    .S(_05960_),
    .X(_01369_));
 sg13g2_mux2_1 _23901_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][10] ),
    .A1(net594),
    .S(net370),
    .X(_01370_));
 sg13g2_mux2_1 _23902_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][11] ),
    .A1(net595),
    .S(net370),
    .X(_01371_));
 sg13g2_mux2_1 _23903_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][1] ),
    .A1(net509),
    .S(_05960_),
    .X(_01372_));
 sg13g2_mux2_1 _23904_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][2] ),
    .A1(net862),
    .S(net370),
    .X(_01373_));
 sg13g2_mux2_1 _23905_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][3] ),
    .A1(net973),
    .S(net370),
    .X(_01374_));
 sg13g2_mux2_1 _23906_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][4] ),
    .A1(net975),
    .S(net370),
    .X(_01375_));
 sg13g2_mux2_1 _23907_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][5] ),
    .A1(net974),
    .S(net370),
    .X(_01376_));
 sg13g2_mux2_1 _23908_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][6] ),
    .A1(net972),
    .S(net370),
    .X(_01377_));
 sg13g2_mux2_1 _23909_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][7] ),
    .A1(net971),
    .S(net370),
    .X(_01378_));
 sg13g2_mux2_1 _23910_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][8] ),
    .A1(net507),
    .S(_05959_),
    .X(_01379_));
 sg13g2_mux2_1 _23911_ (.A0(\cpu.genblk1.mmu.r_vtop_d[28][9] ),
    .A1(net508),
    .S(_05959_),
    .X(_01380_));
 sg13g2_buf_1 _23912_ (.A(_03624_),
    .X(_05961_));
 sg13g2_nor2_1 _23913_ (.A(_05869_),
    .B(_05957_),
    .Y(_05962_));
 sg13g2_buf_1 _23914_ (.A(_05962_),
    .X(_05963_));
 sg13g2_buf_1 _23915_ (.A(_05963_),
    .X(_05964_));
 sg13g2_mux2_1 _23916_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][0] ),
    .A1(net506),
    .S(_05964_),
    .X(_01381_));
 sg13g2_mux2_1 _23917_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][10] ),
    .A1(net594),
    .S(net285),
    .X(_01382_));
 sg13g2_mux2_1 _23918_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][11] ),
    .A1(net595),
    .S(net285),
    .X(_01383_));
 sg13g2_mux2_1 _23919_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][1] ),
    .A1(net509),
    .S(_05964_),
    .X(_01384_));
 sg13g2_buf_1 _23920_ (.A(net1000),
    .X(_05965_));
 sg13g2_mux2_1 _23921_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][2] ),
    .A1(net861),
    .S(net285),
    .X(_01385_));
 sg13g2_mux2_1 _23922_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][3] ),
    .A1(net973),
    .S(net285),
    .X(_01386_));
 sg13g2_mux2_1 _23923_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][4] ),
    .A1(net975),
    .S(net285),
    .X(_01387_));
 sg13g2_mux2_1 _23924_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][5] ),
    .A1(net974),
    .S(net285),
    .X(_01388_));
 sg13g2_mux2_1 _23925_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][6] ),
    .A1(net972),
    .S(net285),
    .X(_01389_));
 sg13g2_mux2_1 _23926_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][7] ),
    .A1(net971),
    .S(net285),
    .X(_01390_));
 sg13g2_mux2_1 _23927_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][8] ),
    .A1(net507),
    .S(_05963_),
    .X(_01391_));
 sg13g2_mux2_1 _23928_ (.A0(\cpu.genblk1.mmu.r_vtop_d[29][9] ),
    .A1(net508),
    .S(_05963_),
    .X(_01392_));
 sg13g2_nor3_1 _23929_ (.A(net746),
    .B(_05836_),
    .C(_05845_),
    .Y(_05966_));
 sg13g2_buf_1 _23930_ (.A(_05966_),
    .X(_05967_));
 sg13g2_buf_1 _23931_ (.A(_05967_),
    .X(_05968_));
 sg13g2_mux2_1 _23932_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][0] ),
    .A1(net506),
    .S(net327),
    .X(_01393_));
 sg13g2_mux2_1 _23933_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][10] ),
    .A1(net594),
    .S(net327),
    .X(_01394_));
 sg13g2_mux2_1 _23934_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][11] ),
    .A1(_05940_),
    .S(net327),
    .X(_01395_));
 sg13g2_mux2_1 _23935_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][1] ),
    .A1(net509),
    .S(net327),
    .X(_01396_));
 sg13g2_mux2_1 _23936_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][2] ),
    .A1(net861),
    .S(net327),
    .X(_01397_));
 sg13g2_mux2_1 _23937_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][3] ),
    .A1(_05946_),
    .S(_05968_),
    .X(_01398_));
 sg13g2_mux2_1 _23938_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][4] ),
    .A1(_05929_),
    .S(net327),
    .X(_01399_));
 sg13g2_mux2_1 _23939_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][5] ),
    .A1(_05930_),
    .S(_05968_),
    .X(_01400_));
 sg13g2_mux2_1 _23940_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][6] ),
    .A1(_05953_),
    .S(net327),
    .X(_01401_));
 sg13g2_mux2_1 _23941_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][7] ),
    .A1(net971),
    .S(net327),
    .X(_01402_));
 sg13g2_mux2_1 _23942_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][8] ),
    .A1(_05955_),
    .S(_05967_),
    .X(_01403_));
 sg13g2_mux2_1 _23943_ (.A0(\cpu.genblk1.mmu.r_vtop_d[2][9] ),
    .A1(net508),
    .S(_05967_),
    .X(_01404_));
 sg13g2_nor3_1 _23944_ (.A(net746),
    .B(net461),
    .C(_05957_),
    .Y(_05969_));
 sg13g2_buf_1 _23945_ (.A(_05969_),
    .X(_05970_));
 sg13g2_buf_1 _23946_ (.A(_05970_),
    .X(_05971_));
 sg13g2_mux2_1 _23947_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][0] ),
    .A1(net506),
    .S(_05971_),
    .X(_01405_));
 sg13g2_mux2_1 _23948_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][10] ),
    .A1(net594),
    .S(net326),
    .X(_01406_));
 sg13g2_mux2_1 _23949_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][11] ),
    .A1(net595),
    .S(net326),
    .X(_01407_));
 sg13g2_mux2_1 _23950_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][1] ),
    .A1(_05936_),
    .S(_05971_),
    .X(_01408_));
 sg13g2_mux2_1 _23951_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][2] ),
    .A1(net861),
    .S(net326),
    .X(_01409_));
 sg13g2_mux2_1 _23952_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][3] ),
    .A1(net973),
    .S(net326),
    .X(_01410_));
 sg13g2_mux2_1 _23953_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][4] ),
    .A1(net975),
    .S(net326),
    .X(_01411_));
 sg13g2_mux2_1 _23954_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][5] ),
    .A1(net974),
    .S(net326),
    .X(_01412_));
 sg13g2_mux2_1 _23955_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][6] ),
    .A1(net972),
    .S(net326),
    .X(_01413_));
 sg13g2_mux2_1 _23956_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][7] ),
    .A1(_05954_),
    .S(net326),
    .X(_01414_));
 sg13g2_mux2_1 _23957_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][8] ),
    .A1(net507),
    .S(_05970_),
    .X(_01415_));
 sg13g2_mux2_1 _23958_ (.A0(\cpu.genblk1.mmu.r_vtop_d[30][9] ),
    .A1(net508),
    .S(_05970_),
    .X(_01416_));
 sg13g2_nor3_1 _23959_ (.A(net867),
    .B(net461),
    .C(_05957_),
    .Y(_05972_));
 sg13g2_buf_1 _23960_ (.A(_05972_),
    .X(_05973_));
 sg13g2_buf_1 _23961_ (.A(_05973_),
    .X(_05974_));
 sg13g2_mux2_1 _23962_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][0] ),
    .A1(net506),
    .S(net325),
    .X(_01417_));
 sg13g2_mux2_1 _23963_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][10] ),
    .A1(net594),
    .S(net325),
    .X(_01418_));
 sg13g2_mux2_1 _23964_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][11] ),
    .A1(net595),
    .S(net325),
    .X(_01419_));
 sg13g2_mux2_1 _23965_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][1] ),
    .A1(_05936_),
    .S(_05974_),
    .X(_01420_));
 sg13g2_mux2_1 _23966_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][2] ),
    .A1(net861),
    .S(_05974_),
    .X(_01421_));
 sg13g2_mux2_1 _23967_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][3] ),
    .A1(net973),
    .S(net325),
    .X(_01422_));
 sg13g2_mux2_1 _23968_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][4] ),
    .A1(_05929_),
    .S(net325),
    .X(_01423_));
 sg13g2_mux2_1 _23969_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][5] ),
    .A1(_05930_),
    .S(net325),
    .X(_01424_));
 sg13g2_mux2_1 _23970_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][6] ),
    .A1(net972),
    .S(net325),
    .X(_01425_));
 sg13g2_mux2_1 _23971_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][7] ),
    .A1(_05954_),
    .S(net325),
    .X(_01426_));
 sg13g2_mux2_1 _23972_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][8] ),
    .A1(net507),
    .S(_05973_),
    .X(_01427_));
 sg13g2_mux2_1 _23973_ (.A0(\cpu.genblk1.mmu.r_vtop_d[31][9] ),
    .A1(net508),
    .S(_05973_),
    .X(_01428_));
 sg13g2_nor3_1 _23974_ (.A(net867),
    .B(_05836_),
    .C(net461),
    .Y(_05975_));
 sg13g2_buf_1 _23975_ (.A(_05975_),
    .X(_05976_));
 sg13g2_buf_1 _23976_ (.A(_05976_),
    .X(_05977_));
 sg13g2_mux2_1 _23977_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][0] ),
    .A1(net506),
    .S(net324),
    .X(_01429_));
 sg13g2_mux2_1 _23978_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][10] ),
    .A1(net594),
    .S(net324),
    .X(_01430_));
 sg13g2_mux2_1 _23979_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][11] ),
    .A1(_05940_),
    .S(net324),
    .X(_01431_));
 sg13g2_mux2_1 _23980_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][1] ),
    .A1(net509),
    .S(net324),
    .X(_01432_));
 sg13g2_mux2_1 _23981_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][2] ),
    .A1(net861),
    .S(net324),
    .X(_01433_));
 sg13g2_mux2_1 _23982_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][3] ),
    .A1(_05946_),
    .S(_05977_),
    .X(_01434_));
 sg13g2_mux2_1 _23983_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][4] ),
    .A1(net996),
    .S(net324),
    .X(_01435_));
 sg13g2_mux2_1 _23984_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][5] ),
    .A1(net995),
    .S(_05977_),
    .X(_01436_));
 sg13g2_mux2_1 _23985_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][6] ),
    .A1(net972),
    .S(net324),
    .X(_01437_));
 sg13g2_mux2_1 _23986_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][7] ),
    .A1(net971),
    .S(net324),
    .X(_01438_));
 sg13g2_mux2_1 _23987_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][8] ),
    .A1(_05955_),
    .S(_05976_),
    .X(_01439_));
 sg13g2_mux2_1 _23988_ (.A0(\cpu.genblk1.mmu.r_vtop_d[3][9] ),
    .A1(_05941_),
    .S(_05976_),
    .X(_01440_));
 sg13g2_nand2_1 _23989_ (.Y(_05978_),
    .A(net1123),
    .B(_05835_));
 sg13g2_nor2_1 _23990_ (.A(_05838_),
    .B(_05978_),
    .Y(_05979_));
 sg13g2_buf_1 _23991_ (.A(_05979_),
    .X(_05980_));
 sg13g2_buf_1 _23992_ (.A(_05980_),
    .X(_05981_));
 sg13g2_mux2_1 _23993_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][0] ),
    .A1(net506),
    .S(net369),
    .X(_01441_));
 sg13g2_mux2_1 _23994_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][10] ),
    .A1(net594),
    .S(net369),
    .X(_01442_));
 sg13g2_mux2_1 _23995_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][11] ),
    .A1(net595),
    .S(net369),
    .X(_01443_));
 sg13g2_mux2_1 _23996_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][1] ),
    .A1(net530),
    .S(net369),
    .X(_01444_));
 sg13g2_mux2_1 _23997_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][2] ),
    .A1(net861),
    .S(net369),
    .X(_01445_));
 sg13g2_mux2_1 _23998_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][3] ),
    .A1(net973),
    .S(net369),
    .X(_01446_));
 sg13g2_mux2_1 _23999_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][4] ),
    .A1(net996),
    .S(net369),
    .X(_01447_));
 sg13g2_mux2_1 _24000_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][5] ),
    .A1(net995),
    .S(_05981_),
    .X(_01448_));
 sg13g2_mux2_1 _24001_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][6] ),
    .A1(net972),
    .S(net369),
    .X(_01449_));
 sg13g2_mux2_1 _24002_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][7] ),
    .A1(net971),
    .S(_05981_),
    .X(_01450_));
 sg13g2_mux2_1 _24003_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][8] ),
    .A1(net507),
    .S(_05980_),
    .X(_01451_));
 sg13g2_mux2_1 _24004_ (.A0(\cpu.genblk1.mmu.r_vtop_d[4][9] ),
    .A1(_05941_),
    .S(_05980_),
    .X(_01452_));
 sg13g2_nor2_1 _24005_ (.A(_05867_),
    .B(_05978_),
    .Y(_05982_));
 sg13g2_buf_2 _24006_ (.A(_05982_),
    .X(_05983_));
 sg13g2_nor2b_1 _24007_ (.A(net462),
    .B_N(_05983_),
    .Y(_05984_));
 sg13g2_buf_1 _24008_ (.A(_05984_),
    .X(_05985_));
 sg13g2_buf_1 _24009_ (.A(_05985_),
    .X(_05986_));
 sg13g2_mux2_1 _24010_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][0] ),
    .A1(net506),
    .S(net323),
    .X(_01453_));
 sg13g2_mux2_1 _24011_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][10] ),
    .A1(_05952_),
    .S(net323),
    .X(_01454_));
 sg13g2_mux2_1 _24012_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][11] ),
    .A1(net617),
    .S(net323),
    .X(_01455_));
 sg13g2_mux2_1 _24013_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][1] ),
    .A1(net530),
    .S(net323),
    .X(_01456_));
 sg13g2_mux2_1 _24014_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][2] ),
    .A1(_05965_),
    .S(net323),
    .X(_01457_));
 sg13g2_mux2_1 _24015_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][3] ),
    .A1(net973),
    .S(net323),
    .X(_01458_));
 sg13g2_mux2_1 _24016_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][4] ),
    .A1(net996),
    .S(net323),
    .X(_01459_));
 sg13g2_mux2_1 _24017_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][5] ),
    .A1(net995),
    .S(_05986_),
    .X(_01460_));
 sg13g2_mux2_1 _24018_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][6] ),
    .A1(net972),
    .S(net323),
    .X(_01461_));
 sg13g2_mux2_1 _24019_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][7] ),
    .A1(net971),
    .S(_05986_),
    .X(_01462_));
 sg13g2_mux2_1 _24020_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][8] ),
    .A1(net507),
    .S(_05985_),
    .X(_01463_));
 sg13g2_mux2_1 _24021_ (.A0(\cpu.genblk1.mmu.r_vtop_d[5][9] ),
    .A1(net536),
    .S(_05985_),
    .X(_01464_));
 sg13g2_nor2_1 _24022_ (.A(net868),
    .B(net746),
    .Y(_05987_));
 sg13g2_and2_1 _24023_ (.A(_05835_),
    .B(_05987_),
    .X(_05988_));
 sg13g2_buf_1 _24024_ (.A(_05988_),
    .X(_05989_));
 sg13g2_nor2b_1 _24025_ (.A(net462),
    .B_N(_05989_),
    .Y(_05990_));
 sg13g2_buf_1 _24026_ (.A(_05990_),
    .X(_05991_));
 sg13g2_buf_1 _24027_ (.A(_05991_),
    .X(_05992_));
 sg13g2_mux2_1 _24028_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][0] ),
    .A1(net506),
    .S(net322),
    .X(_01465_));
 sg13g2_mux2_1 _24029_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][10] ),
    .A1(_05952_),
    .S(net322),
    .X(_01466_));
 sg13g2_mux2_1 _24030_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][11] ),
    .A1(net617),
    .S(net322),
    .X(_01467_));
 sg13g2_mux2_1 _24031_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][1] ),
    .A1(net530),
    .S(net322),
    .X(_01468_));
 sg13g2_mux2_1 _24032_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][2] ),
    .A1(net861),
    .S(net322),
    .X(_01469_));
 sg13g2_mux2_1 _24033_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][3] ),
    .A1(net997),
    .S(_05992_),
    .X(_01470_));
 sg13g2_mux2_1 _24034_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][4] ),
    .A1(net996),
    .S(net322),
    .X(_01471_));
 sg13g2_mux2_1 _24035_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][5] ),
    .A1(_03081_),
    .S(_05992_),
    .X(_01472_));
 sg13g2_mux2_1 _24036_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][6] ),
    .A1(_05953_),
    .S(net322),
    .X(_01473_));
 sg13g2_mux2_1 _24037_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][7] ),
    .A1(net971),
    .S(net322),
    .X(_01474_));
 sg13g2_mux2_1 _24038_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][8] ),
    .A1(net507),
    .S(_05991_),
    .X(_01475_));
 sg13g2_mux2_1 _24039_ (.A0(\cpu.genblk1.mmu.r_vtop_d[6][9] ),
    .A1(net536),
    .S(_05991_),
    .X(_01476_));
 sg13g2_and2_1 _24040_ (.A(_05819_),
    .B(_05835_),
    .X(_05993_));
 sg13g2_buf_2 _24041_ (.A(_05993_),
    .X(_05994_));
 sg13g2_nor2b_1 _24042_ (.A(_05845_),
    .B_N(_05994_),
    .Y(_05995_));
 sg13g2_buf_1 _24043_ (.A(_05995_),
    .X(_05996_));
 sg13g2_buf_1 _24044_ (.A(_05996_),
    .X(_05997_));
 sg13g2_mux2_1 _24045_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][0] ),
    .A1(_05961_),
    .S(net321),
    .X(_01477_));
 sg13g2_mux2_1 _24046_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][10] ),
    .A1(_03615_),
    .S(net321),
    .X(_01478_));
 sg13g2_mux2_1 _24047_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][11] ),
    .A1(net617),
    .S(net321),
    .X(_01479_));
 sg13g2_mux2_1 _24048_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][1] ),
    .A1(net530),
    .S(net321),
    .X(_01480_));
 sg13g2_mux2_1 _24049_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][2] ),
    .A1(net861),
    .S(net321),
    .X(_01481_));
 sg13g2_mux2_1 _24050_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][3] ),
    .A1(net997),
    .S(net321),
    .X(_01482_));
 sg13g2_mux2_1 _24051_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][4] ),
    .A1(_03079_),
    .S(net321),
    .X(_01483_));
 sg13g2_mux2_1 _24052_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][5] ),
    .A1(_03081_),
    .S(_05997_),
    .X(_01484_));
 sg13g2_mux2_1 _24053_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][6] ),
    .A1(net999),
    .S(net321),
    .X(_01485_));
 sg13g2_mux2_1 _24054_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][7] ),
    .A1(net998),
    .S(_05997_),
    .X(_01486_));
 sg13g2_mux2_1 _24055_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][8] ),
    .A1(_03611_),
    .S(_05996_),
    .X(_01487_));
 sg13g2_mux2_1 _24056_ (.A0(\cpu.genblk1.mmu.r_vtop_d[7][9] ),
    .A1(net536),
    .S(_05996_),
    .X(_01488_));
 sg13g2_nor3_1 _24057_ (.A(_05873_),
    .B(_05850_),
    .C(_05885_),
    .Y(_05998_));
 sg13g2_buf_1 _24058_ (.A(_05998_),
    .X(_05999_));
 sg13g2_buf_1 _24059_ (.A(_05999_),
    .X(_06000_));
 sg13g2_mux2_1 _24060_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][0] ),
    .A1(_05961_),
    .S(net320),
    .X(_01489_));
 sg13g2_mux2_1 _24061_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][10] ),
    .A1(net618),
    .S(net320),
    .X(_01490_));
 sg13g2_mux2_1 _24062_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][11] ),
    .A1(_03617_),
    .S(net320),
    .X(_01491_));
 sg13g2_mux2_1 _24063_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][1] ),
    .A1(_03642_),
    .S(net320),
    .X(_01492_));
 sg13g2_mux2_1 _24064_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][2] ),
    .A1(_05965_),
    .S(net320),
    .X(_01493_));
 sg13g2_mux2_1 _24065_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][3] ),
    .A1(_03077_),
    .S(net320),
    .X(_01494_));
 sg13g2_mux2_1 _24066_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][4] ),
    .A1(net996),
    .S(_06000_),
    .X(_01495_));
 sg13g2_mux2_1 _24067_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][5] ),
    .A1(net995),
    .S(net320),
    .X(_01496_));
 sg13g2_mux2_1 _24068_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][6] ),
    .A1(net999),
    .S(net320),
    .X(_01497_));
 sg13g2_mux2_1 _24069_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][7] ),
    .A1(net998),
    .S(_06000_),
    .X(_01498_));
 sg13g2_mux2_1 _24070_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][8] ),
    .A1(net537),
    .S(_05999_),
    .X(_01499_));
 sg13g2_mux2_1 _24071_ (.A0(\cpu.genblk1.mmu.r_vtop_d[8][9] ),
    .A1(_03613_),
    .S(_05999_),
    .X(_01500_));
 sg13g2_nor3_1 _24072_ (.A(_05820_),
    .B(_05850_),
    .C(_05869_),
    .Y(_06001_));
 sg13g2_buf_1 _24073_ (.A(_06001_),
    .X(_06002_));
 sg13g2_buf_1 _24074_ (.A(_06002_),
    .X(_06003_));
 sg13g2_mux2_1 _24075_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][0] ),
    .A1(net616),
    .S(net284),
    .X(_01501_));
 sg13g2_mux2_1 _24076_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][10] ),
    .A1(net618),
    .S(net284),
    .X(_01502_));
 sg13g2_mux2_1 _24077_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][11] ),
    .A1(_03617_),
    .S(net284),
    .X(_01503_));
 sg13g2_mux2_1 _24078_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][1] ),
    .A1(_03642_),
    .S(net284),
    .X(_01504_));
 sg13g2_mux2_1 _24079_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][2] ),
    .A1(_03057_),
    .S(net284),
    .X(_01505_));
 sg13g2_mux2_1 _24080_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][3] ),
    .A1(_03077_),
    .S(net284),
    .X(_01506_));
 sg13g2_mux2_1 _24081_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][4] ),
    .A1(net996),
    .S(net284),
    .X(_01507_));
 sg13g2_mux2_1 _24082_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][5] ),
    .A1(net995),
    .S(_06003_),
    .X(_01508_));
 sg13g2_mux2_1 _24083_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][6] ),
    .A1(_03068_),
    .S(net284),
    .X(_01509_));
 sg13g2_mux2_1 _24084_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][7] ),
    .A1(_03070_),
    .S(_06003_),
    .X(_01510_));
 sg13g2_mux2_1 _24085_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][8] ),
    .A1(_03611_),
    .S(_06002_),
    .X(_01511_));
 sg13g2_mux2_1 _24086_ (.A0(\cpu.genblk1.mmu.r_vtop_d[9][9] ),
    .A1(_03613_),
    .S(_06002_),
    .X(_01512_));
 sg13g2_and2_1 _24087_ (.A(_05832_),
    .B(_05835_),
    .X(_06004_));
 sg13g2_buf_1 _24088_ (.A(_06004_),
    .X(_06005_));
 sg13g2_nand2_1 _24089_ (.Y(_06006_),
    .A(net1162),
    .B(_05794_));
 sg13g2_nor2_1 _24090_ (.A(_11058_),
    .B(_06006_),
    .Y(_06007_));
 sg13g2_buf_1 _24091_ (.A(_06007_),
    .X(_06008_));
 sg13g2_and2_1 _24092_ (.A(_05808_),
    .B(_06008_),
    .X(_06009_));
 sg13g2_buf_1 _24093_ (.A(_06009_),
    .X(_06010_));
 sg13g2_nand2_1 _24094_ (.Y(_06011_),
    .A(_06005_),
    .B(_06010_));
 sg13g2_buf_2 _24095_ (.A(_06011_),
    .X(_06012_));
 sg13g2_buf_1 _24096_ (.A(_06012_),
    .X(_06013_));
 sg13g2_nand2_1 _24097_ (.Y(_06014_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][0] ),
    .B(_06012_));
 sg13g2_o21ai_1 _24098_ (.B1(_06014_),
    .Y(_01513_),
    .A1(net522),
    .A2(net241));
 sg13g2_mux2_1 _24099_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][10] ),
    .S(net241),
    .X(_01514_));
 sg13g2_mux2_1 _24100_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][11] ),
    .S(net241),
    .X(_01515_));
 sg13g2_nand2_1 _24101_ (.Y(_06015_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][1] ),
    .B(_06012_));
 sg13g2_o21ai_1 _24102_ (.B1(_06015_),
    .Y(_01516_),
    .A1(net674),
    .A2(net241));
 sg13g2_mux2_1 _24103_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][2] ),
    .S(net241),
    .X(_01517_));
 sg13g2_nand2_1 _24104_ (.Y(_06016_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][3] ),
    .B(_06012_));
 sg13g2_o21ai_1 _24105_ (.B1(_06016_),
    .Y(_01518_),
    .A1(net753),
    .A2(net241));
 sg13g2_nand2_1 _24106_ (.Y(_06017_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][4] ),
    .B(_06012_));
 sg13g2_o21ai_1 _24107_ (.B1(_06017_),
    .Y(_01519_),
    .A1(net752),
    .A2(_06013_));
 sg13g2_nand2_1 _24108_ (.Y(_06018_),
    .A(\cpu.genblk1.mmu.r_vtop_i[0][5] ),
    .B(_06012_));
 sg13g2_o21ai_1 _24109_ (.B1(_06018_),
    .Y(_01520_),
    .A1(net751),
    .A2(_06013_));
 sg13g2_mux2_1 _24110_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][6] ),
    .S(net241),
    .X(_01521_));
 sg13g2_mux2_1 _24111_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][7] ),
    .S(net241),
    .X(_01522_));
 sg13g2_mux2_1 _24112_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][8] ),
    .S(_06012_),
    .X(_01523_));
 sg13g2_mux2_1 _24113_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[0][9] ),
    .S(_06012_),
    .X(_01524_));
 sg13g2_buf_1 _24114_ (.A(_06008_),
    .X(_06019_));
 sg13g2_nand2_1 _24115_ (.Y(_06020_),
    .A(_05851_),
    .B(net407));
 sg13g2_buf_2 _24116_ (.A(_06020_),
    .X(_06021_));
 sg13g2_buf_1 _24117_ (.A(_06021_),
    .X(_06022_));
 sg13g2_nand2_1 _24118_ (.Y(_06023_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][0] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24119_ (.B1(_06023_),
    .Y(_01525_),
    .A1(net522),
    .A2(net283));
 sg13g2_mux2_1 _24120_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][10] ),
    .S(_06022_),
    .X(_01526_));
 sg13g2_mux2_1 _24121_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][11] ),
    .S(net283),
    .X(_01527_));
 sg13g2_nand2_1 _24122_ (.Y(_06024_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][1] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24123_ (.B1(_06024_),
    .Y(_01528_),
    .A1(_03051_),
    .A2(net283));
 sg13g2_mux2_1 _24124_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][2] ),
    .S(net283),
    .X(_01529_));
 sg13g2_nand2_1 _24125_ (.Y(_06025_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][3] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24126_ (.B1(_06025_),
    .Y(_01530_),
    .A1(_03060_),
    .A2(net283));
 sg13g2_nand2_1 _24127_ (.Y(_06026_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][4] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24128_ (.B1(_06026_),
    .Y(_01531_),
    .A1(_03063_),
    .A2(net283));
 sg13g2_nand2_1 _24129_ (.Y(_06027_),
    .A(\cpu.genblk1.mmu.r_vtop_i[10][5] ),
    .B(_06021_));
 sg13g2_o21ai_1 _24130_ (.B1(_06027_),
    .Y(_01532_),
    .A1(_03066_),
    .A2(net283));
 sg13g2_mux2_1 _24131_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][6] ),
    .S(net283),
    .X(_01533_));
 sg13g2_mux2_1 _24132_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][7] ),
    .S(_06022_),
    .X(_01534_));
 sg13g2_mux2_1 _24133_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][8] ),
    .S(_06021_),
    .X(_01535_));
 sg13g2_mux2_1 _24134_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[10][9] ),
    .S(_06021_),
    .X(_01536_));
 sg13g2_nand2_1 _24135_ (.Y(_06028_),
    .A(_05857_),
    .B(net407));
 sg13g2_buf_2 _24136_ (.A(_06028_),
    .X(_06029_));
 sg13g2_buf_1 _24137_ (.A(_06029_),
    .X(_06030_));
 sg13g2_nand2_1 _24138_ (.Y(_06031_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][0] ),
    .B(_06029_));
 sg13g2_o21ai_1 _24139_ (.B1(_06031_),
    .Y(_01537_),
    .A1(net522),
    .A2(net282));
 sg13g2_mux2_1 _24140_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][10] ),
    .S(_06030_),
    .X(_01538_));
 sg13g2_mux2_1 _24141_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][11] ),
    .S(net282),
    .X(_01539_));
 sg13g2_nand2_1 _24142_ (.Y(_06032_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][1] ),
    .B(_06029_));
 sg13g2_o21ai_1 _24143_ (.B1(_06032_),
    .Y(_01540_),
    .A1(_03051_),
    .A2(net282));
 sg13g2_mux2_1 _24144_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][2] ),
    .S(net282),
    .X(_01541_));
 sg13g2_nand2_1 _24145_ (.Y(_06033_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][3] ),
    .B(_06029_));
 sg13g2_o21ai_1 _24146_ (.B1(_06033_),
    .Y(_01542_),
    .A1(_03060_),
    .A2(net282));
 sg13g2_nand2_1 _24147_ (.Y(_06034_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][4] ),
    .B(_06029_));
 sg13g2_o21ai_1 _24148_ (.B1(_06034_),
    .Y(_01543_),
    .A1(_03063_),
    .A2(net282));
 sg13g2_nand2_1 _24149_ (.Y(_06035_),
    .A(\cpu.genblk1.mmu.r_vtop_i[11][5] ),
    .B(_06029_));
 sg13g2_o21ai_1 _24150_ (.B1(_06035_),
    .Y(_01544_),
    .A1(_03066_),
    .A2(net282));
 sg13g2_mux2_1 _24151_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][6] ),
    .S(net282),
    .X(_01545_));
 sg13g2_mux2_1 _24152_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][7] ),
    .S(_06030_),
    .X(_01546_));
 sg13g2_mux2_1 _24153_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][8] ),
    .S(_06029_),
    .X(_01547_));
 sg13g2_mux2_1 _24154_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[11][9] ),
    .S(_06029_),
    .X(_01548_));
 sg13g2_nor2_2 _24155_ (.A(_05832_),
    .B(_05850_),
    .Y(_06036_));
 sg13g2_nand2_1 _24156_ (.Y(_06037_),
    .A(_06036_),
    .B(_06010_));
 sg13g2_buf_2 _24157_ (.A(_06037_),
    .X(_06038_));
 sg13g2_buf_1 _24158_ (.A(_06038_),
    .X(_06039_));
 sg13g2_nand2_1 _24159_ (.Y(_06040_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][0] ),
    .B(_06038_));
 sg13g2_o21ai_1 _24160_ (.B1(_06040_),
    .Y(_01549_),
    .A1(net522),
    .A2(net240));
 sg13g2_mux2_1 _24161_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][10] ),
    .S(_06039_),
    .X(_01550_));
 sg13g2_mux2_1 _24162_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][11] ),
    .S(net240),
    .X(_01551_));
 sg13g2_nand2_1 _24163_ (.Y(_06041_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][1] ),
    .B(_06038_));
 sg13g2_o21ai_1 _24164_ (.B1(_06041_),
    .Y(_01552_),
    .A1(net674),
    .A2(net240));
 sg13g2_mux2_1 _24165_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][2] ),
    .S(net240),
    .X(_01553_));
 sg13g2_nand2_1 _24166_ (.Y(_06042_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][3] ),
    .B(_06038_));
 sg13g2_o21ai_1 _24167_ (.B1(_06042_),
    .Y(_01554_),
    .A1(net753),
    .A2(net240));
 sg13g2_nand2_1 _24168_ (.Y(_06043_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][4] ),
    .B(_06038_));
 sg13g2_o21ai_1 _24169_ (.B1(_06043_),
    .Y(_01555_),
    .A1(net752),
    .A2(net240));
 sg13g2_nand2_1 _24170_ (.Y(_06044_),
    .A(\cpu.genblk1.mmu.r_vtop_i[12][5] ),
    .B(_06038_));
 sg13g2_o21ai_1 _24171_ (.B1(_06044_),
    .Y(_01556_),
    .A1(net751),
    .A2(net240));
 sg13g2_mux2_1 _24172_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][6] ),
    .S(net240),
    .X(_01557_));
 sg13g2_mux2_1 _24173_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][7] ),
    .S(_06039_),
    .X(_01558_));
 sg13g2_mux2_1 _24174_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][8] ),
    .S(_06038_),
    .X(_01559_));
 sg13g2_mux2_1 _24175_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[12][9] ),
    .S(_06038_),
    .X(_01560_));
 sg13g2_nor3_1 _24176_ (.A(_11058_),
    .B(_05867_),
    .C(_06006_),
    .Y(_06045_));
 sg13g2_buf_2 _24177_ (.A(_06045_),
    .X(_06046_));
 sg13g2_nand2_1 _24178_ (.Y(_06047_),
    .A(_06036_),
    .B(_06046_));
 sg13g2_buf_2 _24179_ (.A(_06047_),
    .X(_06048_));
 sg13g2_buf_1 _24180_ (.A(_06048_),
    .X(_06049_));
 sg13g2_nand2_1 _24181_ (.Y(_06050_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][0] ),
    .B(_06048_));
 sg13g2_o21ai_1 _24182_ (.B1(_06050_),
    .Y(_01561_),
    .A1(net522),
    .A2(net319));
 sg13g2_mux2_1 _24183_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][10] ),
    .S(_06049_),
    .X(_01562_));
 sg13g2_mux2_1 _24184_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][11] ),
    .S(net319),
    .X(_01563_));
 sg13g2_nand2_1 _24185_ (.Y(_06051_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][1] ),
    .B(_06048_));
 sg13g2_o21ai_1 _24186_ (.B1(_06051_),
    .Y(_01564_),
    .A1(net674),
    .A2(net319));
 sg13g2_mux2_1 _24187_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][2] ),
    .S(net319),
    .X(_01565_));
 sg13g2_nand2_1 _24188_ (.Y(_06052_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][3] ),
    .B(_06048_));
 sg13g2_o21ai_1 _24189_ (.B1(_06052_),
    .Y(_01566_),
    .A1(net753),
    .A2(net319));
 sg13g2_nand2_1 _24190_ (.Y(_06053_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][4] ),
    .B(_06048_));
 sg13g2_o21ai_1 _24191_ (.B1(_06053_),
    .Y(_01567_),
    .A1(net752),
    .A2(net319));
 sg13g2_nand2_1 _24192_ (.Y(_06054_),
    .A(\cpu.genblk1.mmu.r_vtop_i[13][5] ),
    .B(_06048_));
 sg13g2_o21ai_1 _24193_ (.B1(_06054_),
    .Y(_01568_),
    .A1(net751),
    .A2(net319));
 sg13g2_mux2_1 _24194_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][6] ),
    .S(net319),
    .X(_01569_));
 sg13g2_mux2_1 _24195_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][7] ),
    .S(_06049_),
    .X(_01570_));
 sg13g2_mux2_1 _24196_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][8] ),
    .S(_06048_),
    .X(_01571_));
 sg13g2_mux2_1 _24197_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[13][9] ),
    .S(_06048_),
    .X(_01572_));
 sg13g2_nor2_2 _24198_ (.A(net980),
    .B(_10799_),
    .Y(_06055_));
 sg13g2_nand3_1 _24199_ (.B(_06036_),
    .C(_06019_),
    .A(_06055_),
    .Y(_06056_));
 sg13g2_buf_2 _24200_ (.A(_06056_),
    .X(_06057_));
 sg13g2_buf_1 _24201_ (.A(_06057_),
    .X(_06058_));
 sg13g2_nand2_1 _24202_ (.Y(_06059_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][0] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24203_ (.B1(_06059_),
    .Y(_01573_),
    .A1(net522),
    .A2(net281));
 sg13g2_mux2_1 _24204_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][10] ),
    .S(net281),
    .X(_01574_));
 sg13g2_mux2_1 _24205_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][11] ),
    .S(net281),
    .X(_01575_));
 sg13g2_nand2_1 _24206_ (.Y(_06060_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][1] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24207_ (.B1(_06060_),
    .Y(_01576_),
    .A1(net674),
    .A2(net281));
 sg13g2_mux2_1 _24208_ (.A0(net754),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][2] ),
    .S(net281),
    .X(_01577_));
 sg13g2_nand2_1 _24209_ (.Y(_06061_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][3] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24210_ (.B1(_06061_),
    .Y(_01578_),
    .A1(net753),
    .A2(net281));
 sg13g2_nand2_1 _24211_ (.Y(_06062_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][4] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24212_ (.B1(_06062_),
    .Y(_01579_),
    .A1(net752),
    .A2(_06058_));
 sg13g2_nand2_1 _24213_ (.Y(_06063_),
    .A(\cpu.genblk1.mmu.r_vtop_i[14][5] ),
    .B(_06057_));
 sg13g2_o21ai_1 _24214_ (.B1(_06063_),
    .Y(_01580_),
    .A1(net751),
    .A2(net281));
 sg13g2_mux2_1 _24215_ (.A0(net886),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][6] ),
    .S(net281),
    .X(_01581_));
 sg13g2_mux2_1 _24216_ (.A0(net885),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][7] ),
    .S(_06058_),
    .X(_01582_));
 sg13g2_mux2_1 _24217_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][8] ),
    .S(_06057_),
    .X(_01583_));
 sg13g2_mux2_1 _24218_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[14][9] ),
    .S(_06057_),
    .X(_01584_));
 sg13g2_buf_1 _24219_ (.A(_06008_),
    .X(_06064_));
 sg13g2_nand3_1 _24220_ (.B(_06036_),
    .C(net406),
    .A(_05806_),
    .Y(_06065_));
 sg13g2_buf_2 _24221_ (.A(_06065_),
    .X(_06066_));
 sg13g2_buf_1 _24222_ (.A(_06066_),
    .X(_06067_));
 sg13g2_nand2_1 _24223_ (.Y(_06068_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][0] ),
    .B(_06066_));
 sg13g2_o21ai_1 _24224_ (.B1(_06068_),
    .Y(_01585_),
    .A1(net522),
    .A2(_06067_));
 sg13g2_mux2_1 _24225_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][10] ),
    .S(net280),
    .X(_01586_));
 sg13g2_mux2_1 _24226_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][11] ),
    .S(net280),
    .X(_01587_));
 sg13g2_buf_1 _24227_ (.A(net755),
    .X(_06069_));
 sg13g2_nand2_1 _24228_ (.Y(_06070_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][1] ),
    .B(_06066_));
 sg13g2_o21ai_1 _24229_ (.B1(_06070_),
    .Y(_01588_),
    .A1(_06069_),
    .A2(net280));
 sg13g2_buf_1 _24230_ (.A(net890),
    .X(_06071_));
 sg13g2_mux2_1 _24231_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][2] ),
    .S(net280),
    .X(_01589_));
 sg13g2_buf_1 _24232_ (.A(net889),
    .X(_06072_));
 sg13g2_nand2_1 _24233_ (.Y(_06073_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][3] ),
    .B(_06066_));
 sg13g2_o21ai_1 _24234_ (.B1(_06073_),
    .Y(_01590_),
    .A1(_06072_),
    .A2(net280));
 sg13g2_buf_1 _24235_ (.A(net888),
    .X(_06074_));
 sg13g2_nand2_1 _24236_ (.Y(_06075_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][4] ),
    .B(_06066_));
 sg13g2_o21ai_1 _24237_ (.B1(_06075_),
    .Y(_01591_),
    .A1(_06074_),
    .A2(net280));
 sg13g2_buf_1 _24238_ (.A(net887),
    .X(_06076_));
 sg13g2_nand2_1 _24239_ (.Y(_06077_),
    .A(\cpu.genblk1.mmu.r_vtop_i[15][5] ),
    .B(_06066_));
 sg13g2_o21ai_1 _24240_ (.B1(_06077_),
    .Y(_01592_),
    .A1(_06076_),
    .A2(_06067_));
 sg13g2_buf_1 _24241_ (.A(net999),
    .X(_06078_));
 sg13g2_mux2_1 _24242_ (.A0(_06078_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][6] ),
    .S(net280),
    .X(_01593_));
 sg13g2_buf_1 _24243_ (.A(net998),
    .X(_06079_));
 sg13g2_mux2_1 _24244_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][7] ),
    .S(net280),
    .X(_01594_));
 sg13g2_mux2_1 _24245_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][8] ),
    .S(_06066_),
    .X(_01595_));
 sg13g2_mux2_1 _24246_ (.A0(net464),
    .A1(\cpu.genblk1.mmu.r_vtop_i[15][9] ),
    .S(_06066_),
    .X(_01596_));
 sg13g2_nor3_2 _24247_ (.A(net980),
    .B(net1124),
    .C(net979),
    .Y(_06080_));
 sg13g2_nand4_1 _24248_ (.B(net1035),
    .C(_06080_),
    .A(net978),
    .Y(_06081_),
    .D(net406));
 sg13g2_buf_2 _24249_ (.A(_06081_),
    .X(_06082_));
 sg13g2_buf_1 _24250_ (.A(_06082_),
    .X(_06083_));
 sg13g2_nand2_1 _24251_ (.Y(_06084_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][0] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24252_ (.B1(_06084_),
    .Y(_01597_),
    .A1(net522),
    .A2(net279));
 sg13g2_mux2_1 _24253_ (.A0(net524),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][10] ),
    .S(net279),
    .X(_01598_));
 sg13g2_mux2_1 _24254_ (.A0(net523),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][11] ),
    .S(net279),
    .X(_01599_));
 sg13g2_nand2_1 _24255_ (.Y(_06085_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][1] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24256_ (.B1(_06085_),
    .Y(_01600_),
    .A1(net662),
    .A2(net279));
 sg13g2_mux2_1 _24257_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][2] ),
    .S(_06083_),
    .X(_01601_));
 sg13g2_nand2_1 _24258_ (.Y(_06086_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][3] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24259_ (.B1(_06086_),
    .Y(_01602_),
    .A1(net744),
    .A2(net279));
 sg13g2_nand2_1 _24260_ (.Y(_06087_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][4] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24261_ (.B1(_06087_),
    .Y(_01603_),
    .A1(net743),
    .A2(net279));
 sg13g2_nand2_1 _24262_ (.Y(_06088_),
    .A(\cpu.genblk1.mmu.r_vtop_i[16][5] ),
    .B(_06082_));
 sg13g2_o21ai_1 _24263_ (.B1(_06088_),
    .Y(_01604_),
    .A1(net742),
    .A2(net279));
 sg13g2_mux2_1 _24264_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][6] ),
    .S(net279),
    .X(_01605_));
 sg13g2_mux2_1 _24265_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][7] ),
    .S(_06083_),
    .X(_01606_));
 sg13g2_mux2_1 _24266_ (.A0(net465),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][8] ),
    .S(_06082_),
    .X(_01607_));
 sg13g2_mux2_1 _24267_ (.A0(_03673_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[16][9] ),
    .S(_06082_),
    .X(_01608_));
 sg13g2_buf_1 _24268_ (.A(net608),
    .X(_06089_));
 sg13g2_nand4_1 _24269_ (.B(net868),
    .C(net1035),
    .A(net978),
    .Y(_06090_),
    .D(_06046_));
 sg13g2_buf_2 _24270_ (.A(_06090_),
    .X(_06091_));
 sg13g2_buf_1 _24271_ (.A(_06091_),
    .X(_06092_));
 sg13g2_nand2_1 _24272_ (.Y(_06093_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][0] ),
    .B(_06091_));
 sg13g2_o21ai_1 _24273_ (.B1(_06093_),
    .Y(_01609_),
    .A1(net505),
    .A2(net318));
 sg13g2_buf_1 _24274_ (.A(net618),
    .X(_06094_));
 sg13g2_mux2_1 _24275_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][10] ),
    .S(_06092_),
    .X(_01610_));
 sg13g2_buf_1 _24276_ (.A(net617),
    .X(_06095_));
 sg13g2_mux2_1 _24277_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][11] ),
    .S(net318),
    .X(_01611_));
 sg13g2_nand2_1 _24278_ (.Y(_06096_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][1] ),
    .B(_06091_));
 sg13g2_o21ai_1 _24279_ (.B1(_06096_),
    .Y(_01612_),
    .A1(net662),
    .A2(net318));
 sg13g2_mux2_1 _24280_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][2] ),
    .S(net318),
    .X(_01613_));
 sg13g2_nand2_1 _24281_ (.Y(_06097_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][3] ),
    .B(_06091_));
 sg13g2_o21ai_1 _24282_ (.B1(_06097_),
    .Y(_01614_),
    .A1(net744),
    .A2(net318));
 sg13g2_nand2_1 _24283_ (.Y(_06098_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][4] ),
    .B(_06091_));
 sg13g2_o21ai_1 _24284_ (.B1(_06098_),
    .Y(_01615_),
    .A1(net743),
    .A2(net318));
 sg13g2_nand2_1 _24285_ (.Y(_06099_),
    .A(\cpu.genblk1.mmu.r_vtop_i[17][5] ),
    .B(_06091_));
 sg13g2_o21ai_1 _24286_ (.B1(_06099_),
    .Y(_01616_),
    .A1(net742),
    .A2(net318));
 sg13g2_mux2_1 _24287_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][6] ),
    .S(net318),
    .X(_01617_));
 sg13g2_mux2_1 _24288_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][7] ),
    .S(_06092_),
    .X(_01618_));
 sg13g2_buf_1 _24289_ (.A(net537),
    .X(_06100_));
 sg13g2_mux2_1 _24290_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][8] ),
    .S(_06091_),
    .X(_01619_));
 sg13g2_buf_1 _24291_ (.A(net536),
    .X(_06101_));
 sg13g2_mux2_1 _24292_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[17][9] ),
    .S(_06091_),
    .X(_01620_));
 sg13g2_nand2_1 _24293_ (.Y(_06102_),
    .A(_05897_),
    .B(net407));
 sg13g2_buf_2 _24294_ (.A(_06102_),
    .X(_06103_));
 sg13g2_buf_1 _24295_ (.A(_06103_),
    .X(_06104_));
 sg13g2_nand2_1 _24296_ (.Y(_06105_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][0] ),
    .B(_06103_));
 sg13g2_o21ai_1 _24297_ (.B1(_06105_),
    .Y(_01621_),
    .A1(net505),
    .A2(net278));
 sg13g2_mux2_1 _24298_ (.A0(_06094_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][10] ),
    .S(_06104_),
    .X(_01622_));
 sg13g2_mux2_1 _24299_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][11] ),
    .S(net278),
    .X(_01623_));
 sg13g2_nand2_1 _24300_ (.Y(_06106_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][1] ),
    .B(_06103_));
 sg13g2_o21ai_1 _24301_ (.B1(_06106_),
    .Y(_01624_),
    .A1(net662),
    .A2(net278));
 sg13g2_mux2_1 _24302_ (.A0(_06071_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][2] ),
    .S(net278),
    .X(_01625_));
 sg13g2_nand2_1 _24303_ (.Y(_06107_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][3] ),
    .B(_06103_));
 sg13g2_o21ai_1 _24304_ (.B1(_06107_),
    .Y(_01626_),
    .A1(net744),
    .A2(net278));
 sg13g2_nand2_1 _24305_ (.Y(_06108_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][4] ),
    .B(_06103_));
 sg13g2_o21ai_1 _24306_ (.B1(_06108_),
    .Y(_01627_),
    .A1(net743),
    .A2(net278));
 sg13g2_nand2_1 _24307_ (.Y(_06109_),
    .A(\cpu.genblk1.mmu.r_vtop_i[18][5] ),
    .B(_06103_));
 sg13g2_o21ai_1 _24308_ (.B1(_06109_),
    .Y(_01628_),
    .A1(net742),
    .A2(net278));
 sg13g2_mux2_1 _24309_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][6] ),
    .S(net278),
    .X(_01629_));
 sg13g2_mux2_1 _24310_ (.A0(_06079_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][7] ),
    .S(_06104_),
    .X(_01630_));
 sg13g2_mux2_1 _24311_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][8] ),
    .S(_06103_),
    .X(_01631_));
 sg13g2_mux2_1 _24312_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[18][9] ),
    .S(_06103_),
    .X(_01632_));
 sg13g2_nand2_1 _24313_ (.Y(_06110_),
    .A(_05906_),
    .B(net407));
 sg13g2_buf_2 _24314_ (.A(_06110_),
    .X(_06111_));
 sg13g2_buf_1 _24315_ (.A(_06111_),
    .X(_06112_));
 sg13g2_nand2_1 _24316_ (.Y(_06113_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][0] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24317_ (.B1(_06113_),
    .Y(_01633_),
    .A1(net505),
    .A2(net277));
 sg13g2_mux2_1 _24318_ (.A0(_06094_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][10] ),
    .S(_06112_),
    .X(_01634_));
 sg13g2_mux2_1 _24319_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][11] ),
    .S(net277),
    .X(_01635_));
 sg13g2_nand2_1 _24320_ (.Y(_06114_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][1] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24321_ (.B1(_06114_),
    .Y(_01636_),
    .A1(net662),
    .A2(net277));
 sg13g2_mux2_1 _24322_ (.A0(_06071_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][2] ),
    .S(_06112_),
    .X(_01637_));
 sg13g2_nand2_1 _24323_ (.Y(_06115_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][3] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24324_ (.B1(_06115_),
    .Y(_01638_),
    .A1(net744),
    .A2(net277));
 sg13g2_nand2_1 _24325_ (.Y(_06116_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][4] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24326_ (.B1(_06116_),
    .Y(_01639_),
    .A1(net743),
    .A2(net277));
 sg13g2_nand2_1 _24327_ (.Y(_06117_),
    .A(\cpu.genblk1.mmu.r_vtop_i[19][5] ),
    .B(_06111_));
 sg13g2_o21ai_1 _24328_ (.B1(_06117_),
    .Y(_01640_),
    .A1(net742),
    .A2(net277));
 sg13g2_mux2_1 _24329_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][6] ),
    .S(net277),
    .X(_01641_));
 sg13g2_mux2_1 _24330_ (.A0(_06079_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][7] ),
    .S(net277),
    .X(_01642_));
 sg13g2_mux2_1 _24331_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][8] ),
    .S(_06111_),
    .X(_01643_));
 sg13g2_mux2_1 _24332_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[19][9] ),
    .S(_06111_),
    .X(_01644_));
 sg13g2_nand2_1 _24333_ (.Y(_06118_),
    .A(_06005_),
    .B(_06046_));
 sg13g2_buf_2 _24334_ (.A(_06118_),
    .X(_06119_));
 sg13g2_buf_1 _24335_ (.A(_06119_),
    .X(_06120_));
 sg13g2_nand2_1 _24336_ (.Y(_06121_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][0] ),
    .B(_06119_));
 sg13g2_o21ai_1 _24337_ (.B1(_06121_),
    .Y(_01645_),
    .A1(_06089_),
    .A2(net317));
 sg13g2_mux2_1 _24338_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][10] ),
    .S(net317),
    .X(_01646_));
 sg13g2_mux2_1 _24339_ (.A0(_06095_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][11] ),
    .S(net317),
    .X(_01647_));
 sg13g2_nand2_1 _24340_ (.Y(_06122_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][1] ),
    .B(_06119_));
 sg13g2_o21ai_1 _24341_ (.B1(_06122_),
    .Y(_01648_),
    .A1(_06069_),
    .A2(net317));
 sg13g2_mux2_1 _24342_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][2] ),
    .S(net317),
    .X(_01649_));
 sg13g2_nand2_1 _24343_ (.Y(_06123_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][3] ),
    .B(_06119_));
 sg13g2_o21ai_1 _24344_ (.B1(_06123_),
    .Y(_01650_),
    .A1(_06072_),
    .A2(net317));
 sg13g2_nand2_1 _24345_ (.Y(_06124_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][4] ),
    .B(_06119_));
 sg13g2_o21ai_1 _24346_ (.B1(_06124_),
    .Y(_01651_),
    .A1(_06074_),
    .A2(_06120_));
 sg13g2_nand2_1 _24347_ (.Y(_06125_),
    .A(\cpu.genblk1.mmu.r_vtop_i[1][5] ),
    .B(_06119_));
 sg13g2_o21ai_1 _24348_ (.B1(_06125_),
    .Y(_01652_),
    .A1(_06076_),
    .A2(_06120_));
 sg13g2_mux2_1 _24349_ (.A0(_06078_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][6] ),
    .S(net317),
    .X(_01653_));
 sg13g2_mux2_1 _24350_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][7] ),
    .S(net317),
    .X(_01654_));
 sg13g2_mux2_1 _24351_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][8] ),
    .S(_06119_),
    .X(_01655_));
 sg13g2_mux2_1 _24352_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[1][9] ),
    .S(_06119_),
    .X(_01656_));
 sg13g2_nor2_2 _24353_ (.A(_05832_),
    .B(_05884_),
    .Y(_06126_));
 sg13g2_nand2_1 _24354_ (.Y(_06127_),
    .A(_06126_),
    .B(_06010_));
 sg13g2_buf_2 _24355_ (.A(_06127_),
    .X(_06128_));
 sg13g2_buf_1 _24356_ (.A(_06128_),
    .X(_06129_));
 sg13g2_nand2_1 _24357_ (.Y(_06130_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][0] ),
    .B(_06128_));
 sg13g2_o21ai_1 _24358_ (.B1(_06130_),
    .Y(_01657_),
    .A1(net505),
    .A2(net239));
 sg13g2_mux2_1 _24359_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][10] ),
    .S(net239),
    .X(_01658_));
 sg13g2_mux2_1 _24360_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][11] ),
    .S(_06129_),
    .X(_01659_));
 sg13g2_nand2_1 _24361_ (.Y(_06131_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][1] ),
    .B(_06128_));
 sg13g2_o21ai_1 _24362_ (.B1(_06131_),
    .Y(_01660_),
    .A1(net662),
    .A2(net239));
 sg13g2_mux2_1 _24363_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][2] ),
    .S(net239),
    .X(_01661_));
 sg13g2_nand2_1 _24364_ (.Y(_06132_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][3] ),
    .B(_06128_));
 sg13g2_o21ai_1 _24365_ (.B1(_06132_),
    .Y(_01662_),
    .A1(net744),
    .A2(net239));
 sg13g2_nand2_1 _24366_ (.Y(_06133_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][4] ),
    .B(_06128_));
 sg13g2_o21ai_1 _24367_ (.B1(_06133_),
    .Y(_01663_),
    .A1(net743),
    .A2(net239));
 sg13g2_nand2_1 _24368_ (.Y(_06134_),
    .A(\cpu.genblk1.mmu.r_vtop_i[20][5] ),
    .B(_06128_));
 sg13g2_o21ai_1 _24369_ (.B1(_06134_),
    .Y(_01664_),
    .A1(net742),
    .A2(net239));
 sg13g2_mux2_1 _24370_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][6] ),
    .S(net239),
    .X(_01665_));
 sg13g2_mux2_1 _24371_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][7] ),
    .S(_06129_),
    .X(_01666_));
 sg13g2_mux2_1 _24372_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][8] ),
    .S(_06128_),
    .X(_01667_));
 sg13g2_mux2_1 _24373_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[20][9] ),
    .S(_06128_),
    .X(_01668_));
 sg13g2_nand2_1 _24374_ (.Y(_06135_),
    .A(_06126_),
    .B(_06046_));
 sg13g2_buf_2 _24375_ (.A(_06135_),
    .X(_06136_));
 sg13g2_buf_1 _24376_ (.A(_06136_),
    .X(_06137_));
 sg13g2_nand2_1 _24377_ (.Y(_06138_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][0] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24378_ (.B1(_06138_),
    .Y(_01669_),
    .A1(net505),
    .A2(net316));
 sg13g2_mux2_1 _24379_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][10] ),
    .S(net316),
    .X(_01670_));
 sg13g2_mux2_1 _24380_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][11] ),
    .S(_06137_),
    .X(_01671_));
 sg13g2_nand2_1 _24381_ (.Y(_06139_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][1] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24382_ (.B1(_06139_),
    .Y(_01672_),
    .A1(net662),
    .A2(net316));
 sg13g2_mux2_1 _24383_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][2] ),
    .S(net316),
    .X(_01673_));
 sg13g2_nand2_1 _24384_ (.Y(_06140_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][3] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24385_ (.B1(_06140_),
    .Y(_01674_),
    .A1(net744),
    .A2(net316));
 sg13g2_nand2_1 _24386_ (.Y(_06141_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][4] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24387_ (.B1(_06141_),
    .Y(_01675_),
    .A1(net743),
    .A2(net316));
 sg13g2_nand2_1 _24388_ (.Y(_06142_),
    .A(\cpu.genblk1.mmu.r_vtop_i[21][5] ),
    .B(_06136_));
 sg13g2_o21ai_1 _24389_ (.B1(_06142_),
    .Y(_01676_),
    .A1(net742),
    .A2(net316));
 sg13g2_mux2_1 _24390_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][6] ),
    .S(net316),
    .X(_01677_));
 sg13g2_mux2_1 _24391_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][7] ),
    .S(_06137_),
    .X(_01678_));
 sg13g2_mux2_1 _24392_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][8] ),
    .S(_06136_),
    .X(_01679_));
 sg13g2_mux2_1 _24393_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[21][9] ),
    .S(_06136_),
    .X(_01680_));
 sg13g2_nand3_1 _24394_ (.B(_06126_),
    .C(net406),
    .A(_06055_),
    .Y(_06143_));
 sg13g2_buf_2 _24395_ (.A(_06143_),
    .X(_06144_));
 sg13g2_buf_1 _24396_ (.A(_06144_),
    .X(_06145_));
 sg13g2_nand2_1 _24397_ (.Y(_06146_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][0] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24398_ (.B1(_06146_),
    .Y(_01681_),
    .A1(net505),
    .A2(net276));
 sg13g2_mux2_1 _24399_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][10] ),
    .S(net276),
    .X(_01682_));
 sg13g2_mux2_1 _24400_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][11] ),
    .S(_06145_),
    .X(_01683_));
 sg13g2_nand2_1 _24401_ (.Y(_06147_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][1] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24402_ (.B1(_06147_),
    .Y(_01684_),
    .A1(net662),
    .A2(net276));
 sg13g2_mux2_1 _24403_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][2] ),
    .S(net276),
    .X(_01685_));
 sg13g2_nand2_1 _24404_ (.Y(_06148_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][3] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24405_ (.B1(_06148_),
    .Y(_01686_),
    .A1(net744),
    .A2(net276));
 sg13g2_nand2_1 _24406_ (.Y(_06149_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][4] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24407_ (.B1(_06149_),
    .Y(_01687_),
    .A1(net743),
    .A2(net276));
 sg13g2_nand2_1 _24408_ (.Y(_06150_),
    .A(\cpu.genblk1.mmu.r_vtop_i[22][5] ),
    .B(_06144_));
 sg13g2_o21ai_1 _24409_ (.B1(_06150_),
    .Y(_01688_),
    .A1(net742),
    .A2(net276));
 sg13g2_mux2_1 _24410_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][6] ),
    .S(net276),
    .X(_01689_));
 sg13g2_mux2_1 _24411_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][7] ),
    .S(_06145_),
    .X(_01690_));
 sg13g2_mux2_1 _24412_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][8] ),
    .S(_06144_),
    .X(_01691_));
 sg13g2_mux2_1 _24413_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[22][9] ),
    .S(_06144_),
    .X(_01692_));
 sg13g2_nand3_1 _24414_ (.B(_06126_),
    .C(net406),
    .A(_05806_),
    .Y(_06151_));
 sg13g2_buf_2 _24415_ (.A(_06151_),
    .X(_06152_));
 sg13g2_buf_1 _24416_ (.A(_06152_),
    .X(_06153_));
 sg13g2_nand2_1 _24417_ (.Y(_06154_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][0] ),
    .B(_06152_));
 sg13g2_o21ai_1 _24418_ (.B1(_06154_),
    .Y(_01693_),
    .A1(net505),
    .A2(net275));
 sg13g2_mux2_1 _24419_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][10] ),
    .S(net275),
    .X(_01694_));
 sg13g2_mux2_1 _24420_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][11] ),
    .S(net275),
    .X(_01695_));
 sg13g2_nand2_1 _24421_ (.Y(_06155_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][1] ),
    .B(_06152_));
 sg13g2_o21ai_1 _24422_ (.B1(_06155_),
    .Y(_01696_),
    .A1(net662),
    .A2(net275));
 sg13g2_mux2_1 _24423_ (.A0(net745),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][2] ),
    .S(net275),
    .X(_01697_));
 sg13g2_nand2_1 _24424_ (.Y(_06156_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][3] ),
    .B(_06152_));
 sg13g2_o21ai_1 _24425_ (.B1(_06156_),
    .Y(_01698_),
    .A1(net744),
    .A2(net275));
 sg13g2_nand2_1 _24426_ (.Y(_06157_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][4] ),
    .B(_06152_));
 sg13g2_o21ai_1 _24427_ (.B1(_06157_),
    .Y(_01699_),
    .A1(net743),
    .A2(_06153_));
 sg13g2_nand2_1 _24428_ (.Y(_06158_),
    .A(\cpu.genblk1.mmu.r_vtop_i[23][5] ),
    .B(_06152_));
 sg13g2_o21ai_1 _24429_ (.B1(_06158_),
    .Y(_01700_),
    .A1(net742),
    .A2(net275));
 sg13g2_mux2_1 _24430_ (.A0(net860),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][6] ),
    .S(net275),
    .X(_01701_));
 sg13g2_mux2_1 _24431_ (.A0(net859),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][7] ),
    .S(_06153_),
    .X(_01702_));
 sg13g2_mux2_1 _24432_ (.A0(net459),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][8] ),
    .S(_06152_),
    .X(_01703_));
 sg13g2_mux2_1 _24433_ (.A0(net458),
    .A1(\cpu.genblk1.mmu.r_vtop_i[23][9] ),
    .S(_06152_),
    .X(_01704_));
 sg13g2_inv_1 _24434_ (.Y(_06159_),
    .A(_05932_));
 sg13g2_nand3_1 _24435_ (.B(_06159_),
    .C(_06064_),
    .A(_06080_),
    .Y(_06160_));
 sg13g2_buf_2 _24436_ (.A(_06160_),
    .X(_06161_));
 sg13g2_buf_1 _24437_ (.A(_06161_),
    .X(_06162_));
 sg13g2_nand2_1 _24438_ (.Y(_06163_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][0] ),
    .B(_06161_));
 sg13g2_o21ai_1 _24439_ (.B1(_06163_),
    .Y(_01705_),
    .A1(net505),
    .A2(net274));
 sg13g2_mux2_1 _24440_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][10] ),
    .S(net274),
    .X(_01706_));
 sg13g2_mux2_1 _24441_ (.A0(net503),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][11] ),
    .S(net274),
    .X(_01707_));
 sg13g2_buf_1 _24442_ (.A(_03050_),
    .X(_06164_));
 sg13g2_nand2_1 _24443_ (.Y(_06165_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][1] ),
    .B(_06161_));
 sg13g2_o21ai_1 _24444_ (.B1(_06165_),
    .Y(_01708_),
    .A1(net661),
    .A2(net274));
 sg13g2_buf_1 _24445_ (.A(net890),
    .X(_06166_));
 sg13g2_mux2_1 _24446_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][2] ),
    .S(net274),
    .X(_01709_));
 sg13g2_buf_1 _24447_ (.A(net889),
    .X(_06167_));
 sg13g2_nand2_1 _24448_ (.Y(_06168_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][3] ),
    .B(_06161_));
 sg13g2_o21ai_1 _24449_ (.B1(_06168_),
    .Y(_01710_),
    .A1(net740),
    .A2(net274));
 sg13g2_buf_1 _24450_ (.A(net888),
    .X(_06169_));
 sg13g2_nand2_1 _24451_ (.Y(_06170_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][4] ),
    .B(_06161_));
 sg13g2_o21ai_1 _24452_ (.B1(_06170_),
    .Y(_01711_),
    .A1(net739),
    .A2(_06162_));
 sg13g2_buf_1 _24453_ (.A(net887),
    .X(_06171_));
 sg13g2_nand2_1 _24454_ (.Y(_06172_),
    .A(\cpu.genblk1.mmu.r_vtop_i[24][5] ),
    .B(_06161_));
 sg13g2_o21ai_1 _24455_ (.B1(_06172_),
    .Y(_01712_),
    .A1(net738),
    .A2(_06162_));
 sg13g2_buf_1 _24456_ (.A(net999),
    .X(_06173_));
 sg13g2_mux2_1 _24457_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][6] ),
    .S(net274),
    .X(_01713_));
 sg13g2_buf_1 _24458_ (.A(net998),
    .X(_06174_));
 sg13g2_mux2_1 _24459_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][7] ),
    .S(net274),
    .X(_01714_));
 sg13g2_mux2_1 _24460_ (.A0(_06100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][8] ),
    .S(_06161_),
    .X(_01715_));
 sg13g2_mux2_1 _24461_ (.A0(_06101_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[24][9] ),
    .S(_06161_),
    .X(_01716_));
 sg13g2_nand3_1 _24462_ (.B(_06159_),
    .C(_06046_),
    .A(net868),
    .Y(_06175_));
 sg13g2_buf_2 _24463_ (.A(_06175_),
    .X(_06176_));
 sg13g2_buf_1 _24464_ (.A(_06176_),
    .X(_06177_));
 sg13g2_nand2_1 _24465_ (.Y(_06178_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][0] ),
    .B(_06176_));
 sg13g2_o21ai_1 _24466_ (.B1(_06178_),
    .Y(_01717_),
    .A1(_06089_),
    .A2(net315));
 sg13g2_mux2_1 _24467_ (.A0(net504),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][10] ),
    .S(net315),
    .X(_01718_));
 sg13g2_mux2_1 _24468_ (.A0(_06095_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][11] ),
    .S(net315),
    .X(_01719_));
 sg13g2_nand2_1 _24469_ (.Y(_06179_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][1] ),
    .B(_06176_));
 sg13g2_o21ai_1 _24470_ (.B1(_06179_),
    .Y(_01720_),
    .A1(net661),
    .A2(net315));
 sg13g2_mux2_1 _24471_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][2] ),
    .S(net315),
    .X(_01721_));
 sg13g2_nand2_1 _24472_ (.Y(_06180_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][3] ),
    .B(_06176_));
 sg13g2_o21ai_1 _24473_ (.B1(_06180_),
    .Y(_01722_),
    .A1(net740),
    .A2(_06177_));
 sg13g2_nand2_1 _24474_ (.Y(_06181_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][4] ),
    .B(_06176_));
 sg13g2_o21ai_1 _24475_ (.B1(_06181_),
    .Y(_01723_),
    .A1(net739),
    .A2(net315));
 sg13g2_nand2_1 _24476_ (.Y(_06182_),
    .A(\cpu.genblk1.mmu.r_vtop_i[25][5] ),
    .B(_06176_));
 sg13g2_o21ai_1 _24477_ (.B1(_06182_),
    .Y(_01724_),
    .A1(net738),
    .A2(_06177_));
 sg13g2_mux2_1 _24478_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][6] ),
    .S(net315),
    .X(_01725_));
 sg13g2_mux2_1 _24479_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][7] ),
    .S(net315),
    .X(_01726_));
 sg13g2_mux2_1 _24480_ (.A0(_06100_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][8] ),
    .S(_06176_),
    .X(_01727_));
 sg13g2_mux2_1 _24481_ (.A0(_06101_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[25][9] ),
    .S(_06176_),
    .X(_01728_));
 sg13g2_buf_1 _24482_ (.A(net608),
    .X(_06183_));
 sg13g2_nand2_1 _24483_ (.Y(_06184_),
    .A(_05942_),
    .B(net407));
 sg13g2_buf_2 _24484_ (.A(_06184_),
    .X(_06185_));
 sg13g2_buf_1 _24485_ (.A(_06185_),
    .X(_06186_));
 sg13g2_nand2_1 _24486_ (.Y(_06187_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][0] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24487_ (.B1(_06187_),
    .Y(_01729_),
    .A1(net502),
    .A2(net273));
 sg13g2_buf_1 _24488_ (.A(net618),
    .X(_06188_));
 sg13g2_mux2_1 _24489_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][10] ),
    .S(net273),
    .X(_01730_));
 sg13g2_buf_1 _24490_ (.A(net617),
    .X(_06189_));
 sg13g2_mux2_1 _24491_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][11] ),
    .S(net273),
    .X(_01731_));
 sg13g2_nand2_1 _24492_ (.Y(_06190_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][1] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24493_ (.B1(_06190_),
    .Y(_01732_),
    .A1(net661),
    .A2(net273));
 sg13g2_mux2_1 _24494_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][2] ),
    .S(net273),
    .X(_01733_));
 sg13g2_nand2_1 _24495_ (.Y(_06191_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][3] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24496_ (.B1(_06191_),
    .Y(_01734_),
    .A1(net740),
    .A2(_06186_));
 sg13g2_nand2_1 _24497_ (.Y(_06192_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][4] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24498_ (.B1(_06192_),
    .Y(_01735_),
    .A1(net739),
    .A2(net273));
 sg13g2_nand2_1 _24499_ (.Y(_06193_),
    .A(\cpu.genblk1.mmu.r_vtop_i[26][5] ),
    .B(_06185_));
 sg13g2_o21ai_1 _24500_ (.B1(_06193_),
    .Y(_01736_),
    .A1(net738),
    .A2(_06186_));
 sg13g2_mux2_1 _24501_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][6] ),
    .S(net273),
    .X(_01737_));
 sg13g2_mux2_1 _24502_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][7] ),
    .S(net273),
    .X(_01738_));
 sg13g2_buf_1 _24503_ (.A(net537),
    .X(_06194_));
 sg13g2_mux2_1 _24504_ (.A0(_06194_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][8] ),
    .S(_06185_),
    .X(_01739_));
 sg13g2_buf_1 _24505_ (.A(net536),
    .X(_06195_));
 sg13g2_mux2_1 _24506_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[26][9] ),
    .S(_06185_),
    .X(_01740_));
 sg13g2_nand2_1 _24507_ (.Y(_06196_),
    .A(_05948_),
    .B(net407));
 sg13g2_buf_2 _24508_ (.A(_06196_),
    .X(_06197_));
 sg13g2_buf_1 _24509_ (.A(_06197_),
    .X(_06198_));
 sg13g2_nand2_1 _24510_ (.Y(_06199_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][0] ),
    .B(_06197_));
 sg13g2_o21ai_1 _24511_ (.B1(_06199_),
    .Y(_01741_),
    .A1(net502),
    .A2(net272));
 sg13g2_mux2_1 _24512_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][10] ),
    .S(net272),
    .X(_01742_));
 sg13g2_mux2_1 _24513_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][11] ),
    .S(net272),
    .X(_01743_));
 sg13g2_nand2_1 _24514_ (.Y(_06200_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][1] ),
    .B(_06197_));
 sg13g2_o21ai_1 _24515_ (.B1(_06200_),
    .Y(_01744_),
    .A1(net661),
    .A2(_06198_));
 sg13g2_mux2_1 _24516_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][2] ),
    .S(net272),
    .X(_01745_));
 sg13g2_nand2_1 _24517_ (.Y(_06201_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][3] ),
    .B(_06197_));
 sg13g2_o21ai_1 _24518_ (.B1(_06201_),
    .Y(_01746_),
    .A1(net740),
    .A2(net272));
 sg13g2_nand2_1 _24519_ (.Y(_06202_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][4] ),
    .B(_06197_));
 sg13g2_o21ai_1 _24520_ (.B1(_06202_),
    .Y(_01747_),
    .A1(net739),
    .A2(_06198_));
 sg13g2_nand2_1 _24521_ (.Y(_06203_),
    .A(\cpu.genblk1.mmu.r_vtop_i[27][5] ),
    .B(_06197_));
 sg13g2_o21ai_1 _24522_ (.B1(_06203_),
    .Y(_01748_),
    .A1(net738),
    .A2(net272));
 sg13g2_mux2_1 _24523_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][6] ),
    .S(net272),
    .X(_01749_));
 sg13g2_mux2_1 _24524_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][7] ),
    .S(net272),
    .X(_01750_));
 sg13g2_mux2_1 _24525_ (.A0(_06194_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][8] ),
    .S(_06197_),
    .X(_01751_));
 sg13g2_mux2_1 _24526_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[27][9] ),
    .S(_06197_),
    .X(_01752_));
 sg13g2_nor2_2 _24527_ (.A(_05832_),
    .B(_05932_),
    .Y(_06204_));
 sg13g2_nand2_1 _24528_ (.Y(_06205_),
    .A(_06204_),
    .B(_06010_));
 sg13g2_buf_2 _24529_ (.A(_06205_),
    .X(_06206_));
 sg13g2_buf_1 _24530_ (.A(_06206_),
    .X(_06207_));
 sg13g2_nand2_1 _24531_ (.Y(_06208_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][0] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24532_ (.B1(_06208_),
    .Y(_01753_),
    .A1(net502),
    .A2(net238));
 sg13g2_mux2_1 _24533_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][10] ),
    .S(net238),
    .X(_01754_));
 sg13g2_mux2_1 _24534_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][11] ),
    .S(net238),
    .X(_01755_));
 sg13g2_nand2_1 _24535_ (.Y(_06209_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][1] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24536_ (.B1(_06209_),
    .Y(_01756_),
    .A1(net661),
    .A2(net238));
 sg13g2_mux2_1 _24537_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][2] ),
    .S(net238),
    .X(_01757_));
 sg13g2_nand2_1 _24538_ (.Y(_06210_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][3] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24539_ (.B1(_06210_),
    .Y(_01758_),
    .A1(net740),
    .A2(net238));
 sg13g2_nand2_1 _24540_ (.Y(_06211_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][4] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24541_ (.B1(_06211_),
    .Y(_01759_),
    .A1(net739),
    .A2(_06207_));
 sg13g2_nand2_1 _24542_ (.Y(_06212_),
    .A(\cpu.genblk1.mmu.r_vtop_i[28][5] ),
    .B(_06206_));
 sg13g2_o21ai_1 _24543_ (.B1(_06212_),
    .Y(_01760_),
    .A1(net738),
    .A2(_06207_));
 sg13g2_mux2_1 _24544_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][6] ),
    .S(net238),
    .X(_01761_));
 sg13g2_mux2_1 _24545_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][7] ),
    .S(net238),
    .X(_01762_));
 sg13g2_mux2_1 _24546_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][8] ),
    .S(_06206_),
    .X(_01763_));
 sg13g2_mux2_1 _24547_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[28][9] ),
    .S(_06206_),
    .X(_01764_));
 sg13g2_nand2_1 _24548_ (.Y(_06213_),
    .A(_06204_),
    .B(_06046_));
 sg13g2_buf_2 _24549_ (.A(_06213_),
    .X(_06214_));
 sg13g2_buf_1 _24550_ (.A(_06214_),
    .X(_06215_));
 sg13g2_nand2_1 _24551_ (.Y(_06216_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][0] ),
    .B(_06214_));
 sg13g2_o21ai_1 _24552_ (.B1(_06216_),
    .Y(_01765_),
    .A1(net502),
    .A2(net314));
 sg13g2_mux2_1 _24553_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][10] ),
    .S(net314),
    .X(_01766_));
 sg13g2_mux2_1 _24554_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][11] ),
    .S(net314),
    .X(_01767_));
 sg13g2_nand2_1 _24555_ (.Y(_06217_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][1] ),
    .B(_06214_));
 sg13g2_o21ai_1 _24556_ (.B1(_06217_),
    .Y(_01768_),
    .A1(net661),
    .A2(net314));
 sg13g2_mux2_1 _24557_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][2] ),
    .S(net314),
    .X(_01769_));
 sg13g2_nand2_1 _24558_ (.Y(_06218_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][3] ),
    .B(_06214_));
 sg13g2_o21ai_1 _24559_ (.B1(_06218_),
    .Y(_01770_),
    .A1(net740),
    .A2(net314));
 sg13g2_nand2_1 _24560_ (.Y(_06219_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][4] ),
    .B(_06214_));
 sg13g2_o21ai_1 _24561_ (.B1(_06219_),
    .Y(_01771_),
    .A1(net739),
    .A2(_06215_));
 sg13g2_nand2_1 _24562_ (.Y(_06220_),
    .A(\cpu.genblk1.mmu.r_vtop_i[29][5] ),
    .B(_06214_));
 sg13g2_o21ai_1 _24563_ (.B1(_06220_),
    .Y(_01772_),
    .A1(net738),
    .A2(_06215_));
 sg13g2_mux2_1 _24564_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][6] ),
    .S(net314),
    .X(_01773_));
 sg13g2_mux2_1 _24565_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][7] ),
    .S(net314),
    .X(_01774_));
 sg13g2_mux2_1 _24566_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][8] ),
    .S(_06214_),
    .X(_01775_));
 sg13g2_mux2_1 _24567_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[29][9] ),
    .S(_06214_),
    .X(_01776_));
 sg13g2_nand3_1 _24568_ (.B(_06005_),
    .C(net406),
    .A(_06055_),
    .Y(_06221_));
 sg13g2_buf_2 _24569_ (.A(_06221_),
    .X(_06222_));
 sg13g2_buf_1 _24570_ (.A(_06222_),
    .X(_06223_));
 sg13g2_nand2_1 _24571_ (.Y(_06224_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][0] ),
    .B(_06222_));
 sg13g2_o21ai_1 _24572_ (.B1(_06224_),
    .Y(_01777_),
    .A1(net502),
    .A2(net271));
 sg13g2_mux2_1 _24573_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][10] ),
    .S(net271),
    .X(_01778_));
 sg13g2_mux2_1 _24574_ (.A0(_06189_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][11] ),
    .S(net271),
    .X(_01779_));
 sg13g2_nand2_1 _24575_ (.Y(_06225_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][1] ),
    .B(_06222_));
 sg13g2_o21ai_1 _24576_ (.B1(_06225_),
    .Y(_01780_),
    .A1(_06164_),
    .A2(net271));
 sg13g2_mux2_1 _24577_ (.A0(_06166_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][2] ),
    .S(net271),
    .X(_01781_));
 sg13g2_nand2_1 _24578_ (.Y(_06226_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][3] ),
    .B(_06222_));
 sg13g2_o21ai_1 _24579_ (.B1(_06226_),
    .Y(_01782_),
    .A1(net740),
    .A2(net271));
 sg13g2_nand2_1 _24580_ (.Y(_06227_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][4] ),
    .B(_06222_));
 sg13g2_o21ai_1 _24581_ (.B1(_06227_),
    .Y(_01783_),
    .A1(_06169_),
    .A2(_06223_));
 sg13g2_nand2_1 _24582_ (.Y(_06228_),
    .A(\cpu.genblk1.mmu.r_vtop_i[2][5] ),
    .B(_06222_));
 sg13g2_o21ai_1 _24583_ (.B1(_06228_),
    .Y(_01784_),
    .A1(_06171_),
    .A2(_06223_));
 sg13g2_mux2_1 _24584_ (.A0(_06173_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][6] ),
    .S(net271),
    .X(_01785_));
 sg13g2_mux2_1 _24585_ (.A0(_06174_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][7] ),
    .S(net271),
    .X(_01786_));
 sg13g2_mux2_1 _24586_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][8] ),
    .S(_06222_),
    .X(_01787_));
 sg13g2_mux2_1 _24587_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[2][9] ),
    .S(_06222_),
    .X(_01788_));
 sg13g2_nand3_1 _24588_ (.B(_06204_),
    .C(net406),
    .A(_06055_),
    .Y(_06229_));
 sg13g2_buf_2 _24589_ (.A(_06229_),
    .X(_06230_));
 sg13g2_buf_1 _24590_ (.A(_06230_),
    .X(_06231_));
 sg13g2_nand2_1 _24591_ (.Y(_06232_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][0] ),
    .B(_06230_));
 sg13g2_o21ai_1 _24592_ (.B1(_06232_),
    .Y(_01789_),
    .A1(net502),
    .A2(net270));
 sg13g2_mux2_1 _24593_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][10] ),
    .S(net270),
    .X(_01790_));
 sg13g2_mux2_1 _24594_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][11] ),
    .S(net270),
    .X(_01791_));
 sg13g2_nand2_1 _24595_ (.Y(_06233_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][1] ),
    .B(_06230_));
 sg13g2_o21ai_1 _24596_ (.B1(_06233_),
    .Y(_01792_),
    .A1(net661),
    .A2(net270));
 sg13g2_mux2_1 _24597_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][2] ),
    .S(net270),
    .X(_01793_));
 sg13g2_nand2_1 _24598_ (.Y(_06234_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][3] ),
    .B(_06230_));
 sg13g2_o21ai_1 _24599_ (.B1(_06234_),
    .Y(_01794_),
    .A1(_06167_),
    .A2(net270));
 sg13g2_nand2_1 _24600_ (.Y(_06235_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][4] ),
    .B(_06230_));
 sg13g2_o21ai_1 _24601_ (.B1(_06235_),
    .Y(_01795_),
    .A1(net739),
    .A2(_06231_));
 sg13g2_nand2_1 _24602_ (.Y(_06236_),
    .A(\cpu.genblk1.mmu.r_vtop_i[30][5] ),
    .B(_06230_));
 sg13g2_o21ai_1 _24603_ (.B1(_06236_),
    .Y(_01796_),
    .A1(net738),
    .A2(_06231_));
 sg13g2_mux2_1 _24604_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][6] ),
    .S(net270),
    .X(_01797_));
 sg13g2_mux2_1 _24605_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][7] ),
    .S(net270),
    .X(_01798_));
 sg13g2_mux2_1 _24606_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][8] ),
    .S(_06230_),
    .X(_01799_));
 sg13g2_mux2_1 _24607_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[30][9] ),
    .S(_06230_),
    .X(_01800_));
 sg13g2_nand3_1 _24608_ (.B(_06204_),
    .C(net406),
    .A(_05806_),
    .Y(_06237_));
 sg13g2_buf_2 _24609_ (.A(_06237_),
    .X(_06238_));
 sg13g2_buf_1 _24610_ (.A(_06238_),
    .X(_06239_));
 sg13g2_nand2_1 _24611_ (.Y(_06240_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][0] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24612_ (.B1(_06240_),
    .Y(_01801_),
    .A1(net502),
    .A2(net269));
 sg13g2_mux2_1 _24613_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][10] ),
    .S(net269),
    .X(_01802_));
 sg13g2_mux2_1 _24614_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][11] ),
    .S(net269),
    .X(_01803_));
 sg13g2_nand2_1 _24615_ (.Y(_06241_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][1] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24616_ (.B1(_06241_),
    .Y(_01804_),
    .A1(net661),
    .A2(net269));
 sg13g2_mux2_1 _24617_ (.A0(net741),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][2] ),
    .S(net269),
    .X(_01805_));
 sg13g2_nand2_1 _24618_ (.Y(_06242_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][3] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24619_ (.B1(_06242_),
    .Y(_01806_),
    .A1(_06167_),
    .A2(net269));
 sg13g2_nand2_1 _24620_ (.Y(_06243_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][4] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24621_ (.B1(_06243_),
    .Y(_01807_),
    .A1(net739),
    .A2(_06239_));
 sg13g2_nand2_1 _24622_ (.Y(_06244_),
    .A(\cpu.genblk1.mmu.r_vtop_i[31][5] ),
    .B(_06238_));
 sg13g2_o21ai_1 _24623_ (.B1(_06244_),
    .Y(_01808_),
    .A1(net738),
    .A2(_06239_));
 sg13g2_mux2_1 _24624_ (.A0(net858),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][6] ),
    .S(net269),
    .X(_01809_));
 sg13g2_mux2_1 _24625_ (.A0(net857),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][7] ),
    .S(net269),
    .X(_01810_));
 sg13g2_mux2_1 _24626_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][8] ),
    .S(_06238_),
    .X(_01811_));
 sg13g2_mux2_1 _24627_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[31][9] ),
    .S(_06238_),
    .X(_01812_));
 sg13g2_nand3_1 _24628_ (.B(_06005_),
    .C(net406),
    .A(_05806_),
    .Y(_06245_));
 sg13g2_buf_2 _24629_ (.A(_06245_),
    .X(_06246_));
 sg13g2_buf_1 _24630_ (.A(_06246_),
    .X(_06247_));
 sg13g2_nand2_1 _24631_ (.Y(_06248_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][0] ),
    .B(_06246_));
 sg13g2_o21ai_1 _24632_ (.B1(_06248_),
    .Y(_01813_),
    .A1(net502),
    .A2(net268));
 sg13g2_mux2_1 _24633_ (.A0(_06188_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][10] ),
    .S(net268),
    .X(_01814_));
 sg13g2_mux2_1 _24634_ (.A0(_06189_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][11] ),
    .S(net268),
    .X(_01815_));
 sg13g2_nand2_1 _24635_ (.Y(_06249_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][1] ),
    .B(_06246_));
 sg13g2_o21ai_1 _24636_ (.B1(_06249_),
    .Y(_01816_),
    .A1(_06164_),
    .A2(net268));
 sg13g2_mux2_1 _24637_ (.A0(_06166_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][2] ),
    .S(net268),
    .X(_01817_));
 sg13g2_nand2_1 _24638_ (.Y(_06250_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][3] ),
    .B(_06246_));
 sg13g2_o21ai_1 _24639_ (.B1(_06250_),
    .Y(_01818_),
    .A1(net740),
    .A2(net268));
 sg13g2_nand2_1 _24640_ (.Y(_06251_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][4] ),
    .B(_06246_));
 sg13g2_o21ai_1 _24641_ (.B1(_06251_),
    .Y(_01819_),
    .A1(_06169_),
    .A2(_06247_));
 sg13g2_nand2_1 _24642_ (.Y(_06252_),
    .A(\cpu.genblk1.mmu.r_vtop_i[3][5] ),
    .B(_06246_));
 sg13g2_o21ai_1 _24643_ (.B1(_06252_),
    .Y(_01820_),
    .A1(_06171_),
    .A2(_06247_));
 sg13g2_mux2_1 _24644_ (.A0(_06173_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][6] ),
    .S(net268),
    .X(_01821_));
 sg13g2_mux2_1 _24645_ (.A0(_06174_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][7] ),
    .S(net268),
    .X(_01822_));
 sg13g2_mux2_1 _24646_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][8] ),
    .S(_06246_),
    .X(_01823_));
 sg13g2_mux2_1 _24647_ (.A0(net456),
    .A1(\cpu.genblk1.mmu.r_vtop_i[3][9] ),
    .S(_06246_),
    .X(_01824_));
 sg13g2_nand2b_1 _24648_ (.Y(_06253_),
    .B(_06010_),
    .A_N(_05978_));
 sg13g2_buf_2 _24649_ (.A(_06253_),
    .X(_06254_));
 sg13g2_buf_1 _24650_ (.A(_06254_),
    .X(_06255_));
 sg13g2_nand2_1 _24651_ (.Y(_06256_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][0] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24652_ (.B1(_06256_),
    .Y(_01825_),
    .A1(_06183_),
    .A2(net237));
 sg13g2_mux2_1 _24653_ (.A0(net501),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][10] ),
    .S(net237),
    .X(_01826_));
 sg13g2_mux2_1 _24654_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][11] ),
    .S(net237),
    .X(_01827_));
 sg13g2_nand2_1 _24655_ (.Y(_06257_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][1] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24656_ (.B1(_06257_),
    .Y(_01828_),
    .A1(net755),
    .A2(net237));
 sg13g2_mux2_1 _24657_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][2] ),
    .S(net237),
    .X(_01829_));
 sg13g2_nand2_1 _24658_ (.Y(_06258_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][3] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24659_ (.B1(_06258_),
    .Y(_01830_),
    .A1(net889),
    .A2(net237));
 sg13g2_nand2_1 _24660_ (.Y(_06259_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][4] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24661_ (.B1(_06259_),
    .Y(_01831_),
    .A1(net888),
    .A2(net237));
 sg13g2_nand2_1 _24662_ (.Y(_06260_),
    .A(\cpu.genblk1.mmu.r_vtop_i[4][5] ),
    .B(_06254_));
 sg13g2_o21ai_1 _24663_ (.B1(_06260_),
    .Y(_01832_),
    .A1(net887),
    .A2(net237));
 sg13g2_mux2_1 _24664_ (.A0(_03083_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][6] ),
    .S(_06255_),
    .X(_01833_));
 sg13g2_mux2_1 _24665_ (.A0(net880),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][7] ),
    .S(_06255_),
    .X(_01834_));
 sg13g2_mux2_1 _24666_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][8] ),
    .S(_06254_),
    .X(_01835_));
 sg13g2_mux2_1 _24667_ (.A0(_06195_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[4][9] ),
    .S(_06254_),
    .X(_01836_));
 sg13g2_nand2_1 _24668_ (.Y(_06261_),
    .A(_05983_),
    .B(net407));
 sg13g2_buf_2 _24669_ (.A(_06261_),
    .X(_06262_));
 sg13g2_buf_1 _24670_ (.A(_06262_),
    .X(_06263_));
 sg13g2_nand2_1 _24671_ (.Y(_06264_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][0] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24672_ (.B1(_06264_),
    .Y(_01837_),
    .A1(_06183_),
    .A2(net267));
 sg13g2_mux2_1 _24673_ (.A0(_06188_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][10] ),
    .S(net267),
    .X(_01838_));
 sg13g2_mux2_1 _24674_ (.A0(net500),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][11] ),
    .S(net267),
    .X(_01839_));
 sg13g2_nand2_1 _24675_ (.Y(_06265_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][1] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24676_ (.B1(_06265_),
    .Y(_01840_),
    .A1(net755),
    .A2(net267));
 sg13g2_mux2_1 _24677_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][2] ),
    .S(net267),
    .X(_01841_));
 sg13g2_nand2_1 _24678_ (.Y(_06266_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][3] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24679_ (.B1(_06266_),
    .Y(_01842_),
    .A1(net889),
    .A2(net267));
 sg13g2_nand2_1 _24680_ (.Y(_06267_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][4] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24681_ (.B1(_06267_),
    .Y(_01843_),
    .A1(net888),
    .A2(net267));
 sg13g2_nand2_1 _24682_ (.Y(_06268_),
    .A(\cpu.genblk1.mmu.r_vtop_i[5][5] ),
    .B(_06262_));
 sg13g2_o21ai_1 _24683_ (.B1(_06268_),
    .Y(_01844_),
    .A1(net887),
    .A2(net267));
 sg13g2_mux2_1 _24684_ (.A0(net881),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][6] ),
    .S(_06263_),
    .X(_01845_));
 sg13g2_mux2_1 _24685_ (.A0(net880),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][7] ),
    .S(_06263_),
    .X(_01846_));
 sg13g2_mux2_1 _24686_ (.A0(net457),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][8] ),
    .S(_06262_),
    .X(_01847_));
 sg13g2_mux2_1 _24687_ (.A0(_06195_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[5][9] ),
    .S(_06262_),
    .X(_01848_));
 sg13g2_nand2_1 _24688_ (.Y(_06269_),
    .A(_05989_),
    .B(net407));
 sg13g2_buf_2 _24689_ (.A(_06269_),
    .X(_06270_));
 sg13g2_buf_1 _24690_ (.A(_06270_),
    .X(_06271_));
 sg13g2_nand2_1 _24691_ (.Y(_06272_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][0] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24692_ (.B1(_06272_),
    .Y(_01849_),
    .A1(net608),
    .A2(net266));
 sg13g2_mux2_1 _24693_ (.A0(net535),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][10] ),
    .S(net266),
    .X(_01850_));
 sg13g2_mux2_1 _24694_ (.A0(net534),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][11] ),
    .S(net266),
    .X(_01851_));
 sg13g2_nand2_1 _24695_ (.Y(_06273_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][1] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24696_ (.B1(_06273_),
    .Y(_01852_),
    .A1(net755),
    .A2(net266));
 sg13g2_mux2_1 _24697_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][2] ),
    .S(net266),
    .X(_01853_));
 sg13g2_nand2_1 _24698_ (.Y(_06274_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][3] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24699_ (.B1(_06274_),
    .Y(_01854_),
    .A1(net889),
    .A2(net266));
 sg13g2_nand2_1 _24700_ (.Y(_06275_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][4] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24701_ (.B1(_06275_),
    .Y(_01855_),
    .A1(_03062_),
    .A2(_06271_));
 sg13g2_nand2_1 _24702_ (.Y(_06276_),
    .A(\cpu.genblk1.mmu.r_vtop_i[6][5] ),
    .B(_06270_));
 sg13g2_o21ai_1 _24703_ (.B1(_06276_),
    .Y(_01856_),
    .A1(net887),
    .A2(net266));
 sg13g2_mux2_1 _24704_ (.A0(net881),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][6] ),
    .S(net266),
    .X(_01857_));
 sg13g2_mux2_1 _24705_ (.A0(net880),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][7] ),
    .S(_06271_),
    .X(_01858_));
 sg13g2_mux2_1 _24706_ (.A0(net468),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][8] ),
    .S(_06270_),
    .X(_01859_));
 sg13g2_mux2_1 _24707_ (.A0(net471),
    .A1(\cpu.genblk1.mmu.r_vtop_i[6][9] ),
    .S(_06270_),
    .X(_01860_));
 sg13g2_nand2_1 _24708_ (.Y(_06277_),
    .A(_05994_),
    .B(_06019_));
 sg13g2_buf_2 _24709_ (.A(_06277_),
    .X(_06278_));
 sg13g2_buf_1 _24710_ (.A(_06278_),
    .X(_06279_));
 sg13g2_nand2_1 _24711_ (.Y(_06280_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][0] ),
    .B(_06278_));
 sg13g2_o21ai_1 _24712_ (.B1(_06280_),
    .Y(_01861_),
    .A1(net608),
    .A2(net265));
 sg13g2_mux2_1 _24713_ (.A0(net535),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][10] ),
    .S(net265),
    .X(_01862_));
 sg13g2_mux2_1 _24714_ (.A0(net534),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][11] ),
    .S(net265),
    .X(_01863_));
 sg13g2_nand2_1 _24715_ (.Y(_06281_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][1] ),
    .B(_06278_));
 sg13g2_o21ai_1 _24716_ (.B1(_06281_),
    .Y(_01864_),
    .A1(net755),
    .A2(net265));
 sg13g2_mux2_1 _24717_ (.A0(net750),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][2] ),
    .S(net265),
    .X(_01865_));
 sg13g2_nand2_1 _24718_ (.Y(_06282_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][3] ),
    .B(_06278_));
 sg13g2_o21ai_1 _24719_ (.B1(_06282_),
    .Y(_01866_),
    .A1(net889),
    .A2(net265));
 sg13g2_nand2_1 _24720_ (.Y(_06283_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][4] ),
    .B(_06278_));
 sg13g2_o21ai_1 _24721_ (.B1(_06283_),
    .Y(_01867_),
    .A1(_03062_),
    .A2(_06279_));
 sg13g2_nand2_1 _24722_ (.Y(_06284_),
    .A(\cpu.genblk1.mmu.r_vtop_i[7][5] ),
    .B(_06278_));
 sg13g2_o21ai_1 _24723_ (.B1(_06284_),
    .Y(_01868_),
    .A1(_03065_),
    .A2(net265));
 sg13g2_mux2_1 _24724_ (.A0(net881),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][6] ),
    .S(net265),
    .X(_01869_));
 sg13g2_mux2_1 _24725_ (.A0(net880),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][7] ),
    .S(_06279_),
    .X(_01870_));
 sg13g2_mux2_1 _24726_ (.A0(net468),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][8] ),
    .S(_06278_),
    .X(_01871_));
 sg13g2_mux2_1 _24727_ (.A0(net471),
    .A1(\cpu.genblk1.mmu.r_vtop_i[7][9] ),
    .S(_06278_),
    .X(_01872_));
 sg13g2_nand3_1 _24728_ (.B(_06080_),
    .C(_06064_),
    .A(_05861_),
    .Y(_06285_));
 sg13g2_buf_2 _24729_ (.A(_06285_),
    .X(_06286_));
 sg13g2_buf_1 _24730_ (.A(_06286_),
    .X(_06287_));
 sg13g2_nand2_1 _24731_ (.Y(_06288_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][0] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24732_ (.B1(_06288_),
    .Y(_01873_),
    .A1(net608),
    .A2(net264));
 sg13g2_mux2_1 _24733_ (.A0(net535),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][10] ),
    .S(_06287_),
    .X(_01874_));
 sg13g2_mux2_1 _24734_ (.A0(net534),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][11] ),
    .S(net264),
    .X(_01875_));
 sg13g2_nand2_1 _24735_ (.Y(_06289_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][1] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24736_ (.B1(_06289_),
    .Y(_01876_),
    .A1(net755),
    .A2(net264));
 sg13g2_mux2_1 _24737_ (.A0(_03075_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][2] ),
    .S(net264),
    .X(_01877_));
 sg13g2_nand2_1 _24738_ (.Y(_06290_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][3] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24739_ (.B1(_06290_),
    .Y(_01878_),
    .A1(_03059_),
    .A2(net264));
 sg13g2_nand2_1 _24740_ (.Y(_06291_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][4] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24741_ (.B1(_06291_),
    .Y(_01879_),
    .A1(net888),
    .A2(net264));
 sg13g2_nand2_1 _24742_ (.Y(_06292_),
    .A(\cpu.genblk1.mmu.r_vtop_i[8][5] ),
    .B(_06286_));
 sg13g2_o21ai_1 _24743_ (.B1(_06292_),
    .Y(_01880_),
    .A1(net887),
    .A2(net264));
 sg13g2_mux2_1 _24744_ (.A0(_03083_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][6] ),
    .S(net264),
    .X(_01881_));
 sg13g2_mux2_1 _24745_ (.A0(_03084_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][7] ),
    .S(_06287_),
    .X(_01882_));
 sg13g2_mux2_1 _24746_ (.A0(net468),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][8] ),
    .S(_06286_),
    .X(_01883_));
 sg13g2_mux2_1 _24747_ (.A0(net471),
    .A1(\cpu.genblk1.mmu.r_vtop_i[8][9] ),
    .S(_06286_),
    .X(_01884_));
 sg13g2_nand3_1 _24748_ (.B(_05861_),
    .C(_06046_),
    .A(net868),
    .Y(_06293_));
 sg13g2_buf_2 _24749_ (.A(_06293_),
    .X(_06294_));
 sg13g2_buf_1 _24750_ (.A(_06294_),
    .X(_06295_));
 sg13g2_nand2_1 _24751_ (.Y(_06296_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][0] ),
    .B(_06294_));
 sg13g2_o21ai_1 _24752_ (.B1(_06296_),
    .Y(_01885_),
    .A1(net608),
    .A2(net313));
 sg13g2_mux2_1 _24753_ (.A0(net535),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][10] ),
    .S(_06295_),
    .X(_01886_));
 sg13g2_mux2_1 _24754_ (.A0(net534),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][11] ),
    .S(net313),
    .X(_01887_));
 sg13g2_nand2_1 _24755_ (.Y(_06297_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][1] ),
    .B(_06294_));
 sg13g2_o21ai_1 _24756_ (.B1(_06297_),
    .Y(_01888_),
    .A1(net755),
    .A2(net313));
 sg13g2_mux2_1 _24757_ (.A0(_03075_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][2] ),
    .S(net313),
    .X(_01889_));
 sg13g2_nand2_1 _24758_ (.Y(_06298_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][3] ),
    .B(_06294_));
 sg13g2_o21ai_1 _24759_ (.B1(_06298_),
    .Y(_01890_),
    .A1(net889),
    .A2(net313));
 sg13g2_nand2_1 _24760_ (.Y(_06299_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][4] ),
    .B(_06294_));
 sg13g2_o21ai_1 _24761_ (.B1(_06299_),
    .Y(_01891_),
    .A1(net888),
    .A2(net313));
 sg13g2_nand2_1 _24762_ (.Y(_06300_),
    .A(\cpu.genblk1.mmu.r_vtop_i[9][5] ),
    .B(_06294_));
 sg13g2_o21ai_1 _24763_ (.B1(_06300_),
    .Y(_01892_),
    .A1(net887),
    .A2(net313));
 sg13g2_mux2_1 _24764_ (.A0(net881),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][6] ),
    .S(net313),
    .X(_01893_));
 sg13g2_mux2_1 _24765_ (.A0(_03084_),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][7] ),
    .S(_06295_),
    .X(_01894_));
 sg13g2_mux2_1 _24766_ (.A0(net468),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][8] ),
    .S(_06294_),
    .X(_01895_));
 sg13g2_mux2_1 _24767_ (.A0(net471),
    .A1(\cpu.genblk1.mmu.r_vtop_i[9][9] ),
    .S(_06294_),
    .X(_01896_));
 sg13g2_mux2_1 _24768_ (.A0(\cpu.genblk1.mmu.r_writeable_d[0] ),
    .A1(_03621_),
    .S(_05840_),
    .X(_01897_));
 sg13g2_buf_1 _24769_ (.A(net533),
    .X(_06301_));
 sg13g2_mux2_1 _24770_ (.A0(\cpu.genblk1.mmu.r_writeable_d[10] ),
    .A1(net455),
    .S(_05853_),
    .X(_01898_));
 sg13g2_mux2_1 _24771_ (.A0(\cpu.genblk1.mmu.r_writeable_d[11] ),
    .A1(net455),
    .S(_05859_),
    .X(_01899_));
 sg13g2_mux2_1 _24772_ (.A0(\cpu.genblk1.mmu.r_writeable_d[12] ),
    .A1(net455),
    .S(_05865_),
    .X(_01900_));
 sg13g2_mux2_1 _24773_ (.A0(\cpu.genblk1.mmu.r_writeable_d[13] ),
    .A1(net455),
    .S(_05871_),
    .X(_01901_));
 sg13g2_mux2_1 _24774_ (.A0(\cpu.genblk1.mmu.r_writeable_d[14] ),
    .A1(_06301_),
    .S(_05875_),
    .X(_01902_));
 sg13g2_mux2_1 _24775_ (.A0(\cpu.genblk1.mmu.r_writeable_d[15] ),
    .A1(_06301_),
    .S(_05880_),
    .X(_01903_));
 sg13g2_mux2_1 _24776_ (.A0(\cpu.genblk1.mmu.r_writeable_d[16] ),
    .A1(net455),
    .S(_05887_),
    .X(_01904_));
 sg13g2_mux2_1 _24777_ (.A0(\cpu.genblk1.mmu.r_writeable_d[17] ),
    .A1(net455),
    .S(_05892_),
    .X(_01905_));
 sg13g2_mux2_1 _24778_ (.A0(\cpu.genblk1.mmu.r_writeable_d[18] ),
    .A1(net455),
    .S(_05899_),
    .X(_01906_));
 sg13g2_mux2_1 _24779_ (.A0(\cpu.genblk1.mmu.r_writeable_d[19] ),
    .A1(net455),
    .S(_05908_),
    .X(_01907_));
 sg13g2_buf_1 _24780_ (.A(net533),
    .X(_06302_));
 sg13g2_mux2_1 _24781_ (.A0(\cpu.genblk1.mmu.r_writeable_d[1] ),
    .A1(_06302_),
    .S(_05912_),
    .X(_01908_));
 sg13g2_mux2_1 _24782_ (.A0(\cpu.genblk1.mmu.r_writeable_d[20] ),
    .A1(net454),
    .S(_05918_),
    .X(_01909_));
 sg13g2_mux2_1 _24783_ (.A0(\cpu.genblk1.mmu.r_writeable_d[21] ),
    .A1(net454),
    .S(_05921_),
    .X(_01910_));
 sg13g2_mux2_1 _24784_ (.A0(\cpu.genblk1.mmu.r_writeable_d[22] ),
    .A1(net454),
    .S(_05924_),
    .X(_01911_));
 sg13g2_mux2_1 _24785_ (.A0(\cpu.genblk1.mmu.r_writeable_d[23] ),
    .A1(net454),
    .S(_05927_),
    .X(_01912_));
 sg13g2_mux2_1 _24786_ (.A0(\cpu.genblk1.mmu.r_writeable_d[24] ),
    .A1(net454),
    .S(_05934_),
    .X(_01913_));
 sg13g2_mux2_1 _24787_ (.A0(\cpu.genblk1.mmu.r_writeable_d[25] ),
    .A1(net454),
    .S(_05938_),
    .X(_01914_));
 sg13g2_mux2_1 _24788_ (.A0(\cpu.genblk1.mmu.r_writeable_d[26] ),
    .A1(net454),
    .S(_05944_),
    .X(_01915_));
 sg13g2_mux2_1 _24789_ (.A0(\cpu.genblk1.mmu.r_writeable_d[27] ),
    .A1(net454),
    .S(_05950_),
    .X(_01916_));
 sg13g2_mux2_1 _24790_ (.A0(\cpu.genblk1.mmu.r_writeable_d[28] ),
    .A1(_06302_),
    .S(_05959_),
    .X(_01917_));
 sg13g2_buf_1 _24791_ (.A(net533),
    .X(_06303_));
 sg13g2_mux2_1 _24792_ (.A0(\cpu.genblk1.mmu.r_writeable_d[29] ),
    .A1(net453),
    .S(_05963_),
    .X(_01918_));
 sg13g2_mux2_1 _24793_ (.A0(\cpu.genblk1.mmu.r_writeable_d[2] ),
    .A1(_06303_),
    .S(_05967_),
    .X(_01919_));
 sg13g2_mux2_1 _24794_ (.A0(\cpu.genblk1.mmu.r_writeable_d[30] ),
    .A1(net453),
    .S(_05970_),
    .X(_01920_));
 sg13g2_mux2_1 _24795_ (.A0(\cpu.genblk1.mmu.r_writeable_d[31] ),
    .A1(net453),
    .S(_05973_),
    .X(_01921_));
 sg13g2_mux2_1 _24796_ (.A0(\cpu.genblk1.mmu.r_writeable_d[3] ),
    .A1(net453),
    .S(_05976_),
    .X(_01922_));
 sg13g2_mux2_1 _24797_ (.A0(\cpu.genblk1.mmu.r_writeable_d[4] ),
    .A1(net453),
    .S(_05980_),
    .X(_01923_));
 sg13g2_mux2_1 _24798_ (.A0(\cpu.genblk1.mmu.r_writeable_d[5] ),
    .A1(net453),
    .S(_05985_),
    .X(_01924_));
 sg13g2_mux2_1 _24799_ (.A0(\cpu.genblk1.mmu.r_writeable_d[6] ),
    .A1(net453),
    .S(_05991_),
    .X(_01925_));
 sg13g2_mux2_1 _24800_ (.A0(\cpu.genblk1.mmu.r_writeable_d[7] ),
    .A1(net453),
    .S(_05996_),
    .X(_01926_));
 sg13g2_mux2_1 _24801_ (.A0(\cpu.genblk1.mmu.r_writeable_d[8] ),
    .A1(_06303_),
    .S(_05999_),
    .X(_01927_));
 sg13g2_mux2_1 _24802_ (.A0(\cpu.genblk1.mmu.r_writeable_d[9] ),
    .A1(_03620_),
    .S(_06002_),
    .X(_01928_));
 sg13g2_buf_1 _24803_ (.A(net1057),
    .X(_06304_));
 sg13g2_nor2b_1 _24804_ (.A(net1000),
    .B_N(_09195_),
    .Y(_06305_));
 sg13g2_and3_1 _24805_ (.X(_06306_),
    .A(net1154),
    .B(_00227_),
    .C(_06305_));
 sg13g2_buf_1 _24806_ (.A(_06306_),
    .X(_06307_));
 sg13g2_and2_1 _24807_ (.A(net1071),
    .B(_06307_),
    .X(_06308_));
 sg13g2_buf_2 _24808_ (.A(_06308_),
    .X(_06309_));
 sg13g2_nand3_1 _24809_ (.B(net340),
    .C(_06309_),
    .A(net869),
    .Y(_06310_));
 sg13g2_buf_2 _24810_ (.A(_06310_),
    .X(_06311_));
 sg13g2_mux2_1 _24811_ (.A0(net856),
    .A1(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .S(_06311_),
    .X(_01945_));
 sg13g2_nand2_1 _24812_ (.Y(_06312_),
    .A(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .B(_06311_));
 sg13g2_o21ai_1 _24813_ (.B1(_06312_),
    .Y(_01946_),
    .A1(net892),
    .A2(_06311_));
 sg13g2_nand2_1 _24814_ (.Y(_06313_),
    .A(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .B(_06311_));
 sg13g2_o21ai_1 _24815_ (.B1(_06313_),
    .Y(_01947_),
    .A1(net757),
    .A2(_06311_));
 sg13g2_nand2_1 _24816_ (.Y(_06314_),
    .A(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .B(_06311_));
 sg13g2_o21ai_1 _24817_ (.B1(_06314_),
    .Y(_01948_),
    .A1(net891),
    .A2(_06311_));
 sg13g2_nand3_1 _24818_ (.B(net374),
    .C(_06309_),
    .A(net869),
    .Y(_06315_));
 sg13g2_buf_2 _24819_ (.A(_06315_),
    .X(_06316_));
 sg13g2_mux2_1 _24820_ (.A0(net981),
    .A1(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .S(_06316_),
    .X(_01949_));
 sg13g2_mux2_1 _24821_ (.A0(net856),
    .A1(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .S(_06316_),
    .X(_01950_));
 sg13g2_nand2_1 _24822_ (.Y(_06317_),
    .A(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .B(_06316_));
 sg13g2_o21ai_1 _24823_ (.B1(_06317_),
    .Y(_01951_),
    .A1(_02743_),
    .A2(_06316_));
 sg13g2_nand2_1 _24824_ (.Y(_06318_),
    .A(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .B(_06316_));
 sg13g2_o21ai_1 _24825_ (.B1(_06318_),
    .Y(_01952_),
    .A1(net757),
    .A2(_06316_));
 sg13g2_nand2_1 _24826_ (.Y(_06319_),
    .A(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .B(_06316_));
 sg13g2_o21ai_1 _24827_ (.B1(_06319_),
    .Y(_01953_),
    .A1(_02749_),
    .A2(_06316_));
 sg13g2_nand2_1 _24828_ (.Y(_06320_),
    .A(_04849_),
    .B(_06309_));
 sg13g2_buf_1 _24829_ (.A(_06320_),
    .X(_06321_));
 sg13g2_buf_1 _24830_ (.A(_06321_),
    .X(_06322_));
 sg13g2_nand2_1 _24831_ (.Y(_06323_),
    .A(_04850_),
    .B(_06322_));
 sg13g2_o21ai_1 _24832_ (.B1(_06323_),
    .Y(_01954_),
    .A1(net761),
    .A2(_06322_));
 sg13g2_buf_1 _24833_ (.A(\cpu.gpio.r_spi_miso_src[0][1] ),
    .X(_06324_));
 sg13g2_nand2_1 _24834_ (.Y(_06325_),
    .A(_06324_),
    .B(net80));
 sg13g2_o21ai_1 _24835_ (.B1(_06325_),
    .Y(_01955_),
    .A1(net759),
    .A2(net80));
 sg13g2_nand2_1 _24836_ (.Y(_06326_),
    .A(\cpu.gpio.r_spi_miso_src[0][2] ),
    .B(_06321_));
 sg13g2_o21ai_1 _24837_ (.B1(_06326_),
    .Y(_01956_),
    .A1(net758),
    .A2(net80));
 sg13g2_buf_1 _24838_ (.A(\cpu.gpio.r_spi_miso_src[0][3] ),
    .X(_06327_));
 sg13g2_mux2_1 _24839_ (.A0(net981),
    .A1(_06327_),
    .S(net80),
    .X(_01957_));
 sg13g2_mux2_1 _24840_ (.A0(net856),
    .A1(_05554_),
    .S(net80),
    .X(_01958_));
 sg13g2_nand2_1 _24841_ (.Y(_06328_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B(_06321_));
 sg13g2_o21ai_1 _24842_ (.B1(_06328_),
    .Y(_01959_),
    .A1(_02743_),
    .A2(net80));
 sg13g2_nand2_1 _24843_ (.Y(_06329_),
    .A(\cpu.gpio.r_spi_miso_src[1][2] ),
    .B(_06321_));
 sg13g2_o21ai_1 _24844_ (.B1(_06329_),
    .Y(_01960_),
    .A1(_02746_),
    .A2(net80));
 sg13g2_buf_1 _24845_ (.A(\cpu.gpio.r_spi_miso_src[1][3] ),
    .X(_06330_));
 sg13g2_nand2_1 _24846_ (.Y(_06331_),
    .A(_06330_),
    .B(_06321_));
 sg13g2_o21ai_1 _24847_ (.B1(_06331_),
    .Y(_01961_),
    .A1(net891),
    .A2(net80));
 sg13g2_nand2_1 _24848_ (.Y(_06332_),
    .A(net413),
    .B(_06309_));
 sg13g2_buf_1 _24849_ (.A(_06332_),
    .X(_06333_));
 sg13g2_buf_1 _24850_ (.A(_06333_),
    .X(_06334_));
 sg13g2_nand2_1 _24851_ (.Y(_06335_),
    .A(_04872_),
    .B(_06334_));
 sg13g2_o21ai_1 _24852_ (.B1(_06335_),
    .Y(_01962_),
    .A1(_12703_),
    .A2(_06334_));
 sg13g2_nand2_1 _24853_ (.Y(_06336_),
    .A(_05341_),
    .B(net79));
 sg13g2_o21ai_1 _24854_ (.B1(_06336_),
    .Y(_01963_),
    .A1(_02727_),
    .A2(net79));
 sg13g2_nand2_1 _24855_ (.Y(_06337_),
    .A(_05421_),
    .B(_06333_));
 sg13g2_o21ai_1 _24856_ (.B1(_06337_),
    .Y(_01964_),
    .A1(_02730_),
    .A2(net79));
 sg13g2_mux2_1 _24857_ (.A0(net981),
    .A1(_05482_),
    .S(net79),
    .X(_01965_));
 sg13g2_mux2_1 _24858_ (.A0(net856),
    .A1(_05558_),
    .S(net79),
    .X(_01966_));
 sg13g2_nand2_1 _24859_ (.Y(_06338_),
    .A(_05622_),
    .B(_06333_));
 sg13g2_o21ai_1 _24860_ (.B1(_06338_),
    .Y(_01967_),
    .A1(net895),
    .A2(net79));
 sg13g2_nand2_1 _24861_ (.Y(_06339_),
    .A(_05664_),
    .B(_06333_));
 sg13g2_o21ai_1 _24862_ (.B1(_06339_),
    .Y(_01968_),
    .A1(_02746_),
    .A2(net79));
 sg13g2_nand2_1 _24863_ (.Y(_06340_),
    .A(_05078_),
    .B(_06333_));
 sg13g2_o21ai_1 _24864_ (.B1(_06340_),
    .Y(_01969_),
    .A1(net893),
    .A2(net79));
 sg13g2_nand2_1 _24865_ (.Y(_06341_),
    .A(_04869_),
    .B(_06309_));
 sg13g2_buf_1 _24866_ (.A(_06341_),
    .X(_06342_));
 sg13g2_buf_1 _24867_ (.A(_06342_),
    .X(_06343_));
 sg13g2_nand2_1 _24868_ (.Y(_06344_),
    .A(_04865_),
    .B(net78));
 sg13g2_o21ai_1 _24869_ (.B1(_06344_),
    .Y(_01970_),
    .A1(net922),
    .A2(net78));
 sg13g2_buf_1 _24870_ (.A(\cpu.gpio.r_src_io[6][1] ),
    .X(_06345_));
 sg13g2_nand2_1 _24871_ (.Y(_06346_),
    .A(_06345_),
    .B(net78));
 sg13g2_o21ai_1 _24872_ (.B1(_06346_),
    .Y(_01971_),
    .A1(_02727_),
    .A2(net78));
 sg13g2_nand2_1 _24873_ (.Y(_06347_),
    .A(\cpu.gpio.r_src_io[6][2] ),
    .B(_06342_));
 sg13g2_o21ai_1 _24874_ (.B1(_06347_),
    .Y(_01972_),
    .A1(_02730_),
    .A2(_06343_));
 sg13g2_mux2_1 _24875_ (.A0(_05781_),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .S(net78),
    .X(_01973_));
 sg13g2_mux2_1 _24876_ (.A0(net856),
    .A1(_05557_),
    .S(net78),
    .X(_01974_));
 sg13g2_buf_1 _24877_ (.A(\cpu.gpio.r_src_io[7][1] ),
    .X(_06348_));
 sg13g2_nand2_1 _24878_ (.Y(_06349_),
    .A(_06348_),
    .B(_06342_));
 sg13g2_o21ai_1 _24879_ (.B1(_06349_),
    .Y(_01975_),
    .A1(net895),
    .A2(_06343_));
 sg13g2_nand2_1 _24880_ (.Y(_06350_),
    .A(\cpu.gpio.r_src_io[7][2] ),
    .B(_06342_));
 sg13g2_o21ai_1 _24881_ (.B1(_06350_),
    .Y(_01976_),
    .A1(net894),
    .A2(net78));
 sg13g2_nand2_1 _24882_ (.Y(_06351_),
    .A(\cpu.gpio.r_src_io[7][3] ),
    .B(_06342_));
 sg13g2_o21ai_1 _24883_ (.B1(_06351_),
    .Y(_01977_),
    .A1(net893),
    .A2(net78));
 sg13g2_nand2b_1 _24884_ (.Y(_06352_),
    .B(_06309_),
    .A_N(_05620_));
 sg13g2_buf_2 _24885_ (.A(_06352_),
    .X(_06353_));
 sg13g2_mux2_1 _24886_ (.A0(net856),
    .A1(_05567_),
    .S(_06353_),
    .X(_01978_));
 sg13g2_buf_1 _24887_ (.A(\cpu.gpio.r_src_o[3][1] ),
    .X(_06354_));
 sg13g2_nand2_1 _24888_ (.Y(_06355_),
    .A(_06354_),
    .B(_06353_));
 sg13g2_o21ai_1 _24889_ (.B1(_06355_),
    .Y(_01979_),
    .A1(net895),
    .A2(_06353_));
 sg13g2_nand2_1 _24890_ (.Y(_06356_),
    .A(\cpu.gpio.r_src_o[3][2] ),
    .B(_06353_));
 sg13g2_o21ai_1 _24891_ (.B1(_06356_),
    .Y(_01980_),
    .A1(net894),
    .A2(_06353_));
 sg13g2_nand2_1 _24892_ (.Y(_06357_),
    .A(\cpu.gpio.r_src_o[3][3] ),
    .B(_06353_));
 sg13g2_o21ai_1 _24893_ (.B1(_06357_),
    .Y(_01981_),
    .A1(net893),
    .A2(_06353_));
 sg13g2_nand2_1 _24894_ (.Y(_06358_),
    .A(_04863_),
    .B(_06309_));
 sg13g2_buf_1 _24895_ (.A(_06358_),
    .X(_06359_));
 sg13g2_buf_1 _24896_ (.A(_06359_),
    .X(_06360_));
 sg13g2_nand2_1 _24897_ (.Y(_06361_),
    .A(_04858_),
    .B(net77));
 sg13g2_o21ai_1 _24898_ (.B1(_06361_),
    .Y(_01982_),
    .A1(net922),
    .A2(net77));
 sg13g2_buf_1 _24899_ (.A(\cpu.gpio.r_src_o[4][1] ),
    .X(_06362_));
 sg13g2_nand2_1 _24900_ (.Y(_06363_),
    .A(_06362_),
    .B(net77));
 sg13g2_o21ai_1 _24901_ (.B1(_06363_),
    .Y(_01983_),
    .A1(net897),
    .A2(net77));
 sg13g2_nand2_1 _24902_ (.Y(_06364_),
    .A(\cpu.gpio.r_src_o[4][2] ),
    .B(_06359_));
 sg13g2_o21ai_1 _24903_ (.B1(_06364_),
    .Y(_01984_),
    .A1(net896),
    .A2(net77));
 sg13g2_mux2_1 _24904_ (.A0(net981),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .S(net77),
    .X(_01985_));
 sg13g2_mux2_1 _24905_ (.A0(_06304_),
    .A1(_05561_),
    .S(net77),
    .X(_01986_));
 sg13g2_buf_1 _24906_ (.A(\cpu.gpio.r_src_o[5][1] ),
    .X(_06365_));
 sg13g2_nand2_1 _24907_ (.Y(_06366_),
    .A(_06365_),
    .B(_06359_));
 sg13g2_o21ai_1 _24908_ (.B1(_06366_),
    .Y(_01987_),
    .A1(net895),
    .A2(_06360_));
 sg13g2_nand2_1 _24909_ (.Y(_06367_),
    .A(\cpu.gpio.r_src_o[5][2] ),
    .B(_06359_));
 sg13g2_o21ai_1 _24910_ (.B1(_06367_),
    .Y(_01988_),
    .A1(net894),
    .A2(net77));
 sg13g2_nand2_1 _24911_ (.Y(_06368_),
    .A(\cpu.gpio.r_src_o[5][3] ),
    .B(_06359_));
 sg13g2_o21ai_1 _24912_ (.B1(_06368_),
    .Y(_01989_),
    .A1(net893),
    .A2(_06360_));
 sg13g2_nand2b_1 _24913_ (.Y(_06369_),
    .B(_06309_),
    .A_N(_05340_));
 sg13g2_buf_2 _24914_ (.A(_06369_),
    .X(_06370_));
 sg13g2_mux2_1 _24915_ (.A0(_06304_),
    .A1(_05559_),
    .S(_06370_),
    .X(_01994_));
 sg13g2_buf_1 _24916_ (.A(\cpu.gpio.r_src_o[7][1] ),
    .X(_06371_));
 sg13g2_nand2_1 _24917_ (.Y(_06372_),
    .A(_06371_),
    .B(_06370_));
 sg13g2_o21ai_1 _24918_ (.B1(_06372_),
    .Y(_01995_),
    .A1(_12261_),
    .A2(_06370_));
 sg13g2_nand2_1 _24919_ (.Y(_06373_),
    .A(\cpu.gpio.r_src_o[7][2] ),
    .B(_06370_));
 sg13g2_o21ai_1 _24920_ (.B1(_06373_),
    .Y(_01996_),
    .A1(_12265_),
    .A2(_06370_));
 sg13g2_nand2_1 _24921_ (.Y(_06374_),
    .A(\cpu.gpio.r_src_o[7][3] ),
    .B(_06370_));
 sg13g2_o21ai_1 _24922_ (.B1(_06374_),
    .Y(_01997_),
    .A1(net893),
    .A2(_06370_));
 sg13g2_buf_1 _24923_ (.A(net1002),
    .X(_06375_));
 sg13g2_and2_1 _24924_ (.A(net719),
    .B(_08572_),
    .X(_06376_));
 sg13g2_buf_4 _24925_ (.X(_06377_),
    .A(_06376_));
 sg13g2_buf_1 _24926_ (.A(_00245_),
    .X(_06378_));
 sg13g2_nor2_1 _24927_ (.A(\cpu.icache.r_offset[2] ),
    .B(_06378_),
    .Y(_06379_));
 sg13g2_buf_2 _24928_ (.A(_06379_),
    .X(_06380_));
 sg13g2_buf_1 _24929_ (.A(\cpu.icache.r_offset[1] ),
    .X(_06381_));
 sg13g2_buf_1 _24930_ (.A(\cpu.icache.r_offset[0] ),
    .X(_06382_));
 sg13g2_nor2b_1 _24931_ (.A(_06381_),
    .B_N(_06382_),
    .Y(_06383_));
 sg13g2_buf_2 _24932_ (.A(_06383_),
    .X(_06384_));
 sg13g2_and2_1 _24933_ (.A(_06380_),
    .B(_06384_),
    .X(_06385_));
 sg13g2_buf_2 _24934_ (.A(_06385_),
    .X(_06386_));
 sg13g2_nand2_2 _24935_ (.Y(_06387_),
    .A(_06377_),
    .B(_06386_));
 sg13g2_mux2_1 _24936_ (.A0(_06375_),
    .A1(\cpu.icache.r_data[0][0] ),
    .S(_06387_),
    .X(_02001_));
 sg13g2_buf_1 _24937_ (.A(_12632_),
    .X(_06388_));
 sg13g2_inv_1 _24938_ (.Y(_06389_),
    .A(_00246_));
 sg13g2_nand2_1 _24939_ (.Y(_06390_),
    .A(_06381_),
    .B(_06382_));
 sg13g2_buf_2 _24940_ (.A(_06390_),
    .X(_06391_));
 sg13g2_nor3_2 _24941_ (.A(_06378_),
    .B(_06389_),
    .C(_06391_),
    .Y(_06392_));
 sg13g2_nand2_2 _24942_ (.Y(_06393_),
    .A(_06377_),
    .B(_06392_));
 sg13g2_mux2_1 _24943_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][10] ),
    .S(_06393_),
    .X(_02002_));
 sg13g2_buf_1 _24944_ (.A(net1003),
    .X(_06394_));
 sg13g2_mux2_1 _24945_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][11] ),
    .S(_06393_),
    .X(_02003_));
 sg13g2_nor2b_1 _24946_ (.A(_06382_),
    .B_N(_06381_),
    .Y(_06395_));
 sg13g2_buf_1 _24947_ (.A(_06395_),
    .X(_06396_));
 sg13g2_and2_1 _24948_ (.A(_06380_),
    .B(_06396_),
    .X(_06397_));
 sg13g2_buf_2 _24949_ (.A(_06397_),
    .X(_06398_));
 sg13g2_nand2_2 _24950_ (.Y(_06399_),
    .A(_06377_),
    .B(_06398_));
 sg13g2_mux2_1 _24951_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][12] ),
    .S(_06399_),
    .X(_02004_));
 sg13g2_buf_1 _24952_ (.A(_12668_),
    .X(_06400_));
 sg13g2_mux2_1 _24953_ (.A0(_06400_),
    .A1(\cpu.icache.r_data[0][13] ),
    .S(_06399_),
    .X(_02005_));
 sg13g2_mux2_1 _24954_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][14] ),
    .S(_06399_),
    .X(_02006_));
 sg13g2_mux2_1 _24955_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][15] ),
    .S(_06399_),
    .X(_02007_));
 sg13g2_nor2_1 _24956_ (.A(_06378_),
    .B(_00246_),
    .Y(_06401_));
 sg13g2_buf_2 _24957_ (.A(_06401_),
    .X(_06402_));
 sg13g2_and2_1 _24958_ (.A(_06384_),
    .B(_06402_),
    .X(_06403_));
 sg13g2_buf_2 _24959_ (.A(_06403_),
    .X(_06404_));
 sg13g2_nand2_2 _24960_ (.Y(_06405_),
    .A(_06377_),
    .B(_06404_));
 sg13g2_mux2_1 _24961_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][16] ),
    .S(_06405_),
    .X(_02008_));
 sg13g2_mux2_1 _24962_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][17] ),
    .S(_06405_),
    .X(_02009_));
 sg13g2_mux2_1 _24963_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][18] ),
    .S(_06405_),
    .X(_02010_));
 sg13g2_mux2_1 _24964_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][19] ),
    .S(_06405_),
    .X(_02011_));
 sg13g2_mux2_1 _24965_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][1] ),
    .S(_06387_),
    .X(_02012_));
 sg13g2_nor2_2 _24966_ (.A(_06381_),
    .B(_06382_),
    .Y(_06406_));
 sg13g2_and2_1 _24967_ (.A(_06402_),
    .B(_06406_),
    .X(_06407_));
 sg13g2_buf_2 _24968_ (.A(_06407_),
    .X(_06408_));
 sg13g2_nand2_2 _24969_ (.Y(_06409_),
    .A(_06377_),
    .B(_06408_));
 sg13g2_mux2_1 _24970_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][20] ),
    .S(_06409_),
    .X(_02013_));
 sg13g2_mux2_1 _24971_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][21] ),
    .S(_06409_),
    .X(_02014_));
 sg13g2_mux2_1 _24972_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][22] ),
    .S(_06409_),
    .X(_02015_));
 sg13g2_mux2_1 _24973_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][23] ),
    .S(_06409_),
    .X(_02016_));
 sg13g2_inv_1 _24974_ (.Y(_06410_),
    .A(\cpu.i_wstrobe_d ));
 sg13g2_nor3_2 _24975_ (.A(_00246_),
    .B(_06410_),
    .C(_06391_),
    .Y(_06411_));
 sg13g2_nand2_1 _24976_ (.Y(_06412_),
    .A(_06377_),
    .B(_06411_));
 sg13g2_buf_1 _24977_ (.A(_06412_),
    .X(_06413_));
 sg13g2_buf_1 _24978_ (.A(net405),
    .X(_06414_));
 sg13g2_mux2_1 _24979_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][24] ),
    .S(net368),
    .X(_02017_));
 sg13g2_mux2_1 _24980_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][25] ),
    .S(net368),
    .X(_02018_));
 sg13g2_mux2_1 _24981_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][26] ),
    .S(_06414_),
    .X(_02019_));
 sg13g2_mux2_1 _24982_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][27] ),
    .S(_06414_),
    .X(_02020_));
 sg13g2_and2_1 _24983_ (.A(_06396_),
    .B(_06402_),
    .X(_06415_));
 sg13g2_buf_2 _24984_ (.A(_06415_),
    .X(_06416_));
 sg13g2_nand2_2 _24985_ (.Y(_06417_),
    .A(_06377_),
    .B(_06416_));
 sg13g2_mux2_1 _24986_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][28] ),
    .S(_06417_),
    .X(_02021_));
 sg13g2_mux2_1 _24987_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][29] ),
    .S(_06417_),
    .X(_02022_));
 sg13g2_mux2_1 _24988_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][2] ),
    .S(_06387_),
    .X(_02023_));
 sg13g2_mux2_1 _24989_ (.A0(_06388_),
    .A1(\cpu.icache.r_data[0][30] ),
    .S(_06417_),
    .X(_02024_));
 sg13g2_mux2_1 _24990_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][31] ),
    .S(_06417_),
    .X(_02025_));
 sg13g2_mux2_1 _24991_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][3] ),
    .S(_06387_),
    .X(_02026_));
 sg13g2_and2_1 _24992_ (.A(_06380_),
    .B(_06406_),
    .X(_06418_));
 sg13g2_buf_2 _24993_ (.A(_06418_),
    .X(_06419_));
 sg13g2_nand2_2 _24994_ (.Y(_06420_),
    .A(_06377_),
    .B(_06419_));
 sg13g2_mux2_1 _24995_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][4] ),
    .S(_06420_),
    .X(_02027_));
 sg13g2_mux2_1 _24996_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][5] ),
    .S(_06420_),
    .X(_02028_));
 sg13g2_mux2_1 _24997_ (.A0(net854),
    .A1(\cpu.icache.r_data[0][6] ),
    .S(_06420_),
    .X(_02029_));
 sg13g2_mux2_1 _24998_ (.A0(net853),
    .A1(\cpu.icache.r_data[0][7] ),
    .S(_06420_),
    .X(_02030_));
 sg13g2_mux2_1 _24999_ (.A0(net855),
    .A1(\cpu.icache.r_data[0][8] ),
    .S(_06393_),
    .X(_02031_));
 sg13g2_mux2_1 _25000_ (.A0(net852),
    .A1(\cpu.icache.r_data[0][9] ),
    .S(_06393_),
    .X(_02032_));
 sg13g2_buf_1 _25001_ (.A(net1002),
    .X(_06421_));
 sg13g2_nand2b_1 _25002_ (.Y(_06422_),
    .B(_08864_),
    .A_N(_08451_));
 sg13g2_buf_4 _25003_ (.X(_06423_),
    .A(_06422_));
 sg13g2_nand2_2 _25004_ (.Y(_06424_),
    .A(_06380_),
    .B(_06384_));
 sg13g2_nor2_2 _25005_ (.A(_06423_),
    .B(_06424_),
    .Y(_06425_));
 sg13g2_mux2_1 _25006_ (.A0(\cpu.icache.r_data[1][0] ),
    .A1(_06421_),
    .S(_06425_),
    .X(_02033_));
 sg13g2_buf_1 _25007_ (.A(net1108),
    .X(_06426_));
 sg13g2_or3_1 _25008_ (.A(_06378_),
    .B(_06389_),
    .C(_06391_),
    .X(_06427_));
 sg13g2_buf_2 _25009_ (.A(_06427_),
    .X(_06428_));
 sg13g2_nor2_2 _25010_ (.A(_06423_),
    .B(_06428_),
    .Y(_06429_));
 sg13g2_mux2_1 _25011_ (.A0(\cpu.icache.r_data[1][10] ),
    .A1(net970),
    .S(_06429_),
    .X(_02034_));
 sg13g2_buf_1 _25012_ (.A(net1003),
    .X(_06430_));
 sg13g2_mux2_1 _25013_ (.A0(\cpu.icache.r_data[1][11] ),
    .A1(net850),
    .S(_06429_),
    .X(_02035_));
 sg13g2_buf_1 _25014_ (.A(net1002),
    .X(_06431_));
 sg13g2_nand2_2 _25015_ (.Y(_06432_),
    .A(_06380_),
    .B(_06396_));
 sg13g2_nor2_2 _25016_ (.A(_06423_),
    .B(_06432_),
    .Y(_06433_));
 sg13g2_mux2_1 _25017_ (.A0(\cpu.icache.r_data[1][12] ),
    .A1(net849),
    .S(_06433_),
    .X(_02036_));
 sg13g2_buf_1 _25018_ (.A(net1109),
    .X(_06434_));
 sg13g2_mux2_1 _25019_ (.A0(\cpu.icache.r_data[1][13] ),
    .A1(net969),
    .S(_06433_),
    .X(_02037_));
 sg13g2_buf_1 _25020_ (.A(net1108),
    .X(_06435_));
 sg13g2_mux2_1 _25021_ (.A0(\cpu.icache.r_data[1][14] ),
    .A1(net968),
    .S(_06433_),
    .X(_02038_));
 sg13g2_buf_1 _25022_ (.A(net1003),
    .X(_06436_));
 sg13g2_mux2_1 _25023_ (.A0(\cpu.icache.r_data[1][15] ),
    .A1(net848),
    .S(_06433_),
    .X(_02039_));
 sg13g2_nand2_2 _25024_ (.Y(_06437_),
    .A(_06384_),
    .B(_06402_));
 sg13g2_nor2_2 _25025_ (.A(_06423_),
    .B(_06437_),
    .Y(_06438_));
 sg13g2_mux2_1 _25026_ (.A0(\cpu.icache.r_data[1][16] ),
    .A1(net849),
    .S(_06438_),
    .X(_02040_));
 sg13g2_buf_1 _25027_ (.A(net1109),
    .X(_06439_));
 sg13g2_mux2_1 _25028_ (.A0(\cpu.icache.r_data[1][17] ),
    .A1(net967),
    .S(_06438_),
    .X(_02041_));
 sg13g2_mux2_1 _25029_ (.A0(\cpu.icache.r_data[1][18] ),
    .A1(net968),
    .S(_06438_),
    .X(_02042_));
 sg13g2_mux2_1 _25030_ (.A0(\cpu.icache.r_data[1][19] ),
    .A1(net848),
    .S(_06438_),
    .X(_02043_));
 sg13g2_mux2_1 _25031_ (.A0(\cpu.icache.r_data[1][1] ),
    .A1(net967),
    .S(_06425_),
    .X(_02044_));
 sg13g2_nand2_2 _25032_ (.Y(_06440_),
    .A(_06402_),
    .B(_06406_));
 sg13g2_nor2_2 _25033_ (.A(_06423_),
    .B(_06440_),
    .Y(_06441_));
 sg13g2_mux2_1 _25034_ (.A0(\cpu.icache.r_data[1][20] ),
    .A1(net849),
    .S(_06441_),
    .X(_02045_));
 sg13g2_mux2_1 _25035_ (.A0(\cpu.icache.r_data[1][21] ),
    .A1(net967),
    .S(_06441_),
    .X(_02046_));
 sg13g2_mux2_1 _25036_ (.A0(\cpu.icache.r_data[1][22] ),
    .A1(net968),
    .S(_06441_),
    .X(_02047_));
 sg13g2_mux2_1 _25037_ (.A0(\cpu.icache.r_data[1][23] ),
    .A1(net848),
    .S(_06441_),
    .X(_02048_));
 sg13g2_nand4_1 _25038_ (.B(_06382_),
    .C(_06389_),
    .A(_06381_),
    .Y(_06442_),
    .D(\cpu.i_wstrobe_d ));
 sg13g2_buf_1 _25039_ (.A(_06442_),
    .X(_06443_));
 sg13g2_nor2_1 _25040_ (.A(_06423_),
    .B(_06443_),
    .Y(_06444_));
 sg13g2_buf_2 _25041_ (.A(_06444_),
    .X(_06445_));
 sg13g2_mux2_1 _25042_ (.A0(\cpu.icache.r_data[1][24] ),
    .A1(net849),
    .S(_06445_),
    .X(_02049_));
 sg13g2_mux2_1 _25043_ (.A0(\cpu.icache.r_data[1][25] ),
    .A1(net967),
    .S(_06445_),
    .X(_02050_));
 sg13g2_mux2_1 _25044_ (.A0(\cpu.icache.r_data[1][26] ),
    .A1(net968),
    .S(_06445_),
    .X(_02051_));
 sg13g2_mux2_1 _25045_ (.A0(\cpu.icache.r_data[1][27] ),
    .A1(net848),
    .S(_06445_),
    .X(_02052_));
 sg13g2_nand2_2 _25046_ (.Y(_06446_),
    .A(_06396_),
    .B(_06402_));
 sg13g2_nor2_2 _25047_ (.A(_06423_),
    .B(_06446_),
    .Y(_06447_));
 sg13g2_mux2_1 _25048_ (.A0(\cpu.icache.r_data[1][28] ),
    .A1(net849),
    .S(_06447_),
    .X(_02053_));
 sg13g2_mux2_1 _25049_ (.A0(\cpu.icache.r_data[1][29] ),
    .A1(net967),
    .S(_06447_),
    .X(_02054_));
 sg13g2_mux2_1 _25050_ (.A0(\cpu.icache.r_data[1][2] ),
    .A1(_06435_),
    .S(_06425_),
    .X(_02055_));
 sg13g2_mux2_1 _25051_ (.A0(\cpu.icache.r_data[1][30] ),
    .A1(_06435_),
    .S(_06447_),
    .X(_02056_));
 sg13g2_mux2_1 _25052_ (.A0(\cpu.icache.r_data[1][31] ),
    .A1(net848),
    .S(_06447_),
    .X(_02057_));
 sg13g2_mux2_1 _25053_ (.A0(\cpu.icache.r_data[1][3] ),
    .A1(_06436_),
    .S(_06425_),
    .X(_02058_));
 sg13g2_nand2_2 _25054_ (.Y(_06448_),
    .A(_06380_),
    .B(_06406_));
 sg13g2_nor2_2 _25055_ (.A(_06423_),
    .B(_06448_),
    .Y(_06449_));
 sg13g2_mux2_1 _25056_ (.A0(\cpu.icache.r_data[1][4] ),
    .A1(net849),
    .S(_06449_),
    .X(_02059_));
 sg13g2_mux2_1 _25057_ (.A0(\cpu.icache.r_data[1][5] ),
    .A1(net967),
    .S(_06449_),
    .X(_02060_));
 sg13g2_mux2_1 _25058_ (.A0(\cpu.icache.r_data[1][6] ),
    .A1(net968),
    .S(_06449_),
    .X(_02061_));
 sg13g2_mux2_1 _25059_ (.A0(\cpu.icache.r_data[1][7] ),
    .A1(_06436_),
    .S(_06449_),
    .X(_02062_));
 sg13g2_mux2_1 _25060_ (.A0(\cpu.icache.r_data[1][8] ),
    .A1(net849),
    .S(_06429_),
    .X(_02063_));
 sg13g2_mux2_1 _25061_ (.A0(\cpu.icache.r_data[1][9] ),
    .A1(net967),
    .S(_06429_),
    .X(_02064_));
 sg13g2_nand2_1 _25062_ (.Y(_06450_),
    .A(net820),
    .B(_08453_));
 sg13g2_buf_4 _25063_ (.X(_06451_),
    .A(_06450_));
 sg13g2_nor2_2 _25064_ (.A(_06451_),
    .B(_06424_),
    .Y(_06452_));
 sg13g2_mux2_1 _25065_ (.A0(\cpu.icache.r_data[2][0] ),
    .A1(_06431_),
    .S(_06452_),
    .X(_02065_));
 sg13g2_nor2_2 _25066_ (.A(_06451_),
    .B(_06428_),
    .Y(_06453_));
 sg13g2_mux2_1 _25067_ (.A0(\cpu.icache.r_data[2][10] ),
    .A1(net968),
    .S(_06453_),
    .X(_02066_));
 sg13g2_mux2_1 _25068_ (.A0(\cpu.icache.r_data[2][11] ),
    .A1(net848),
    .S(_06453_),
    .X(_02067_));
 sg13g2_nor2_2 _25069_ (.A(_06451_),
    .B(_06432_),
    .Y(_06454_));
 sg13g2_mux2_1 _25070_ (.A0(\cpu.icache.r_data[2][12] ),
    .A1(_06431_),
    .S(_06454_),
    .X(_02068_));
 sg13g2_mux2_1 _25071_ (.A0(\cpu.icache.r_data[2][13] ),
    .A1(_06439_),
    .S(_06454_),
    .X(_02069_));
 sg13g2_mux2_1 _25072_ (.A0(\cpu.icache.r_data[2][14] ),
    .A1(net968),
    .S(_06454_),
    .X(_02070_));
 sg13g2_mux2_1 _25073_ (.A0(\cpu.icache.r_data[2][15] ),
    .A1(net848),
    .S(_06454_),
    .X(_02071_));
 sg13g2_nor2_2 _25074_ (.A(_06451_),
    .B(_06437_),
    .Y(_06455_));
 sg13g2_mux2_1 _25075_ (.A0(\cpu.icache.r_data[2][16] ),
    .A1(net849),
    .S(_06455_),
    .X(_02072_));
 sg13g2_mux2_1 _25076_ (.A0(\cpu.icache.r_data[2][17] ),
    .A1(_06439_),
    .S(_06455_),
    .X(_02073_));
 sg13g2_mux2_1 _25077_ (.A0(\cpu.icache.r_data[2][18] ),
    .A1(net968),
    .S(_06455_),
    .X(_02074_));
 sg13g2_mux2_1 _25078_ (.A0(\cpu.icache.r_data[2][19] ),
    .A1(net848),
    .S(_06455_),
    .X(_02075_));
 sg13g2_mux2_1 _25079_ (.A0(\cpu.icache.r_data[2][1] ),
    .A1(net967),
    .S(_06452_),
    .X(_02076_));
 sg13g2_buf_1 _25080_ (.A(net1002),
    .X(_06456_));
 sg13g2_nor2_2 _25081_ (.A(_06451_),
    .B(_06440_),
    .Y(_06457_));
 sg13g2_mux2_1 _25082_ (.A0(\cpu.icache.r_data[2][20] ),
    .A1(net847),
    .S(_06457_),
    .X(_02077_));
 sg13g2_buf_1 _25083_ (.A(_12207_),
    .X(_06458_));
 sg13g2_mux2_1 _25084_ (.A0(\cpu.icache.r_data[2][21] ),
    .A1(net966),
    .S(_06457_),
    .X(_02078_));
 sg13g2_buf_1 _25085_ (.A(_12214_),
    .X(_06459_));
 sg13g2_mux2_1 _25086_ (.A0(\cpu.icache.r_data[2][22] ),
    .A1(net965),
    .S(_06457_),
    .X(_02079_));
 sg13g2_buf_1 _25087_ (.A(net1003),
    .X(_06460_));
 sg13g2_mux2_1 _25088_ (.A0(\cpu.icache.r_data[2][23] ),
    .A1(net846),
    .S(_06457_),
    .X(_02080_));
 sg13g2_nor2_1 _25089_ (.A(_06451_),
    .B(_06443_),
    .Y(_06461_));
 sg13g2_buf_2 _25090_ (.A(_06461_),
    .X(_06462_));
 sg13g2_mux2_1 _25091_ (.A0(\cpu.icache.r_data[2][24] ),
    .A1(net847),
    .S(_06462_),
    .X(_02081_));
 sg13g2_mux2_1 _25092_ (.A0(\cpu.icache.r_data[2][25] ),
    .A1(net966),
    .S(_06462_),
    .X(_02082_));
 sg13g2_mux2_1 _25093_ (.A0(\cpu.icache.r_data[2][26] ),
    .A1(net965),
    .S(_06462_),
    .X(_02083_));
 sg13g2_mux2_1 _25094_ (.A0(\cpu.icache.r_data[2][27] ),
    .A1(net846),
    .S(_06462_),
    .X(_02084_));
 sg13g2_nor2_2 _25095_ (.A(_06451_),
    .B(_06446_),
    .Y(_06463_));
 sg13g2_mux2_1 _25096_ (.A0(\cpu.icache.r_data[2][28] ),
    .A1(_06456_),
    .S(_06463_),
    .X(_02085_));
 sg13g2_mux2_1 _25097_ (.A0(\cpu.icache.r_data[2][29] ),
    .A1(net966),
    .S(_06463_),
    .X(_02086_));
 sg13g2_mux2_1 _25098_ (.A0(\cpu.icache.r_data[2][2] ),
    .A1(_06459_),
    .S(_06452_),
    .X(_02087_));
 sg13g2_mux2_1 _25099_ (.A0(\cpu.icache.r_data[2][30] ),
    .A1(_06459_),
    .S(_06463_),
    .X(_02088_));
 sg13g2_mux2_1 _25100_ (.A0(\cpu.icache.r_data[2][31] ),
    .A1(_06460_),
    .S(_06463_),
    .X(_02089_));
 sg13g2_mux2_1 _25101_ (.A0(\cpu.icache.r_data[2][3] ),
    .A1(_06460_),
    .S(_06452_),
    .X(_02090_));
 sg13g2_nor2_2 _25102_ (.A(_06451_),
    .B(_06448_),
    .Y(_06464_));
 sg13g2_mux2_1 _25103_ (.A0(\cpu.icache.r_data[2][4] ),
    .A1(net847),
    .S(_06464_),
    .X(_02091_));
 sg13g2_mux2_1 _25104_ (.A0(\cpu.icache.r_data[2][5] ),
    .A1(net966),
    .S(_06464_),
    .X(_02092_));
 sg13g2_mux2_1 _25105_ (.A0(\cpu.icache.r_data[2][6] ),
    .A1(net965),
    .S(_06464_),
    .X(_02093_));
 sg13g2_mux2_1 _25106_ (.A0(\cpu.icache.r_data[2][7] ),
    .A1(net846),
    .S(_06464_),
    .X(_02094_));
 sg13g2_mux2_1 _25107_ (.A0(\cpu.icache.r_data[2][8] ),
    .A1(net847),
    .S(_06453_),
    .X(_02095_));
 sg13g2_mux2_1 _25108_ (.A0(\cpu.icache.r_data[2][9] ),
    .A1(net966),
    .S(_06453_),
    .X(_02096_));
 sg13g2_nand2_2 _25109_ (.Y(_06465_),
    .A(net472),
    .B(_06386_));
 sg13g2_mux2_1 _25110_ (.A0(_06375_),
    .A1(\cpu.icache.r_data[3][0] ),
    .S(_06465_),
    .X(_02097_));
 sg13g2_and2_1 _25111_ (.A(net472),
    .B(_06392_),
    .X(_06466_));
 sg13g2_buf_1 _25112_ (.A(_06466_),
    .X(_06467_));
 sg13g2_mux2_1 _25113_ (.A0(\cpu.icache.r_data[3][10] ),
    .A1(net965),
    .S(_06467_),
    .X(_02098_));
 sg13g2_mux2_1 _25114_ (.A0(\cpu.icache.r_data[3][11] ),
    .A1(net846),
    .S(_06467_),
    .X(_02099_));
 sg13g2_nand2_2 _25115_ (.Y(_06468_),
    .A(net472),
    .B(_06398_));
 sg13g2_mux2_1 _25116_ (.A0(net855),
    .A1(\cpu.icache.r_data[3][12] ),
    .S(_06468_),
    .X(_02100_));
 sg13g2_mux2_1 _25117_ (.A0(net852),
    .A1(\cpu.icache.r_data[3][13] ),
    .S(_06468_),
    .X(_02101_));
 sg13g2_mux2_1 _25118_ (.A0(net854),
    .A1(\cpu.icache.r_data[3][14] ),
    .S(_06468_),
    .X(_02102_));
 sg13g2_mux2_1 _25119_ (.A0(_06394_),
    .A1(\cpu.icache.r_data[3][15] ),
    .S(_06468_),
    .X(_02103_));
 sg13g2_buf_1 _25120_ (.A(_02950_),
    .X(_06469_));
 sg13g2_nand2_2 _25121_ (.Y(_06470_),
    .A(_03213_),
    .B(_06404_));
 sg13g2_mux2_1 _25122_ (.A0(net845),
    .A1(\cpu.icache.r_data[3][16] ),
    .S(_06470_),
    .X(_02104_));
 sg13g2_mux2_1 _25123_ (.A0(_06400_),
    .A1(\cpu.icache.r_data[3][17] ),
    .S(_06470_),
    .X(_02105_));
 sg13g2_mux2_1 _25124_ (.A0(_06388_),
    .A1(\cpu.icache.r_data[3][18] ),
    .S(_06470_),
    .X(_02106_));
 sg13g2_mux2_1 _25125_ (.A0(_06394_),
    .A1(\cpu.icache.r_data[3][19] ),
    .S(_06470_),
    .X(_02107_));
 sg13g2_buf_1 _25126_ (.A(_12668_),
    .X(_06471_));
 sg13g2_mux2_1 _25127_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][1] ),
    .S(_06465_),
    .X(_02108_));
 sg13g2_nand2_2 _25128_ (.Y(_06472_),
    .A(net472),
    .B(_06408_));
 sg13g2_mux2_1 _25129_ (.A0(net845),
    .A1(\cpu.icache.r_data[3][20] ),
    .S(_06472_),
    .X(_02109_));
 sg13g2_mux2_1 _25130_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][21] ),
    .S(_06472_),
    .X(_02110_));
 sg13g2_buf_1 _25131_ (.A(_12632_),
    .X(_06473_));
 sg13g2_mux2_1 _25132_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][22] ),
    .S(_06472_),
    .X(_02111_));
 sg13g2_buf_1 _25133_ (.A(_02921_),
    .X(_06474_));
 sg13g2_mux2_1 _25134_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][23] ),
    .S(_06472_),
    .X(_02112_));
 sg13g2_nand2_1 _25135_ (.Y(_06475_),
    .A(net472),
    .B(_06411_));
 sg13g2_buf_1 _25136_ (.A(_06475_),
    .X(_06476_));
 sg13g2_buf_1 _25137_ (.A(_06476_),
    .X(_06477_));
 sg13g2_mux2_1 _25138_ (.A0(net845),
    .A1(\cpu.icache.r_data[3][24] ),
    .S(net312),
    .X(_02113_));
 sg13g2_mux2_1 _25139_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][25] ),
    .S(net312),
    .X(_02114_));
 sg13g2_mux2_1 _25140_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][26] ),
    .S(_06477_),
    .X(_02115_));
 sg13g2_mux2_1 _25141_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][27] ),
    .S(_06477_),
    .X(_02116_));
 sg13g2_nand2_2 _25142_ (.Y(_06478_),
    .A(_03213_),
    .B(_06416_));
 sg13g2_mux2_1 _25143_ (.A0(net845),
    .A1(\cpu.icache.r_data[3][28] ),
    .S(_06478_),
    .X(_02117_));
 sg13g2_mux2_1 _25144_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][29] ),
    .S(_06478_),
    .X(_02118_));
 sg13g2_mux2_1 _25145_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][2] ),
    .S(_06465_),
    .X(_02119_));
 sg13g2_mux2_1 _25146_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][30] ),
    .S(_06478_),
    .X(_02120_));
 sg13g2_mux2_1 _25147_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][31] ),
    .S(_06478_),
    .X(_02121_));
 sg13g2_mux2_1 _25148_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][3] ),
    .S(_06465_),
    .X(_02122_));
 sg13g2_nand2_2 _25149_ (.Y(_06479_),
    .A(net472),
    .B(_06419_));
 sg13g2_mux2_1 _25150_ (.A0(net845),
    .A1(\cpu.icache.r_data[3][4] ),
    .S(_06479_),
    .X(_02123_));
 sg13g2_mux2_1 _25151_ (.A0(net844),
    .A1(\cpu.icache.r_data[3][5] ),
    .S(_06479_),
    .X(_02124_));
 sg13g2_mux2_1 _25152_ (.A0(net843),
    .A1(\cpu.icache.r_data[3][6] ),
    .S(_06479_),
    .X(_02125_));
 sg13g2_mux2_1 _25153_ (.A0(net842),
    .A1(\cpu.icache.r_data[3][7] ),
    .S(_06479_),
    .X(_02126_));
 sg13g2_mux2_1 _25154_ (.A0(\cpu.icache.r_data[3][8] ),
    .A1(net847),
    .S(_06467_),
    .X(_02127_));
 sg13g2_mux2_1 _25155_ (.A0(\cpu.icache.r_data[3][9] ),
    .A1(net966),
    .S(_06467_),
    .X(_02128_));
 sg13g2_nand2_2 _25156_ (.Y(_06480_),
    .A(net619),
    .B(_06386_));
 sg13g2_mux2_1 _25157_ (.A0(_06469_),
    .A1(\cpu.icache.r_data[4][0] ),
    .S(_06480_),
    .X(_02129_));
 sg13g2_and2_1 _25158_ (.A(net619),
    .B(_06392_),
    .X(_06481_));
 sg13g2_buf_1 _25159_ (.A(_06481_),
    .X(_06482_));
 sg13g2_mux2_1 _25160_ (.A0(\cpu.icache.r_data[4][10] ),
    .A1(net965),
    .S(_06482_),
    .X(_02130_));
 sg13g2_mux2_1 _25161_ (.A0(\cpu.icache.r_data[4][11] ),
    .A1(net846),
    .S(_06482_),
    .X(_02131_));
 sg13g2_nand2_2 _25162_ (.Y(_06483_),
    .A(net619),
    .B(_06398_));
 sg13g2_mux2_1 _25163_ (.A0(_06469_),
    .A1(\cpu.icache.r_data[4][12] ),
    .S(_06483_),
    .X(_02132_));
 sg13g2_mux2_1 _25164_ (.A0(net844),
    .A1(\cpu.icache.r_data[4][13] ),
    .S(_06483_),
    .X(_02133_));
 sg13g2_mux2_1 _25165_ (.A0(net843),
    .A1(\cpu.icache.r_data[4][14] ),
    .S(_06483_),
    .X(_02134_));
 sg13g2_mux2_1 _25166_ (.A0(net842),
    .A1(\cpu.icache.r_data[4][15] ),
    .S(_06483_),
    .X(_02135_));
 sg13g2_nand2_2 _25167_ (.Y(_06484_),
    .A(_03248_),
    .B(_06404_));
 sg13g2_mux2_1 _25168_ (.A0(net845),
    .A1(\cpu.icache.r_data[4][16] ),
    .S(_06484_),
    .X(_02136_));
 sg13g2_mux2_1 _25169_ (.A0(net844),
    .A1(\cpu.icache.r_data[4][17] ),
    .S(_06484_),
    .X(_02137_));
 sg13g2_mux2_1 _25170_ (.A0(net843),
    .A1(\cpu.icache.r_data[4][18] ),
    .S(_06484_),
    .X(_02138_));
 sg13g2_mux2_1 _25171_ (.A0(net842),
    .A1(\cpu.icache.r_data[4][19] ),
    .S(_06484_),
    .X(_02139_));
 sg13g2_mux2_1 _25172_ (.A0(_06471_),
    .A1(\cpu.icache.r_data[4][1] ),
    .S(_06480_),
    .X(_02140_));
 sg13g2_nand2_2 _25173_ (.Y(_06485_),
    .A(net619),
    .B(_06408_));
 sg13g2_mux2_1 _25174_ (.A0(net845),
    .A1(\cpu.icache.r_data[4][20] ),
    .S(_06485_),
    .X(_02141_));
 sg13g2_mux2_1 _25175_ (.A0(net844),
    .A1(\cpu.icache.r_data[4][21] ),
    .S(_06485_),
    .X(_02142_));
 sg13g2_mux2_1 _25176_ (.A0(net843),
    .A1(\cpu.icache.r_data[4][22] ),
    .S(_06485_),
    .X(_02143_));
 sg13g2_mux2_1 _25177_ (.A0(net842),
    .A1(\cpu.icache.r_data[4][23] ),
    .S(_06485_),
    .X(_02144_));
 sg13g2_and2_1 _25178_ (.A(net619),
    .B(_06411_),
    .X(_06486_));
 sg13g2_buf_2 _25179_ (.A(_06486_),
    .X(_06487_));
 sg13g2_mux2_1 _25180_ (.A0(\cpu.icache.r_data[4][24] ),
    .A1(net847),
    .S(_06487_),
    .X(_02145_));
 sg13g2_mux2_1 _25181_ (.A0(\cpu.icache.r_data[4][25] ),
    .A1(net966),
    .S(_06487_),
    .X(_02146_));
 sg13g2_mux2_1 _25182_ (.A0(\cpu.icache.r_data[4][26] ),
    .A1(net965),
    .S(_06487_),
    .X(_02147_));
 sg13g2_mux2_1 _25183_ (.A0(\cpu.icache.r_data[4][27] ),
    .A1(net846),
    .S(_06487_),
    .X(_02148_));
 sg13g2_nand2_2 _25184_ (.Y(_06488_),
    .A(_03248_),
    .B(_06416_));
 sg13g2_mux2_1 _25185_ (.A0(net845),
    .A1(\cpu.icache.r_data[4][28] ),
    .S(_06488_),
    .X(_02149_));
 sg13g2_mux2_1 _25186_ (.A0(_06471_),
    .A1(\cpu.icache.r_data[4][29] ),
    .S(_06488_),
    .X(_02150_));
 sg13g2_mux2_1 _25187_ (.A0(_06473_),
    .A1(\cpu.icache.r_data[4][2] ),
    .S(_06480_),
    .X(_02151_));
 sg13g2_mux2_1 _25188_ (.A0(_06473_),
    .A1(\cpu.icache.r_data[4][30] ),
    .S(_06488_),
    .X(_02152_));
 sg13g2_mux2_1 _25189_ (.A0(_06474_),
    .A1(\cpu.icache.r_data[4][31] ),
    .S(_06488_),
    .X(_02153_));
 sg13g2_mux2_1 _25190_ (.A0(_06474_),
    .A1(\cpu.icache.r_data[4][3] ),
    .S(_06480_),
    .X(_02154_));
 sg13g2_nand2_2 _25191_ (.Y(_06489_),
    .A(net619),
    .B(_06419_));
 sg13g2_mux2_1 _25192_ (.A0(net851),
    .A1(\cpu.icache.r_data[4][4] ),
    .S(_06489_),
    .X(_02155_));
 sg13g2_mux2_1 _25193_ (.A0(net969),
    .A1(\cpu.icache.r_data[4][5] ),
    .S(_06489_),
    .X(_02156_));
 sg13g2_mux2_1 _25194_ (.A0(net970),
    .A1(\cpu.icache.r_data[4][6] ),
    .S(_06489_),
    .X(_02157_));
 sg13g2_mux2_1 _25195_ (.A0(net850),
    .A1(\cpu.icache.r_data[4][7] ),
    .S(_06489_),
    .X(_02158_));
 sg13g2_mux2_1 _25196_ (.A0(\cpu.icache.r_data[4][8] ),
    .A1(net847),
    .S(_06482_),
    .X(_02159_));
 sg13g2_mux2_1 _25197_ (.A0(\cpu.icache.r_data[4][9] ),
    .A1(net966),
    .S(_06482_),
    .X(_02160_));
 sg13g2_nand2_1 _25198_ (.Y(_06490_),
    .A(net1076),
    .B(_08864_));
 sg13g2_buf_4 _25199_ (.X(_06491_),
    .A(_06490_));
 sg13g2_nor2_2 _25200_ (.A(_06491_),
    .B(_06424_),
    .Y(_06492_));
 sg13g2_mux2_1 _25201_ (.A0(\cpu.icache.r_data[5][0] ),
    .A1(net847),
    .S(_06492_),
    .X(_02161_));
 sg13g2_nor2_2 _25202_ (.A(_06491_),
    .B(_06428_),
    .Y(_06493_));
 sg13g2_mux2_1 _25203_ (.A0(\cpu.icache.r_data[5][10] ),
    .A1(net965),
    .S(_06493_),
    .X(_02162_));
 sg13g2_mux2_1 _25204_ (.A0(\cpu.icache.r_data[5][11] ),
    .A1(net846),
    .S(_06493_),
    .X(_02163_));
 sg13g2_nor2_2 _25205_ (.A(_06491_),
    .B(_06432_),
    .Y(_06494_));
 sg13g2_mux2_1 _25206_ (.A0(\cpu.icache.r_data[5][12] ),
    .A1(_06456_),
    .S(_06494_),
    .X(_02164_));
 sg13g2_mux2_1 _25207_ (.A0(\cpu.icache.r_data[5][13] ),
    .A1(_06458_),
    .S(_06494_),
    .X(_02165_));
 sg13g2_mux2_1 _25208_ (.A0(\cpu.icache.r_data[5][14] ),
    .A1(net965),
    .S(_06494_),
    .X(_02166_));
 sg13g2_mux2_1 _25209_ (.A0(\cpu.icache.r_data[5][15] ),
    .A1(net846),
    .S(_06494_),
    .X(_02167_));
 sg13g2_buf_2 _25210_ (.A(net1113),
    .X(_06495_));
 sg13g2_nor2_2 _25211_ (.A(_06491_),
    .B(_06437_),
    .Y(_06496_));
 sg13g2_mux2_1 _25212_ (.A0(\cpu.icache.r_data[5][16] ),
    .A1(net964),
    .S(_06496_),
    .X(_02168_));
 sg13g2_mux2_1 _25213_ (.A0(\cpu.icache.r_data[5][17] ),
    .A1(_06458_),
    .S(_06496_),
    .X(_02169_));
 sg13g2_buf_1 _25214_ (.A(_12214_),
    .X(_06497_));
 sg13g2_mux2_1 _25215_ (.A0(\cpu.icache.r_data[5][18] ),
    .A1(net963),
    .S(_06496_),
    .X(_02170_));
 sg13g2_buf_2 _25216_ (.A(net1107),
    .X(_06498_));
 sg13g2_mux2_1 _25217_ (.A0(\cpu.icache.r_data[5][19] ),
    .A1(net962),
    .S(_06496_),
    .X(_02171_));
 sg13g2_buf_1 _25218_ (.A(_12207_),
    .X(_06499_));
 sg13g2_mux2_1 _25219_ (.A0(\cpu.icache.r_data[5][1] ),
    .A1(net961),
    .S(_06492_),
    .X(_02172_));
 sg13g2_nor2_2 _25220_ (.A(_06491_),
    .B(_06440_),
    .Y(_06500_));
 sg13g2_mux2_1 _25221_ (.A0(\cpu.icache.r_data[5][20] ),
    .A1(net964),
    .S(_06500_),
    .X(_02173_));
 sg13g2_mux2_1 _25222_ (.A0(\cpu.icache.r_data[5][21] ),
    .A1(net961),
    .S(_06500_),
    .X(_02174_));
 sg13g2_mux2_1 _25223_ (.A0(\cpu.icache.r_data[5][22] ),
    .A1(net963),
    .S(_06500_),
    .X(_02175_));
 sg13g2_mux2_1 _25224_ (.A0(\cpu.icache.r_data[5][23] ),
    .A1(net962),
    .S(_06500_),
    .X(_02176_));
 sg13g2_nor2_1 _25225_ (.A(_06491_),
    .B(_06443_),
    .Y(_06501_));
 sg13g2_buf_2 _25226_ (.A(_06501_),
    .X(_06502_));
 sg13g2_mux2_1 _25227_ (.A0(\cpu.icache.r_data[5][24] ),
    .A1(net964),
    .S(_06502_),
    .X(_02177_));
 sg13g2_mux2_1 _25228_ (.A0(\cpu.icache.r_data[5][25] ),
    .A1(net961),
    .S(_06502_),
    .X(_02178_));
 sg13g2_mux2_1 _25229_ (.A0(\cpu.icache.r_data[5][26] ),
    .A1(net963),
    .S(_06502_),
    .X(_02179_));
 sg13g2_mux2_1 _25230_ (.A0(\cpu.icache.r_data[5][27] ),
    .A1(net962),
    .S(_06502_),
    .X(_02180_));
 sg13g2_nor2_2 _25231_ (.A(_06491_),
    .B(_06446_),
    .Y(_06503_));
 sg13g2_mux2_1 _25232_ (.A0(\cpu.icache.r_data[5][28] ),
    .A1(net964),
    .S(_06503_),
    .X(_02181_));
 sg13g2_mux2_1 _25233_ (.A0(\cpu.icache.r_data[5][29] ),
    .A1(net961),
    .S(_06503_),
    .X(_02182_));
 sg13g2_mux2_1 _25234_ (.A0(\cpu.icache.r_data[5][2] ),
    .A1(_06497_),
    .S(_06492_),
    .X(_02183_));
 sg13g2_mux2_1 _25235_ (.A0(\cpu.icache.r_data[5][30] ),
    .A1(net963),
    .S(_06503_),
    .X(_02184_));
 sg13g2_mux2_1 _25236_ (.A0(\cpu.icache.r_data[5][31] ),
    .A1(net962),
    .S(_06503_),
    .X(_02185_));
 sg13g2_mux2_1 _25237_ (.A0(\cpu.icache.r_data[5][3] ),
    .A1(net962),
    .S(_06492_),
    .X(_02186_));
 sg13g2_nor2_2 _25238_ (.A(_06491_),
    .B(_06448_),
    .Y(_06504_));
 sg13g2_mux2_1 _25239_ (.A0(\cpu.icache.r_data[5][4] ),
    .A1(net964),
    .S(_06504_),
    .X(_02187_));
 sg13g2_mux2_1 _25240_ (.A0(\cpu.icache.r_data[5][5] ),
    .A1(net961),
    .S(_06504_),
    .X(_02188_));
 sg13g2_mux2_1 _25241_ (.A0(\cpu.icache.r_data[5][6] ),
    .A1(net963),
    .S(_06504_),
    .X(_02189_));
 sg13g2_mux2_1 _25242_ (.A0(\cpu.icache.r_data[5][7] ),
    .A1(net962),
    .S(_06504_),
    .X(_02190_));
 sg13g2_mux2_1 _25243_ (.A0(\cpu.icache.r_data[5][8] ),
    .A1(net964),
    .S(_06493_),
    .X(_02191_));
 sg13g2_mux2_1 _25244_ (.A0(\cpu.icache.r_data[5][9] ),
    .A1(net961),
    .S(_06493_),
    .X(_02192_));
 sg13g2_nand2_2 _25245_ (.Y(_06505_),
    .A(net570),
    .B(_06386_));
 sg13g2_mux2_1 _25246_ (.A0(_06421_),
    .A1(\cpu.icache.r_data[6][0] ),
    .S(_06505_),
    .X(_02193_));
 sg13g2_nand2_2 _25247_ (.Y(_06506_),
    .A(net570),
    .B(_06392_));
 sg13g2_mux2_1 _25248_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][10] ),
    .S(_06506_),
    .X(_02194_));
 sg13g2_mux2_1 _25249_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][11] ),
    .S(_06506_),
    .X(_02195_));
 sg13g2_nand2_2 _25250_ (.Y(_06507_),
    .A(net570),
    .B(_06398_));
 sg13g2_mux2_1 _25251_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][12] ),
    .S(_06507_),
    .X(_02196_));
 sg13g2_mux2_1 _25252_ (.A0(_06434_),
    .A1(\cpu.icache.r_data[6][13] ),
    .S(_06507_),
    .X(_02197_));
 sg13g2_mux2_1 _25253_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][14] ),
    .S(_06507_),
    .X(_02198_));
 sg13g2_mux2_1 _25254_ (.A0(_06430_),
    .A1(\cpu.icache.r_data[6][15] ),
    .S(_06507_),
    .X(_02199_));
 sg13g2_nand2_2 _25255_ (.Y(_06508_),
    .A(net570),
    .B(_06404_));
 sg13g2_mux2_1 _25256_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][16] ),
    .S(_06508_),
    .X(_02200_));
 sg13g2_mux2_1 _25257_ (.A0(_06434_),
    .A1(\cpu.icache.r_data[6][17] ),
    .S(_06508_),
    .X(_02201_));
 sg13g2_mux2_1 _25258_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][18] ),
    .S(_06508_),
    .X(_02202_));
 sg13g2_mux2_1 _25259_ (.A0(_06430_),
    .A1(\cpu.icache.r_data[6][19] ),
    .S(_06508_),
    .X(_02203_));
 sg13g2_mux2_1 _25260_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][1] ),
    .S(_06505_),
    .X(_02204_));
 sg13g2_nand2_2 _25261_ (.Y(_06509_),
    .A(net570),
    .B(_06408_));
 sg13g2_mux2_1 _25262_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][20] ),
    .S(_06509_),
    .X(_02205_));
 sg13g2_mux2_1 _25263_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][21] ),
    .S(_06509_),
    .X(_02206_));
 sg13g2_mux2_1 _25264_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][22] ),
    .S(_06509_),
    .X(_02207_));
 sg13g2_mux2_1 _25265_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][23] ),
    .S(_06509_),
    .X(_02208_));
 sg13g2_nand2_1 _25266_ (.Y(_06510_),
    .A(net570),
    .B(_06411_));
 sg13g2_buf_2 _25267_ (.A(_06510_),
    .X(_06511_));
 sg13g2_mux2_1 _25268_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][24] ),
    .S(_06511_),
    .X(_02209_));
 sg13g2_mux2_1 _25269_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][25] ),
    .S(_06511_),
    .X(_02210_));
 sg13g2_mux2_1 _25270_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][26] ),
    .S(_06511_),
    .X(_02211_));
 sg13g2_mux2_1 _25271_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][27] ),
    .S(_06511_),
    .X(_02212_));
 sg13g2_nand2_2 _25272_ (.Y(_06512_),
    .A(_08620_),
    .B(_06416_));
 sg13g2_mux2_1 _25273_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][28] ),
    .S(_06512_),
    .X(_02213_));
 sg13g2_mux2_1 _25274_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][29] ),
    .S(_06512_),
    .X(_02214_));
 sg13g2_mux2_1 _25275_ (.A0(_06426_),
    .A1(\cpu.icache.r_data[6][2] ),
    .S(_06505_),
    .X(_02215_));
 sg13g2_mux2_1 _25276_ (.A0(_06426_),
    .A1(\cpu.icache.r_data[6][30] ),
    .S(_06512_),
    .X(_02216_));
 sg13g2_mux2_1 _25277_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][31] ),
    .S(_06512_),
    .X(_02217_));
 sg13g2_mux2_1 _25278_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][3] ),
    .S(_06505_),
    .X(_02218_));
 sg13g2_nand2_2 _25279_ (.Y(_06513_),
    .A(_08620_),
    .B(_06419_));
 sg13g2_mux2_1 _25280_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][4] ),
    .S(_06513_),
    .X(_02219_));
 sg13g2_mux2_1 _25281_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][5] ),
    .S(_06513_),
    .X(_02220_));
 sg13g2_mux2_1 _25282_ (.A0(net970),
    .A1(\cpu.icache.r_data[6][6] ),
    .S(_06513_),
    .X(_02221_));
 sg13g2_mux2_1 _25283_ (.A0(net850),
    .A1(\cpu.icache.r_data[6][7] ),
    .S(_06513_),
    .X(_02222_));
 sg13g2_mux2_1 _25284_ (.A0(net851),
    .A1(\cpu.icache.r_data[6][8] ),
    .S(_06506_),
    .X(_02223_));
 sg13g2_mux2_1 _25285_ (.A0(net969),
    .A1(\cpu.icache.r_data[6][9] ),
    .S(_06506_),
    .X(_02224_));
 sg13g2_nand2_1 _25286_ (.Y(_06514_),
    .A(_08525_),
    .B(_08598_));
 sg13g2_buf_4 _25287_ (.X(_06515_),
    .A(_06514_));
 sg13g2_nor2_2 _25288_ (.A(_06515_),
    .B(_06424_),
    .Y(_06516_));
 sg13g2_mux2_1 _25289_ (.A0(\cpu.icache.r_data[7][0] ),
    .A1(_06495_),
    .S(_06516_),
    .X(_02225_));
 sg13g2_nor2_2 _25290_ (.A(_06515_),
    .B(_06428_),
    .Y(_06517_));
 sg13g2_mux2_1 _25291_ (.A0(\cpu.icache.r_data[7][10] ),
    .A1(net963),
    .S(_06517_),
    .X(_02226_));
 sg13g2_mux2_1 _25292_ (.A0(\cpu.icache.r_data[7][11] ),
    .A1(net962),
    .S(_06517_),
    .X(_02227_));
 sg13g2_nor2_2 _25293_ (.A(_06515_),
    .B(_06432_),
    .Y(_06518_));
 sg13g2_mux2_1 _25294_ (.A0(\cpu.icache.r_data[7][12] ),
    .A1(net964),
    .S(_06518_),
    .X(_02228_));
 sg13g2_mux2_1 _25295_ (.A0(\cpu.icache.r_data[7][13] ),
    .A1(_06499_),
    .S(_06518_),
    .X(_02229_));
 sg13g2_mux2_1 _25296_ (.A0(\cpu.icache.r_data[7][14] ),
    .A1(net963),
    .S(_06518_),
    .X(_02230_));
 sg13g2_mux2_1 _25297_ (.A0(\cpu.icache.r_data[7][15] ),
    .A1(_06498_),
    .S(_06518_),
    .X(_02231_));
 sg13g2_nor2_2 _25298_ (.A(_06515_),
    .B(_06437_),
    .Y(_06519_));
 sg13g2_mux2_1 _25299_ (.A0(\cpu.icache.r_data[7][16] ),
    .A1(_06495_),
    .S(_06519_),
    .X(_02232_));
 sg13g2_mux2_1 _25300_ (.A0(\cpu.icache.r_data[7][17] ),
    .A1(net961),
    .S(_06519_),
    .X(_02233_));
 sg13g2_mux2_1 _25301_ (.A0(\cpu.icache.r_data[7][18] ),
    .A1(_06497_),
    .S(_06519_),
    .X(_02234_));
 sg13g2_mux2_1 _25302_ (.A0(\cpu.icache.r_data[7][19] ),
    .A1(_06498_),
    .S(_06519_),
    .X(_02235_));
 sg13g2_mux2_1 _25303_ (.A0(\cpu.icache.r_data[7][1] ),
    .A1(net961),
    .S(_06516_),
    .X(_02236_));
 sg13g2_nor2_2 _25304_ (.A(_06515_),
    .B(_06440_),
    .Y(_06520_));
 sg13g2_mux2_1 _25305_ (.A0(\cpu.icache.r_data[7][20] ),
    .A1(net964),
    .S(_06520_),
    .X(_02237_));
 sg13g2_mux2_1 _25306_ (.A0(\cpu.icache.r_data[7][21] ),
    .A1(_06499_),
    .S(_06520_),
    .X(_02238_));
 sg13g2_mux2_1 _25307_ (.A0(\cpu.icache.r_data[7][22] ),
    .A1(net963),
    .S(_06520_),
    .X(_02239_));
 sg13g2_mux2_1 _25308_ (.A0(\cpu.icache.r_data[7][23] ),
    .A1(net962),
    .S(_06520_),
    .X(_02240_));
 sg13g2_nor2_1 _25309_ (.A(_06515_),
    .B(_06443_),
    .Y(_06521_));
 sg13g2_buf_2 _25310_ (.A(_06521_),
    .X(_06522_));
 sg13g2_mux2_1 _25311_ (.A0(\cpu.icache.r_data[7][24] ),
    .A1(net1023),
    .S(_06522_),
    .X(_02241_));
 sg13g2_mux2_1 _25312_ (.A0(\cpu.icache.r_data[7][25] ),
    .A1(net1018),
    .S(_06522_),
    .X(_02242_));
 sg13g2_mux2_1 _25313_ (.A0(\cpu.icache.r_data[7][26] ),
    .A1(net1027),
    .S(_06522_),
    .X(_02243_));
 sg13g2_mux2_1 _25314_ (.A0(\cpu.icache.r_data[7][27] ),
    .A1(net1026),
    .S(_06522_),
    .X(_02244_));
 sg13g2_nor2_2 _25315_ (.A(_06515_),
    .B(_06446_),
    .Y(_06523_));
 sg13g2_mux2_1 _25316_ (.A0(\cpu.icache.r_data[7][28] ),
    .A1(net1023),
    .S(_06523_),
    .X(_02245_));
 sg13g2_mux2_1 _25317_ (.A0(\cpu.icache.r_data[7][29] ),
    .A1(net1018),
    .S(_06523_),
    .X(_02246_));
 sg13g2_mux2_1 _25318_ (.A0(\cpu.icache.r_data[7][2] ),
    .A1(net1027),
    .S(_06516_),
    .X(_02247_));
 sg13g2_mux2_1 _25319_ (.A0(\cpu.icache.r_data[7][30] ),
    .A1(_12168_),
    .S(_06523_),
    .X(_02248_));
 sg13g2_mux2_1 _25320_ (.A0(\cpu.icache.r_data[7][31] ),
    .A1(net1026),
    .S(_06523_),
    .X(_02249_));
 sg13g2_mux2_1 _25321_ (.A0(\cpu.icache.r_data[7][3] ),
    .A1(_12185_),
    .S(_06516_),
    .X(_02250_));
 sg13g2_nor2_2 _25322_ (.A(_06515_),
    .B(_06448_),
    .Y(_06524_));
 sg13g2_mux2_1 _25323_ (.A0(\cpu.icache.r_data[7][4] ),
    .A1(_12251_),
    .S(_06524_),
    .X(_02251_));
 sg13g2_mux2_1 _25324_ (.A0(\cpu.icache.r_data[7][5] ),
    .A1(_12335_),
    .S(_06524_),
    .X(_02252_));
 sg13g2_mux2_1 _25325_ (.A0(\cpu.icache.r_data[7][6] ),
    .A1(_12168_),
    .S(_06524_),
    .X(_02253_));
 sg13g2_mux2_1 _25326_ (.A0(\cpu.icache.r_data[7][7] ),
    .A1(_12185_),
    .S(_06524_),
    .X(_02254_));
 sg13g2_mux2_1 _25327_ (.A0(\cpu.icache.r_data[7][8] ),
    .A1(_12251_),
    .S(_06517_),
    .X(_02255_));
 sg13g2_mux2_1 _25328_ (.A0(\cpu.icache.r_data[7][9] ),
    .A1(_12335_),
    .S(_06517_),
    .X(_02256_));
 sg13g2_mux2_1 _25329_ (.A0(net988),
    .A1(\cpu.icache.r_tag[0][5] ),
    .S(net368),
    .X(_02260_));
 sg13g2_buf_1 _25330_ (.A(net405),
    .X(_06525_));
 sg13g2_buf_1 _25331_ (.A(_06412_),
    .X(_06526_));
 sg13g2_nand2_1 _25332_ (.Y(_06527_),
    .A(\cpu.icache.r_tag[0][15] ),
    .B(net404));
 sg13g2_o21ai_1 _25333_ (.B1(_06527_),
    .Y(_02261_),
    .A1(_08733_),
    .A2(_06525_));
 sg13g2_nand2_1 _25334_ (.Y(_06528_),
    .A(\cpu.icache.r_tag[0][16] ),
    .B(_06526_));
 sg13g2_o21ai_1 _25335_ (.B1(_06528_),
    .Y(_02262_),
    .A1(net396),
    .A2(net366));
 sg13g2_nand2_1 _25336_ (.Y(_06529_),
    .A(\cpu.icache.r_tag[0][17] ),
    .B(net404));
 sg13g2_o21ai_1 _25337_ (.B1(_06529_),
    .Y(_02263_),
    .A1(net395),
    .A2(net366));
 sg13g2_nand2_1 _25338_ (.Y(_06530_),
    .A(\cpu.icache.r_tag[0][18] ),
    .B(net404));
 sg13g2_o21ai_1 _25339_ (.B1(_06530_),
    .Y(_02264_),
    .A1(net447),
    .A2(net366));
 sg13g2_nand2_1 _25340_ (.Y(_06531_),
    .A(\cpu.icache.r_tag[0][19] ),
    .B(_06526_));
 sg13g2_o21ai_1 _25341_ (.B1(_06531_),
    .Y(_02265_),
    .A1(net392),
    .A2(net366));
 sg13g2_nand2_1 _25342_ (.Y(_06532_),
    .A(\cpu.icache.r_tag[0][20] ),
    .B(net404));
 sg13g2_o21ai_1 _25343_ (.B1(_06532_),
    .Y(_02266_),
    .A1(net393),
    .A2(net366));
 sg13g2_nand2_1 _25344_ (.Y(_06533_),
    .A(\cpu.icache.r_tag[0][21] ),
    .B(net405));
 sg13g2_o21ai_1 _25345_ (.B1(_06533_),
    .Y(_02267_),
    .A1(net398),
    .A2(net366));
 sg13g2_nand2_1 _25346_ (.Y(_06534_),
    .A(\cpu.icache.r_tag[0][22] ),
    .B(net405));
 sg13g2_o21ai_1 _25347_ (.B1(_06534_),
    .Y(_02268_),
    .A1(net397),
    .A2(net366));
 sg13g2_nand2_1 _25348_ (.Y(_06535_),
    .A(\cpu.icache.r_tag[0][23] ),
    .B(net405));
 sg13g2_o21ai_1 _25349_ (.B1(_06535_),
    .Y(_02269_),
    .A1(net496),
    .A2(net366));
 sg13g2_mux2_1 _25350_ (.A0(net987),
    .A1(\cpu.icache.r_tag[0][6] ),
    .S(net404),
    .X(_02270_));
 sg13g2_mux2_1 _25351_ (.A0(net986),
    .A1(\cpu.icache.r_tag[0][7] ),
    .S(net404),
    .X(_02271_));
 sg13g2_nand2_1 _25352_ (.Y(_06536_),
    .A(\cpu.icache.r_tag[0][8] ),
    .B(net405));
 sg13g2_o21ai_1 _25353_ (.B1(_06536_),
    .Y(_02272_),
    .A1(net990),
    .A2(net368));
 sg13g2_mux2_1 _25354_ (.A0(net985),
    .A1(\cpu.icache.r_tag[0][9] ),
    .S(net404),
    .X(_02273_));
 sg13g2_mux2_1 _25355_ (.A0(net984),
    .A1(\cpu.icache.r_tag[0][10] ),
    .S(net404),
    .X(_02274_));
 sg13g2_nand2_1 _25356_ (.Y(_06537_),
    .A(\cpu.icache.r_tag[0][11] ),
    .B(net405));
 sg13g2_o21ai_1 _25357_ (.B1(_06537_),
    .Y(_02275_),
    .A1(net989),
    .A2(net368));
 sg13g2_nand2_1 _25358_ (.Y(_06538_),
    .A(\cpu.icache.r_tag[0][12] ),
    .B(_06413_));
 sg13g2_o21ai_1 _25359_ (.B1(_06538_),
    .Y(_02276_),
    .A1(net399),
    .A2(net368));
 sg13g2_nand2_1 _25360_ (.Y(_06539_),
    .A(\cpu.icache.r_tag[0][13] ),
    .B(_06413_));
 sg13g2_o21ai_1 _25361_ (.B1(_06539_),
    .Y(_02277_),
    .A1(net400),
    .A2(net368));
 sg13g2_nand2_1 _25362_ (.Y(_06540_),
    .A(\cpu.icache.r_tag[0][14] ),
    .B(net405));
 sg13g2_o21ai_1 _25363_ (.B1(_06540_),
    .Y(_02278_),
    .A1(net394),
    .A2(net368));
 sg13g2_nor2b_1 _25364_ (.A(_06391_),
    .B_N(_06402_),
    .Y(_06541_));
 sg13g2_buf_1 _25365_ (.A(_06541_),
    .X(_06542_));
 sg13g2_nand2_1 _25366_ (.Y(_06543_),
    .A(net495),
    .B(_06542_));
 sg13g2_buf_1 _25367_ (.A(_06543_),
    .X(_06544_));
 sg13g2_buf_1 _25368_ (.A(_06544_),
    .X(_06545_));
 sg13g2_mux2_1 _25369_ (.A0(net988),
    .A1(\cpu.icache.r_tag[1][5] ),
    .S(net311),
    .X(_02279_));
 sg13g2_buf_1 _25370_ (.A(_06544_),
    .X(_06546_));
 sg13g2_nand2_1 _25371_ (.Y(_06547_),
    .A(\cpu.icache.r_tag[1][15] ),
    .B(net311));
 sg13g2_o21ai_1 _25372_ (.B1(_06547_),
    .Y(_02280_),
    .A1(net448),
    .A2(_06546_));
 sg13g2_buf_1 _25373_ (.A(_06544_),
    .X(_06548_));
 sg13g2_nand2_1 _25374_ (.Y(_06549_),
    .A(\cpu.icache.r_tag[1][16] ),
    .B(net309));
 sg13g2_o21ai_1 _25375_ (.B1(_06549_),
    .Y(_02281_),
    .A1(net396),
    .A2(net310));
 sg13g2_nand2_1 _25376_ (.Y(_06550_),
    .A(\cpu.icache.r_tag[1][17] ),
    .B(_06548_));
 sg13g2_o21ai_1 _25377_ (.B1(_06550_),
    .Y(_02282_),
    .A1(net395),
    .A2(net310));
 sg13g2_nand2_1 _25378_ (.Y(_06551_),
    .A(\cpu.icache.r_tag[1][18] ),
    .B(net309));
 sg13g2_o21ai_1 _25379_ (.B1(_06551_),
    .Y(_02283_),
    .A1(_08757_),
    .A2(_06546_));
 sg13g2_nand2_1 _25380_ (.Y(_06552_),
    .A(\cpu.icache.r_tag[1][19] ),
    .B(net309));
 sg13g2_o21ai_1 _25381_ (.B1(_06552_),
    .Y(_02284_),
    .A1(net392),
    .A2(net310));
 sg13g2_nand2_1 _25382_ (.Y(_06553_),
    .A(\cpu.icache.r_tag[1][20] ),
    .B(net309));
 sg13g2_o21ai_1 _25383_ (.B1(_06553_),
    .Y(_02285_),
    .A1(net393),
    .A2(net310));
 sg13g2_nand2_1 _25384_ (.Y(_06554_),
    .A(\cpu.icache.r_tag[1][21] ),
    .B(_06548_));
 sg13g2_o21ai_1 _25385_ (.B1(_06554_),
    .Y(_02286_),
    .A1(net398),
    .A2(net310));
 sg13g2_nand2_1 _25386_ (.Y(_06555_),
    .A(\cpu.icache.r_tag[1][22] ),
    .B(net309));
 sg13g2_o21ai_1 _25387_ (.B1(_06555_),
    .Y(_02287_),
    .A1(net397),
    .A2(net310));
 sg13g2_nand2_1 _25388_ (.Y(_06556_),
    .A(\cpu.icache.r_tag[1][23] ),
    .B(net309));
 sg13g2_o21ai_1 _25389_ (.B1(_06556_),
    .Y(_02288_),
    .A1(net496),
    .A2(net310));
 sg13g2_mux2_1 _25390_ (.A0(net987),
    .A1(\cpu.icache.r_tag[1][6] ),
    .S(net311),
    .X(_02289_));
 sg13g2_mux2_1 _25391_ (.A0(net986),
    .A1(\cpu.icache.r_tag[1][7] ),
    .S(net311),
    .X(_02290_));
 sg13g2_nand2_1 _25392_ (.Y(_06557_),
    .A(\cpu.icache.r_tag[1][8] ),
    .B(net309));
 sg13g2_o21ai_1 _25393_ (.B1(_06557_),
    .Y(_02291_),
    .A1(net990),
    .A2(net310));
 sg13g2_mux2_1 _25394_ (.A0(net985),
    .A1(\cpu.icache.r_tag[1][9] ),
    .S(net311),
    .X(_02292_));
 sg13g2_mux2_1 _25395_ (.A0(net984),
    .A1(\cpu.icache.r_tag[1][10] ),
    .S(net311),
    .X(_02293_));
 sg13g2_nand2_1 _25396_ (.Y(_06558_),
    .A(\cpu.icache.r_tag[1][11] ),
    .B(net309));
 sg13g2_o21ai_1 _25397_ (.B1(_06558_),
    .Y(_02294_),
    .A1(net989),
    .A2(net311));
 sg13g2_nand2_1 _25398_ (.Y(_06559_),
    .A(\cpu.icache.r_tag[1][12] ),
    .B(_06544_));
 sg13g2_o21ai_1 _25399_ (.B1(_06559_),
    .Y(_02295_),
    .A1(net399),
    .A2(net311));
 sg13g2_nand2_1 _25400_ (.Y(_06560_),
    .A(\cpu.icache.r_tag[1][13] ),
    .B(_06544_));
 sg13g2_o21ai_1 _25401_ (.B1(_06560_),
    .Y(_02296_),
    .A1(net400),
    .A2(_06545_));
 sg13g2_nand2_1 _25402_ (.Y(_06561_),
    .A(\cpu.icache.r_tag[1][14] ),
    .B(_06544_));
 sg13g2_o21ai_1 _25403_ (.B1(_06561_),
    .Y(_02297_),
    .A1(net394),
    .A2(_06545_));
 sg13g2_nand2_1 _25404_ (.Y(_06562_),
    .A(net494),
    .B(_06542_));
 sg13g2_buf_1 _25405_ (.A(_06562_),
    .X(_06563_));
 sg13g2_buf_1 _25406_ (.A(_06563_),
    .X(_06564_));
 sg13g2_mux2_1 _25407_ (.A0(net988),
    .A1(\cpu.icache.r_tag[2][5] ),
    .S(net308),
    .X(_02298_));
 sg13g2_buf_1 _25408_ (.A(_06563_),
    .X(_06565_));
 sg13g2_nand2_1 _25409_ (.Y(_06566_),
    .A(\cpu.icache.r_tag[2][15] ),
    .B(_06564_));
 sg13g2_o21ai_1 _25410_ (.B1(_06566_),
    .Y(_02299_),
    .A1(net448),
    .A2(net307));
 sg13g2_buf_1 _25411_ (.A(_06563_),
    .X(_06567_));
 sg13g2_nand2_1 _25412_ (.Y(_06568_),
    .A(\cpu.icache.r_tag[2][16] ),
    .B(net306));
 sg13g2_o21ai_1 _25413_ (.B1(_06568_),
    .Y(_02300_),
    .A1(net396),
    .A2(net307));
 sg13g2_nand2_1 _25414_ (.Y(_06569_),
    .A(\cpu.icache.r_tag[2][17] ),
    .B(net306));
 sg13g2_o21ai_1 _25415_ (.B1(_06569_),
    .Y(_02301_),
    .A1(net395),
    .A2(net307));
 sg13g2_nand2_1 _25416_ (.Y(_06570_),
    .A(\cpu.icache.r_tag[2][18] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25417_ (.B1(_06570_),
    .Y(_02302_),
    .A1(net447),
    .A2(net307));
 sg13g2_nand2_1 _25418_ (.Y(_06571_),
    .A(\cpu.icache.r_tag[2][19] ),
    .B(net306));
 sg13g2_o21ai_1 _25419_ (.B1(_06571_),
    .Y(_02303_),
    .A1(_08712_),
    .A2(_06565_));
 sg13g2_nand2_1 _25420_ (.Y(_06572_),
    .A(\cpu.icache.r_tag[2][20] ),
    .B(net306));
 sg13g2_o21ai_1 _25421_ (.B1(_06572_),
    .Y(_02304_),
    .A1(_08692_),
    .A2(net307));
 sg13g2_nand2_1 _25422_ (.Y(_06573_),
    .A(\cpu.icache.r_tag[2][21] ),
    .B(net306));
 sg13g2_o21ai_1 _25423_ (.B1(_06573_),
    .Y(_02305_),
    .A1(net398),
    .A2(net307));
 sg13g2_nand2_1 _25424_ (.Y(_06574_),
    .A(\cpu.icache.r_tag[2][22] ),
    .B(net306));
 sg13g2_o21ai_1 _25425_ (.B1(_06574_),
    .Y(_02306_),
    .A1(net397),
    .A2(net307));
 sg13g2_nand2_1 _25426_ (.Y(_06575_),
    .A(\cpu.icache.r_tag[2][23] ),
    .B(net306));
 sg13g2_o21ai_1 _25427_ (.B1(_06575_),
    .Y(_02307_),
    .A1(net496),
    .A2(net307));
 sg13g2_mux2_1 _25428_ (.A0(net987),
    .A1(\cpu.icache.r_tag[2][6] ),
    .S(net308),
    .X(_02308_));
 sg13g2_mux2_1 _25429_ (.A0(net986),
    .A1(\cpu.icache.r_tag[2][7] ),
    .S(net308),
    .X(_02309_));
 sg13g2_nand2_1 _25430_ (.Y(_06576_),
    .A(\cpu.icache.r_tag[2][8] ),
    .B(net306));
 sg13g2_o21ai_1 _25431_ (.B1(_06576_),
    .Y(_02310_),
    .A1(net990),
    .A2(_06565_));
 sg13g2_mux2_1 _25432_ (.A0(net985),
    .A1(\cpu.icache.r_tag[2][9] ),
    .S(net308),
    .X(_02311_));
 sg13g2_mux2_1 _25433_ (.A0(net984),
    .A1(\cpu.icache.r_tag[2][10] ),
    .S(net308),
    .X(_02312_));
 sg13g2_nand2_1 _25434_ (.Y(_06577_),
    .A(\cpu.icache.r_tag[2][11] ),
    .B(_06567_));
 sg13g2_o21ai_1 _25435_ (.B1(_06577_),
    .Y(_02313_),
    .A1(net989),
    .A2(net308));
 sg13g2_nand2_1 _25436_ (.Y(_06578_),
    .A(\cpu.icache.r_tag[2][12] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25437_ (.B1(_06578_),
    .Y(_02314_),
    .A1(net399),
    .A2(net308));
 sg13g2_nand2_1 _25438_ (.Y(_06579_),
    .A(\cpu.icache.r_tag[2][13] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25439_ (.B1(_06579_),
    .Y(_02315_),
    .A1(net400),
    .A2(net308));
 sg13g2_nand2_1 _25440_ (.Y(_06580_),
    .A(\cpu.icache.r_tag[2][14] ),
    .B(_06563_));
 sg13g2_o21ai_1 _25441_ (.B1(_06580_),
    .Y(_02316_),
    .A1(net394),
    .A2(_06564_));
 sg13g2_mux2_1 _25442_ (.A0(net988),
    .A1(\cpu.icache.r_tag[3][5] ),
    .S(net312),
    .X(_02317_));
 sg13g2_buf_1 _25443_ (.A(net367),
    .X(_06581_));
 sg13g2_buf_1 _25444_ (.A(_06475_),
    .X(_06582_));
 sg13g2_nand2_1 _25445_ (.Y(_06583_),
    .A(\cpu.icache.r_tag[3][15] ),
    .B(net365));
 sg13g2_o21ai_1 _25446_ (.B1(_06583_),
    .Y(_02318_),
    .A1(net448),
    .A2(net305));
 sg13g2_nand2_1 _25447_ (.Y(_06584_),
    .A(\cpu.icache.r_tag[3][16] ),
    .B(net365));
 sg13g2_o21ai_1 _25448_ (.B1(_06584_),
    .Y(_02319_),
    .A1(net396),
    .A2(net305));
 sg13g2_nand2_1 _25449_ (.Y(_06585_),
    .A(\cpu.icache.r_tag[3][17] ),
    .B(net365));
 sg13g2_o21ai_1 _25450_ (.B1(_06585_),
    .Y(_02320_),
    .A1(net395),
    .A2(_06581_));
 sg13g2_nand2_1 _25451_ (.Y(_06586_),
    .A(\cpu.icache.r_tag[3][18] ),
    .B(net365));
 sg13g2_o21ai_1 _25452_ (.B1(_06586_),
    .Y(_02321_),
    .A1(net447),
    .A2(net305));
 sg13g2_nand2_1 _25453_ (.Y(_06587_),
    .A(\cpu.icache.r_tag[3][19] ),
    .B(net365));
 sg13g2_o21ai_1 _25454_ (.B1(_06587_),
    .Y(_02322_),
    .A1(net392),
    .A2(_06581_));
 sg13g2_nand2_1 _25455_ (.Y(_06588_),
    .A(\cpu.icache.r_tag[3][20] ),
    .B(net365));
 sg13g2_o21ai_1 _25456_ (.B1(_06588_),
    .Y(_02323_),
    .A1(net393),
    .A2(net305));
 sg13g2_nand2_1 _25457_ (.Y(_06589_),
    .A(\cpu.icache.r_tag[3][21] ),
    .B(net367));
 sg13g2_o21ai_1 _25458_ (.B1(_06589_),
    .Y(_02324_),
    .A1(net398),
    .A2(net305));
 sg13g2_nand2_1 _25459_ (.Y(_06590_),
    .A(\cpu.icache.r_tag[3][22] ),
    .B(net367));
 sg13g2_o21ai_1 _25460_ (.B1(_06590_),
    .Y(_02325_),
    .A1(net397),
    .A2(net305));
 sg13g2_nand2_1 _25461_ (.Y(_06591_),
    .A(\cpu.icache.r_tag[3][23] ),
    .B(net367));
 sg13g2_o21ai_1 _25462_ (.B1(_06591_),
    .Y(_02326_),
    .A1(net496),
    .A2(net305));
 sg13g2_mux2_1 _25463_ (.A0(net987),
    .A1(\cpu.icache.r_tag[3][6] ),
    .S(net365),
    .X(_02327_));
 sg13g2_mux2_1 _25464_ (.A0(net986),
    .A1(\cpu.icache.r_tag[3][7] ),
    .S(net365),
    .X(_02328_));
 sg13g2_nand2_1 _25465_ (.Y(_06592_),
    .A(\cpu.icache.r_tag[3][8] ),
    .B(net367));
 sg13g2_o21ai_1 _25466_ (.B1(_06592_),
    .Y(_02329_),
    .A1(net990),
    .A2(net312));
 sg13g2_mux2_1 _25467_ (.A0(net985),
    .A1(\cpu.icache.r_tag[3][9] ),
    .S(_06582_),
    .X(_02330_));
 sg13g2_mux2_1 _25468_ (.A0(net984),
    .A1(\cpu.icache.r_tag[3][10] ),
    .S(_06582_),
    .X(_02331_));
 sg13g2_nand2_1 _25469_ (.Y(_06593_),
    .A(\cpu.icache.r_tag[3][11] ),
    .B(net367));
 sg13g2_o21ai_1 _25470_ (.B1(_06593_),
    .Y(_02332_),
    .A1(net989),
    .A2(net312));
 sg13g2_nand2_1 _25471_ (.Y(_06594_),
    .A(\cpu.icache.r_tag[3][12] ),
    .B(net367));
 sg13g2_o21ai_1 _25472_ (.B1(_06594_),
    .Y(_02333_),
    .A1(net399),
    .A2(net312));
 sg13g2_nand2_1 _25473_ (.Y(_06595_),
    .A(\cpu.icache.r_tag[3][13] ),
    .B(net367));
 sg13g2_o21ai_1 _25474_ (.B1(_06595_),
    .Y(_02334_),
    .A1(net400),
    .A2(net312));
 sg13g2_nand2_1 _25475_ (.Y(_06596_),
    .A(\cpu.icache.r_tag[3][14] ),
    .B(_06476_));
 sg13g2_o21ai_1 _25476_ (.B1(_06596_),
    .Y(_02335_),
    .A1(net394),
    .A2(net312));
 sg13g2_nand2_1 _25477_ (.Y(_06597_),
    .A(net619),
    .B(_06542_));
 sg13g2_buf_1 _25478_ (.A(_06597_),
    .X(_06598_));
 sg13g2_buf_1 _25479_ (.A(_06598_),
    .X(_06599_));
 sg13g2_mux2_1 _25480_ (.A0(net988),
    .A1(\cpu.icache.r_tag[4][5] ),
    .S(net403),
    .X(_02336_));
 sg13g2_buf_1 _25481_ (.A(_06598_),
    .X(_06600_));
 sg13g2_nand2_1 _25482_ (.Y(_06601_),
    .A(\cpu.icache.r_tag[4][15] ),
    .B(_06599_));
 sg13g2_o21ai_1 _25483_ (.B1(_06601_),
    .Y(_02337_),
    .A1(net448),
    .A2(net402));
 sg13g2_buf_1 _25484_ (.A(_06598_),
    .X(_06602_));
 sg13g2_nand2_1 _25485_ (.Y(_06603_),
    .A(\cpu.icache.r_tag[4][16] ),
    .B(net401));
 sg13g2_o21ai_1 _25486_ (.B1(_06603_),
    .Y(_02338_),
    .A1(net396),
    .A2(net402));
 sg13g2_nand2_1 _25487_ (.Y(_06604_),
    .A(\cpu.icache.r_tag[4][17] ),
    .B(net401));
 sg13g2_o21ai_1 _25488_ (.B1(_06604_),
    .Y(_02339_),
    .A1(net395),
    .A2(net402));
 sg13g2_nand2_1 _25489_ (.Y(_06605_),
    .A(\cpu.icache.r_tag[4][18] ),
    .B(_06602_));
 sg13g2_o21ai_1 _25490_ (.B1(_06605_),
    .Y(_02340_),
    .A1(net447),
    .A2(_06600_));
 sg13g2_nand2_1 _25491_ (.Y(_06606_),
    .A(\cpu.icache.r_tag[4][19] ),
    .B(net401));
 sg13g2_o21ai_1 _25492_ (.B1(_06606_),
    .Y(_02341_),
    .A1(net392),
    .A2(net402));
 sg13g2_nand2_1 _25493_ (.Y(_06607_),
    .A(\cpu.icache.r_tag[4][20] ),
    .B(net401));
 sg13g2_o21ai_1 _25494_ (.B1(_06607_),
    .Y(_02342_),
    .A1(net393),
    .A2(net402));
 sg13g2_nand2_1 _25495_ (.Y(_06608_),
    .A(\cpu.icache.r_tag[4][21] ),
    .B(net401));
 sg13g2_o21ai_1 _25496_ (.B1(_06608_),
    .Y(_02343_),
    .A1(net398),
    .A2(net402));
 sg13g2_nand2_1 _25497_ (.Y(_06609_),
    .A(\cpu.icache.r_tag[4][22] ),
    .B(net401));
 sg13g2_o21ai_1 _25498_ (.B1(_06609_),
    .Y(_02344_),
    .A1(_08591_),
    .A2(net402));
 sg13g2_nand2_1 _25499_ (.Y(_06610_),
    .A(\cpu.icache.r_tag[4][23] ),
    .B(net401));
 sg13g2_o21ai_1 _25500_ (.B1(_06610_),
    .Y(_02345_),
    .A1(net496),
    .A2(_06600_));
 sg13g2_mux2_1 _25501_ (.A0(net987),
    .A1(\cpu.icache.r_tag[4][6] ),
    .S(net403),
    .X(_02346_));
 sg13g2_mux2_1 _25502_ (.A0(net986),
    .A1(\cpu.icache.r_tag[4][7] ),
    .S(net403),
    .X(_02347_));
 sg13g2_nand2_1 _25503_ (.Y(_06611_),
    .A(\cpu.icache.r_tag[4][8] ),
    .B(net401));
 sg13g2_o21ai_1 _25504_ (.B1(_06611_),
    .Y(_02348_),
    .A1(net990),
    .A2(net402));
 sg13g2_mux2_1 _25505_ (.A0(net985),
    .A1(\cpu.icache.r_tag[4][9] ),
    .S(net403),
    .X(_02349_));
 sg13g2_mux2_1 _25506_ (.A0(net984),
    .A1(\cpu.icache.r_tag[4][10] ),
    .S(net403),
    .X(_02350_));
 sg13g2_nand2_1 _25507_ (.Y(_06612_),
    .A(\cpu.icache.r_tag[4][11] ),
    .B(_06602_));
 sg13g2_o21ai_1 _25508_ (.B1(_06612_),
    .Y(_02351_),
    .A1(net989),
    .A2(net403));
 sg13g2_nand2_1 _25509_ (.Y(_06613_),
    .A(\cpu.icache.r_tag[4][12] ),
    .B(_06598_));
 sg13g2_o21ai_1 _25510_ (.B1(_06613_),
    .Y(_02352_),
    .A1(net399),
    .A2(net403));
 sg13g2_nand2_1 _25511_ (.Y(_06614_),
    .A(\cpu.icache.r_tag[4][13] ),
    .B(_06598_));
 sg13g2_o21ai_1 _25512_ (.B1(_06614_),
    .Y(_02353_),
    .A1(net400),
    .A2(net403));
 sg13g2_nand2_1 _25513_ (.Y(_06615_),
    .A(\cpu.icache.r_tag[4][14] ),
    .B(_06598_));
 sg13g2_o21ai_1 _25514_ (.B1(_06615_),
    .Y(_02354_),
    .A1(net394),
    .A2(_06599_));
 sg13g2_nand2_1 _25515_ (.Y(_06616_),
    .A(net571),
    .B(_06542_));
 sg13g2_buf_1 _25516_ (.A(_06616_),
    .X(_06617_));
 sg13g2_buf_1 _25517_ (.A(_06617_),
    .X(_06618_));
 sg13g2_mux2_1 _25518_ (.A0(net988),
    .A1(\cpu.icache.r_tag[5][5] ),
    .S(net364),
    .X(_02355_));
 sg13g2_buf_1 _25519_ (.A(_06617_),
    .X(_06619_));
 sg13g2_nand2_1 _25520_ (.Y(_06620_),
    .A(\cpu.icache.r_tag[5][15] ),
    .B(net364));
 sg13g2_o21ai_1 _25521_ (.B1(_06620_),
    .Y(_02356_),
    .A1(net448),
    .A2(net363));
 sg13g2_buf_1 _25522_ (.A(_06617_),
    .X(_06621_));
 sg13g2_nand2_1 _25523_ (.Y(_06622_),
    .A(\cpu.icache.r_tag[5][16] ),
    .B(net362));
 sg13g2_o21ai_1 _25524_ (.B1(_06622_),
    .Y(_02357_),
    .A1(net396),
    .A2(net363));
 sg13g2_nand2_1 _25525_ (.Y(_06623_),
    .A(\cpu.icache.r_tag[5][17] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25526_ (.B1(_06623_),
    .Y(_02358_),
    .A1(net395),
    .A2(_06619_));
 sg13g2_nand2_1 _25527_ (.Y(_06624_),
    .A(\cpu.icache.r_tag[5][18] ),
    .B(net362));
 sg13g2_o21ai_1 _25528_ (.B1(_06624_),
    .Y(_02359_),
    .A1(net447),
    .A2(net363));
 sg13g2_nand2_1 _25529_ (.Y(_06625_),
    .A(\cpu.icache.r_tag[5][19] ),
    .B(net362));
 sg13g2_o21ai_1 _25530_ (.B1(_06625_),
    .Y(_02360_),
    .A1(net392),
    .A2(net363));
 sg13g2_nand2_1 _25531_ (.Y(_06626_),
    .A(\cpu.icache.r_tag[5][20] ),
    .B(net362));
 sg13g2_o21ai_1 _25532_ (.B1(_06626_),
    .Y(_02361_),
    .A1(net393),
    .A2(net363));
 sg13g2_nand2_1 _25533_ (.Y(_06627_),
    .A(\cpu.icache.r_tag[5][21] ),
    .B(net362));
 sg13g2_o21ai_1 _25534_ (.B1(_06627_),
    .Y(_02362_),
    .A1(net398),
    .A2(net363));
 sg13g2_nand2_1 _25535_ (.Y(_06628_),
    .A(\cpu.icache.r_tag[5][22] ),
    .B(net362));
 sg13g2_o21ai_1 _25536_ (.B1(_06628_),
    .Y(_02363_),
    .A1(net397),
    .A2(net363));
 sg13g2_nand2_1 _25537_ (.Y(_06629_),
    .A(\cpu.icache.r_tag[5][23] ),
    .B(net362));
 sg13g2_o21ai_1 _25538_ (.B1(_06629_),
    .Y(_02364_),
    .A1(net496),
    .A2(_06619_));
 sg13g2_mux2_1 _25539_ (.A0(net987),
    .A1(\cpu.icache.r_tag[5][6] ),
    .S(net364),
    .X(_02365_));
 sg13g2_mux2_1 _25540_ (.A0(net986),
    .A1(\cpu.icache.r_tag[5][7] ),
    .S(net364),
    .X(_02366_));
 sg13g2_nand2_1 _25541_ (.Y(_06630_),
    .A(\cpu.icache.r_tag[5][8] ),
    .B(net362));
 sg13g2_o21ai_1 _25542_ (.B1(_06630_),
    .Y(_02367_),
    .A1(net990),
    .A2(net363));
 sg13g2_mux2_1 _25543_ (.A0(net985),
    .A1(\cpu.icache.r_tag[5][9] ),
    .S(net364),
    .X(_02368_));
 sg13g2_mux2_1 _25544_ (.A0(net984),
    .A1(\cpu.icache.r_tag[5][10] ),
    .S(net364),
    .X(_02369_));
 sg13g2_nand2_1 _25545_ (.Y(_06631_),
    .A(\cpu.icache.r_tag[5][11] ),
    .B(_06621_));
 sg13g2_o21ai_1 _25546_ (.B1(_06631_),
    .Y(_02370_),
    .A1(net989),
    .A2(net364));
 sg13g2_nand2_1 _25547_ (.Y(_06632_),
    .A(\cpu.icache.r_tag[5][12] ),
    .B(_06617_));
 sg13g2_o21ai_1 _25548_ (.B1(_06632_),
    .Y(_02371_),
    .A1(net399),
    .A2(net364));
 sg13g2_nand2_1 _25549_ (.Y(_06633_),
    .A(\cpu.icache.r_tag[5][13] ),
    .B(_06617_));
 sg13g2_o21ai_1 _25550_ (.B1(_06633_),
    .Y(_02372_),
    .A1(net400),
    .A2(_06618_));
 sg13g2_nand2_1 _25551_ (.Y(_06634_),
    .A(\cpu.icache.r_tag[5][14] ),
    .B(_06617_));
 sg13g2_o21ai_1 _25552_ (.B1(_06634_),
    .Y(_02373_),
    .A1(net394),
    .A2(_06618_));
 sg13g2_nand2_1 _25553_ (.Y(_06635_),
    .A(net570),
    .B(_06542_));
 sg13g2_buf_1 _25554_ (.A(_06635_),
    .X(_06636_));
 sg13g2_buf_1 _25555_ (.A(_06636_),
    .X(_06637_));
 sg13g2_mux2_1 _25556_ (.A0(_04577_),
    .A1(\cpu.icache.r_tag[6][5] ),
    .S(net361),
    .X(_02374_));
 sg13g2_buf_1 _25557_ (.A(_06636_),
    .X(_06638_));
 sg13g2_nand2_1 _25558_ (.Y(_06639_),
    .A(\cpu.icache.r_tag[6][15] ),
    .B(_06637_));
 sg13g2_o21ai_1 _25559_ (.B1(_06639_),
    .Y(_02375_),
    .A1(net448),
    .A2(net360));
 sg13g2_buf_1 _25560_ (.A(_06636_),
    .X(_06640_));
 sg13g2_nand2_1 _25561_ (.Y(_06641_),
    .A(\cpu.icache.r_tag[6][16] ),
    .B(net359));
 sg13g2_o21ai_1 _25562_ (.B1(_06641_),
    .Y(_02376_),
    .A1(net396),
    .A2(net360));
 sg13g2_nand2_1 _25563_ (.Y(_06642_),
    .A(\cpu.icache.r_tag[6][17] ),
    .B(net359));
 sg13g2_o21ai_1 _25564_ (.B1(_06642_),
    .Y(_02377_),
    .A1(net395),
    .A2(net360));
 sg13g2_nand2_1 _25565_ (.Y(_06643_),
    .A(\cpu.icache.r_tag[6][18] ),
    .B(net359));
 sg13g2_o21ai_1 _25566_ (.B1(_06643_),
    .Y(_02378_),
    .A1(net447),
    .A2(_06638_));
 sg13g2_nand2_1 _25567_ (.Y(_06644_),
    .A(\cpu.icache.r_tag[6][19] ),
    .B(net359));
 sg13g2_o21ai_1 _25568_ (.B1(_06644_),
    .Y(_02379_),
    .A1(net392),
    .A2(net360));
 sg13g2_nand2_1 _25569_ (.Y(_06645_),
    .A(\cpu.icache.r_tag[6][20] ),
    .B(net359));
 sg13g2_o21ai_1 _25570_ (.B1(_06645_),
    .Y(_02380_),
    .A1(net393),
    .A2(net360));
 sg13g2_nand2_1 _25571_ (.Y(_06646_),
    .A(\cpu.icache.r_tag[6][21] ),
    .B(net359));
 sg13g2_o21ai_1 _25572_ (.B1(_06646_),
    .Y(_02381_),
    .A1(_08563_),
    .A2(net360));
 sg13g2_nand2_1 _25573_ (.Y(_06647_),
    .A(\cpu.icache.r_tag[6][22] ),
    .B(net359));
 sg13g2_o21ai_1 _25574_ (.B1(_06647_),
    .Y(_02382_),
    .A1(net397),
    .A2(net360));
 sg13g2_nand2_1 _25575_ (.Y(_06648_),
    .A(\cpu.icache.r_tag[6][23] ),
    .B(net359));
 sg13g2_o21ai_1 _25576_ (.B1(_06648_),
    .Y(_02383_),
    .A1(net496),
    .A2(net360));
 sg13g2_mux2_1 _25577_ (.A0(_04611_),
    .A1(\cpu.icache.r_tag[6][6] ),
    .S(net361),
    .X(_02384_));
 sg13g2_mux2_1 _25578_ (.A0(_04639_),
    .A1(\cpu.icache.r_tag[6][7] ),
    .S(net361),
    .X(_02385_));
 sg13g2_nand2_1 _25579_ (.Y(_06649_),
    .A(\cpu.icache.r_tag[6][8] ),
    .B(_06640_));
 sg13g2_o21ai_1 _25580_ (.B1(_06649_),
    .Y(_02386_),
    .A1(_04222_),
    .A2(_06638_));
 sg13g2_mux2_1 _25581_ (.A0(_04713_),
    .A1(\cpu.icache.r_tag[6][9] ),
    .S(net361),
    .X(_02387_));
 sg13g2_mux2_1 _25582_ (.A0(_04750_),
    .A1(\cpu.icache.r_tag[6][10] ),
    .S(net361),
    .X(_02388_));
 sg13g2_nand2_1 _25583_ (.Y(_06650_),
    .A(\cpu.icache.r_tag[6][11] ),
    .B(_06640_));
 sg13g2_o21ai_1 _25584_ (.B1(_06650_),
    .Y(_02389_),
    .A1(net989),
    .A2(net361));
 sg13g2_nand2_1 _25585_ (.Y(_06651_),
    .A(\cpu.icache.r_tag[6][12] ),
    .B(_06636_));
 sg13g2_o21ai_1 _25586_ (.B1(_06651_),
    .Y(_02390_),
    .A1(net399),
    .A2(_06637_));
 sg13g2_nand2_1 _25587_ (.Y(_06652_),
    .A(\cpu.icache.r_tag[6][13] ),
    .B(_06636_));
 sg13g2_o21ai_1 _25588_ (.B1(_06652_),
    .Y(_02391_),
    .A1(net400),
    .A2(net361));
 sg13g2_nand2_1 _25589_ (.Y(_06653_),
    .A(\cpu.icache.r_tag[6][14] ),
    .B(_06636_));
 sg13g2_o21ai_1 _25590_ (.B1(_06653_),
    .Y(_02392_),
    .A1(net394),
    .A2(net361));
 sg13g2_nand2_1 _25591_ (.Y(_06654_),
    .A(_08523_),
    .B(_06542_));
 sg13g2_buf_1 _25592_ (.A(_06654_),
    .X(_06655_));
 sg13g2_buf_1 _25593_ (.A(_06655_),
    .X(_06656_));
 sg13g2_mux2_1 _25594_ (.A0(_04577_),
    .A1(\cpu.icache.r_tag[7][5] ),
    .S(net452),
    .X(_02393_));
 sg13g2_buf_1 _25595_ (.A(_06655_),
    .X(_06657_));
 sg13g2_nand2_1 _25596_ (.Y(_06658_),
    .A(\cpu.icache.r_tag[7][15] ),
    .B(_06656_));
 sg13g2_o21ai_1 _25597_ (.B1(_06658_),
    .Y(_02394_),
    .A1(net448),
    .A2(_06657_));
 sg13g2_buf_1 _25598_ (.A(_06655_),
    .X(_06659_));
 sg13g2_nand2_1 _25599_ (.Y(_06660_),
    .A(\cpu.icache.r_tag[7][16] ),
    .B(net450));
 sg13g2_o21ai_1 _25600_ (.B1(_06660_),
    .Y(_02395_),
    .A1(net396),
    .A2(net451));
 sg13g2_nand2_1 _25601_ (.Y(_06661_),
    .A(\cpu.icache.r_tag[7][17] ),
    .B(net450));
 sg13g2_o21ai_1 _25602_ (.B1(_06661_),
    .Y(_02396_),
    .A1(_08646_),
    .A2(net451));
 sg13g2_nand2_1 _25603_ (.Y(_06662_),
    .A(\cpu.icache.r_tag[7][18] ),
    .B(_06659_));
 sg13g2_o21ai_1 _25604_ (.B1(_06662_),
    .Y(_02397_),
    .A1(net447),
    .A2(net451));
 sg13g2_nand2_1 _25605_ (.Y(_06663_),
    .A(\cpu.icache.r_tag[7][19] ),
    .B(net450));
 sg13g2_o21ai_1 _25606_ (.B1(_06663_),
    .Y(_02398_),
    .A1(net392),
    .A2(net451));
 sg13g2_nand2_1 _25607_ (.Y(_06664_),
    .A(\cpu.icache.r_tag[7][20] ),
    .B(net450));
 sg13g2_o21ai_1 _25608_ (.B1(_06664_),
    .Y(_02399_),
    .A1(net393),
    .A2(net451));
 sg13g2_nand2_1 _25609_ (.Y(_06665_),
    .A(\cpu.icache.r_tag[7][21] ),
    .B(net450));
 sg13g2_o21ai_1 _25610_ (.B1(_06665_),
    .Y(_02400_),
    .A1(net398),
    .A2(net451));
 sg13g2_nand2_1 _25611_ (.Y(_06666_),
    .A(\cpu.icache.r_tag[7][22] ),
    .B(net450));
 sg13g2_o21ai_1 _25612_ (.B1(_06666_),
    .Y(_02401_),
    .A1(net397),
    .A2(net451));
 sg13g2_nand2_1 _25613_ (.Y(_06667_),
    .A(\cpu.icache.r_tag[7][23] ),
    .B(net450));
 sg13g2_o21ai_1 _25614_ (.B1(_06667_),
    .Y(_02402_),
    .A1(_08777_),
    .A2(net451));
 sg13g2_mux2_1 _25615_ (.A0(_04611_),
    .A1(\cpu.icache.r_tag[7][6] ),
    .S(net452),
    .X(_02403_));
 sg13g2_mux2_1 _25616_ (.A0(_04639_),
    .A1(\cpu.icache.r_tag[7][7] ),
    .S(net452),
    .X(_02404_));
 sg13g2_nand2_1 _25617_ (.Y(_06668_),
    .A(\cpu.icache.r_tag[7][8] ),
    .B(_06659_));
 sg13g2_o21ai_1 _25618_ (.B1(_06668_),
    .Y(_02405_),
    .A1(_04222_),
    .A2(_06657_));
 sg13g2_mux2_1 _25619_ (.A0(_04713_),
    .A1(\cpu.icache.r_tag[7][9] ),
    .S(net452),
    .X(_02406_));
 sg13g2_mux2_1 _25620_ (.A0(_04750_),
    .A1(\cpu.icache.r_tag[7][10] ),
    .S(net452),
    .X(_02407_));
 sg13g2_nand2_1 _25621_ (.Y(_06669_),
    .A(\cpu.icache.r_tag[7][11] ),
    .B(net450));
 sg13g2_o21ai_1 _25622_ (.B1(_06669_),
    .Y(_02408_),
    .A1(_04280_),
    .A2(net452));
 sg13g2_nand2_1 _25623_ (.Y(_06670_),
    .A(\cpu.icache.r_tag[7][12] ),
    .B(_06655_));
 sg13g2_o21ai_1 _25624_ (.B1(_06670_),
    .Y(_02409_),
    .A1(_08511_),
    .A2(net452));
 sg13g2_nand2_1 _25625_ (.Y(_06671_),
    .A(\cpu.icache.r_tag[7][13] ),
    .B(_06655_));
 sg13g2_o21ai_1 _25626_ (.B1(_06671_),
    .Y(_02410_),
    .A1(_08447_),
    .A2(_06656_));
 sg13g2_nand2_1 _25627_ (.Y(_06672_),
    .A(\cpu.icache.r_tag[7][14] ),
    .B(_06655_));
 sg13g2_o21ai_1 _25628_ (.B1(_06672_),
    .Y(_02411_),
    .A1(_08670_),
    .A2(net452));
 sg13g2_buf_1 _25629_ (.A(_09968_),
    .X(_06673_));
 sg13g2_buf_1 _25630_ (.A(net960),
    .X(_06674_));
 sg13g2_and2_1 _25631_ (.A(net234),
    .B(_05146_),
    .X(_06675_));
 sg13g2_buf_2 _25632_ (.A(_06675_),
    .X(_06676_));
 sg13g2_buf_1 _25633_ (.A(_06676_),
    .X(_06677_));
 sg13g2_mux2_1 _25634_ (.A0(\cpu.intr.r_clock_cmp[0] ),
    .A1(_06674_),
    .S(net128),
    .X(_02421_));
 sg13g2_mux2_1 _25635_ (.A0(\cpu.intr.r_clock_cmp[10] ),
    .A1(_10091_),
    .S(net128),
    .X(_02422_));
 sg13g2_mux2_1 _25636_ (.A0(\cpu.intr.r_clock_cmp[11] ),
    .A1(_10098_),
    .S(net128),
    .X(_02423_));
 sg13g2_mux2_1 _25637_ (.A0(\cpu.intr.r_clock_cmp[12] ),
    .A1(_10103_),
    .S(net128),
    .X(_02424_));
 sg13g2_mux2_1 _25638_ (.A0(\cpu.intr.r_clock_cmp[13] ),
    .A1(_10108_),
    .S(net128),
    .X(_02425_));
 sg13g2_mux2_1 _25639_ (.A0(\cpu.intr.r_clock_cmp[14] ),
    .A1(_10114_),
    .S(_06677_),
    .X(_02426_));
 sg13g2_mux2_1 _25640_ (.A0(\cpu.intr.r_clock_cmp[15] ),
    .A1(_10122_),
    .S(_06677_),
    .X(_02427_));
 sg13g2_nor2_1 _25641_ (.A(_09898_),
    .B(_05477_),
    .Y(_06678_));
 sg13g2_buf_2 _25642_ (.A(_06678_),
    .X(_06679_));
 sg13g2_buf_1 _25643_ (.A(_06679_),
    .X(_06680_));
 sg13g2_mux2_1 _25644_ (.A0(\cpu.intr.r_clock_cmp[16] ),
    .A1(_06674_),
    .S(net163),
    .X(_02428_));
 sg13g2_mux2_1 _25645_ (.A0(\cpu.intr.r_clock_cmp[17] ),
    .A1(net1060),
    .S(net163),
    .X(_02429_));
 sg13g2_mux2_1 _25646_ (.A0(\cpu.intr.r_clock_cmp[18] ),
    .A1(net921),
    .S(net163),
    .X(_02430_));
 sg13g2_mux2_1 _25647_ (.A0(\cpu.intr.r_clock_cmp[19] ),
    .A1(net981),
    .S(net163),
    .X(_02431_));
 sg13g2_mux2_1 _25648_ (.A0(\cpu.intr.r_clock_cmp[1] ),
    .A1(net1060),
    .S(net128),
    .X(_02432_));
 sg13g2_mux2_1 _25649_ (.A0(\cpu.intr.r_clock_cmp[20] ),
    .A1(_12259_),
    .S(net163),
    .X(_02433_));
 sg13g2_mux2_1 _25650_ (.A0(\cpu.intr.r_clock_cmp[21] ),
    .A1(_10063_),
    .S(net163),
    .X(_02434_));
 sg13g2_mux2_1 _25651_ (.A0(\cpu.intr.r_clock_cmp[22] ),
    .A1(net1053),
    .S(net163),
    .X(_02435_));
 sg13g2_mux2_1 _25652_ (.A0(\cpu.intr.r_clock_cmp[23] ),
    .A1(_10016_),
    .S(net163),
    .X(_02436_));
 sg13g2_mux2_1 _25653_ (.A0(\cpu.intr.r_clock_cmp[24] ),
    .A1(_10081_),
    .S(_06680_),
    .X(_02437_));
 sg13g2_mux2_1 _25654_ (.A0(\cpu.intr.r_clock_cmp[25] ),
    .A1(_10086_),
    .S(_06680_),
    .X(_02438_));
 sg13g2_mux2_1 _25655_ (.A0(\cpu.intr.r_clock_cmp[26] ),
    .A1(_10091_),
    .S(_06679_),
    .X(_02439_));
 sg13g2_mux2_1 _25656_ (.A0(\cpu.intr.r_clock_cmp[27] ),
    .A1(_10098_),
    .S(_06679_),
    .X(_02440_));
 sg13g2_mux2_1 _25657_ (.A0(\cpu.intr.r_clock_cmp[28] ),
    .A1(_10103_),
    .S(_06679_),
    .X(_02441_));
 sg13g2_mux2_1 _25658_ (.A0(\cpu.intr.r_clock_cmp[29] ),
    .A1(_10108_),
    .S(_06679_),
    .X(_02442_));
 sg13g2_mux2_1 _25659_ (.A0(\cpu.intr.r_clock_cmp[2] ),
    .A1(net921),
    .S(net128),
    .X(_02443_));
 sg13g2_mux2_1 _25660_ (.A0(\cpu.intr.r_clock_cmp[30] ),
    .A1(_10114_),
    .S(_06679_),
    .X(_02444_));
 sg13g2_mux2_1 _25661_ (.A0(\cpu.intr.r_clock_cmp[31] ),
    .A1(_10122_),
    .S(_06679_),
    .X(_02445_));
 sg13g2_mux2_1 _25662_ (.A0(\cpu.intr.r_clock_cmp[3] ),
    .A1(net981),
    .S(net128),
    .X(_02446_));
 sg13g2_mux2_1 _25663_ (.A0(\cpu.intr.r_clock_cmp[4] ),
    .A1(net1022),
    .S(_06676_),
    .X(_02447_));
 sg13g2_mux2_1 _25664_ (.A0(\cpu.intr.r_clock_cmp[5] ),
    .A1(_10063_),
    .S(_06676_),
    .X(_02448_));
 sg13g2_mux2_1 _25665_ (.A0(\cpu.intr.r_clock_cmp[6] ),
    .A1(_10069_),
    .S(_06676_),
    .X(_02449_));
 sg13g2_mux2_1 _25666_ (.A0(\cpu.intr.r_clock_cmp[7] ),
    .A1(_10016_),
    .S(_06676_),
    .X(_02450_));
 sg13g2_mux2_1 _25667_ (.A0(\cpu.intr.r_clock_cmp[8] ),
    .A1(_10081_),
    .S(_06676_),
    .X(_02451_));
 sg13g2_mux2_1 _25668_ (.A0(\cpu.intr.r_clock_cmp[9] ),
    .A1(_10086_),
    .S(_06676_),
    .X(_02452_));
 sg13g2_and2_1 _25669_ (.A(_10021_),
    .B(net341),
    .X(_06681_));
 sg13g2_buf_2 _25670_ (.A(_06681_),
    .X(_06682_));
 sg13g2_buf_1 _25671_ (.A(_06682_),
    .X(_06683_));
 sg13g2_mux2_1 _25672_ (.A0(\cpu.intr.r_timer_reload[0] ),
    .A1(net841),
    .S(net127),
    .X(_02476_));
 sg13g2_mux2_1 _25673_ (.A0(\cpu.intr.r_timer_reload[10] ),
    .A1(_10091_),
    .S(net127),
    .X(_02477_));
 sg13g2_mux2_1 _25674_ (.A0(\cpu.intr.r_timer_reload[11] ),
    .A1(_10098_),
    .S(net127),
    .X(_02478_));
 sg13g2_mux2_1 _25675_ (.A0(\cpu.intr.r_timer_reload[12] ),
    .A1(_10103_),
    .S(net127),
    .X(_02479_));
 sg13g2_mux2_1 _25676_ (.A0(\cpu.intr.r_timer_reload[13] ),
    .A1(_10108_),
    .S(net127),
    .X(_02480_));
 sg13g2_mux2_1 _25677_ (.A0(\cpu.intr.r_timer_reload[14] ),
    .A1(_10114_),
    .S(_06683_),
    .X(_02481_));
 sg13g2_mux2_1 _25678_ (.A0(\cpu.intr.r_timer_reload[15] ),
    .A1(_10122_),
    .S(_06683_),
    .X(_02482_));
 sg13g2_mux2_1 _25679_ (.A0(\cpu.intr.r_timer_reload[16] ),
    .A1(net841),
    .S(net184),
    .X(_02483_));
 sg13g2_mux2_1 _25680_ (.A0(\cpu.intr.r_timer_reload[17] ),
    .A1(net1060),
    .S(net184),
    .X(_02484_));
 sg13g2_mux2_1 _25681_ (.A0(\cpu.intr.r_timer_reload[18] ),
    .A1(net921),
    .S(net184),
    .X(_02485_));
 sg13g2_inv_1 _25682_ (.Y(_06684_),
    .A(\cpu.intr.r_timer_reload[19] ));
 sg13g2_o21ai_1 _25683_ (.B1(_09994_),
    .Y(_02486_),
    .A1(_06684_),
    .A2(net185));
 sg13g2_mux2_1 _25684_ (.A0(\cpu.intr.r_timer_reload[1] ),
    .A1(net1060),
    .S(net127),
    .X(_02487_));
 sg13g2_o21ai_1 _25685_ (.B1(_10001_),
    .Y(_02488_),
    .A1(_09995_),
    .A2(_09972_));
 sg13g2_inv_1 _25686_ (.Y(_06685_),
    .A(\cpu.intr.r_timer_reload[21] ));
 sg13g2_o21ai_1 _25687_ (.B1(_10006_),
    .Y(_02489_),
    .A1(_06685_),
    .A2(net185));
 sg13g2_inv_1 _25688_ (.Y(_06686_),
    .A(\cpu.intr.r_timer_reload[22] ));
 sg13g2_o21ai_1 _25689_ (.B1(_10011_),
    .Y(_02490_),
    .A1(_06686_),
    .A2(net185));
 sg13g2_mux2_1 _25690_ (.A0(\cpu.intr.r_timer_reload[23] ),
    .A1(net1056),
    .S(_09973_),
    .X(_02491_));
 sg13g2_mux2_1 _25691_ (.A0(\cpu.intr.r_timer_reload[2] ),
    .A1(net921),
    .S(net127),
    .X(_02492_));
 sg13g2_mux2_1 _25692_ (.A0(\cpu.intr.r_timer_reload[3] ),
    .A1(net1024),
    .S(net127),
    .X(_02493_));
 sg13g2_mux2_1 _25693_ (.A0(\cpu.intr.r_timer_reload[4] ),
    .A1(_12259_),
    .S(_06682_),
    .X(_02494_));
 sg13g2_mux2_1 _25694_ (.A0(\cpu.intr.r_timer_reload[5] ),
    .A1(net1054),
    .S(_06682_),
    .X(_02495_));
 sg13g2_mux2_1 _25695_ (.A0(\cpu.intr.r_timer_reload[6] ),
    .A1(net1053),
    .S(_06682_),
    .X(_02496_));
 sg13g2_mux2_1 _25696_ (.A0(\cpu.intr.r_timer_reload[7] ),
    .A1(net1056),
    .S(_06682_),
    .X(_02497_));
 sg13g2_mux2_1 _25697_ (.A0(\cpu.intr.r_timer_reload[8] ),
    .A1(_10081_),
    .S(_06682_),
    .X(_02498_));
 sg13g2_mux2_1 _25698_ (.A0(\cpu.intr.r_timer_reload[9] ),
    .A1(_10086_),
    .S(_06682_),
    .X(_02499_));
 sg13g2_inv_1 _25699_ (.Y(_06687_),
    .A(_09763_));
 sg13g2_nor4_2 _25700_ (.A(_12018_),
    .B(_12015_),
    .C(_09782_),
    .Y(_06688_),
    .D(_12016_));
 sg13g2_nor3_1 _25701_ (.A(_12038_),
    .B(_12019_),
    .C(_12039_),
    .Y(_06689_));
 sg13g2_nand2_1 _25702_ (.Y(_06690_),
    .A(_06688_),
    .B(_06689_));
 sg13g2_nor3_1 _25703_ (.A(_09770_),
    .B(_09761_),
    .C(_06690_),
    .Y(_06691_));
 sg13g2_nand3_1 _25704_ (.B(_12021_),
    .C(_06691_),
    .A(_09760_),
    .Y(_06692_));
 sg13g2_buf_1 _25705_ (.A(_06692_),
    .X(_06693_));
 sg13g2_inv_1 _25706_ (.Y(_06694_),
    .A(_09832_));
 sg13g2_and2_1 _25707_ (.A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_09795_),
    .X(_06695_));
 sg13g2_a221oi_1 _25708_ (.B2(\cpu.qspi.r_read_delay[0][0] ),
    .C1(_06695_),
    .B1(_09800_),
    .A1(\cpu.qspi.r_read_delay[2][0] ),
    .Y(_06696_),
    .A2(_09798_));
 sg13g2_or4_1 _25709_ (.A(_09769_),
    .B(_09781_),
    .C(net1148),
    .D(net1149),
    .X(_06697_));
 sg13g2_buf_1 _25710_ (.A(_06697_),
    .X(_06698_));
 sg13g2_a221oi_1 _25711_ (.B2(_06698_),
    .C1(_09779_),
    .B1(_00181_),
    .A1(net1147),
    .Y(_06699_),
    .A2(_06687_));
 sg13g2_o21ai_1 _25712_ (.B1(_06699_),
    .Y(_06700_),
    .A1(_06694_),
    .A2(_06696_));
 sg13g2_nor2_1 _25713_ (.A(net28),
    .B(_06700_),
    .Y(_06701_));
 sg13g2_a21oi_1 _25714_ (.A1(_06687_),
    .A2(net28),
    .Y(_02500_),
    .B1(_06701_));
 sg13g2_nor3_1 _25715_ (.A(_09832_),
    .B(net1147),
    .C(_06698_),
    .Y(_06702_));
 sg13g2_nor2_1 _25716_ (.A(net1147),
    .B(_06698_),
    .Y(_06703_));
 sg13g2_xor2_1 _25717_ (.B(_09764_),
    .A(_09763_),
    .X(_06704_));
 sg13g2_nor2_1 _25718_ (.A(_06703_),
    .B(_06704_),
    .Y(_06705_));
 sg13g2_a22oi_1 _25719_ (.Y(_06706_),
    .B1(_09795_),
    .B2(\cpu.qspi.r_read_delay[1][1] ),
    .A2(_09798_),
    .A1(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_nand2_1 _25720_ (.Y(_06707_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_09800_));
 sg13g2_a21oi_1 _25721_ (.A1(_06706_),
    .A2(_06707_),
    .Y(_06708_),
    .B1(_06694_));
 sg13g2_nor4_1 _25722_ (.A(_09779_),
    .B(_06702_),
    .C(_06705_),
    .D(_06708_),
    .Y(_06709_));
 sg13g2_nand2_1 _25723_ (.Y(_06710_),
    .A(_09764_),
    .B(net28));
 sg13g2_o21ai_1 _25724_ (.B1(_06710_),
    .Y(_02501_),
    .A1(net28),
    .A2(_06709_));
 sg13g2_a22oi_1 _25725_ (.Y(_06711_),
    .B1(_09795_),
    .B2(\cpu.qspi.r_read_delay[1][2] ),
    .A2(_09798_),
    .A1(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_nand2_1 _25726_ (.Y(_06712_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_09800_));
 sg13g2_a21oi_1 _25727_ (.A1(_06711_),
    .A2(_06712_),
    .Y(_06713_),
    .B1(_06694_));
 sg13g2_nor2_1 _25728_ (.A(_09763_),
    .B(_09764_),
    .Y(_06714_));
 sg13g2_xor2_1 _25729_ (.B(_06714_),
    .A(_00182_),
    .X(_06715_));
 sg13g2_mux2_1 _25730_ (.A0(_06698_),
    .A1(net799),
    .S(net1147),
    .X(_06716_));
 sg13g2_a22oi_1 _25731_ (.Y(_06717_),
    .B1(_06715_),
    .B2(_06716_),
    .A2(_06703_),
    .A1(_09832_));
 sg13g2_nor3_1 _25732_ (.A(_09779_),
    .B(_06713_),
    .C(_06717_),
    .Y(_06718_));
 sg13g2_nand2_1 _25733_ (.Y(_06719_),
    .A(_09765_),
    .B(_06693_));
 sg13g2_o21ai_1 _25734_ (.B1(_06719_),
    .Y(_02502_),
    .A1(net28),
    .A2(_06718_));
 sg13g2_a21oi_1 _25735_ (.A1(net1147),
    .A2(_09776_),
    .Y(_06720_),
    .B1(_06698_));
 sg13g2_inv_1 _25736_ (.Y(_06721_),
    .A(_06720_));
 sg13g2_a22oi_1 _25737_ (.Y(_06722_),
    .B1(_09795_),
    .B2(\cpu.qspi.r_read_delay[1][3] ),
    .A2(_09798_),
    .A1(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_nand2_1 _25738_ (.Y(_06723_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_09800_));
 sg13g2_nand2_1 _25739_ (.Y(_06724_),
    .A(_06722_),
    .B(_06723_));
 sg13g2_a22oi_1 _25740_ (.Y(_06725_),
    .B1(_06724_),
    .B2(_09832_),
    .A2(_06721_),
    .A1(_09766_));
 sg13g2_inv_1 _25741_ (.Y(_06726_),
    .A(_09765_));
 sg13g2_a21oi_1 _25742_ (.A1(_06726_),
    .A2(_06714_),
    .Y(_06727_),
    .B1(_06720_));
 sg13g2_o21ai_1 _25743_ (.B1(\cpu.qspi.r_count[3] ),
    .Y(_06728_),
    .A1(net28),
    .A2(_06727_));
 sg13g2_o21ai_1 _25744_ (.B1(_06728_),
    .Y(_02503_),
    .A1(net28),
    .A2(_06725_));
 sg13g2_or2_1 _25745_ (.X(_06729_),
    .B(_09766_),
    .A(_00244_));
 sg13g2_a21oi_1 _25746_ (.A1(_09776_),
    .A2(_06729_),
    .Y(_06730_),
    .B1(_06720_));
 sg13g2_mux2_1 _25747_ (.A0(_06730_),
    .A1(\cpu.qspi.r_count[4] ),
    .S(net28),
    .X(_02504_));
 sg13g2_and2_1 _25748_ (.A(_09895_),
    .B(_06305_),
    .X(_06731_));
 sg13g2_buf_2 _25749_ (.A(_06731_),
    .X(_06732_));
 sg13g2_and2_1 _25750_ (.A(_09181_),
    .B(_06732_),
    .X(_06733_));
 sg13g2_buf_1 _25751_ (.A(_06733_),
    .X(_06734_));
 sg13g2_nand2_1 _25752_ (.Y(_06735_),
    .A(net841),
    .B(_06734_));
 sg13g2_nand2_1 _25753_ (.Y(_06736_),
    .A(_09181_),
    .B(_06732_));
 sg13g2_buf_1 _25754_ (.A(_06736_),
    .X(_06737_));
 sg13g2_nand2_1 _25755_ (.Y(_06738_),
    .A(\cpu.qspi.r_read_delay[0][0] ),
    .B(_06737_));
 sg13g2_a21oi_1 _25756_ (.A1(_06735_),
    .A2(_06738_),
    .Y(_02515_),
    .B1(net637));
 sg13g2_nand2_1 _25757_ (.Y(_06739_),
    .A(_09979_),
    .B(_06734_));
 sg13g2_nand2_1 _25758_ (.Y(_06740_),
    .A(\cpu.qspi.r_read_delay[0][1] ),
    .B(_06737_));
 sg13g2_a21oi_1 _25759_ (.A1(_06739_),
    .A2(_06740_),
    .Y(_02516_),
    .B1(net637));
 sg13g2_nand2_1 _25760_ (.Y(_06741_),
    .A(_09986_),
    .B(_06734_));
 sg13g2_nand2_1 _25761_ (.Y(_06742_),
    .A(\cpu.qspi.r_read_delay[0][2] ),
    .B(_06737_));
 sg13g2_nand3_1 _25762_ (.B(_06741_),
    .C(_06742_),
    .A(net663),
    .Y(_02517_));
 sg13g2_nand2_1 _25763_ (.Y(_06743_),
    .A(net1058),
    .B(_06734_));
 sg13g2_nand2_1 _25764_ (.Y(_06744_),
    .A(\cpu.qspi.r_read_delay[0][3] ),
    .B(_06737_));
 sg13g2_buf_1 _25765_ (.A(_09772_),
    .X(_06745_));
 sg13g2_a21oi_1 _25766_ (.A1(_06743_),
    .A2(_06744_),
    .Y(_02518_),
    .B1(net593));
 sg13g2_and2_1 _25767_ (.A(_04915_),
    .B(_06732_),
    .X(_06746_));
 sg13g2_buf_1 _25768_ (.A(_06746_),
    .X(_06747_));
 sg13g2_nand2_1 _25769_ (.Y(_06748_),
    .A(net841),
    .B(_06747_));
 sg13g2_nand2_1 _25770_ (.Y(_06749_),
    .A(_04915_),
    .B(_06732_));
 sg13g2_buf_1 _25771_ (.A(_06749_),
    .X(_06750_));
 sg13g2_nand2_1 _25772_ (.Y(_06751_),
    .A(\cpu.qspi.r_read_delay[1][0] ),
    .B(_06750_));
 sg13g2_a21oi_1 _25773_ (.A1(_06748_),
    .A2(_06751_),
    .Y(_02519_),
    .B1(net593));
 sg13g2_nand2_1 _25774_ (.Y(_06752_),
    .A(_09979_),
    .B(_06747_));
 sg13g2_nand2_1 _25775_ (.Y(_06753_),
    .A(\cpu.qspi.r_read_delay[1][1] ),
    .B(_06750_));
 sg13g2_a21oi_1 _25776_ (.A1(_06752_),
    .A2(_06753_),
    .Y(_02520_),
    .B1(net593));
 sg13g2_nand2_1 _25777_ (.Y(_06754_),
    .A(_09986_),
    .B(_06747_));
 sg13g2_nand2_1 _25778_ (.Y(_06755_),
    .A(\cpu.qspi.r_read_delay[1][2] ),
    .B(_06750_));
 sg13g2_nand3_1 _25779_ (.B(_06754_),
    .C(_06755_),
    .A(net663),
    .Y(_02521_));
 sg13g2_nand2_1 _25780_ (.Y(_06756_),
    .A(net1058),
    .B(_06747_));
 sg13g2_nand2_1 _25781_ (.Y(_06757_),
    .A(\cpu.qspi.r_read_delay[1][3] ),
    .B(_06750_));
 sg13g2_a21oi_1 _25782_ (.A1(_06756_),
    .A2(_06757_),
    .Y(_02522_),
    .B1(net593));
 sg13g2_nor2b_1 _25783_ (.A(_04861_),
    .B_N(_06732_),
    .Y(_06758_));
 sg13g2_buf_1 _25784_ (.A(_06758_),
    .X(_06759_));
 sg13g2_nand2_1 _25785_ (.Y(_06760_),
    .A(_06673_),
    .B(_06759_));
 sg13g2_nand2b_1 _25786_ (.Y(_06761_),
    .B(_06732_),
    .A_N(_04861_));
 sg13g2_buf_1 _25787_ (.A(_06761_),
    .X(_06762_));
 sg13g2_nand2_1 _25788_ (.Y(_06763_),
    .A(\cpu.qspi.r_read_delay[2][0] ),
    .B(_06762_));
 sg13g2_a21oi_1 _25789_ (.A1(_06760_),
    .A2(_06763_),
    .Y(_02523_),
    .B1(net593));
 sg13g2_nand2_1 _25790_ (.Y(_06764_),
    .A(net1055),
    .B(_06759_));
 sg13g2_nand2_1 _25791_ (.Y(_06765_),
    .A(\cpu.qspi.r_read_delay[2][1] ),
    .B(_06762_));
 sg13g2_a21oi_1 _25792_ (.A1(_06764_),
    .A2(_06765_),
    .Y(_02524_),
    .B1(net593));
 sg13g2_nand2_1 _25793_ (.Y(_06766_),
    .A(_09985_),
    .B(_06759_));
 sg13g2_nand2_1 _25794_ (.Y(_06767_),
    .A(\cpu.qspi.r_read_delay[2][2] ),
    .B(_06762_));
 sg13g2_nand3_1 _25795_ (.B(_06766_),
    .C(_06767_),
    .A(net663),
    .Y(_02525_));
 sg13g2_nand2_1 _25796_ (.Y(_06768_),
    .A(_09993_),
    .B(_06759_));
 sg13g2_nand2_1 _25797_ (.Y(_06769_),
    .A(\cpu.qspi.r_read_delay[2][3] ),
    .B(_06762_));
 sg13g2_a21oi_1 _25798_ (.A1(_06768_),
    .A2(_06769_),
    .Y(_02526_),
    .B1(net593));
 sg13g2_inv_1 _25799_ (.Y(_06770_),
    .A(_06689_));
 sg13g2_nor4_1 _25800_ (.A(_09781_),
    .B(_09779_),
    .C(net1149),
    .D(_06770_),
    .Y(_06771_));
 sg13g2_nor2b_1 _25801_ (.A(\cpu.qspi.r_state[12] ),
    .B_N(_06688_),
    .Y(_06772_));
 sg13g2_and3_1 _25802_ (.X(_06773_),
    .A(_09784_),
    .B(_06771_),
    .C(_06772_));
 sg13g2_buf_1 _25803_ (.A(_06773_),
    .X(_06774_));
 sg13g2_xnor2_1 _25804_ (.Y(_06775_),
    .A(_09778_),
    .B(_09803_));
 sg13g2_buf_1 _25805_ (.A(_08273_),
    .X(_06776_));
 sg13g2_buf_1 _25806_ (.A(_09744_),
    .X(_06777_));
 sg13g2_mux2_1 _25807_ (.A0(_09451_),
    .A1(_09441_),
    .S(net126),
    .X(_06778_));
 sg13g2_nor2_1 _25808_ (.A(net959),
    .B(_06778_),
    .Y(_06779_));
 sg13g2_a21oi_1 _25809_ (.A1(net959),
    .A2(_08511_),
    .Y(_06780_),
    .B1(_06779_));
 sg13g2_o21ai_1 _25810_ (.B1(_09782_),
    .Y(_06781_),
    .A1(net1164),
    .A2(_09740_));
 sg13g2_nand2b_1 _25811_ (.Y(_06782_),
    .B(_06781_),
    .A_N(_12018_));
 sg13g2_inv_1 _25812_ (.Y(_06783_),
    .A(_09762_));
 sg13g2_buf_1 _25813_ (.A(\cpu.qspi.r_state[0] ),
    .X(_06784_));
 sg13g2_nand2_1 _25814_ (.Y(_06785_),
    .A(net1159),
    .B(net1164));
 sg13g2_o21ai_1 _25815_ (.B1(_06785_),
    .Y(_06786_),
    .A1(net1164),
    .A2(_12076_));
 sg13g2_a221oi_1 _25816_ (.B2(_12039_),
    .C1(_06774_),
    .B1(_06786_),
    .A1(_06783_),
    .Y(_06787_),
    .A2(_06784_));
 sg13g2_nand2b_1 _25817_ (.Y(_06788_),
    .B(net1114),
    .A_N(_12127_));
 sg13g2_nand2_1 _25818_ (.Y(_06789_),
    .A(_12149_),
    .B(_05012_));
 sg13g2_nand2b_1 _25819_ (.Y(_06790_),
    .B(net1114),
    .A_N(_04983_));
 sg13g2_nand3_1 _25820_ (.B(_06789_),
    .C(_06790_),
    .A(net1025),
    .Y(_06791_));
 sg13g2_o21ai_1 _25821_ (.B1(_06791_),
    .Y(_06792_),
    .A1(_05522_),
    .A2(_06788_));
 sg13g2_nand2_1 _25822_ (.Y(_06793_),
    .A(_12127_),
    .B(_04994_));
 sg13g2_o21ai_1 _25823_ (.B1(_06793_),
    .Y(_06794_),
    .A1(_12127_),
    .A2(_05197_));
 sg13g2_mux2_1 _25824_ (.A0(_05204_),
    .A1(_05002_),
    .S(_12127_),
    .X(_06795_));
 sg13g2_a22oi_1 _25825_ (.Y(_06796_),
    .B1(_06795_),
    .B2(net1028),
    .A2(_06794_),
    .A1(net1114));
 sg13g2_mux2_1 _25826_ (.A0(_06792_),
    .A1(_06796_),
    .S(net1112),
    .X(_06797_));
 sg13g2_o21ai_1 _25827_ (.B1(_06797_),
    .Y(_06798_),
    .A1(net1021),
    .A2(net1028));
 sg13g2_inv_1 _25828_ (.Y(_06799_),
    .A(_12149_));
 sg13g2_nor2_1 _25829_ (.A(_06799_),
    .B(_12252_),
    .Y(_06800_));
 sg13g2_nor2_2 _25830_ (.A(net1114),
    .B(_06800_),
    .Y(_06801_));
 sg13g2_nand2b_1 _25831_ (.Y(_06802_),
    .B(_06801_),
    .A_N(_05515_));
 sg13g2_nand3_1 _25832_ (.B(_06798_),
    .C(_06802_),
    .A(net1149),
    .Y(_06803_));
 sg13g2_nand3b_1 _25833_ (.B(_06787_),
    .C(_06803_),
    .Y(_06804_),
    .A_N(_06782_));
 sg13g2_a21oi_1 _25834_ (.A1(_12019_),
    .A2(_06780_),
    .Y(_06805_),
    .B1(_06804_));
 sg13g2_mux2_1 _25835_ (.A0(_09394_),
    .A1(net390),
    .S(_09744_),
    .X(_06806_));
 sg13g2_nand2_1 _25836_ (.Y(_06807_),
    .A(net950),
    .B(_06806_));
 sg13g2_o21ai_1 _25837_ (.B1(_06807_),
    .Y(_06808_),
    .A1(net950),
    .A2(_08619_));
 sg13g2_buf_1 _25838_ (.A(_09744_),
    .X(_06809_));
 sg13g2_nor2_1 _25839_ (.A(_09583_),
    .B(net126),
    .Y(_06810_));
 sg13g2_a21oi_1 _25840_ (.A1(_00227_),
    .A2(net125),
    .Y(_06811_),
    .B1(_06810_));
 sg13g2_mux2_1 _25841_ (.A0(_04673_),
    .A1(_06811_),
    .S(net950),
    .X(_06812_));
 sg13g2_a22oi_1 _25842_ (.Y(_06813_),
    .B1(_06812_),
    .B2(_12015_),
    .A2(_06808_),
    .A1(_12038_));
 sg13g2_nand2_1 _25843_ (.Y(_06814_),
    .A(_06687_),
    .B(_09764_));
 sg13g2_mux2_1 _25844_ (.A0(_06814_),
    .A1(_09764_),
    .S(_09778_),
    .X(_06815_));
 sg13g2_nand2_1 _25845_ (.Y(_06816_),
    .A(net1148),
    .B(_09762_));
 sg13g2_a21o_1 _25846_ (.A2(_06816_),
    .A1(_00181_),
    .B1(_09764_),
    .X(_06817_));
 sg13g2_o21ai_1 _25847_ (.B1(_06817_),
    .Y(_06818_),
    .A1(net1148),
    .A2(_06815_));
 sg13g2_nand3_1 _25848_ (.B(_09763_),
    .C(_09762_),
    .A(net1148),
    .Y(_06819_));
 sg13g2_o21ai_1 _25849_ (.B1(_06819_),
    .Y(_06820_),
    .A1(_09762_),
    .A2(_06814_));
 sg13g2_nand2b_1 _25850_ (.Y(_06821_),
    .B(_09778_),
    .A_N(_09764_));
 sg13g2_a21oi_1 _25851_ (.A1(_06814_),
    .A2(_06821_),
    .Y(_06822_),
    .B1(net1148));
 sg13g2_nor3_1 _25852_ (.A(_09765_),
    .B(_06820_),
    .C(_06822_),
    .Y(_06823_));
 sg13g2_a21o_1 _25853_ (.A2(_06818_),
    .A1(_09765_),
    .B1(_06823_),
    .X(_06824_));
 sg13g2_o21ai_1 _25854_ (.B1(_06824_),
    .Y(_06825_),
    .A1(_09781_),
    .A2(net1148));
 sg13g2_and3_1 _25855_ (.X(_06826_),
    .A(_06805_),
    .B(_06813_),
    .C(_06825_));
 sg13g2_a21oi_1 _25856_ (.A1(_06774_),
    .A2(_06775_),
    .Y(_06827_),
    .B1(_06826_));
 sg13g2_and2_1 _25857_ (.A(\cpu.qspi.r_mask[1] ),
    .B(_09795_),
    .X(_06828_));
 sg13g2_a221oi_1 _25858_ (.B2(\cpu.qspi.r_mask[0] ),
    .C1(_06828_),
    .B1(_09800_),
    .A1(\cpu.qspi.r_mask[2] ),
    .Y(_06829_),
    .A2(_09798_));
 sg13g2_nand2_1 _25859_ (.Y(_06830_),
    .A(_12018_),
    .B(_06829_));
 sg13g2_nor3_2 _25860_ (.A(_09769_),
    .B(_09770_),
    .C(_09761_),
    .Y(_06831_));
 sg13g2_nor2_1 _25861_ (.A(_09832_),
    .B(\cpu.qspi.r_state[14] ),
    .Y(_06832_));
 sg13g2_nand4_1 _25862_ (.B(_06830_),
    .C(_06831_),
    .A(_09760_),
    .Y(_06833_),
    .D(_06832_));
 sg13g2_buf_1 _25863_ (.A(_06833_),
    .X(_06834_));
 sg13g2_mux2_1 _25864_ (.A0(_06827_),
    .A1(net11),
    .S(_06834_),
    .X(_02531_));
 sg13g2_buf_1 _25865_ (.A(net959),
    .X(_06835_));
 sg13g2_mux2_1 _25866_ (.A0(_09595_),
    .A1(_00229_),
    .S(net125),
    .X(_06836_));
 sg13g2_nand2_1 _25867_ (.Y(_06837_),
    .A(net840),
    .B(_10277_));
 sg13g2_o21ai_1 _25868_ (.B1(_06837_),
    .Y(_06838_),
    .A1(net840),
    .A2(_06836_));
 sg13g2_nand2_1 _25869_ (.Y(_06839_),
    .A(_12015_),
    .B(_06838_));
 sg13g2_mux2_1 _25870_ (.A0(_09464_),
    .A1(_09479_),
    .S(net126),
    .X(_06840_));
 sg13g2_nor2_1 _25871_ (.A(net959),
    .B(_06840_),
    .Y(_06841_));
 sg13g2_a21oi_1 _25872_ (.A1(net840),
    .A2(_08447_),
    .Y(_06842_),
    .B1(_06841_));
 sg13g2_a22oi_1 _25873_ (.Y(_06843_),
    .B1(_05238_),
    .B2(_12150_),
    .A2(_05230_),
    .A1(net1021));
 sg13g2_nand3_1 _25874_ (.B(net1028),
    .C(_05321_),
    .A(net1025),
    .Y(_06844_));
 sg13g2_o21ai_1 _25875_ (.B1(_06844_),
    .Y(_06845_),
    .A1(_12195_),
    .A2(_06843_));
 sg13g2_nor2b_1 _25876_ (.A(_06845_),
    .B_N(net1112),
    .Y(_06846_));
 sg13g2_a22oi_1 _25877_ (.Y(_06847_),
    .B1(_05314_),
    .B2(net1021),
    .A2(_05304_),
    .A1(net1028));
 sg13g2_nand2_1 _25878_ (.Y(_06848_),
    .A(net1025),
    .B(_06847_));
 sg13g2_a21oi_1 _25879_ (.A1(_06788_),
    .A2(_06848_),
    .Y(_06849_),
    .B1(net1112));
 sg13g2_a22oi_1 _25880_ (.Y(_06850_),
    .B1(_05601_),
    .B2(_12252_),
    .A2(_05327_),
    .A1(_12129_));
 sg13g2_nand2_1 _25881_ (.Y(_06851_),
    .A(net1021),
    .B(_06850_));
 sg13g2_o21ai_1 _25882_ (.B1(_06851_),
    .Y(_06852_),
    .A1(net1021),
    .A2(_06799_));
 sg13g2_o21ai_1 _25883_ (.B1(_06852_),
    .Y(_06853_),
    .A1(_06846_),
    .A2(_06849_));
 sg13g2_a21oi_1 _25884_ (.A1(_05591_),
    .A2(_06801_),
    .Y(_06854_),
    .B1(_12020_));
 sg13g2_a221oi_1 _25885_ (.B2(_06854_),
    .C1(_06782_),
    .B1(_06853_),
    .A1(_12019_),
    .Y(_06855_),
    .A2(_06842_));
 sg13g2_buf_1 _25886_ (.A(net950),
    .X(_06856_));
 sg13g2_mux2_1 _25887_ (.A0(_09372_),
    .A1(net391),
    .S(net125),
    .X(_06857_));
 sg13g2_nand2_1 _25888_ (.Y(_06858_),
    .A(net737),
    .B(_06857_));
 sg13g2_o21ai_1 _25889_ (.B1(_06858_),
    .Y(_06859_),
    .A1(net737),
    .A2(_08646_));
 sg13g2_nor2_1 _25890_ (.A(_09573_),
    .B(net125),
    .Y(_06860_));
 sg13g2_a21oi_1 _25891_ (.A1(_09564_),
    .A2(net125),
    .Y(_06861_),
    .B1(_06860_));
 sg13g2_nand2b_1 _25892_ (.Y(_06862_),
    .B(_06835_),
    .A_N(_10507_));
 sg13g2_o21ai_1 _25893_ (.B1(_06862_),
    .Y(_06863_),
    .A1(net840),
    .A2(_06861_));
 sg13g2_a22oi_1 _25894_ (.Y(_06864_),
    .B1(_06863_),
    .B2(_12039_),
    .A2(_06859_),
    .A1(_12038_));
 sg13g2_nand2b_1 _25895_ (.Y(_06865_),
    .B(_06774_),
    .A_N(_09803_));
 sg13g2_nand4_1 _25896_ (.B(_06855_),
    .C(_06864_),
    .A(_06839_),
    .Y(_06866_),
    .D(_06865_));
 sg13g2_mux2_1 _25897_ (.A0(_06866_),
    .A1(net12),
    .S(_06834_),
    .X(_02532_));
 sg13g2_inv_1 _25898_ (.Y(_06867_),
    .A(_00223_));
 sg13g2_mux2_1 _25899_ (.A0(_09497_),
    .A1(_06867_),
    .S(_06809_),
    .X(_06868_));
 sg13g2_mux2_1 _25900_ (.A0(_10434_),
    .A1(_06868_),
    .S(net737),
    .X(_06869_));
 sg13g2_mux2_1 _25901_ (.A0(_05261_),
    .A1(_05124_),
    .S(_12195_),
    .X(_06870_));
 sg13g2_a22oi_1 _25902_ (.Y(_06871_),
    .B1(_06870_),
    .B2(_12151_),
    .A2(_05398_),
    .A1(_12153_));
 sg13g2_nor2b_1 _25903_ (.A(_06871_),
    .B_N(net1021),
    .Y(_06872_));
 sg13g2_a22oi_1 _25904_ (.Y(_06873_),
    .B1(_05269_),
    .B2(_12196_),
    .A2(_05134_),
    .A1(_12129_));
 sg13g2_nor2_1 _25905_ (.A(_06799_),
    .B(_06873_),
    .Y(_06874_));
 sg13g2_nand2b_1 _25906_ (.Y(_06875_),
    .B(_05695_),
    .A_N(net1025));
 sg13g2_nand3b_1 _25907_ (.B(net1028),
    .C(net1025),
    .Y(_06876_),
    .A_N(_05391_));
 sg13g2_a21oi_1 _25908_ (.A1(_06875_),
    .A2(_06876_),
    .Y(_06877_),
    .B1(net1112));
 sg13g2_nor3_1 _25909_ (.A(_06872_),
    .B(_06874_),
    .C(_06877_),
    .Y(_06878_));
 sg13g2_nand2_1 _25910_ (.Y(_06879_),
    .A(_05704_),
    .B(_06801_));
 sg13g2_o21ai_1 _25911_ (.B1(_06879_),
    .Y(_06880_),
    .A1(_06801_),
    .A2(_06878_));
 sg13g2_nor2_1 _25912_ (.A(_09522_),
    .B(net126),
    .Y(_06881_));
 sg13g2_a21oi_1 _25913_ (.A1(_09539_),
    .A2(net125),
    .Y(_06882_),
    .B1(_06881_));
 sg13g2_nand2b_1 _25914_ (.Y(_06883_),
    .B(net959),
    .A_N(_08670_));
 sg13g2_o21ai_1 _25915_ (.B1(_06883_),
    .Y(_06884_),
    .A1(net959),
    .A2(_06882_));
 sg13g2_mux2_1 _25916_ (.A0(_08866_),
    .A1(_12122_),
    .S(net950),
    .X(_06885_));
 sg13g2_nor2_1 _25917_ (.A(_12018_),
    .B(_06774_),
    .Y(_06886_));
 sg13g2_o21ai_1 _25918_ (.B1(_06886_),
    .Y(_06887_),
    .A1(_00183_),
    .A2(_06885_));
 sg13g2_a221oi_1 _25919_ (.B2(_12019_),
    .C1(_06887_),
    .B1(_06884_),
    .A1(_09774_),
    .Y(_06888_),
    .A2(_06880_));
 sg13g2_mux2_1 _25920_ (.A0(_09664_),
    .A1(net445),
    .S(_06777_),
    .X(_06889_));
 sg13g2_nand2_1 _25921_ (.Y(_06890_),
    .A(net950),
    .B(_06889_));
 sg13g2_o21ai_1 _25922_ (.B1(_06890_),
    .Y(_06891_),
    .A1(net737),
    .A2(_08757_));
 sg13g2_inv_1 _25923_ (.Y(_06892_),
    .A(_00231_));
 sg13g2_mux2_1 _25924_ (.A0(_09489_),
    .A1(_06892_),
    .S(net126),
    .X(_06893_));
 sg13g2_nor2_1 _25925_ (.A(net950),
    .B(_10136_),
    .Y(_06894_));
 sg13g2_a21o_1 _25926_ (.A2(_06893_),
    .A1(net737),
    .B1(_06894_),
    .X(_06895_));
 sg13g2_a22oi_1 _25927_ (.Y(_06896_),
    .B1(_06895_),
    .B2(_12015_),
    .A2(_06891_),
    .A1(_12038_));
 sg13g2_nand2_1 _25928_ (.Y(_06897_),
    .A(_06888_),
    .B(_06896_));
 sg13g2_a21oi_1 _25929_ (.A1(_12039_),
    .A2(_06869_),
    .Y(_06898_),
    .B1(_06897_));
 sg13g2_o21ai_1 _25930_ (.B1(_06774_),
    .Y(_06899_),
    .A1(_09778_),
    .A2(_09803_));
 sg13g2_nand2b_1 _25931_ (.Y(_06900_),
    .B(_06899_),
    .A_N(_06834_));
 sg13g2_nand2_1 _25932_ (.Y(_06901_),
    .A(net13),
    .B(_06834_));
 sg13g2_o21ai_1 _25933_ (.B1(_06901_),
    .Y(_02533_),
    .A1(_06898_),
    .A2(_06900_));
 sg13g2_mux2_1 _25934_ (.A0(_09561_),
    .A1(_09541_),
    .S(net126),
    .X(_06902_));
 sg13g2_nor2_1 _25935_ (.A(net959),
    .B(_06902_),
    .Y(_06903_));
 sg13g2_a21oi_1 _25936_ (.A1(net840),
    .A2(_10411_),
    .Y(_06904_),
    .B1(_06903_));
 sg13g2_mux2_1 _25937_ (.A0(_09713_),
    .A1(net442),
    .S(_06777_),
    .X(_06905_));
 sg13g2_nor2_1 _25938_ (.A(_06776_),
    .B(_06905_),
    .Y(_06906_));
 sg13g2_a21oi_1 _25939_ (.A1(_06835_),
    .A2(_08733_),
    .Y(_06907_),
    .B1(_06906_));
 sg13g2_a22oi_1 _25940_ (.Y(_06908_),
    .B1(_06907_),
    .B2(_12019_),
    .A2(_06904_),
    .A1(_12039_));
 sg13g2_mux2_1 _25941_ (.A0(_09419_),
    .A1(_09412_),
    .S(net126),
    .X(_06909_));
 sg13g2_nand2_1 _25942_ (.Y(_06910_),
    .A(net737),
    .B(_06909_));
 sg13g2_o21ai_1 _25943_ (.B1(_06910_),
    .Y(_06911_),
    .A1(net737),
    .A2(_08712_));
 sg13g2_nor2_1 _25944_ (.A(_09620_),
    .B(net126),
    .Y(_06912_));
 sg13g2_a21oi_1 _25945_ (.A1(_09789_),
    .A2(net125),
    .Y(_06913_),
    .B1(_06912_));
 sg13g2_nand2_1 _25946_ (.Y(_06914_),
    .A(net737),
    .B(_06913_));
 sg13g2_nand3b_1 _25947_ (.B(_12016_),
    .C(_09788_),
    .Y(_06915_),
    .A_N(_09787_));
 sg13g2_a21oi_1 _25948_ (.A1(_09790_),
    .A2(_06914_),
    .Y(_06916_),
    .B1(_06915_));
 sg13g2_a21oi_1 _25949_ (.A1(_12038_),
    .A2(_06911_),
    .Y(_06917_),
    .B1(_06916_));
 sg13g2_mux2_1 _25950_ (.A0(_05051_),
    .A1(_05174_),
    .S(net1025),
    .X(_06918_));
 sg13g2_a22oi_1 _25951_ (.Y(_06919_),
    .B1(_06918_),
    .B2(net1112),
    .A2(_05459_),
    .A1(_12153_));
 sg13g2_mux4_1 _25952_ (.S0(net1112),
    .A0(_05041_),
    .A1(_05057_),
    .A2(_05466_),
    .A3(_05182_),
    .S1(net1025),
    .X(_06920_));
 sg13g2_a22oi_1 _25953_ (.Y(_06921_),
    .B1(_06920_),
    .B2(net1021),
    .A2(_06801_),
    .A1(_05034_));
 sg13g2_o21ai_1 _25954_ (.B1(_06921_),
    .Y(_06922_),
    .A1(_06799_),
    .A2(_06919_));
 sg13g2_inv_1 _25955_ (.Y(_06923_),
    .A(_00183_));
 sg13g2_mux2_1 _25956_ (.A0(_03622_),
    .A1(net649),
    .S(net959),
    .X(_06924_));
 sg13g2_a21oi_1 _25957_ (.A1(_06923_),
    .A2(_06924_),
    .Y(_06925_),
    .B1(_09782_));
 sg13g2_nand2_1 _25958_ (.Y(_06926_),
    .A(_06886_),
    .B(_06925_));
 sg13g2_a21oi_1 _25959_ (.A1(net1149),
    .A2(_06922_),
    .Y(_06927_),
    .B1(_06926_));
 sg13g2_nor2b_1 _25960_ (.A(_00233_),
    .B_N(net125),
    .Y(_06928_));
 sg13g2_nor2_1 _25961_ (.A(_09508_),
    .B(_06809_),
    .Y(_06929_));
 sg13g2_nor3_1 _25962_ (.A(_06776_),
    .B(_06928_),
    .C(_06929_),
    .Y(_06930_));
 sg13g2_a21oi_1 _25963_ (.A1(net840),
    .A2(_10319_),
    .Y(_06931_),
    .B1(_06930_));
 sg13g2_nand2_1 _25964_ (.Y(_06932_),
    .A(_12015_),
    .B(_06931_));
 sg13g2_and4_1 _25965_ (.A(_06908_),
    .B(_06917_),
    .C(_06927_),
    .D(_06932_),
    .X(_06933_));
 sg13g2_nand2_1 _25966_ (.Y(_06934_),
    .A(net14),
    .B(_06834_));
 sg13g2_o21ai_1 _25967_ (.B1(_06934_),
    .Y(_02534_),
    .A1(_06900_),
    .A2(_06933_));
 sg13g2_buf_1 _25968_ (.A(_12086_),
    .X(_06935_));
 sg13g2_nor2b_1 _25969_ (.A(_09171_),
    .B_N(_09197_),
    .Y(_06936_));
 sg13g2_nand2_1 _25970_ (.Y(_06937_),
    .A(net900),
    .B(_06936_));
 sg13g2_nor3_1 _25971_ (.A(_06935_),
    .B(net668),
    .C(_06937_),
    .Y(_06938_));
 sg13g2_buf_4 _25972_ (.X(_06939_),
    .A(_06938_));
 sg13g2_mux2_1 _25973_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(net841),
    .S(_06939_),
    .X(_02539_));
 sg13g2_mux2_1 _25974_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(net1060),
    .S(_06939_),
    .X(_02540_));
 sg13g2_mux2_1 _25975_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(net921),
    .S(_06939_),
    .X(_02541_));
 sg13g2_mux2_1 _25976_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(net1024),
    .S(_06939_),
    .X(_02542_));
 sg13g2_mux2_1 _25977_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(net1022),
    .S(_06939_),
    .X(_02543_));
 sg13g2_mux2_1 _25978_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(net1054),
    .S(_06939_),
    .X(_02544_));
 sg13g2_mux2_1 _25979_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(net1053),
    .S(_06939_),
    .X(_02545_));
 sg13g2_mux2_1 _25980_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(net1056),
    .S(_06939_),
    .X(_02546_));
 sg13g2_and2_1 _25981_ (.A(net900),
    .B(_06936_),
    .X(_06940_));
 sg13g2_nand3_1 _25982_ (.B(_04915_),
    .C(_06940_),
    .A(_12086_),
    .Y(_06941_));
 sg13g2_buf_1 _25983_ (.A(_06941_),
    .X(_06942_));
 sg13g2_buf_1 _25984_ (.A(_06942_),
    .X(_06943_));
 sg13g2_nand2_1 _25985_ (.Y(_06944_),
    .A(\cpu.spi.r_clk_count[1][0] ),
    .B(net85));
 sg13g2_o21ai_1 _25986_ (.B1(_06944_),
    .Y(_02547_),
    .A1(net922),
    .A2(net85));
 sg13g2_nand2_1 _25987_ (.Y(_06945_),
    .A(\cpu.spi.r_clk_count[1][1] ),
    .B(_06943_));
 sg13g2_o21ai_1 _25988_ (.B1(_06945_),
    .Y(_02548_),
    .A1(net897),
    .A2(_06943_));
 sg13g2_nand2_1 _25989_ (.Y(_06946_),
    .A(\cpu.spi.r_clk_count[1][2] ),
    .B(_06942_));
 sg13g2_o21ai_1 _25990_ (.B1(_06946_),
    .Y(_02549_),
    .A1(net896),
    .A2(net85));
 sg13g2_mux2_1 _25991_ (.A0(net981),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net85),
    .X(_02550_));
 sg13g2_mux2_1 _25992_ (.A0(net856),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(net85),
    .X(_02551_));
 sg13g2_nand2_1 _25993_ (.Y(_06947_),
    .A(\cpu.spi.r_clk_count[1][5] ),
    .B(_06942_));
 sg13g2_o21ai_1 _25994_ (.B1(_06947_),
    .Y(_02552_),
    .A1(net895),
    .A2(net85));
 sg13g2_nand2_1 _25995_ (.Y(_06948_),
    .A(\cpu.spi.r_clk_count[1][6] ),
    .B(_06942_));
 sg13g2_o21ai_1 _25996_ (.B1(_06948_),
    .Y(_02553_),
    .A1(net894),
    .A2(net85));
 sg13g2_nand2_1 _25997_ (.Y(_06949_),
    .A(\cpu.spi.r_clk_count[1][7] ),
    .B(_06942_));
 sg13g2_o21ai_1 _25998_ (.B1(_06949_),
    .Y(_02554_),
    .A1(net893),
    .A2(net85));
 sg13g2_nand3_1 _25999_ (.B(_04915_),
    .C(_06936_),
    .A(_12080_),
    .Y(_06950_));
 sg13g2_buf_1 _26000_ (.A(_06950_),
    .X(_06951_));
 sg13g2_buf_1 _26001_ (.A(_06951_),
    .X(_06952_));
 sg13g2_nand2_1 _26002_ (.Y(_06953_),
    .A(_04950_),
    .B(net98));
 sg13g2_o21ai_1 _26003_ (.B1(_06953_),
    .Y(_02555_),
    .A1(net922),
    .A2(net98));
 sg13g2_nand2_1 _26004_ (.Y(_06954_),
    .A(_05370_),
    .B(net98));
 sg13g2_o21ai_1 _26005_ (.B1(_06954_),
    .Y(_02556_),
    .A1(net897),
    .A2(net98));
 sg13g2_nand2_1 _26006_ (.Y(_06955_),
    .A(_05427_),
    .B(_06951_));
 sg13g2_o21ai_1 _26007_ (.B1(_06955_),
    .Y(_02557_),
    .A1(net896),
    .A2(_06952_));
 sg13g2_mux2_1 _26008_ (.A0(net981),
    .A1(_05472_),
    .S(net98),
    .X(_02558_));
 sg13g2_mux2_1 _26009_ (.A0(net856),
    .A1(_05533_),
    .S(net98),
    .X(_02559_));
 sg13g2_nand2_1 _26010_ (.Y(_06956_),
    .A(_05606_),
    .B(_06951_));
 sg13g2_o21ai_1 _26011_ (.B1(_06956_),
    .Y(_02560_),
    .A1(net895),
    .A2(net98));
 sg13g2_nand2_1 _26012_ (.Y(_06957_),
    .A(_05681_),
    .B(_06951_));
 sg13g2_o21ai_1 _26013_ (.B1(_06957_),
    .Y(_02561_),
    .A1(net894),
    .A2(_06952_));
 sg13g2_nand2_1 _26014_ (.Y(_06958_),
    .A(_05103_),
    .B(_06951_));
 sg13g2_o21ai_1 _26015_ (.B1(_06958_),
    .Y(_02562_),
    .A1(net893),
    .A2(net98));
 sg13g2_mux2_1 _26016_ (.A0(\cpu.spi.r_clk_count[0][0] ),
    .A1(\cpu.spi.r_clk_count[1][0] ),
    .S(net677),
    .X(_06959_));
 sg13g2_nand2_1 _26017_ (.Y(_06960_),
    .A(net679),
    .B(_04950_));
 sg13g2_nand2_1 _26018_ (.Y(_06961_),
    .A(net677),
    .B(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_nand3_1 _26019_ (.B(_06960_),
    .C(_06961_),
    .A(net678),
    .Y(_06962_));
 sg13g2_o21ai_1 _26020_ (.B1(_06962_),
    .Y(_06963_),
    .A1(net620),
    .A2(_06959_));
 sg13g2_buf_2 _26021_ (.A(_00218_),
    .X(_06964_));
 sg13g2_nor4_1 _26022_ (.A(\cpu.spi.r_state[5] ),
    .B(net1150),
    .C(_09263_),
    .D(_12044_),
    .Y(_06965_));
 sg13g2_buf_1 _26023_ (.A(_06965_),
    .X(_06966_));
 sg13g2_nand2_1 _26024_ (.Y(_06967_),
    .A(_06964_),
    .B(net660));
 sg13g2_buf_2 _26025_ (.A(_06967_),
    .X(_06968_));
 sg13g2_buf_1 _26026_ (.A(_06968_),
    .X(_06969_));
 sg13g2_buf_1 _26027_ (.A(_09261_),
    .X(_06970_));
 sg13g2_buf_1 _26028_ (.A(net1119),
    .X(_06971_));
 sg13g2_mux2_1 _26029_ (.A0(_00294_),
    .A1(_00295_),
    .S(net958),
    .X(_06972_));
 sg13g2_nand2b_1 _26030_ (.Y(_06973_),
    .B(net1032),
    .A_N(_04950_));
 sg13g2_nand2b_1 _26031_ (.Y(_06974_),
    .B(_00295_),
    .A_N(_12054_));
 sg13g2_nand3_1 _26032_ (.B(_06973_),
    .C(_06974_),
    .A(_12064_),
    .Y(_06975_));
 sg13g2_o21ai_1 _26033_ (.B1(_06975_),
    .Y(_06976_),
    .A1(net772),
    .A2(_06972_));
 sg13g2_nor2_1 _26034_ (.A(_09230_),
    .B(net157),
    .Y(_06977_));
 sg13g2_a21oi_1 _26035_ (.A1(net111),
    .A2(_06976_),
    .Y(_06978_),
    .B1(_06977_));
 sg13g2_nor2_1 _26036_ (.A(_09230_),
    .B(_06966_),
    .Y(_06979_));
 sg13g2_o21ai_1 _26037_ (.B1(_06979_),
    .Y(_06980_),
    .A1(net352),
    .A2(_06976_));
 sg13g2_o21ai_1 _26038_ (.B1(_06980_),
    .Y(_06981_),
    .A1(_06970_),
    .A2(_06978_));
 sg13g2_nand2_1 _26039_ (.Y(_06982_),
    .A(net449),
    .B(_06981_));
 sg13g2_o21ai_1 _26040_ (.B1(_06982_),
    .Y(_06983_),
    .A1(_06963_),
    .A2(_06969_));
 sg13g2_and2_1 _26041_ (.A(_09300_),
    .B(net660),
    .X(_06984_));
 sg13g2_nor2_1 _26042_ (.A(_06964_),
    .B(net353),
    .Y(_06985_));
 sg13g2_nor2_1 _26043_ (.A(_09185_),
    .B(_09239_),
    .Y(_06986_));
 sg13g2_o21ai_1 _26044_ (.B1(_09302_),
    .Y(_06987_),
    .A1(_09202_),
    .A2(_06986_));
 sg13g2_a221oi_1 _26045_ (.B2(_09244_),
    .C1(_06987_),
    .B1(_06985_),
    .A1(_06964_),
    .Y(_06988_),
    .A2(_06984_));
 sg13g2_buf_1 _26046_ (.A(_06988_),
    .X(_06989_));
 sg13g2_mux2_1 _26047_ (.A0(_09230_),
    .A1(_06983_),
    .S(net67),
    .X(_02563_));
 sg13g2_nand2b_1 _26048_ (.Y(_06990_),
    .B(net770),
    .A_N(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_o21ai_1 _26049_ (.B1(_06990_),
    .Y(_06991_),
    .A1(net677),
    .A2(_05370_));
 sg13g2_mux2_1 _26050_ (.A0(\cpu.spi.r_clk_count[0][1] ),
    .A1(\cpu.spi.r_clk_count[1][1] ),
    .S(net770),
    .X(_06992_));
 sg13g2_nor2_1 _26051_ (.A(net769),
    .B(_06992_),
    .Y(_06993_));
 sg13g2_a21oi_1 _26052_ (.A1(net769),
    .A2(_06991_),
    .Y(_06994_),
    .B1(_06993_));
 sg13g2_nor2_1 _26053_ (.A(net449),
    .B(_06994_),
    .Y(_06995_));
 sg13g2_buf_1 _26054_ (.A(net839),
    .X(_06996_));
 sg13g2_mux2_1 _26055_ (.A0(_00299_),
    .A1(_00300_),
    .S(_06971_),
    .X(_06997_));
 sg13g2_nand2b_1 _26056_ (.Y(_06998_),
    .B(net958),
    .A_N(_05370_));
 sg13g2_nand2b_1 _26057_ (.Y(_06999_),
    .B(_00300_),
    .A_N(net1033));
 sg13g2_nand3_1 _26058_ (.B(_06998_),
    .C(_06999_),
    .A(net901),
    .Y(_07000_));
 sg13g2_o21ai_1 _26059_ (.B1(_07000_),
    .Y(_07001_),
    .A1(net772),
    .A2(_06997_));
 sg13g2_nor2_1 _26060_ (.A(net111),
    .B(_09232_),
    .Y(_07002_));
 sg13g2_a21oi_1 _26061_ (.A1(net111),
    .A2(_07001_),
    .Y(_07003_),
    .B1(_07002_));
 sg13g2_nand2_1 _26062_ (.Y(_07004_),
    .A(_09230_),
    .B(\cpu.spi.r_count[1] ));
 sg13g2_a21oi_1 _26063_ (.A1(_09232_),
    .A2(_07004_),
    .Y(_07005_),
    .B1(_06966_));
 sg13g2_o21ai_1 _26064_ (.B1(_07005_),
    .Y(_07006_),
    .A1(_09249_),
    .A2(_07001_));
 sg13g2_and2_1 _26065_ (.A(_06968_),
    .B(_07006_),
    .X(_07007_));
 sg13g2_o21ai_1 _26066_ (.B1(_07007_),
    .Y(_07008_),
    .A1(net736),
    .A2(_07003_));
 sg13g2_nand2_1 _26067_ (.Y(_07009_),
    .A(net67),
    .B(_07008_));
 sg13g2_o21ai_1 _26068_ (.B1(_09230_),
    .Y(_07010_),
    .A1(_06968_),
    .A2(_06994_));
 sg13g2_o21ai_1 _26069_ (.B1(net67),
    .Y(_07011_),
    .A1(_09202_),
    .A2(_07010_));
 sg13g2_nand2_1 _26070_ (.Y(_07012_),
    .A(\cpu.spi.r_count[1] ),
    .B(_07011_));
 sg13g2_o21ai_1 _26071_ (.B1(_07012_),
    .Y(_02564_),
    .A1(_06995_),
    .A2(_07009_));
 sg13g2_mux2_1 _26072_ (.A0(\cpu.spi.r_clk_count[0][2] ),
    .A1(\cpu.spi.r_clk_count[1][2] ),
    .S(net592),
    .X(_07013_));
 sg13g2_nand2_1 _26073_ (.Y(_07014_),
    .A(net679),
    .B(_05427_));
 sg13g2_nand2_1 _26074_ (.Y(_07015_),
    .A(net592),
    .B(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_nand3_1 _26075_ (.B(_07014_),
    .C(_07015_),
    .A(net678),
    .Y(_07016_));
 sg13g2_o21ai_1 _26076_ (.B1(_07016_),
    .Y(_07017_),
    .A1(net620),
    .A2(_07013_));
 sg13g2_mux2_1 _26077_ (.A0(_00096_),
    .A1(_00097_),
    .S(net958),
    .X(_07018_));
 sg13g2_nand2b_1 _26078_ (.Y(_07019_),
    .B(net1032),
    .A_N(_05427_));
 sg13g2_nand2b_1 _26079_ (.Y(_07020_),
    .B(_00097_),
    .A_N(net1033));
 sg13g2_nand3_1 _26080_ (.B(_07019_),
    .C(_07020_),
    .A(net901),
    .Y(_07021_));
 sg13g2_o21ai_1 _26081_ (.B1(_07021_),
    .Y(_07022_),
    .A1(net772),
    .A2(_07018_));
 sg13g2_xor2_1 _26082_ (.B(_09232_),
    .A(_09229_),
    .X(_07023_));
 sg13g2_nor2_1 _26083_ (.A(net157),
    .B(_07023_),
    .Y(_07024_));
 sg13g2_a21oi_1 _26084_ (.A1(net111),
    .A2(_07022_),
    .Y(_07025_),
    .B1(_07024_));
 sg13g2_nor2_1 _26085_ (.A(net660),
    .B(_07023_),
    .Y(_07026_));
 sg13g2_o21ai_1 _26086_ (.B1(_07026_),
    .Y(_07027_),
    .A1(net352),
    .A2(_07022_));
 sg13g2_o21ai_1 _26087_ (.B1(_07027_),
    .Y(_07028_),
    .A1(net839),
    .A2(_07025_));
 sg13g2_nand2_1 _26088_ (.Y(_07029_),
    .A(net449),
    .B(_07028_));
 sg13g2_o21ai_1 _26089_ (.B1(_07029_),
    .Y(_07030_),
    .A1(net449),
    .A2(_07017_));
 sg13g2_mux2_1 _26090_ (.A0(_09229_),
    .A1(_07030_),
    .S(net67),
    .X(_02565_));
 sg13g2_mux2_1 _26091_ (.A0(\cpu.spi.r_clk_count[0][3] ),
    .A1(\cpu.spi.r_clk_count[1][3] ),
    .S(net592),
    .X(_07031_));
 sg13g2_nand2_1 _26092_ (.Y(_07032_),
    .A(net679),
    .B(_05472_));
 sg13g2_nand2_1 _26093_ (.Y(_07033_),
    .A(net592),
    .B(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_nand3_1 _26094_ (.B(_07032_),
    .C(_07033_),
    .A(net678),
    .Y(_07034_));
 sg13g2_o21ai_1 _26095_ (.B1(_07034_),
    .Y(_07035_),
    .A1(net620),
    .A2(_07031_));
 sg13g2_mux2_1 _26096_ (.A0(_00107_),
    .A1(_00108_),
    .S(net958),
    .X(_07036_));
 sg13g2_nand2b_1 _26097_ (.Y(_07037_),
    .B(net1032),
    .A_N(_05472_));
 sg13g2_nand2b_1 _26098_ (.Y(_07038_),
    .B(_00108_),
    .A_N(net1033));
 sg13g2_nand3_1 _26099_ (.B(_07037_),
    .C(_07038_),
    .A(net901),
    .Y(_07039_));
 sg13g2_o21ai_1 _26100_ (.B1(_07039_),
    .Y(_07040_),
    .A1(net772),
    .A2(_07036_));
 sg13g2_nor2_1 _26101_ (.A(_09229_),
    .B(_09232_),
    .Y(_07041_));
 sg13g2_xnor2_1 _26102_ (.Y(_07042_),
    .A(\cpu.spi.r_count[3] ),
    .B(_07041_));
 sg13g2_nor2_1 _26103_ (.A(net157),
    .B(_07042_),
    .Y(_07043_));
 sg13g2_a21oi_1 _26104_ (.A1(net111),
    .A2(_07040_),
    .Y(_07044_),
    .B1(_07043_));
 sg13g2_nor2_1 _26105_ (.A(net660),
    .B(_07042_),
    .Y(_07045_));
 sg13g2_o21ai_1 _26106_ (.B1(_07045_),
    .Y(_07046_),
    .A1(net352),
    .A2(_07040_));
 sg13g2_o21ai_1 _26107_ (.B1(_07046_),
    .Y(_07047_),
    .A1(net839),
    .A2(_07044_));
 sg13g2_nand2_1 _26108_ (.Y(_07048_),
    .A(net449),
    .B(_07047_));
 sg13g2_o21ai_1 _26109_ (.B1(_07048_),
    .Y(_07049_),
    .A1(net449),
    .A2(_07035_));
 sg13g2_mux2_1 _26110_ (.A0(\cpu.spi.r_count[3] ),
    .A1(_07049_),
    .S(net67),
    .X(_02566_));
 sg13g2_mux2_1 _26111_ (.A0(\cpu.spi.r_clk_count[0][4] ),
    .A1(\cpu.spi.r_clk_count[1][4] ),
    .S(_06935_),
    .X(_07050_));
 sg13g2_nand2_1 _26112_ (.Y(_07051_),
    .A(net679),
    .B(_05533_));
 sg13g2_nand2_1 _26113_ (.Y(_07052_),
    .A(net592),
    .B(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_nand3_1 _26114_ (.B(_07051_),
    .C(_07052_),
    .A(net678),
    .Y(_07053_));
 sg13g2_o21ai_1 _26115_ (.B1(_07053_),
    .Y(_07054_),
    .A1(net620),
    .A2(_07050_));
 sg13g2_mux2_1 _26116_ (.A0(_00118_),
    .A1(_00119_),
    .S(net958),
    .X(_07055_));
 sg13g2_nand2b_1 _26117_ (.Y(_07056_),
    .B(net1032),
    .A_N(_05533_));
 sg13g2_nand2b_1 _26118_ (.Y(_07057_),
    .B(_00119_),
    .A_N(net1033));
 sg13g2_nand3_1 _26119_ (.B(_07056_),
    .C(_07057_),
    .A(net901),
    .Y(_07058_));
 sg13g2_o21ai_1 _26120_ (.B1(_07058_),
    .Y(_07059_),
    .A1(net772),
    .A2(_07055_));
 sg13g2_xnor2_1 _26121_ (.Y(_07060_),
    .A(\cpu.spi.r_count[4] ),
    .B(_09233_));
 sg13g2_nor2_1 _26122_ (.A(net157),
    .B(_07060_),
    .Y(_07061_));
 sg13g2_a21oi_1 _26123_ (.A1(net111),
    .A2(_07059_),
    .Y(_07062_),
    .B1(_07061_));
 sg13g2_nor2_1 _26124_ (.A(net660),
    .B(_07060_),
    .Y(_07063_));
 sg13g2_o21ai_1 _26125_ (.B1(_07063_),
    .Y(_07064_),
    .A1(net352),
    .A2(_07059_));
 sg13g2_o21ai_1 _26126_ (.B1(_07064_),
    .Y(_07065_),
    .A1(net839),
    .A2(_07062_));
 sg13g2_nand2_1 _26127_ (.Y(_07066_),
    .A(_06968_),
    .B(_07065_));
 sg13g2_o21ai_1 _26128_ (.B1(_07066_),
    .Y(_07067_),
    .A1(net449),
    .A2(_07054_));
 sg13g2_mux2_1 _26129_ (.A0(\cpu.spi.r_count[4] ),
    .A1(_07067_),
    .S(net67),
    .X(_02567_));
 sg13g2_mux2_1 _26130_ (.A0(\cpu.spi.r_clk_count[0][5] ),
    .A1(\cpu.spi.r_clk_count[1][5] ),
    .S(net592),
    .X(_07068_));
 sg13g2_nand2_1 _26131_ (.Y(_07069_),
    .A(net679),
    .B(_05606_));
 sg13g2_nand2_1 _26132_ (.Y(_07070_),
    .A(net592),
    .B(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_nand3_1 _26133_ (.B(_07069_),
    .C(_07070_),
    .A(net678),
    .Y(_07071_));
 sg13g2_o21ai_1 _26134_ (.B1(_07071_),
    .Y(_07072_),
    .A1(net620),
    .A2(_07068_));
 sg13g2_mux2_1 _26135_ (.A0(_00125_),
    .A1(_00126_),
    .S(net958),
    .X(_07073_));
 sg13g2_nand2b_1 _26136_ (.Y(_07074_),
    .B(net1032),
    .A_N(_05606_));
 sg13g2_nand2b_1 _26137_ (.Y(_07075_),
    .B(_00126_),
    .A_N(net1033));
 sg13g2_nand3_1 _26138_ (.B(_07074_),
    .C(_07075_),
    .A(net901),
    .Y(_07076_));
 sg13g2_o21ai_1 _26139_ (.B1(_07076_),
    .Y(_07077_),
    .A1(net772),
    .A2(_07073_));
 sg13g2_xnor2_1 _26140_ (.Y(_07078_),
    .A(\cpu.spi.r_count[5] ),
    .B(_09234_));
 sg13g2_nor2_1 _26141_ (.A(net157),
    .B(_07078_),
    .Y(_07079_));
 sg13g2_a21oi_1 _26142_ (.A1(net111),
    .A2(_07077_),
    .Y(_07080_),
    .B1(_07079_));
 sg13g2_nor2_1 _26143_ (.A(net660),
    .B(_07078_),
    .Y(_07081_));
 sg13g2_o21ai_1 _26144_ (.B1(_07081_),
    .Y(_07082_),
    .A1(net352),
    .A2(_07077_));
 sg13g2_o21ai_1 _26145_ (.B1(_07082_),
    .Y(_07083_),
    .A1(net839),
    .A2(_07080_));
 sg13g2_nand2_1 _26146_ (.Y(_07084_),
    .A(_06968_),
    .B(_07083_));
 sg13g2_o21ai_1 _26147_ (.B1(_07084_),
    .Y(_07085_),
    .A1(net449),
    .A2(_07072_));
 sg13g2_mux2_1 _26148_ (.A0(\cpu.spi.r_count[5] ),
    .A1(_07085_),
    .S(net67),
    .X(_02568_));
 sg13g2_mux2_1 _26149_ (.A0(\cpu.spi.r_clk_count[0][6] ),
    .A1(\cpu.spi.r_clk_count[1][6] ),
    .S(net677),
    .X(_07086_));
 sg13g2_nand2_1 _26150_ (.Y(_07087_),
    .A(net679),
    .B(_05681_));
 sg13g2_nand2_1 _26151_ (.Y(_07088_),
    .A(net592),
    .B(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_nand3_1 _26152_ (.B(_07087_),
    .C(_07088_),
    .A(net678),
    .Y(_07089_));
 sg13g2_o21ai_1 _26153_ (.B1(_07089_),
    .Y(_07090_),
    .A1(net620),
    .A2(_07086_));
 sg13g2_mux2_1 _26154_ (.A0(_00137_),
    .A1(_00138_),
    .S(net958),
    .X(_07091_));
 sg13g2_nand2b_1 _26155_ (.Y(_07092_),
    .B(net958),
    .A_N(_05681_));
 sg13g2_nand2b_1 _26156_ (.Y(_07093_),
    .B(_00138_),
    .A_N(net1033));
 sg13g2_nand3_1 _26157_ (.B(_07092_),
    .C(_07093_),
    .A(net901),
    .Y(_07094_));
 sg13g2_o21ai_1 _26158_ (.B1(_07094_),
    .Y(_07095_),
    .A1(net772),
    .A2(_07091_));
 sg13g2_xnor2_1 _26159_ (.Y(_07096_),
    .A(\cpu.spi.r_count[6] ),
    .B(_09235_));
 sg13g2_nor2_1 _26160_ (.A(net157),
    .B(_07096_),
    .Y(_07097_));
 sg13g2_a21oi_1 _26161_ (.A1(net157),
    .A2(_07095_),
    .Y(_07098_),
    .B1(_07097_));
 sg13g2_nor2_1 _26162_ (.A(net660),
    .B(_07096_),
    .Y(_07099_));
 sg13g2_o21ai_1 _26163_ (.B1(_07099_),
    .Y(_07100_),
    .A1(net352),
    .A2(_07095_));
 sg13g2_o21ai_1 _26164_ (.B1(_07100_),
    .Y(_07101_),
    .A1(net839),
    .A2(_07098_));
 sg13g2_nand2_1 _26165_ (.Y(_07102_),
    .A(_06968_),
    .B(_07101_));
 sg13g2_o21ai_1 _26166_ (.B1(_07102_),
    .Y(_07103_),
    .A1(_06969_),
    .A2(_07090_));
 sg13g2_mux2_1 _26167_ (.A0(\cpu.spi.r_count[6] ),
    .A1(_07103_),
    .S(_06989_),
    .X(_02569_));
 sg13g2_nand2b_1 _26168_ (.Y(_07104_),
    .B(net770),
    .A_N(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_o21ai_1 _26169_ (.B1(_07104_),
    .Y(_07105_),
    .A1(net770),
    .A2(_05103_));
 sg13g2_mux2_1 _26170_ (.A0(\cpu.spi.r_clk_count[0][7] ),
    .A1(\cpu.spi.r_clk_count[1][7] ),
    .S(net770),
    .X(_07106_));
 sg13g2_nor2_1 _26171_ (.A(net769),
    .B(_07106_),
    .Y(_07107_));
 sg13g2_a21oi_1 _26172_ (.A1(net769),
    .A2(_07105_),
    .Y(_07108_),
    .B1(_07107_));
 sg13g2_nor2_1 _26173_ (.A(_06968_),
    .B(_07108_),
    .Y(_07109_));
 sg13g2_nor3_1 _26174_ (.A(_09202_),
    .B(_09237_),
    .C(_07109_),
    .Y(_07110_));
 sg13g2_nand2b_1 _26175_ (.Y(_07111_),
    .B(_06989_),
    .A_N(_07110_));
 sg13g2_nand2b_1 _26176_ (.Y(_07112_),
    .B(net1119),
    .A_N(_00150_));
 sg13g2_o21ai_1 _26177_ (.B1(_07112_),
    .Y(_07113_),
    .A1(net1033),
    .A2(_00149_));
 sg13g2_nor2b_1 _26178_ (.A(_05103_),
    .B_N(net1119),
    .Y(_07114_));
 sg13g2_nor2b_1 _26179_ (.A(net1119),
    .B_N(_00150_),
    .Y(_07115_));
 sg13g2_nor3_1 _26180_ (.A(_12051_),
    .B(_07114_),
    .C(_07115_),
    .Y(_07116_));
 sg13g2_a21oi_1 _26181_ (.A1(_12051_),
    .A2(_07113_),
    .Y(_07117_),
    .B1(_07116_));
 sg13g2_nor2_1 _26182_ (.A(_09244_),
    .B(net353),
    .Y(_07118_));
 sg13g2_a21oi_1 _26183_ (.A1(net111),
    .A2(_07117_),
    .Y(_07119_),
    .B1(_07118_));
 sg13g2_nor2_1 _26184_ (.A(_09228_),
    .B(_07117_),
    .Y(_07120_));
 sg13g2_nor2b_1 _26185_ (.A(_09237_),
    .B_N(_09228_),
    .Y(_07121_));
 sg13g2_a21oi_1 _26186_ (.A1(_09237_),
    .A2(_07120_),
    .Y(_07122_),
    .B1(_07121_));
 sg13g2_o21ai_1 _26187_ (.B1(_06968_),
    .Y(_07123_),
    .A1(net660),
    .A2(_07122_));
 sg13g2_a21oi_1 _26188_ (.A1(net1031),
    .A2(_07119_),
    .Y(_07124_),
    .B1(_07123_));
 sg13g2_nor2_1 _26189_ (.A(_07109_),
    .B(_07124_),
    .Y(_07125_));
 sg13g2_a22oi_1 _26190_ (.Y(_07126_),
    .B1(_07125_),
    .B2(net67),
    .A2(_07111_),
    .A1(_09228_));
 sg13g2_inv_1 _26191_ (.Y(_02570_),
    .A(_07126_));
 sg13g2_mux4_1 _26192_ (.S0(_04850_),
    .A0(_09137_),
    .A1(_09145_),
    .A2(_09151_),
    .A3(_09139_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07127_));
 sg13g2_nand2_1 _26193_ (.Y(_07128_),
    .A(_09132_),
    .B(_04850_));
 sg13g2_nand2b_1 _26194_ (.Y(_07129_),
    .B(_09131_),
    .A_N(_04850_));
 sg13g2_nand3_1 _26195_ (.B(_07128_),
    .C(_07129_),
    .A(_06327_),
    .Y(_07130_));
 sg13g2_o21ai_1 _26196_ (.B1(_07130_),
    .Y(_07131_),
    .A1(_06327_),
    .A2(_07127_));
 sg13g2_mux2_1 _26197_ (.A0(_09141_),
    .A1(_09142_),
    .S(_04850_),
    .X(_07132_));
 sg13g2_inv_1 _26198_ (.Y(_07133_),
    .A(_00102_));
 sg13g2_o21ai_1 _26199_ (.B1(_07133_),
    .Y(_07134_),
    .A1(_06324_),
    .A2(_07132_));
 sg13g2_mux4_1 _26200_ (.S0(_04850_),
    .A0(_09149_),
    .A1(_09126_),
    .A2(_09147_),
    .A3(_09128_),
    .S1(\cpu.gpio.r_spi_miso_src[0][2] ),
    .X(_07135_));
 sg13g2_nor3_1 _26201_ (.A(_06324_),
    .B(_06327_),
    .C(_07135_),
    .Y(_07136_));
 sg13g2_a221oi_1 _26202_ (.B2(_06327_),
    .C1(_07136_),
    .B1(_07134_),
    .A1(_06324_),
    .Y(_07137_),
    .A2(_07131_));
 sg13g2_inv_1 _26203_ (.Y(_07138_),
    .A(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_mux4_1 _26204_ (.S0(_05554_),
    .A0(_09149_),
    .A1(_09126_),
    .A2(_09147_),
    .A3(_09128_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07139_));
 sg13g2_nand2_1 _26205_ (.Y(_07140_),
    .A(_09142_),
    .B(_05554_));
 sg13g2_nand2b_1 _26206_ (.Y(_07141_),
    .B(_09141_),
    .A_N(_05554_));
 sg13g2_nand3_1 _26207_ (.B(_07140_),
    .C(_07141_),
    .A(_06330_),
    .Y(_07142_));
 sg13g2_o21ai_1 _26208_ (.B1(_07142_),
    .Y(_07143_),
    .A1(_06330_),
    .A2(_07139_));
 sg13g2_nand2b_1 _26209_ (.Y(_07144_),
    .B(_05554_),
    .A_N(_09132_));
 sg13g2_o21ai_1 _26210_ (.B1(_07144_),
    .Y(_07145_),
    .A1(_09131_),
    .A2(_05554_));
 sg13g2_a21o_1 _26211_ (.A2(_07145_),
    .A1(\cpu.gpio.r_spi_miso_src[1][1] ),
    .B1(_00143_),
    .X(_07146_));
 sg13g2_mux4_1 _26212_ (.S0(_05554_),
    .A0(_09137_),
    .A1(_09145_),
    .A2(_09151_),
    .A3(_09139_),
    .S1(\cpu.gpio.r_spi_miso_src[1][2] ),
    .X(_07147_));
 sg13g2_nor3_1 _26213_ (.A(_07138_),
    .B(_06330_),
    .C(_07147_),
    .Y(_07148_));
 sg13g2_a221oi_1 _26214_ (.B2(_06330_),
    .C1(_07148_),
    .B1(_07146_),
    .A1(_07138_),
    .Y(_07149_),
    .A2(_07143_));
 sg13g2_mux2_1 _26215_ (.A0(_07137_),
    .A1(_07149_),
    .S(_12060_),
    .X(_07150_));
 sg13g2_nor3_1 _26216_ (.A(_09251_),
    .B(_09254_),
    .C(_12108_),
    .Y(_07151_));
 sg13g2_nand3_1 _26217_ (.B(_09254_),
    .C(net553),
    .A(_09251_),
    .Y(_07152_));
 sg13g2_nand2b_1 _26218_ (.Y(_07153_),
    .B(_07152_),
    .A_N(_07151_));
 sg13g2_nand3_1 _26219_ (.B(net353),
    .C(_07153_),
    .A(net933),
    .Y(_07154_));
 sg13g2_buf_4 _26220_ (.X(_07155_),
    .A(_07154_));
 sg13g2_mux2_1 _26221_ (.A0(_07150_),
    .A1(_09217_),
    .S(_07155_),
    .X(_02574_));
 sg13g2_mux2_1 _26222_ (.A0(_09217_),
    .A1(_09216_),
    .S(_07155_),
    .X(_02575_));
 sg13g2_mux2_1 _26223_ (.A0(_09216_),
    .A1(_09220_),
    .S(_07155_),
    .X(_02576_));
 sg13g2_mux2_1 _26224_ (.A0(_09220_),
    .A1(_09215_),
    .S(_07155_),
    .X(_02577_));
 sg13g2_mux2_1 _26225_ (.A0(_09215_),
    .A1(_09222_),
    .S(_07155_),
    .X(_02578_));
 sg13g2_mux2_1 _26226_ (.A0(_09222_),
    .A1(_09221_),
    .S(_07155_),
    .X(_02579_));
 sg13g2_mux2_1 _26227_ (.A0(_09221_),
    .A1(_09223_),
    .S(_07155_),
    .X(_02580_));
 sg13g2_mux2_1 _26228_ (.A0(_09223_),
    .A1(\cpu.spi.r_in[7] ),
    .S(_07155_),
    .X(_02581_));
 sg13g2_nor4_2 _26229_ (.A(net533),
    .B(net566),
    .C(net616),
    .Y(_07156_),
    .D(_06937_));
 sg13g2_mux2_1 _26230_ (.A0(\cpu.spi.r_mode[0][0] ),
    .A1(net841),
    .S(_07156_),
    .X(_02583_));
 sg13g2_mux2_1 _26231_ (.A0(_12066_),
    .A1(net1060),
    .S(_07156_),
    .X(_02584_));
 sg13g2_nand3_1 _26232_ (.B(_09181_),
    .C(_06940_),
    .A(net616),
    .Y(_07157_));
 sg13g2_buf_1 _26233_ (.A(_07157_),
    .X(_07158_));
 sg13g2_nand2_1 _26234_ (.Y(_07159_),
    .A(\cpu.spi.r_mode[1][0] ),
    .B(_07158_));
 sg13g2_o21ai_1 _26235_ (.B1(_07159_),
    .Y(_02585_),
    .A1(net922),
    .A2(_07158_));
 sg13g2_nand2_1 _26236_ (.Y(_07160_),
    .A(_12071_),
    .B(_07158_));
 sg13g2_o21ai_1 _26237_ (.B1(_07160_),
    .Y(_02586_),
    .A1(net897),
    .A2(_07158_));
 sg13g2_nand3_1 _26238_ (.B(_12080_),
    .C(_06936_),
    .A(_09181_),
    .Y(_07161_));
 sg13g2_buf_1 _26239_ (.A(_07161_),
    .X(_07162_));
 sg13g2_nand2_1 _26240_ (.Y(_07163_),
    .A(\cpu.spi.r_mode[2][0] ),
    .B(_07162_));
 sg13g2_o21ai_1 _26241_ (.B1(_07163_),
    .Y(_02587_),
    .A1(net922),
    .A2(_07162_));
 sg13g2_nand2_1 _26242_ (.Y(_07164_),
    .A(_12067_),
    .B(_07162_));
 sg13g2_o21ai_1 _26243_ (.B1(_07164_),
    .Y(_02588_),
    .A1(net897),
    .A2(_07162_));
 sg13g2_nor3_1 _26244_ (.A(_09200_),
    .B(_09265_),
    .C(_12050_),
    .Y(_07165_));
 sg13g2_a21oi_1 _26245_ (.A1(net1150),
    .A2(_12112_),
    .Y(_07166_),
    .B1(_07165_));
 sg13g2_nand4_1 _26246_ (.B(_09302_),
    .C(_12116_),
    .A(_09202_),
    .Y(_07167_),
    .D(_07166_));
 sg13g2_buf_1 _26247_ (.A(_07167_),
    .X(_07168_));
 sg13g2_nand2b_1 _26248_ (.Y(_07169_),
    .B(_00216_),
    .A_N(net553));
 sg13g2_nor2_1 _26249_ (.A(_06970_),
    .B(_06964_),
    .Y(_07170_));
 sg13g2_a221oi_1 _26250_ (.B2(_07170_),
    .C1(net768),
    .B1(_07169_),
    .A1(net736),
    .Y(_07171_),
    .A2(net960));
 sg13g2_nand2_1 _26251_ (.Y(_07172_),
    .A(\cpu.spi.r_out[0] ),
    .B(net76));
 sg13g2_o21ai_1 _26252_ (.B1(_07172_),
    .Y(_02589_),
    .A1(net76),
    .A2(_07171_));
 sg13g2_mux2_1 _26253_ (.A0(_00176_),
    .A1(_00216_),
    .S(net553),
    .X(_07173_));
 sg13g2_nor2_1 _26254_ (.A(_09200_),
    .B(_12050_),
    .Y(_07174_));
 sg13g2_buf_2 _26255_ (.A(_07174_),
    .X(_07175_));
 sg13g2_a22oi_1 _26256_ (.Y(_07176_),
    .B1(_07175_),
    .B2(_09978_),
    .A2(net768),
    .A1(\cpu.spi.r_out[0] ));
 sg13g2_o21ai_1 _26257_ (.B1(_07176_),
    .Y(_07177_),
    .A1(net736),
    .A2(_07173_));
 sg13g2_mux2_1 _26258_ (.A0(_07177_),
    .A1(\cpu.spi.r_out[1] ),
    .S(net76),
    .X(_02590_));
 sg13g2_mux2_1 _26259_ (.A0(_00177_),
    .A1(_00176_),
    .S(net553),
    .X(_07178_));
 sg13g2_a22oi_1 _26260_ (.Y(_07179_),
    .B1(_07175_),
    .B2(net1059),
    .A2(net768),
    .A1(\cpu.spi.r_out[1] ));
 sg13g2_o21ai_1 _26261_ (.B1(_07179_),
    .Y(_07180_),
    .A1(net736),
    .A2(_07178_));
 sg13g2_mux2_1 _26262_ (.A0(_07180_),
    .A1(\cpu.spi.r_out[2] ),
    .S(net76),
    .X(_02591_));
 sg13g2_mux2_1 _26263_ (.A0(_00280_),
    .A1(_00177_),
    .S(net553),
    .X(_07181_));
 sg13g2_a22oi_1 _26264_ (.Y(_07182_),
    .B1(_07175_),
    .B2(net1144),
    .A2(net768),
    .A1(\cpu.spi.r_out[2] ));
 sg13g2_o21ai_1 _26265_ (.B1(_07182_),
    .Y(_07183_),
    .A1(net736),
    .A2(_07181_));
 sg13g2_mux2_1 _26266_ (.A0(_07183_),
    .A1(\cpu.spi.r_out[3] ),
    .S(net76),
    .X(_02592_));
 sg13g2_mux2_1 _26267_ (.A0(_00178_),
    .A1(_00280_),
    .S(net553),
    .X(_07184_));
 sg13g2_a22oi_1 _26268_ (.Y(_07185_),
    .B1(_07175_),
    .B2(_09999_),
    .A2(net768),
    .A1(\cpu.spi.r_out[3] ));
 sg13g2_o21ai_1 _26269_ (.B1(_07185_),
    .Y(_07186_),
    .A1(net736),
    .A2(_07184_));
 sg13g2_mux2_1 _26270_ (.A0(_07186_),
    .A1(\cpu.spi.r_out[4] ),
    .S(_07168_),
    .X(_02593_));
 sg13g2_mux2_1 _26271_ (.A0(_00179_),
    .A1(_00178_),
    .S(net553),
    .X(_07187_));
 sg13g2_a22oi_1 _26272_ (.Y(_07188_),
    .B1(_07175_),
    .B2(_10005_),
    .A2(_12097_),
    .A1(\cpu.spi.r_out[4] ));
 sg13g2_o21ai_1 _26273_ (.B1(_07188_),
    .Y(_07189_),
    .A1(net736),
    .A2(_07187_));
 sg13g2_mux2_1 _26274_ (.A0(_07189_),
    .A1(\cpu.spi.r_out[5] ),
    .S(net76),
    .X(_02594_));
 sg13g2_buf_1 _26275_ (.A(_00180_),
    .X(_07190_));
 sg13g2_mux2_1 _26276_ (.A0(_07190_),
    .A1(_00179_),
    .S(_12109_),
    .X(_07191_));
 sg13g2_a22oi_1 _26277_ (.Y(_07192_),
    .B1(_07175_),
    .B2(_10010_),
    .A2(net768),
    .A1(\cpu.spi.r_out[5] ));
 sg13g2_o21ai_1 _26278_ (.B1(_07192_),
    .Y(_07193_),
    .A1(_06996_),
    .A2(_07191_));
 sg13g2_mux2_1 _26279_ (.A0(_07193_),
    .A1(\cpu.spi.r_out[6] ),
    .S(net76),
    .X(_02595_));
 sg13g2_buf_1 _26280_ (.A(_00274_),
    .X(_07194_));
 sg13g2_mux2_1 _26281_ (.A0(_07194_),
    .A1(_07190_),
    .S(_12109_),
    .X(_07195_));
 sg13g2_a22oi_1 _26282_ (.Y(_07196_),
    .B1(_07175_),
    .B2(_10015_),
    .A2(net768),
    .A1(\cpu.spi.r_out[6] ));
 sg13g2_o21ai_1 _26283_ (.B1(_07196_),
    .Y(_07197_),
    .A1(_06996_),
    .A2(_07195_));
 sg13g2_mux2_1 _26284_ (.A0(_07197_),
    .A1(\cpu.spi.r_out[7] ),
    .S(net76),
    .X(_02596_));
 sg13g2_nand2_1 _26285_ (.Y(_07198_),
    .A(_12051_),
    .B(_09267_));
 sg13g2_o21ai_1 _26286_ (.B1(_07198_),
    .Y(_02599_),
    .A1(_03677_),
    .A2(_09267_));
 sg13g2_nand2_1 _26287_ (.Y(_07199_),
    .A(net1032),
    .B(_09267_));
 sg13g2_o21ai_1 _26288_ (.B1(_07199_),
    .Y(_02600_),
    .A1(_03050_),
    .A2(_09267_));
 sg13g2_mux2_1 _26289_ (.A0(\cpu.spi.r_src[0] ),
    .A1(net921),
    .S(_07156_),
    .X(_02601_));
 sg13g2_nand2_1 _26290_ (.Y(_07200_),
    .A(\cpu.spi.r_src[1] ),
    .B(_07158_));
 sg13g2_o21ai_1 _26291_ (.B1(_07200_),
    .Y(_02602_),
    .A1(net896),
    .A2(_07158_));
 sg13g2_nand2_1 _26292_ (.Y(_07201_),
    .A(_12056_),
    .B(_07162_));
 sg13g2_o21ai_1 _26293_ (.B1(_07201_),
    .Y(_02603_),
    .A1(net896),
    .A2(_07162_));
 sg13g2_and2_1 _26294_ (.A(_09197_),
    .B(_05105_),
    .X(_07202_));
 sg13g2_buf_4 _26295_ (.X(_07203_),
    .A(_07202_));
 sg13g2_mux2_1 _26296_ (.A0(\cpu.spi.r_timeout[0] ),
    .A1(net841),
    .S(_07203_),
    .X(_02604_));
 sg13g2_mux2_1 _26297_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(net1060),
    .S(_07203_),
    .X(_02605_));
 sg13g2_mux2_1 _26298_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(net921),
    .S(_07203_),
    .X(_02606_));
 sg13g2_mux2_1 _26299_ (.A0(\cpu.spi.r_timeout[3] ),
    .A1(net1024),
    .S(_07203_),
    .X(_02607_));
 sg13g2_mux2_1 _26300_ (.A0(\cpu.spi.r_timeout[4] ),
    .A1(net1022),
    .S(_07203_),
    .X(_02608_));
 sg13g2_mux2_1 _26301_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(net1054),
    .S(_07203_),
    .X(_02609_));
 sg13g2_mux2_1 _26302_ (.A0(\cpu.spi.r_timeout[6] ),
    .A1(net1053),
    .S(_07203_),
    .X(_02610_));
 sg13g2_mux2_1 _26303_ (.A0(\cpu.spi.r_timeout[7] ),
    .A1(net1056),
    .S(_07203_),
    .X(_02611_));
 sg13g2_inv_1 _26304_ (.Y(_07204_),
    .A(\cpu.spi.r_timeout_count[0] ));
 sg13g2_nor2_1 _26305_ (.A(_09251_),
    .B(net1152),
    .Y(_07205_));
 sg13g2_a21oi_1 _26306_ (.A1(net1152),
    .A2(_09199_),
    .Y(_07206_),
    .B1(_07205_));
 sg13g2_nor2_1 _26307_ (.A(_09227_),
    .B(_09249_),
    .Y(_07207_));
 sg13g2_nor2_1 _26308_ (.A(_09251_),
    .B(_07207_),
    .Y(_07208_));
 sg13g2_nor4_1 _26309_ (.A(_00219_),
    .B(_09206_),
    .C(_09227_),
    .D(_09249_),
    .Y(_07209_));
 sg13g2_nor4_1 _26310_ (.A(net929),
    .B(_07206_),
    .C(_07208_),
    .D(_07209_),
    .Y(_07210_));
 sg13g2_buf_2 _26311_ (.A(_07210_),
    .X(_07211_));
 sg13g2_buf_1 _26312_ (.A(_07211_),
    .X(_07212_));
 sg13g2_mux2_1 _26313_ (.A0(_00277_),
    .A1(\cpu.spi.r_timeout[0] ),
    .S(net1031),
    .X(_07213_));
 sg13g2_nand2_1 _26314_ (.Y(_07214_),
    .A(net75),
    .B(_07213_));
 sg13g2_o21ai_1 _26315_ (.B1(_07214_),
    .Y(_02612_),
    .A1(_07204_),
    .A2(net75));
 sg13g2_o21ai_1 _26316_ (.B1(_07212_),
    .Y(_07215_),
    .A1(_07204_),
    .A2(net1066));
 sg13g2_nor2_1 _26317_ (.A(\cpu.spi.r_timeout_count[0] ),
    .B(\cpu.spi.r_timeout_count[1] ),
    .Y(_07216_));
 sg13g2_mux2_1 _26318_ (.A0(\cpu.spi.r_timeout[1] ),
    .A1(_07216_),
    .S(net736),
    .X(_07217_));
 sg13g2_a22oi_1 _26319_ (.Y(_07218_),
    .B1(_07217_),
    .B2(_07212_),
    .A2(_07215_),
    .A1(\cpu.spi.r_timeout_count[1] ));
 sg13g2_inv_1 _26320_ (.Y(_02613_),
    .A(_07218_));
 sg13g2_o21ai_1 _26321_ (.B1(_07211_),
    .Y(_07219_),
    .A1(net1066),
    .A2(_07216_));
 sg13g2_mux2_1 _26322_ (.A0(\cpu.spi.r_timeout[2] ),
    .A1(_09207_),
    .S(net839),
    .X(_07220_));
 sg13g2_a22oi_1 _26323_ (.Y(_07221_),
    .B1(_07220_),
    .B2(net75),
    .A2(_07219_),
    .A1(\cpu.spi.r_timeout_count[2] ));
 sg13g2_inv_1 _26324_ (.Y(_02614_),
    .A(_07221_));
 sg13g2_o21ai_1 _26325_ (.B1(_07211_),
    .Y(_07222_),
    .A1(net1066),
    .A2(_09207_));
 sg13g2_nand2b_1 _26326_ (.Y(_07223_),
    .B(_09207_),
    .A_N(\cpu.spi.r_timeout_count[3] ));
 sg13g2_nand2_1 _26327_ (.Y(_07224_),
    .A(net1031),
    .B(\cpu.spi.r_timeout[3] ));
 sg13g2_o21ai_1 _26328_ (.B1(_07224_),
    .Y(_07225_),
    .A1(net1066),
    .A2(_07223_));
 sg13g2_a22oi_1 _26329_ (.Y(_07226_),
    .B1(_07225_),
    .B2(net75),
    .A2(_07222_),
    .A1(\cpu.spi.r_timeout_count[3] ));
 sg13g2_inv_1 _26330_ (.Y(_02615_),
    .A(_07226_));
 sg13g2_o21ai_1 _26331_ (.B1(_07211_),
    .Y(_07227_),
    .A1(net1066),
    .A2(_09208_));
 sg13g2_nand2_1 _26332_ (.Y(_07228_),
    .A(net1031),
    .B(\cpu.spi.r_timeout[4] ));
 sg13g2_o21ai_1 _26333_ (.B1(_07228_),
    .Y(_07229_),
    .A1(net1066),
    .A2(_09209_));
 sg13g2_a22oi_1 _26334_ (.Y(_07230_),
    .B1(_07229_),
    .B2(net75),
    .A2(_07227_),
    .A1(\cpu.spi.r_timeout_count[4] ));
 sg13g2_inv_1 _26335_ (.Y(_02616_),
    .A(_07230_));
 sg13g2_nor2_1 _26336_ (.A(\cpu.spi.r_timeout_count[4] ),
    .B(_07223_),
    .Y(_07231_));
 sg13g2_o21ai_1 _26337_ (.B1(_07211_),
    .Y(_07232_),
    .A1(net1066),
    .A2(_07231_));
 sg13g2_mux2_1 _26338_ (.A0(\cpu.spi.r_timeout[5] ),
    .A1(_09210_),
    .S(net839),
    .X(_07233_));
 sg13g2_a22oi_1 _26339_ (.Y(_07234_),
    .B1(_07233_),
    .B2(net75),
    .A2(_07232_),
    .A1(\cpu.spi.r_timeout_count[5] ));
 sg13g2_inv_1 _26340_ (.Y(_02617_),
    .A(_07234_));
 sg13g2_o21ai_1 _26341_ (.B1(_07211_),
    .Y(_07235_),
    .A1(net1031),
    .A2(_09210_));
 sg13g2_nand2_1 _26342_ (.Y(_07236_),
    .A(net1031),
    .B(\cpu.spi.r_timeout[6] ));
 sg13g2_o21ai_1 _26343_ (.B1(_07236_),
    .Y(_07237_),
    .A1(_09243_),
    .A2(_09212_));
 sg13g2_a22oi_1 _26344_ (.Y(_07238_),
    .B1(_07237_),
    .B2(net75),
    .A2(_07235_),
    .A1(\cpu.spi.r_timeout_count[6] ));
 sg13g2_inv_1 _26345_ (.Y(_02618_),
    .A(_07238_));
 sg13g2_inv_1 _26346_ (.Y(_07239_),
    .A(_09212_));
 sg13g2_o21ai_1 _26347_ (.B1(_07211_),
    .Y(_07240_),
    .A1(net1031),
    .A2(_07239_));
 sg13g2_nor3_1 _26348_ (.A(\cpu.spi.r_timeout_count[7] ),
    .B(net1031),
    .C(_09212_),
    .Y(_07241_));
 sg13g2_a21o_1 _26349_ (.A2(\cpu.spi.r_timeout[7] ),
    .A1(net1066),
    .B1(_07241_),
    .X(_07242_));
 sg13g2_a22oi_1 _26350_ (.Y(_07243_),
    .B1(_07242_),
    .B2(net75),
    .A2(_07240_),
    .A1(\cpu.spi.r_timeout_count[7] ));
 sg13g2_inv_1 _26351_ (.Y(_02619_),
    .A(_07243_));
 sg13g2_buf_1 _26352_ (.A(\cpu.uart.r_rcnt[0] ),
    .X(_07244_));
 sg13g2_nor2_1 _26353_ (.A(_07244_),
    .B(\cpu.uart.r_rcnt[1] ),
    .Y(_07245_));
 sg13g2_nand2_1 _26354_ (.Y(_07246_),
    .A(net349),
    .B(_07245_));
 sg13g2_nor2_1 _26355_ (.A(net929),
    .B(_07246_),
    .Y(_07247_));
 sg13g2_buf_2 _26356_ (.A(\cpu.uart.r_rstate[3] ),
    .X(_07248_));
 sg13g2_buf_1 _26357_ (.A(_07248_),
    .X(_07249_));
 sg13g2_buf_1 _26358_ (.A(\cpu.uart.r_rstate[1] ),
    .X(_07250_));
 sg13g2_buf_1 _26359_ (.A(\cpu.uart.r_rstate[2] ),
    .X(_07251_));
 sg13g2_buf_1 _26360_ (.A(_07251_),
    .X(_07252_));
 sg13g2_nor2_2 _26361_ (.A(net1099),
    .B(net956),
    .Y(_07253_));
 sg13g2_buf_2 _26362_ (.A(\cpu.uart.r_rstate[0] ),
    .X(_07254_));
 sg13g2_inv_1 _26363_ (.Y(_07255_),
    .A(_07254_));
 sg13g2_nand3_1 _26364_ (.B(net957),
    .C(_07253_),
    .A(_07255_),
    .Y(_07256_));
 sg13g2_o21ai_1 _26365_ (.B1(_07256_),
    .Y(_07257_),
    .A1(net957),
    .A2(_07253_));
 sg13g2_and2_1 _26366_ (.A(_07247_),
    .B(_07257_),
    .X(_07258_));
 sg13g2_buf_2 _26367_ (.A(_07258_),
    .X(_07259_));
 sg13g2_mux2_1 _26368_ (.A0(\cpu.uart.r_ib[0] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(_07259_),
    .X(_02632_));
 sg13g2_mux2_1 _26369_ (.A0(\cpu.uart.r_ib[1] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(_07259_),
    .X(_02633_));
 sg13g2_mux2_1 _26370_ (.A0(\cpu.uart.r_ib[2] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(_07259_),
    .X(_02634_));
 sg13g2_mux2_1 _26371_ (.A0(\cpu.uart.r_ib[3] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(_07259_),
    .X(_02635_));
 sg13g2_mux2_1 _26372_ (.A0(\cpu.uart.r_ib[4] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(_07259_),
    .X(_02636_));
 sg13g2_mux2_1 _26373_ (.A0(\cpu.uart.r_ib[5] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(_07259_),
    .X(_02637_));
 sg13g2_xor2_1 _26374_ (.B(\cpu.uart.r_r ),
    .A(\cpu.uart.r_r_invert ),
    .X(_07260_));
 sg13g2_mux2_1 _26375_ (.A0(\cpu.uart.r_ib[6] ),
    .A1(_07260_),
    .S(_07259_),
    .X(_02638_));
 sg13g2_and4_1 _26376_ (.A(_07254_),
    .B(_07249_),
    .C(_07247_),
    .D(_07253_),
    .X(_07261_));
 sg13g2_buf_1 _26377_ (.A(_07261_),
    .X(_07262_));
 sg13g2_mux2_1 _26378_ (.A0(\cpu.uart.r_in[0] ),
    .A1(\cpu.uart.r_ib[0] ),
    .S(net188),
    .X(_02639_));
 sg13g2_mux2_1 _26379_ (.A0(\cpu.uart.r_in[1] ),
    .A1(\cpu.uart.r_ib[1] ),
    .S(net188),
    .X(_02640_));
 sg13g2_mux2_1 _26380_ (.A0(\cpu.uart.r_in[2] ),
    .A1(\cpu.uart.r_ib[2] ),
    .S(net188),
    .X(_02641_));
 sg13g2_mux2_1 _26381_ (.A0(\cpu.uart.r_in[3] ),
    .A1(\cpu.uart.r_ib[3] ),
    .S(net188),
    .X(_02642_));
 sg13g2_mux2_1 _26382_ (.A0(\cpu.uart.r_in[4] ),
    .A1(\cpu.uart.r_ib[4] ),
    .S(net188),
    .X(_02643_));
 sg13g2_mux2_1 _26383_ (.A0(\cpu.uart.r_in[5] ),
    .A1(\cpu.uart.r_ib[5] ),
    .S(net188),
    .X(_02644_));
 sg13g2_mux2_1 _26384_ (.A0(\cpu.uart.r_in[6] ),
    .A1(\cpu.uart.r_ib[6] ),
    .S(net188),
    .X(_02645_));
 sg13g2_mux2_1 _26385_ (.A0(\cpu.uart.r_in[7] ),
    .A1(_07260_),
    .S(_07262_),
    .X(_02646_));
 sg13g2_nor2_1 _26386_ (.A(_09165_),
    .B(net1154),
    .Y(_07263_));
 sg13g2_and3_1 _26387_ (.X(_07264_),
    .A(net899),
    .B(_07263_),
    .C(_06305_));
 sg13g2_buf_1 _26388_ (.A(_07264_),
    .X(_07265_));
 sg13g2_buf_1 _26389_ (.A(\cpu.uart.r_xstate[2] ),
    .X(_07266_));
 sg13g2_a21oi_1 _26390_ (.A1(net517),
    .A2(_07265_),
    .Y(_07267_),
    .B1(net1098));
 sg13g2_nand3_1 _26391_ (.B(_07263_),
    .C(_06305_),
    .A(net899),
    .Y(_07268_));
 sg13g2_buf_1 _26392_ (.A(_07268_),
    .X(_07269_));
 sg13g2_buf_1 _26393_ (.A(\cpu.uart.r_xstate[3] ),
    .X(_07270_));
 sg13g2_buf_1 _26394_ (.A(\cpu.uart.r_xstate[1] ),
    .X(_07271_));
 sg13g2_buf_1 _26395_ (.A(_07271_),
    .X(_07272_));
 sg13g2_buf_1 _26396_ (.A(\cpu.uart.r_xstate[0] ),
    .X(_07273_));
 sg13g2_nor2_1 _26397_ (.A(net955),
    .B(_07273_),
    .Y(_07274_));
 sg13g2_nand2b_1 _26398_ (.Y(_07275_),
    .B(_07274_),
    .A_N(net1097));
 sg13g2_and2_1 _26399_ (.A(_07271_),
    .B(_07273_),
    .X(_07276_));
 sg13g2_buf_1 _26400_ (.A(_07276_),
    .X(_07277_));
 sg13g2_nand2_2 _26401_ (.Y(_07278_),
    .A(net1097),
    .B(_07277_));
 sg13g2_o21ai_1 _26402_ (.B1(_07278_),
    .Y(_07279_),
    .A1(_07269_),
    .A2(_07275_));
 sg13g2_buf_1 _26403_ (.A(\cpu.uart.r_xcnt[0] ),
    .X(_07280_));
 sg13g2_nor2_1 _26404_ (.A(_07280_),
    .B(\cpu.uart.r_xcnt[1] ),
    .Y(_07281_));
 sg13g2_nand2_1 _26405_ (.Y(_07282_),
    .A(_09857_),
    .B(_07281_));
 sg13g2_buf_1 _26406_ (.A(_07282_),
    .X(_07283_));
 sg13g2_a21o_1 _26407_ (.A2(_07283_),
    .A1(net1097),
    .B1(net955),
    .X(_07284_));
 sg13g2_a21oi_1 _26408_ (.A1(_07278_),
    .A2(_07284_),
    .Y(_07285_),
    .B1(net1098));
 sg13g2_nor2_1 _26409_ (.A(net1097),
    .B(_07283_),
    .Y(_07286_));
 sg13g2_buf_1 _26410_ (.A(_07273_),
    .X(_07287_));
 sg13g2_nor3_1 _26411_ (.A(net955),
    .B(net1097),
    .C(net1098),
    .Y(_07288_));
 sg13g2_o21ai_1 _26412_ (.B1(_07288_),
    .Y(_07289_),
    .A1(net954),
    .A2(_07269_));
 sg13g2_o21ai_1 _26413_ (.B1(_07289_),
    .Y(_07290_),
    .A1(_07285_),
    .A2(_07286_));
 sg13g2_or2_1 _26414_ (.X(_07291_),
    .B(_07290_),
    .A(net929));
 sg13g2_a21o_1 _26415_ (.A2(_07279_),
    .A1(_07267_),
    .B1(_07291_),
    .X(_07292_));
 sg13g2_buf_2 _26416_ (.A(_07292_),
    .X(_07293_));
 sg13g2_buf_1 _26417_ (.A(_07293_),
    .X(_07294_));
 sg13g2_buf_1 _26418_ (.A(net1098),
    .X(_07295_));
 sg13g2_nor2_1 _26419_ (.A(net955),
    .B(net953),
    .Y(_07296_));
 sg13g2_xnor2_1 _26420_ (.Y(_07297_),
    .A(net1097),
    .B(_07296_));
 sg13g2_buf_1 _26421_ (.A(_07297_),
    .X(_07298_));
 sg13g2_buf_1 _26422_ (.A(_07298_),
    .X(_07299_));
 sg13g2_nor2_1 _26423_ (.A(_09969_),
    .B(net591),
    .Y(_07300_));
 sg13g2_a21oi_1 _26424_ (.A1(\cpu.uart.r_out[1] ),
    .A2(net591),
    .Y(_07301_),
    .B1(_07300_));
 sg13g2_buf_1 _26425_ (.A(\cpu.uart.r_out[0] ),
    .X(_07302_));
 sg13g2_nand2_1 _26426_ (.Y(_07303_),
    .A(_07302_),
    .B(net66));
 sg13g2_o21ai_1 _26427_ (.B1(_07303_),
    .Y(_02647_),
    .A1(net66),
    .A2(_07301_));
 sg13g2_nor2_1 _26428_ (.A(net897),
    .B(_07299_),
    .Y(_07304_));
 sg13g2_a21oi_1 _26429_ (.A1(\cpu.uart.r_out[2] ),
    .A2(_07299_),
    .Y(_07305_),
    .B1(_07304_));
 sg13g2_nand2_1 _26430_ (.Y(_07306_),
    .A(\cpu.uart.r_out[1] ),
    .B(net66));
 sg13g2_o21ai_1 _26431_ (.B1(_07306_),
    .Y(_02648_),
    .A1(_07294_),
    .A2(_07305_));
 sg13g2_nor2_1 _26432_ (.A(_12175_),
    .B(_07298_),
    .Y(_07307_));
 sg13g2_a21oi_1 _26433_ (.A1(\cpu.uart.r_out[3] ),
    .A2(net591),
    .Y(_07308_),
    .B1(_07307_));
 sg13g2_nand2_1 _26434_ (.Y(_07309_),
    .A(\cpu.uart.r_out[2] ),
    .B(_07293_));
 sg13g2_o21ai_1 _26435_ (.B1(_07309_),
    .Y(_02649_),
    .A1(_07294_),
    .A2(_07308_));
 sg13g2_nor2b_1 _26436_ (.A(_07298_),
    .B_N(net1144),
    .Y(_07310_));
 sg13g2_a21oi_1 _26437_ (.A1(\cpu.uart.r_out[4] ),
    .A2(net591),
    .Y(_07311_),
    .B1(_07310_));
 sg13g2_nand2_1 _26438_ (.Y(_07312_),
    .A(\cpu.uart.r_out[3] ),
    .B(_07293_));
 sg13g2_o21ai_1 _26439_ (.B1(_07312_),
    .Y(_02650_),
    .A1(net66),
    .A2(_07311_));
 sg13g2_nor2b_1 _26440_ (.A(_07298_),
    .B_N(_09999_),
    .Y(_07313_));
 sg13g2_a21oi_1 _26441_ (.A1(\cpu.uart.r_out[5] ),
    .A2(net591),
    .Y(_07314_),
    .B1(_07313_));
 sg13g2_nand2_1 _26442_ (.Y(_07315_),
    .A(\cpu.uart.r_out[4] ),
    .B(_07293_));
 sg13g2_o21ai_1 _26443_ (.B1(_07315_),
    .Y(_02651_),
    .A1(net66),
    .A2(_07314_));
 sg13g2_nor2_1 _26444_ (.A(_12202_),
    .B(_07298_),
    .Y(_07316_));
 sg13g2_a21oi_1 _26445_ (.A1(\cpu.uart.r_out[6] ),
    .A2(net591),
    .Y(_07317_),
    .B1(_07316_));
 sg13g2_nand2_1 _26446_ (.Y(_07318_),
    .A(\cpu.uart.r_out[5] ),
    .B(_07293_));
 sg13g2_o21ai_1 _26447_ (.B1(_07318_),
    .Y(_02652_),
    .A1(net66),
    .A2(_07317_));
 sg13g2_nor2_1 _26448_ (.A(_12210_),
    .B(_07298_),
    .Y(_07319_));
 sg13g2_a21oi_1 _26449_ (.A1(\cpu.uart.r_out[7] ),
    .A2(net591),
    .Y(_07320_),
    .B1(_07319_));
 sg13g2_nand2_1 _26450_ (.Y(_07321_),
    .A(\cpu.uart.r_out[6] ),
    .B(_07293_));
 sg13g2_o21ai_1 _26451_ (.B1(_07321_),
    .Y(_02653_),
    .A1(net66),
    .A2(_07320_));
 sg13g2_nor3_1 _26452_ (.A(_07194_),
    .B(_07293_),
    .C(net591),
    .Y(_07322_));
 sg13g2_a21o_1 _26453_ (.A2(net66),
    .A1(\cpu.uart.r_out[7] ),
    .B1(_07322_),
    .X(_02654_));
 sg13g2_nand2_1 _26454_ (.Y(_07323_),
    .A(net1099),
    .B(_07248_));
 sg13g2_inv_1 _26455_ (.Y(_07324_),
    .A(_07323_));
 sg13g2_nor4_1 _26456_ (.A(net1099),
    .B(_07251_),
    .C(_07248_),
    .D(_09857_),
    .Y(_07325_));
 sg13g2_o21ai_1 _26457_ (.B1(_07254_),
    .Y(_07326_),
    .A1(_07324_),
    .A2(_07325_));
 sg13g2_nor4_1 _26458_ (.A(_07254_),
    .B(_07250_),
    .C(_07251_),
    .D(_07248_),
    .Y(_07327_));
 sg13g2_nand2b_1 _26459_ (.Y(_07328_),
    .B(_09885_),
    .A_N(_09847_));
 sg13g2_a21o_1 _26460_ (.A2(_07328_),
    .A1(net1099),
    .B1(_07251_),
    .X(_07329_));
 sg13g2_a22oi_1 _26461_ (.Y(_07330_),
    .B1(_07329_),
    .B2(_07248_),
    .A2(_07327_),
    .A1(_07260_));
 sg13g2_nand2_1 _26462_ (.Y(_07331_),
    .A(_07326_),
    .B(_07330_));
 sg13g2_nor2b_1 _26463_ (.A(_07248_),
    .B_N(_07260_),
    .Y(_07332_));
 sg13g2_nor2_1 _26464_ (.A(_07255_),
    .B(net1099),
    .Y(_07333_));
 sg13g2_a22oi_1 _26465_ (.Y(_07334_),
    .B1(_07332_),
    .B2(_07333_),
    .A2(_07324_),
    .A1(_07255_));
 sg13g2_nor3_1 _26466_ (.A(net956),
    .B(_07246_),
    .C(_07334_),
    .Y(_07335_));
 sg13g2_xor2_1 _26467_ (.B(_07253_),
    .A(_07249_),
    .X(_07336_));
 sg13g2_o21ai_1 _26468_ (.B1(net1071),
    .Y(_07337_),
    .A1(net349),
    .A2(_07336_));
 sg13g2_nor3_2 _26469_ (.A(_07331_),
    .B(_07335_),
    .C(_07337_),
    .Y(_07338_));
 sg13g2_and2_1 _26470_ (.A(_07254_),
    .B(net1099),
    .X(_07339_));
 sg13g2_buf_1 _26471_ (.A(_07339_),
    .X(_07340_));
 sg13g2_o21ai_1 _26472_ (.B1(net957),
    .Y(_07341_),
    .A1(net956),
    .A2(_07340_));
 sg13g2_nor2b_1 _26473_ (.A(_07327_),
    .B_N(_07341_),
    .Y(_07342_));
 sg13g2_nand3_1 _26474_ (.B(_07338_),
    .C(_07342_),
    .A(_07244_),
    .Y(_07343_));
 sg13g2_o21ai_1 _26475_ (.B1(_07343_),
    .Y(_07344_),
    .A1(_07244_),
    .A2(_07338_));
 sg13g2_inv_1 _26476_ (.Y(_02657_),
    .A(_07344_));
 sg13g2_nand2_1 _26477_ (.Y(_07345_),
    .A(_07244_),
    .B(_07342_));
 sg13g2_nand2_1 _26478_ (.Y(_07346_),
    .A(_07338_),
    .B(_07345_));
 sg13g2_nand2_1 _26479_ (.Y(_07347_),
    .A(\cpu.uart.r_rcnt[1] ),
    .B(_07346_));
 sg13g2_nand3_1 _26480_ (.B(_07338_),
    .C(_07342_),
    .A(_07245_),
    .Y(_07348_));
 sg13g2_nand2_1 _26481_ (.Y(_02658_),
    .A(_07347_),
    .B(_07348_));
 sg13g2_buf_1 _26482_ (.A(\cpu.gpio.genblk1[3].srcs_o[1] ),
    .X(_07349_));
 sg13g2_buf_1 _26483_ (.A(_07270_),
    .X(_07350_));
 sg13g2_a21oi_1 _26484_ (.A1(net952),
    .A2(_04969_),
    .Y(_07351_),
    .B1(net953));
 sg13g2_nor2b_1 _26485_ (.A(_07302_),
    .B_N(_04969_),
    .Y(_07352_));
 sg13g2_a21oi_1 _26486_ (.A1(_07302_),
    .A2(_07351_),
    .Y(_07353_),
    .B1(_07352_));
 sg13g2_nor2_1 _26487_ (.A(net955),
    .B(_07353_),
    .Y(_07354_));
 sg13g2_xnor2_1 _26488_ (.Y(_07355_),
    .A(_07302_),
    .B(_04969_));
 sg13g2_nand3_1 _26489_ (.B(_07295_),
    .C(_04969_),
    .A(net952),
    .Y(_07356_));
 sg13g2_o21ai_1 _26490_ (.B1(_07356_),
    .Y(_07357_),
    .A1(_07350_),
    .A2(_07355_));
 sg13g2_inv_1 _26491_ (.Y(_07358_),
    .A(_07271_));
 sg13g2_or2_1 _26492_ (.X(_07359_),
    .B(net1098),
    .A(\cpu.uart.r_xstate[3] ));
 sg13g2_buf_1 _26493_ (.A(_07359_),
    .X(_07360_));
 sg13g2_nand2_2 _26494_ (.Y(_07361_),
    .A(_07270_),
    .B(net1098));
 sg13g2_a21o_1 _26495_ (.A2(_07361_),
    .A1(_07360_),
    .B1(_07273_),
    .X(_07362_));
 sg13g2_buf_1 _26496_ (.A(_07362_),
    .X(_07363_));
 sg13g2_o21ai_1 _26497_ (.B1(_07363_),
    .Y(_07364_),
    .A1(_04969_),
    .A2(_07360_));
 sg13g2_a21oi_1 _26498_ (.A1(_07358_),
    .A2(_07364_),
    .Y(_07365_),
    .B1(net929));
 sg13g2_o21ai_1 _26499_ (.B1(_07365_),
    .Y(_07366_),
    .A1(_07354_),
    .A2(_07357_));
 sg13g2_nor2b_1 _26500_ (.A(net1098),
    .B_N(net1097),
    .Y(_07367_));
 sg13g2_nor2_1 _26501_ (.A(_07358_),
    .B(_07367_),
    .Y(_07368_));
 sg13g2_a21oi_1 _26502_ (.A1(_07358_),
    .A2(_07363_),
    .Y(_07369_),
    .B1(_07368_));
 sg13g2_o21ai_1 _26503_ (.B1(_00273_),
    .Y(_07370_),
    .A1(net815),
    .A2(_07369_));
 sg13g2_nand2_1 _26504_ (.Y(_07371_),
    .A(_07366_),
    .B(_07370_));
 sg13g2_and4_1 _26505_ (.A(net517),
    .B(_07265_),
    .C(_07277_),
    .D(_07367_),
    .X(_07372_));
 sg13g2_buf_1 _26506_ (.A(_07372_),
    .X(_07373_));
 sg13g2_o21ai_1 _26507_ (.B1(_07363_),
    .Y(_07374_),
    .A1(_07328_),
    .A2(_07360_));
 sg13g2_and2_1 _26508_ (.A(_07358_),
    .B(_07374_),
    .X(_07375_));
 sg13g2_a21oi_1 _26509_ (.A1(_07278_),
    .A2(_07283_),
    .Y(_07376_),
    .B1(net1098));
 sg13g2_nor3_1 _26510_ (.A(_07286_),
    .B(_07375_),
    .C(_07376_),
    .Y(_07377_));
 sg13g2_o21ai_1 _26511_ (.B1(net933),
    .Y(_07378_),
    .A1(_07373_),
    .A2(_07377_));
 sg13g2_mux2_1 _26512_ (.A0(net1096),
    .A1(_07371_),
    .S(_07378_),
    .X(_02663_));
 sg13g2_o21ai_1 _26513_ (.B1(net349),
    .Y(_07379_),
    .A1(net954),
    .A2(net952));
 sg13g2_o21ai_1 _26514_ (.B1(_07361_),
    .Y(_07380_),
    .A1(net954),
    .A2(net349));
 sg13g2_and2_1 _26515_ (.A(net1097),
    .B(_07266_),
    .X(_07381_));
 sg13g2_buf_1 _26516_ (.A(_07381_),
    .X(_07382_));
 sg13g2_a21oi_1 _26517_ (.A1(net954),
    .A2(_07382_),
    .Y(_07383_),
    .B1(net929));
 sg13g2_o21ai_1 _26518_ (.B1(_07383_),
    .Y(_07384_),
    .A1(net952),
    .A2(_09858_));
 sg13g2_a221oi_1 _26519_ (.B2(net955),
    .C1(_07384_),
    .B1(_07380_),
    .A1(_07296_),
    .Y(_07385_),
    .A2(_07379_));
 sg13g2_nand2b_1 _26520_ (.Y(_07386_),
    .B(_09858_),
    .A_N(_07281_));
 sg13g2_nand2_1 _26521_ (.Y(_07387_),
    .A(net955),
    .B(net954));
 sg13g2_nor2_1 _26522_ (.A(net953),
    .B(_07387_),
    .Y(_07388_));
 sg13g2_a21oi_1 _26523_ (.A1(net953),
    .A2(_07274_),
    .Y(_07389_),
    .B1(_07388_));
 sg13g2_nor2b_1 _26524_ (.A(_07389_),
    .B_N(net952),
    .Y(_07390_));
 sg13g2_o21ai_1 _26525_ (.B1(_07390_),
    .Y(_07391_),
    .A1(_07373_),
    .A2(_07386_));
 sg13g2_nand2_1 _26526_ (.Y(_07392_),
    .A(_07385_),
    .B(_07391_));
 sg13g2_nor2_1 _26527_ (.A(_07274_),
    .B(_07361_),
    .Y(_07393_));
 sg13g2_nor2_1 _26528_ (.A(_07288_),
    .B(_07393_),
    .Y(_07394_));
 sg13g2_nand3_1 _26529_ (.B(_07391_),
    .C(_07394_),
    .A(_07385_),
    .Y(_07395_));
 sg13g2_nand2_1 _26530_ (.Y(_07396_),
    .A(_07280_),
    .B(_07395_));
 sg13g2_o21ai_1 _26531_ (.B1(_07396_),
    .Y(_02666_),
    .A1(_07280_),
    .A2(_07392_));
 sg13g2_a21o_1 _26532_ (.A2(_07394_),
    .A1(_07280_),
    .B1(_07392_),
    .X(_07397_));
 sg13g2_o21ai_1 _26533_ (.B1(\cpu.uart.r_xcnt[1] ),
    .Y(_07398_),
    .A1(_07280_),
    .A2(_07395_));
 sg13g2_o21ai_1 _26534_ (.B1(_07398_),
    .Y(_02667_),
    .A1(\cpu.uart.r_xcnt[1] ),
    .A2(_07397_));
 sg13g2_nor2_1 _26535_ (.A(net694),
    .B(_10023_),
    .Y(_07399_));
 sg13g2_buf_2 _26536_ (.A(_07399_),
    .X(_07400_));
 sg13g2_buf_1 _26537_ (.A(_07400_),
    .X(_07401_));
 sg13g2_or2_1 _26538_ (.X(_07402_),
    .B(_10111_),
    .A(_10118_));
 sg13g2_or2_1 _26539_ (.X(_07403_),
    .B(_07402_),
    .A(_10077_));
 sg13g2_nor2_1 _26540_ (.A(_10117_),
    .B(_07403_),
    .Y(_07404_));
 sg13g2_and2_1 _26541_ (.A(_04919_),
    .B(_07404_),
    .X(_07405_));
 sg13g2_buf_1 _26542_ (.A(_07405_),
    .X(_07406_));
 sg13g2_nor2_1 _26543_ (.A(net636),
    .B(_10023_),
    .Y(_07407_));
 sg13g2_buf_1 _26544_ (.A(_07407_),
    .X(_07408_));
 sg13g2_buf_1 _26545_ (.A(_07408_),
    .X(_07409_));
 sg13g2_nor2_1 _26546_ (.A(_10033_),
    .B(_07404_),
    .Y(_07410_));
 sg13g2_nor2_1 _26547_ (.A(net83),
    .B(_07410_),
    .Y(_07411_));
 sg13g2_nor2_1 _26548_ (.A(_04919_),
    .B(_07411_),
    .Y(_07412_));
 sg13g2_a221oi_1 _26549_ (.B2(net153),
    .C1(_07412_),
    .B1(_07406_),
    .A1(_09970_),
    .Y(_02453_),
    .A2(net84));
 sg13g2_nor2_1 _26550_ (.A(_10033_),
    .B(_07406_),
    .Y(_07413_));
 sg13g2_or2_1 _26551_ (.X(_07414_),
    .B(_07413_),
    .A(net83));
 sg13g2_inv_1 _26552_ (.Y(_07415_),
    .A(_05359_));
 sg13g2_nand2_1 _26553_ (.Y(_07416_),
    .A(_05359_),
    .B(_07406_));
 sg13g2_nor2_1 _26554_ (.A(net183),
    .B(_07416_),
    .Y(_07417_));
 sg13g2_a221oi_1 _26555_ (.B2(_07415_),
    .C1(_07417_),
    .B1(_07414_),
    .A1(_12236_),
    .Y(_02454_),
    .A2(net84));
 sg13g2_a21oi_1 _26556_ (.A1(net153),
    .A2(_07416_),
    .Y(_07418_),
    .B1(_07408_));
 sg13g2_nor2_1 _26557_ (.A(_05408_),
    .B(_07418_),
    .Y(_07419_));
 sg13g2_a221oi_1 _26558_ (.B2(_05408_),
    .C1(_07419_),
    .B1(_07417_),
    .A1(net896),
    .Y(_02455_),
    .A2(net84));
 sg13g2_inv_1 _26559_ (.Y(_07420_),
    .A(_05495_));
 sg13g2_nand4_1 _26560_ (.B(_04919_),
    .C(_05359_),
    .A(_10116_),
    .Y(_07421_),
    .D(_05408_));
 sg13g2_or2_1 _26561_ (.X(_07422_),
    .B(_07421_),
    .A(_10120_));
 sg13g2_a21oi_1 _26562_ (.A1(net153),
    .A2(_07422_),
    .Y(_07423_),
    .B1(net83));
 sg13g2_nor2_1 _26563_ (.A(net183),
    .B(_07422_),
    .Y(_07424_));
 sg13g2_a22oi_1 _26564_ (.Y(_07425_),
    .B1(_07424_),
    .B2(_07420_),
    .A2(_07400_),
    .A1(net1058));
 sg13g2_o21ai_1 _26565_ (.B1(_07425_),
    .Y(_02456_),
    .A1(_07420_),
    .A2(_07423_));
 sg13g2_nor2_1 _26566_ (.A(_07403_),
    .B(_07421_),
    .Y(_07426_));
 sg13g2_buf_1 _26567_ (.A(_07426_),
    .X(_07427_));
 sg13g2_a21oi_1 _26568_ (.A1(_05495_),
    .A2(_07427_),
    .Y(_07428_),
    .B1(net183));
 sg13g2_o21ai_1 _26569_ (.B1(_05542_),
    .Y(_07429_),
    .A1(net83),
    .A2(_07428_));
 sg13g2_and2_1 _26570_ (.A(_10023_),
    .B(_07427_),
    .X(_07430_));
 sg13g2_buf_1 _26571_ (.A(_07430_),
    .X(_07431_));
 sg13g2_nor2_1 _26572_ (.A(_07420_),
    .B(_05542_),
    .Y(_07432_));
 sg13g2_a22oi_1 _26573_ (.Y(_07433_),
    .B1(_07431_),
    .B2(_07432_),
    .A2(net84),
    .A1(net1057));
 sg13g2_nand2_1 _26574_ (.Y(_02457_),
    .A(_07429_),
    .B(_07433_));
 sg13g2_and3_1 _26575_ (.X(_07434_),
    .A(_05495_),
    .B(_05542_),
    .C(_05636_));
 sg13g2_buf_1 _26576_ (.A(_07434_),
    .X(_07435_));
 sg13g2_nor2_1 _26577_ (.A(_10120_),
    .B(_07421_),
    .Y(_07436_));
 sg13g2_nand3_1 _26578_ (.B(_05542_),
    .C(_07436_),
    .A(_05495_),
    .Y(_07437_));
 sg13g2_a21oi_1 _26579_ (.A1(net153),
    .A2(_07437_),
    .Y(_07438_),
    .B1(_07408_));
 sg13g2_nor2_1 _26580_ (.A(_05636_),
    .B(_07438_),
    .Y(_07439_));
 sg13g2_a221oi_1 _26581_ (.B2(_07435_),
    .C1(_07439_),
    .B1(_07424_),
    .A1(net895),
    .Y(_02458_),
    .A2(net84));
 sg13g2_and2_1 _26582_ (.A(_05659_),
    .B(_07435_),
    .X(_07440_));
 sg13g2_buf_1 _26583_ (.A(_07440_),
    .X(_07441_));
 sg13g2_a21oi_1 _26584_ (.A1(_07427_),
    .A2(_07435_),
    .Y(_07442_),
    .B1(_10033_));
 sg13g2_nor2_1 _26585_ (.A(net83),
    .B(_07442_),
    .Y(_07443_));
 sg13g2_nor2_1 _26586_ (.A(_05659_),
    .B(_07443_),
    .Y(_07444_));
 sg13g2_a221oi_1 _26587_ (.B2(_07441_),
    .C1(_07444_),
    .B1(_07431_),
    .A1(net894),
    .Y(_02459_),
    .A2(net84));
 sg13g2_and2_1 _26588_ (.A(_05067_),
    .B(_07441_),
    .X(_07445_));
 sg13g2_buf_1 _26589_ (.A(_07445_),
    .X(_07446_));
 sg13g2_a21oi_1 _26590_ (.A1(_07436_),
    .A2(_07441_),
    .Y(_07447_),
    .B1(_10033_));
 sg13g2_nor2_1 _26591_ (.A(_07408_),
    .B(_07447_),
    .Y(_07448_));
 sg13g2_nor2_1 _26592_ (.A(_05067_),
    .B(_07448_),
    .Y(_07449_));
 sg13g2_a221oi_1 _26593_ (.B2(_07446_),
    .C1(_07449_),
    .B1(_07424_),
    .A1(_12269_),
    .Y(_02460_),
    .A2(net84));
 sg13g2_a21oi_1 _26594_ (.A1(_07427_),
    .A2(_07446_),
    .Y(_07450_),
    .B1(_10034_));
 sg13g2_o21ai_1 _26595_ (.B1(_05727_),
    .Y(_07451_),
    .A1(_07409_),
    .A2(_07450_));
 sg13g2_nor2b_1 _26596_ (.A(_05727_),
    .B_N(_07446_),
    .Y(_07452_));
 sg13g2_a22oi_1 _26597_ (.Y(_07453_),
    .B1(_07431_),
    .B2(_07452_),
    .A2(_07400_),
    .A1(_10081_));
 sg13g2_nand2_1 _26598_ (.Y(_02461_),
    .A(_07451_),
    .B(_07453_));
 sg13g2_inv_1 _26599_ (.Y(_07454_),
    .A(_05740_));
 sg13g2_nand3_1 _26600_ (.B(_07427_),
    .C(_07446_),
    .A(_05727_),
    .Y(_07455_));
 sg13g2_a21oi_1 _26601_ (.A1(_10024_),
    .A2(_07455_),
    .Y(_07456_),
    .B1(net83));
 sg13g2_nor2_2 _26602_ (.A(_10033_),
    .B(_07455_),
    .Y(_07457_));
 sg13g2_a22oi_1 _26603_ (.Y(_07458_),
    .B1(_07457_),
    .B2(_07454_),
    .A2(_07400_),
    .A1(_10086_));
 sg13g2_o21ai_1 _26604_ (.B1(_07458_),
    .Y(_02462_),
    .A1(_07454_),
    .A2(_07456_));
 sg13g2_and3_1 _26605_ (.X(_07459_),
    .A(_05727_),
    .B(_07427_),
    .C(_07446_));
 sg13g2_buf_1 _26606_ (.A(_07459_),
    .X(_07460_));
 sg13g2_a21oi_1 _26607_ (.A1(_05740_),
    .A2(_07460_),
    .Y(_07461_),
    .B1(net183));
 sg13g2_o21ai_1 _26608_ (.B1(_05142_),
    .Y(_07462_),
    .A1(net83),
    .A2(_07461_));
 sg13g2_nor2_1 _26609_ (.A(_07454_),
    .B(_05142_),
    .Y(_07463_));
 sg13g2_a22oi_1 _26610_ (.Y(_07464_),
    .B1(_07457_),
    .B2(_07463_),
    .A2(_07400_),
    .A1(_10091_));
 sg13g2_nand2_1 _26611_ (.Y(_02463_),
    .A(_07462_),
    .B(_07464_));
 sg13g2_and3_1 _26612_ (.X(_07465_),
    .A(_05727_),
    .B(_07436_),
    .C(_07446_));
 sg13g2_buf_1 _26613_ (.A(_07465_),
    .X(_07466_));
 sg13g2_and4_1 _26614_ (.A(_05740_),
    .B(_05142_),
    .C(_05165_),
    .D(_07466_),
    .X(_07467_));
 sg13g2_nand3_1 _26615_ (.B(_05142_),
    .C(_07466_),
    .A(_05740_),
    .Y(_07468_));
 sg13g2_a21oi_1 _26616_ (.A1(net153),
    .A2(_07468_),
    .Y(_07469_),
    .B1(_07408_));
 sg13g2_nor2_1 _26617_ (.A(_05165_),
    .B(_07469_),
    .Y(_07470_));
 sg13g2_a221oi_1 _26618_ (.B2(net153),
    .C1(_07470_),
    .B1(_07467_),
    .A1(_05761_),
    .Y(_02464_),
    .A2(net84));
 sg13g2_and4_1 _26619_ (.A(_05740_),
    .B(_05142_),
    .C(_05165_),
    .D(_05208_),
    .X(_07471_));
 sg13g2_buf_1 _26620_ (.A(_07471_),
    .X(_07472_));
 sg13g2_nand4_1 _26621_ (.B(_05142_),
    .C(_05165_),
    .A(_05740_),
    .Y(_07473_),
    .D(_07460_));
 sg13g2_a21oi_1 _26622_ (.A1(_10023_),
    .A2(_07473_),
    .Y(_07474_),
    .B1(_07408_));
 sg13g2_nor2_1 _26623_ (.A(_05208_),
    .B(_07474_),
    .Y(_07475_));
 sg13g2_a221oi_1 _26624_ (.B2(_07472_),
    .C1(_07475_),
    .B1(_07457_),
    .A1(_12192_),
    .Y(_02465_),
    .A2(_07401_));
 sg13g2_nand2_1 _26625_ (.Y(_07476_),
    .A(_07466_),
    .B(_07472_));
 sg13g2_a21oi_1 _26626_ (.A1(_10024_),
    .A2(_07476_),
    .Y(_07477_),
    .B1(net83));
 sg13g2_nand2b_1 _26627_ (.Y(_07478_),
    .B(_07477_),
    .A_N(_05222_));
 sg13g2_o21ai_1 _26628_ (.B1(_05222_),
    .Y(_07479_),
    .A1(net183),
    .A2(_07476_));
 sg13g2_a22oi_1 _26629_ (.Y(_02466_),
    .B1(_07478_),
    .B2(_07479_),
    .A2(_07401_),
    .A1(_12203_));
 sg13g2_and2_1 _26630_ (.A(_05222_),
    .B(_07472_),
    .X(_07480_));
 sg13g2_buf_1 _26631_ (.A(_07480_),
    .X(_07481_));
 sg13g2_a21oi_1 _26632_ (.A1(_07460_),
    .A2(_07481_),
    .Y(_07482_),
    .B1(_10034_));
 sg13g2_o21ai_1 _26633_ (.B1(_05272_),
    .Y(_07483_),
    .A1(_07409_),
    .A2(_07482_));
 sg13g2_nor2b_1 _26634_ (.A(_05272_),
    .B_N(_07481_),
    .Y(_07484_));
 sg13g2_a22oi_1 _26635_ (.Y(_07485_),
    .B1(_07457_),
    .B2(_07484_),
    .A2(_07400_),
    .A1(_10114_));
 sg13g2_nand2_1 _26636_ (.Y(_02467_),
    .A(_07483_),
    .B(_07485_));
 sg13g2_nand3_1 _26637_ (.B(_07466_),
    .C(_07481_),
    .A(_05272_),
    .Y(_07486_));
 sg13g2_a21o_1 _26638_ (.A2(_07486_),
    .A1(_10023_),
    .B1(_07408_),
    .X(_07487_));
 sg13g2_nor3_1 _26639_ (.A(_05282_),
    .B(net183),
    .C(_07486_),
    .Y(_07488_));
 sg13g2_a221oi_1 _26640_ (.B2(_05282_),
    .C1(_07488_),
    .B1(_07487_),
    .A1(_10122_),
    .Y(_07489_),
    .A2(_07400_));
 sg13g2_inv_1 _26641_ (.Y(_02468_),
    .A(_07489_));
 sg13g2_nor2_1 _26642_ (.A(\cpu.r_clk_invert ),
    .B(net714),
    .Y(_07490_));
 sg13g2_a21oi_1 _26643_ (.A1(_09139_),
    .A2(net714),
    .Y(_02535_),
    .B1(_07490_));
 sg13g2_nand2b_1 _26644_ (.Y(_07491_),
    .B(_09105_),
    .A_N(\cpu.d_flush_all ));
 sg13g2_buf_2 _26645_ (.A(_07491_),
    .X(_07492_));
 sg13g2_nor2b_1 _26646_ (.A(\cpu.dcache.r_valid[0] ),
    .B_N(net432),
    .Y(_07493_));
 sg13g2_nand4_1 _26647_ (.B(_03012_),
    .C(_12296_),
    .A(_09303_),
    .Y(_07494_),
    .D(_12129_));
 sg13g2_buf_2 _26648_ (.A(_07494_),
    .X(_07495_));
 sg13g2_nor2_1 _26649_ (.A(net625),
    .B(_07495_),
    .Y(_07496_));
 sg13g2_nor3_1 _26650_ (.A(_07492_),
    .B(_07493_),
    .C(_07496_),
    .Y(_00732_));
 sg13g2_nor2_1 _26651_ (.A(\cpu.dcache.r_valid[1] ),
    .B(net476),
    .Y(_07497_));
 sg13g2_nor2_1 _26652_ (.A(_12339_),
    .B(_07495_),
    .Y(_07498_));
 sg13g2_nor3_1 _26653_ (.A(_07492_),
    .B(_07497_),
    .C(_07498_),
    .Y(_00733_));
 sg13g2_nor2_1 _26654_ (.A(\cpu.dcache.r_valid[2] ),
    .B(_12518_),
    .Y(_07499_));
 sg13g2_nor2_1 _26655_ (.A(_12457_),
    .B(_07495_),
    .Y(_07500_));
 sg13g2_nor3_1 _26656_ (.A(_07492_),
    .B(_07499_),
    .C(_07500_),
    .Y(_00734_));
 sg13g2_nor2_1 _26657_ (.A(\cpu.dcache.r_valid[3] ),
    .B(net343),
    .Y(_07501_));
 sg13g2_nor2_1 _26658_ (.A(_12566_),
    .B(_07495_),
    .Y(_07502_));
 sg13g2_nor3_1 _26659_ (.A(_07492_),
    .B(_07501_),
    .C(_07502_),
    .Y(_00735_));
 sg13g2_a21oi_1 _26660_ (.A1(_10019_),
    .A2(_12274_),
    .Y(_07503_),
    .B1(\cpu.dcache.r_valid[4] ));
 sg13g2_nor2_1 _26661_ (.A(net484),
    .B(_07495_),
    .Y(_07504_));
 sg13g2_nor3_1 _26662_ (.A(_07492_),
    .B(_07503_),
    .C(_07504_),
    .Y(_00736_));
 sg13g2_nor2_1 _26663_ (.A(\cpu.dcache.r_valid[5] ),
    .B(net550),
    .Y(_07505_));
 sg13g2_nor2_1 _26664_ (.A(net760),
    .B(_07495_),
    .Y(_07506_));
 sg13g2_nor3_1 _26665_ (.A(_07492_),
    .B(_07505_),
    .C(_07506_),
    .Y(_00737_));
 sg13g2_nor2_1 _26666_ (.A(\cpu.dcache.r_valid[6] ),
    .B(_02861_),
    .Y(_07507_));
 sg13g2_nor2_1 _26667_ (.A(net756),
    .B(_07495_),
    .Y(_07508_));
 sg13g2_nor3_1 _26668_ (.A(_07492_),
    .B(_07507_),
    .C(_07508_),
    .Y(_00738_));
 sg13g2_nor2_1 _26669_ (.A(\cpu.dcache.r_valid[7] ),
    .B(net295),
    .Y(_07509_));
 sg13g2_nor2_1 _26670_ (.A(net381),
    .B(_07495_),
    .Y(_07510_));
 sg13g2_nor3_1 _26671_ (.A(_07492_),
    .B(_07509_),
    .C(_07510_),
    .Y(_00739_));
 sg13g2_nand3_1 _26672_ (.B(_10146_),
    .C(_04769_),
    .A(_11431_),
    .Y(_07511_));
 sg13g2_buf_1 _26673_ (.A(_07511_),
    .X(_07512_));
 sg13g2_nand2_1 _26674_ (.Y(_07513_),
    .A(_08274_),
    .B(net499));
 sg13g2_o21ai_1 _26675_ (.B1(_07513_),
    .Y(_07514_),
    .A1(_03677_),
    .A2(net499));
 sg13g2_and3_1 _26676_ (.X(_00787_),
    .A(net292),
    .B(net680),
    .C(_07514_));
 sg13g2_and4_1 _26677_ (.A(_03571_),
    .B(_11168_),
    .C(\cpu.dec.do_flush_all ),
    .D(_09288_),
    .X(_00919_));
 sg13g2_and4_1 _26678_ (.A(net993),
    .B(_10589_),
    .C(\cpu.dec.do_flush_all ),
    .D(net814),
    .X(_00937_));
 sg13g2_a21oi_1 _26679_ (.A1(_11011_),
    .A2(_09160_),
    .Y(_07515_),
    .B1(_09280_));
 sg13g2_nand2_1 _26680_ (.Y(_07516_),
    .A(_06856_),
    .B(_09280_));
 sg13g2_o21ai_1 _26681_ (.B1(_07516_),
    .Y(_07517_),
    .A1(_08419_),
    .A2(_07515_));
 sg13g2_nand2_1 _26682_ (.Y(_07518_),
    .A(net773),
    .B(net683));
 sg13g2_nor3_1 _26683_ (.A(_11619_),
    .B(_09280_),
    .C(_07518_),
    .Y(_07519_));
 sg13g2_nand3_1 _26684_ (.B(net1071),
    .C(_07519_),
    .A(net993),
    .Y(_07520_));
 sg13g2_mux2_1 _26685_ (.A0(_10580_),
    .A1(_09158_),
    .S(_07520_),
    .X(_07521_));
 sg13g2_nand2_1 _26686_ (.Y(_07522_),
    .A(net499),
    .B(_07521_));
 sg13g2_o21ai_1 _26687_ (.B1(_07522_),
    .Y(_07523_),
    .A1(_10984_),
    .A2(net499));
 sg13g2_and3_1 _26688_ (.X(_00938_),
    .A(_12014_),
    .B(_07517_),
    .C(_07523_));
 sg13g2_nand2_1 _26689_ (.Y(_07524_),
    .A(_08355_),
    .B(net814));
 sg13g2_nor2_1 _26690_ (.A(_00291_),
    .B(_07524_),
    .Y(_07525_));
 sg13g2_nand4_1 _26691_ (.B(_09162_),
    .C(_09734_),
    .A(net350),
    .Y(_07526_),
    .D(_09737_));
 sg13g2_a22oi_1 _26692_ (.Y(_07527_),
    .B1(_12274_),
    .B2(net1071),
    .A2(_07526_),
    .A1(_09303_));
 sg13g2_a21oi_1 _26693_ (.A1(_11635_),
    .A2(_07527_),
    .Y(_07528_),
    .B1(_08355_));
 sg13g2_nor2_1 _26694_ (.A(_09259_),
    .B(_07528_),
    .Y(_07529_));
 sg13g2_o21ai_1 _26695_ (.B1(_07529_),
    .Y(_07530_),
    .A1(_08268_),
    .A2(_07525_));
 sg13g2_and3_1 _26696_ (.X(_07531_),
    .A(net877),
    .B(_08290_),
    .C(_04832_));
 sg13g2_o21ai_1 _26697_ (.B1(_07531_),
    .Y(_07532_),
    .A1(\cpu.ex.c_mult[0] ),
    .A2(net246));
 sg13g2_nor2b_1 _26698_ (.A(_07530_),
    .B_N(_07532_),
    .Y(_01056_));
 sg13g2_nand2_1 _26699_ (.Y(_07533_),
    .A(_04832_),
    .B(_07525_));
 sg13g2_a22oi_1 _26700_ (.Y(_07534_),
    .B1(_07525_),
    .B2(_08375_),
    .A2(_07529_),
    .A1(_08267_));
 sg13g2_o21ai_1 _26701_ (.B1(_07534_),
    .Y(_01057_),
    .A1(_04811_),
    .A2(_07533_));
 sg13g2_inv_1 _26702_ (.Y(_07535_),
    .A(\cpu.icache.r_valid[0] ));
 sg13g2_nand2b_1 _26703_ (.Y(_07536_),
    .B(net933),
    .A_N(\cpu.ex.i_flush_all ));
 sg13g2_buf_2 _26704_ (.A(_07536_),
    .X(_07537_));
 sg13g2_a21oi_1 _26705_ (.A1(_07535_),
    .A2(_06525_),
    .Y(_02412_),
    .B1(_07537_));
 sg13g2_nor2_1 _26706_ (.A(\cpu.icache.r_valid[1] ),
    .B(_06445_),
    .Y(_07538_));
 sg13g2_nor2_1 _26707_ (.A(_07537_),
    .B(_07538_),
    .Y(_02413_));
 sg13g2_nor2_1 _26708_ (.A(\cpu.icache.r_valid[2] ),
    .B(_06462_),
    .Y(_07539_));
 sg13g2_nor2_1 _26709_ (.A(_07537_),
    .B(_07539_),
    .Y(_02414_));
 sg13g2_inv_1 _26710_ (.Y(_07540_),
    .A(\cpu.icache.r_valid[3] ));
 sg13g2_a21oi_1 _26711_ (.A1(_07540_),
    .A2(net305),
    .Y(_02415_),
    .B1(_07537_));
 sg13g2_nor2_1 _26712_ (.A(\cpu.icache.r_valid[4] ),
    .B(_06487_),
    .Y(_07541_));
 sg13g2_nor2_1 _26713_ (.A(_07537_),
    .B(_07541_),
    .Y(_02416_));
 sg13g2_nor2_1 _26714_ (.A(\cpu.icache.r_valid[5] ),
    .B(_06502_),
    .Y(_07542_));
 sg13g2_nor2_1 _26715_ (.A(_07537_),
    .B(_07542_),
    .Y(_02417_));
 sg13g2_inv_1 _26716_ (.Y(_07543_),
    .A(\cpu.icache.r_valid[6] ));
 sg13g2_a21oi_1 _26717_ (.A1(_07543_),
    .A2(_06511_),
    .Y(_02418_),
    .B1(_07537_));
 sg13g2_nor2_1 _26718_ (.A(\cpu.icache.r_valid[7] ),
    .B(_06522_),
    .Y(_07544_));
 sg13g2_nor2_1 _26719_ (.A(_07537_),
    .B(_07544_),
    .Y(_02419_));
 sg13g2_nand3_1 _26720_ (.B(net234),
    .C(net409),
    .A(net1144),
    .Y(_07545_));
 sg13g2_and2_1 _26721_ (.A(net234),
    .B(_04931_),
    .X(_07546_));
 sg13g2_buf_1 _26722_ (.A(_07546_),
    .X(_07547_));
 sg13g2_a22oi_1 _26723_ (.Y(_07548_),
    .B1(_07547_),
    .B2(net1009),
    .A2(_07545_),
    .A1(_09118_));
 sg13g2_nor2_1 _26724_ (.A(net647),
    .B(_07548_),
    .Y(_00308_));
 sg13g2_nor2_1 _26725_ (.A(_03012_),
    .B(_12148_),
    .Y(_07549_));
 sg13g2_nor2b_1 _26726_ (.A(_07549_),
    .B_N(_00306_),
    .Y(_00577_));
 sg13g2_nor2_1 _26727_ (.A(_12153_),
    .B(_12196_),
    .Y(_07550_));
 sg13g2_nor2_1 _26728_ (.A(_07549_),
    .B(_07550_),
    .Y(_00578_));
 sg13g2_xnor2_1 _26729_ (.Y(_07551_),
    .A(_06799_),
    .B(_12129_));
 sg13g2_nor2_1 _26730_ (.A(_07549_),
    .B(_07551_),
    .Y(_00579_));
 sg13g2_mux2_1 _26731_ (.A0(net418),
    .A1(_08424_),
    .S(_07512_),
    .X(_07552_));
 sg13g2_and2_1 _26732_ (.A(_09107_),
    .B(_07552_),
    .X(_00788_));
 sg13g2_a21oi_2 _26733_ (.B1(net247),
    .Y(_07553_),
    .A2(_11624_),
    .A1(_11617_));
 sg13g2_and2_1 _26734_ (.A(net825),
    .B(_07553_),
    .X(_07554_));
 sg13g2_nor2b_1 _26735_ (.A(_10994_),
    .B_N(_07519_),
    .Y(_07555_));
 sg13g2_o21ai_1 _26736_ (.B1(_09104_),
    .Y(_07556_),
    .A1(net825),
    .A2(_07555_));
 sg13g2_nand2b_1 _26737_ (.Y(_07557_),
    .B(_07556_),
    .A_N(_03666_));
 sg13g2_nand2_1 _26738_ (.Y(_07558_),
    .A(_10994_),
    .B(_07557_));
 sg13g2_o21ai_1 _26739_ (.B1(_07558_),
    .Y(_07559_),
    .A1(_10984_),
    .A2(_07557_));
 sg13g2_nor2_1 _26740_ (.A(_07553_),
    .B(_07559_),
    .Y(_07560_));
 sg13g2_o21ai_1 _26741_ (.B1(_09812_),
    .Y(_00789_),
    .A1(_07554_),
    .A2(_07560_));
 sg13g2_nand2_1 _26742_ (.Y(_07561_),
    .A(_10402_),
    .B(net499));
 sg13g2_o21ai_1 _26743_ (.B1(_07561_),
    .Y(_07562_),
    .A1(net889),
    .A2(net499));
 sg13g2_and2_1 _26744_ (.A(_09107_),
    .B(_07562_),
    .X(_00790_));
 sg13g2_nor2_1 _26745_ (.A(_06856_),
    .B(_03397_),
    .Y(_07563_));
 sg13g2_nor4_1 _26746_ (.A(\cpu.ex.r_branch_stall ),
    .B(_11616_),
    .C(_03558_),
    .D(_07524_),
    .Y(_07564_));
 sg13g2_nor3_1 _26747_ (.A(_03729_),
    .B(_07528_),
    .C(_07564_),
    .Y(_07565_));
 sg13g2_nand2_1 _26748_ (.Y(_07566_),
    .A(_08377_),
    .B(_11618_));
 sg13g2_o21ai_1 _26749_ (.B1(_05024_),
    .Y(_07567_),
    .A1(_07565_),
    .A2(_07566_));
 sg13g2_nor2_1 _26750_ (.A(net840),
    .B(_07567_),
    .Y(_07568_));
 sg13g2_o21ai_1 _26751_ (.B1(_09812_),
    .Y(_00935_),
    .A1(_07563_),
    .A2(_07568_));
 sg13g2_nand2_1 _26752_ (.Y(_07569_),
    .A(_09303_),
    .B(_09280_));
 sg13g2_nand3_1 _26753_ (.B(\cpu.dec.do_flush_write ),
    .C(_12024_),
    .A(net993),
    .Y(_07570_));
 sg13g2_a21oi_1 _26754_ (.A1(_07569_),
    .A2(_07570_),
    .Y(_00936_),
    .B1(net593));
 sg13g2_nand2_1 _26755_ (.Y(_07571_),
    .A(\cpu.dec.io ),
    .B(_12024_));
 sg13g2_nand2_1 _26756_ (.Y(_07572_),
    .A(_03011_),
    .B(_09280_));
 sg13g2_a21oi_1 _26757_ (.A1(_07571_),
    .A2(_07572_),
    .Y(_00939_),
    .B1(_06745_));
 sg13g2_nor2b_1 _26758_ (.A(_09158_),
    .B_N(_07553_),
    .Y(_07573_));
 sg13g2_nand2_1 _26759_ (.Y(_07574_),
    .A(_10580_),
    .B(net499));
 sg13g2_o21ai_1 _26760_ (.B1(_07574_),
    .Y(_07575_),
    .A1(_10039_),
    .A2(net499));
 sg13g2_nor2_1 _26761_ (.A(_07553_),
    .B(_07575_),
    .Y(_07576_));
 sg13g2_nor3_1 _26762_ (.A(_09260_),
    .B(_07573_),
    .C(_07576_),
    .Y(_00986_));
 sg13g2_buf_1 _26763_ (.A(net815),
    .X(_07577_));
 sg13g2_buf_1 _26764_ (.A(_07577_),
    .X(_07578_));
 sg13g2_a22oi_1 _26765_ (.Y(_07579_),
    .B1(_11637_),
    .B2(net1081),
    .A2(_12024_),
    .A1(_11616_));
 sg13g2_nor2_1 _26766_ (.A(_07578_),
    .B(_07579_),
    .Y(_00987_));
 sg13g2_and2_1 _26767_ (.A(_10984_),
    .B(_05796_),
    .X(_07580_));
 sg13g2_buf_2 _26768_ (.A(_07580_),
    .X(_07581_));
 sg13g2_nand2_1 _26769_ (.Y(_07582_),
    .A(_03622_),
    .B(_07581_));
 sg13g2_o21ai_1 _26770_ (.B1(_07582_),
    .Y(_07583_),
    .A1(_11058_),
    .A2(_07581_));
 sg13g2_nand2_1 _26771_ (.Y(_07584_),
    .A(net292),
    .B(_07583_));
 sg13g2_a21oi_1 _26772_ (.A1(_11617_),
    .A2(_07584_),
    .Y(_01062_),
    .B1(_06745_));
 sg13g2_nand2_1 _26773_ (.Y(_07585_),
    .A(_03620_),
    .B(_07581_));
 sg13g2_o21ai_1 _26774_ (.B1(_07585_),
    .Y(_07586_),
    .A1(_05848_),
    .A2(_07581_));
 sg13g2_nor2_1 _26775_ (.A(net708),
    .B(net292),
    .Y(_07587_));
 sg13g2_a21oi_1 _26776_ (.A1(net292),
    .A2(_07586_),
    .Y(_07588_),
    .B1(_07587_));
 sg13g2_nor2_1 _26777_ (.A(net590),
    .B(_07588_),
    .Y(_01063_));
 sg13g2_mux2_1 _26778_ (.A0(\cpu.ex.mmu_read[1] ),
    .A1(_10028_),
    .S(_07581_),
    .X(_07589_));
 sg13g2_nand2_1 _26779_ (.Y(_07590_),
    .A(net498),
    .B(_07589_));
 sg13g2_buf_1 _26780_ (.A(_09772_),
    .X(_07591_));
 sg13g2_a21oi_1 _26781_ (.A1(net358),
    .A2(_07590_),
    .Y(_01064_),
    .B1(_07591_));
 sg13g2_nor2_1 _26782_ (.A(net978),
    .B(_05807_),
    .Y(_07592_));
 sg13g2_nor2_1 _26783_ (.A(net1124),
    .B(net1123),
    .Y(_07593_));
 sg13g2_and3_1 _26784_ (.X(_07594_),
    .A(net1035),
    .B(net1100),
    .C(_07593_));
 sg13g2_buf_1 _26785_ (.A(_07594_),
    .X(_07595_));
 sg13g2_and2_1 _26786_ (.A(_07592_),
    .B(_07595_),
    .X(_07596_));
 sg13g2_buf_1 _26787_ (.A(_07596_),
    .X(_07597_));
 sg13g2_nor2b_1 _26788_ (.A(_00249_),
    .B_N(_05794_),
    .Y(_07598_));
 sg13g2_o21ai_1 _26789_ (.B1(_07598_),
    .Y(_07599_),
    .A1(_10984_),
    .A2(_00247_));
 sg13g2_a21oi_1 _26790_ (.A1(_05793_),
    .A2(_07599_),
    .Y(_07600_),
    .B1(_08419_));
 sg13g2_nand2_1 _26791_ (.Y(_07601_),
    .A(_05793_),
    .B(_07600_));
 sg13g2_buf_1 _26792_ (.A(_07601_),
    .X(_07602_));
 sg13g2_a21oi_1 _26793_ (.A1(_03447_),
    .A2(_11168_),
    .Y(_07603_),
    .B1(_05793_));
 sg13g2_nor2b_1 _26794_ (.A(_07603_),
    .B_N(_07600_),
    .Y(_07604_));
 sg13g2_buf_2 _26795_ (.A(_07604_),
    .X(_07605_));
 sg13g2_o21ai_1 _26796_ (.B1(_07605_),
    .Y(_07606_),
    .A1(_07597_),
    .A2(net162));
 sg13g2_nor2_1 _26797_ (.A(net694),
    .B(_07601_),
    .Y(_07607_));
 sg13g2_buf_2 _26798_ (.A(_07607_),
    .X(_07608_));
 sg13g2_buf_1 _26799_ (.A(_07608_),
    .X(_07609_));
 sg13g2_a22oi_1 _26800_ (.Y(_07610_),
    .B1(_07609_),
    .B2(_07597_),
    .A2(_07606_),
    .A1(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_nor2_1 _26801_ (.A(net590),
    .B(_07610_),
    .Y(_01065_));
 sg13g2_nor3_1 _26802_ (.A(net979),
    .B(_12140_),
    .C(net746),
    .Y(_07611_));
 sg13g2_buf_2 _26803_ (.A(_07611_),
    .X(_07612_));
 sg13g2_a21oi_1 _26804_ (.A1(net1100),
    .A2(_07593_),
    .Y(_07613_),
    .B1(_11336_));
 sg13g2_a21oi_1 _26805_ (.A1(net980),
    .A2(_07595_),
    .Y(_07614_),
    .B1(_07613_));
 sg13g2_nand2_1 _26806_ (.Y(_07615_),
    .A(_05895_),
    .B(_07595_));
 sg13g2_o21ai_1 _26807_ (.B1(_07615_),
    .Y(_07616_),
    .A1(_05833_),
    .A2(_07614_));
 sg13g2_buf_1 _26808_ (.A(_07616_),
    .X(_07617_));
 sg13g2_nor2b_2 _26809_ (.A(_07602_),
    .B_N(_07617_),
    .Y(_07618_));
 sg13g2_buf_1 _26810_ (.A(net162),
    .X(_07619_));
 sg13g2_buf_1 _26811_ (.A(_07605_),
    .X(_07620_));
 sg13g2_o21ai_1 _26812_ (.B1(net123),
    .Y(_07621_),
    .A1(_05851_),
    .A2(net124));
 sg13g2_a22oi_1 _26813_ (.Y(_07622_),
    .B1(_07621_),
    .B2(\cpu.genblk1.mmu.r_valid_d[10] ),
    .A2(_07618_),
    .A1(_07612_));
 sg13g2_nor2_1 _26814_ (.A(net590),
    .B(_07622_),
    .Y(_01066_));
 sg13g2_o21ai_1 _26815_ (.B1(net123),
    .Y(_07623_),
    .A1(_05857_),
    .A2(_07619_));
 sg13g2_a22oi_1 _26816_ (.Y(_07624_),
    .B1(_07623_),
    .B2(\cpu.genblk1.mmu.r_valid_d[11] ),
    .A2(_07608_),
    .A1(_05857_));
 sg13g2_nor2_1 _26817_ (.A(net590),
    .B(_07624_),
    .Y(_01067_));
 sg13g2_nand2_1 _26818_ (.Y(_07625_),
    .A(net979),
    .B(_12161_));
 sg13g2_nor3_1 _26819_ (.A(net980),
    .B(net1124),
    .C(_07625_),
    .Y(_07626_));
 sg13g2_buf_2 _26820_ (.A(_07626_),
    .X(_07627_));
 sg13g2_buf_1 _26821_ (.A(net162),
    .X(_07628_));
 sg13g2_nor2_1 _26822_ (.A(net1123),
    .B(net867),
    .Y(_07629_));
 sg13g2_nor3_1 _26823_ (.A(net980),
    .B(_10798_),
    .C(_05815_),
    .Y(_07630_));
 sg13g2_o21ai_1 _26824_ (.B1(net1100),
    .Y(_07631_),
    .A1(_07629_),
    .A2(_07630_));
 sg13g2_buf_1 _26825_ (.A(_07631_),
    .X(_07632_));
 sg13g2_nor2b_1 _26826_ (.A(_07632_),
    .B_N(_07617_),
    .Y(_07633_));
 sg13g2_o21ai_1 _26827_ (.B1(net123),
    .Y(_07634_),
    .A1(net122),
    .A2(_07633_));
 sg13g2_a22oi_1 _26828_ (.Y(_07635_),
    .B1(_07634_),
    .B2(\cpu.genblk1.mmu.r_valid_d[12] ),
    .A2(_07627_),
    .A1(_07618_));
 sg13g2_nor2_1 _26829_ (.A(net590),
    .B(_07635_),
    .Y(_01068_));
 sg13g2_nor2_1 _26830_ (.A(_05815_),
    .B(_05867_),
    .Y(_07636_));
 sg13g2_and2_1 _26831_ (.A(_07617_),
    .B(_07636_),
    .X(_07637_));
 sg13g2_buf_1 _26832_ (.A(_07637_),
    .X(_07638_));
 sg13g2_o21ai_1 _26833_ (.B1(net123),
    .Y(_07639_),
    .A1(net122),
    .A2(_07638_));
 sg13g2_a22oi_1 _26834_ (.Y(_07640_),
    .B1(_07639_),
    .B2(\cpu.genblk1.mmu.r_valid_d[13] ),
    .A2(_07638_),
    .A1(_07609_));
 sg13g2_nor2_1 _26835_ (.A(net590),
    .B(_07640_),
    .Y(_01069_));
 sg13g2_nor2_1 _26836_ (.A(net746),
    .B(_07625_),
    .Y(_07641_));
 sg13g2_buf_2 _26837_ (.A(_07641_),
    .X(_07642_));
 sg13g2_and2_1 _26838_ (.A(_05987_),
    .B(_07617_),
    .X(_07643_));
 sg13g2_o21ai_1 _26839_ (.B1(_07620_),
    .Y(_07644_),
    .A1(_07628_),
    .A2(_07643_));
 sg13g2_a22oi_1 _26840_ (.Y(_07645_),
    .B1(_07644_),
    .B2(\cpu.genblk1.mmu.r_valid_d[14] ),
    .A2(_07642_),
    .A1(_07618_));
 sg13g2_nor2_1 _26841_ (.A(net590),
    .B(_07645_),
    .Y(_01070_));
 sg13g2_and2_1 _26842_ (.A(_05819_),
    .B(_07617_),
    .X(_07646_));
 sg13g2_buf_1 _26843_ (.A(_07646_),
    .X(_07647_));
 sg13g2_o21ai_1 _26844_ (.B1(net123),
    .Y(_07648_),
    .A1(_07628_),
    .A2(_07647_));
 sg13g2_a22oi_1 _26845_ (.Y(_07649_),
    .B1(_07648_),
    .B2(\cpu.genblk1.mmu.r_valid_d[15] ),
    .A2(_07647_),
    .A1(net97));
 sg13g2_nor2_1 _26846_ (.A(_07578_),
    .B(_07649_),
    .Y(_01071_));
 sg13g2_a21oi_1 _26847_ (.A1(_05797_),
    .A2(_05835_),
    .Y(_07650_),
    .B1(_12140_));
 sg13g2_and2_1 _26848_ (.A(_06080_),
    .B(_07650_),
    .X(_07651_));
 sg13g2_buf_2 _26849_ (.A(_07651_),
    .X(_07652_));
 sg13g2_nand2_1 _26850_ (.Y(_07653_),
    .A(net1123),
    .B(_05806_));
 sg13g2_o21ai_1 _26851_ (.B1(_07653_),
    .Y(_07654_),
    .A1(_05835_),
    .A2(_05885_));
 sg13g2_nand2_1 _26852_ (.Y(_07655_),
    .A(net1100),
    .B(_07654_));
 sg13g2_nor2b_1 _26853_ (.A(_07655_),
    .B_N(_07617_),
    .Y(_07656_));
 sg13g2_a21oi_1 _26854_ (.A1(_03447_),
    .A2(_10551_),
    .Y(_07657_),
    .B1(_05793_));
 sg13g2_nor2b_1 _26855_ (.A(_07657_),
    .B_N(_07600_),
    .Y(_07658_));
 sg13g2_buf_2 _26856_ (.A(_07658_),
    .X(_07659_));
 sg13g2_buf_1 _26857_ (.A(_07659_),
    .X(_07660_));
 sg13g2_o21ai_1 _26858_ (.B1(net121),
    .Y(_07661_),
    .A1(net122),
    .A2(_07656_));
 sg13g2_a22oi_1 _26859_ (.Y(_07662_),
    .B1(_07661_),
    .B2(\cpu.genblk1.mmu.r_valid_d[16] ),
    .A2(_07652_),
    .A1(_07618_));
 sg13g2_nor2_1 _26860_ (.A(net590),
    .B(_07662_),
    .Y(_01072_));
 sg13g2_buf_1 _26861_ (.A(_07577_),
    .X(_07663_));
 sg13g2_nor2_1 _26862_ (.A(net979),
    .B(_05867_),
    .Y(_07664_));
 sg13g2_nand2b_1 _26863_ (.Y(_07665_),
    .B(net980),
    .A_N(net1100));
 sg13g2_a21oi_1 _26864_ (.A1(_07593_),
    .A2(_07665_),
    .Y(_07666_),
    .B1(_10743_));
 sg13g2_nor2_1 _26865_ (.A(net1125),
    .B(net1100),
    .Y(_07667_));
 sg13g2_a22oi_1 _26866_ (.Y(_07668_),
    .B1(_07667_),
    .B2(_07592_),
    .A2(_06159_),
    .A1(net1100));
 sg13g2_nor2b_1 _26867_ (.A(_07668_),
    .B_N(_07593_),
    .Y(_07669_));
 sg13g2_a21o_1 _26868_ (.A2(_07666_),
    .A1(_05833_),
    .B1(_07669_),
    .X(_07670_));
 sg13g2_buf_1 _26869_ (.A(_07670_),
    .X(_07671_));
 sg13g2_and2_1 _26870_ (.A(_07664_),
    .B(_07671_),
    .X(_07672_));
 sg13g2_buf_1 _26871_ (.A(_07672_),
    .X(_07673_));
 sg13g2_o21ai_1 _26872_ (.B1(net121),
    .Y(_07674_),
    .A1(net122),
    .A2(_07673_));
 sg13g2_a22oi_1 _26873_ (.Y(_07675_),
    .B1(_07674_),
    .B2(\cpu.genblk1.mmu.r_valid_d[17] ),
    .A2(_07673_),
    .A1(net97));
 sg13g2_nor2_1 _26874_ (.A(_07663_),
    .B(_07675_),
    .Y(_01073_));
 sg13g2_nor2b_1 _26875_ (.A(net162),
    .B_N(_07671_),
    .Y(_07676_));
 sg13g2_o21ai_1 _26876_ (.B1(net121),
    .Y(_07677_),
    .A1(_05897_),
    .A2(net124));
 sg13g2_a22oi_1 _26877_ (.Y(_07678_),
    .B1(_07677_),
    .B2(\cpu.genblk1.mmu.r_valid_d[18] ),
    .A2(_07676_),
    .A1(_07612_));
 sg13g2_nor2_1 _26878_ (.A(net588),
    .B(_07678_),
    .Y(_01074_));
 sg13g2_o21ai_1 _26879_ (.B1(net121),
    .Y(_07679_),
    .A1(_05906_),
    .A2(net124));
 sg13g2_a22oi_1 _26880_ (.Y(_07680_),
    .B1(_07679_),
    .B2(\cpu.genblk1.mmu.r_valid_d[19] ),
    .A2(_07608_),
    .A1(_05906_));
 sg13g2_nor2_1 _26881_ (.A(net588),
    .B(_07680_),
    .Y(_01075_));
 sg13g2_a22oi_1 _26882_ (.Y(_07681_),
    .B1(_05895_),
    .B2(_07667_),
    .A2(_05861_),
    .A1(net1100));
 sg13g2_nor2b_1 _26883_ (.A(_07681_),
    .B_N(_07593_),
    .Y(_07682_));
 sg13g2_a21oi_1 _26884_ (.A1(_05848_),
    .A2(_07666_),
    .Y(_07683_),
    .B1(_07682_));
 sg13g2_buf_2 _26885_ (.A(_07683_),
    .X(_07684_));
 sg13g2_nor2b_1 _26886_ (.A(_07684_),
    .B_N(_07664_),
    .Y(_07685_));
 sg13g2_o21ai_1 _26887_ (.B1(net123),
    .Y(_07686_),
    .A1(net122),
    .A2(_07685_));
 sg13g2_a22oi_1 _26888_ (.Y(_07687_),
    .B1(_07686_),
    .B2(\cpu.genblk1.mmu.r_valid_d[1] ),
    .A2(_07685_),
    .A1(net97));
 sg13g2_nor2_1 _26889_ (.A(net588),
    .B(_07687_),
    .Y(_01076_));
 sg13g2_nor2b_1 _26890_ (.A(_07632_),
    .B_N(_07671_),
    .Y(_07688_));
 sg13g2_o21ai_1 _26891_ (.B1(net121),
    .Y(_07689_),
    .A1(net122),
    .A2(_07688_));
 sg13g2_a22oi_1 _26892_ (.Y(_07690_),
    .B1(_07689_),
    .B2(\cpu.genblk1.mmu.r_valid_d[20] ),
    .A2(_07676_),
    .A1(_07627_));
 sg13g2_nor2_1 _26893_ (.A(net588),
    .B(_07690_),
    .Y(_01077_));
 sg13g2_and2_1 _26894_ (.A(_07636_),
    .B(_07671_),
    .X(_07691_));
 sg13g2_buf_1 _26895_ (.A(_07691_),
    .X(_07692_));
 sg13g2_o21ai_1 _26896_ (.B1(_07660_),
    .Y(_07693_),
    .A1(net122),
    .A2(_07692_));
 sg13g2_a22oi_1 _26897_ (.Y(_07694_),
    .B1(_07693_),
    .B2(\cpu.genblk1.mmu.r_valid_d[21] ),
    .A2(_07692_),
    .A1(net97));
 sg13g2_nor2_1 _26898_ (.A(_07663_),
    .B(_07694_),
    .Y(_01078_));
 sg13g2_and2_1 _26899_ (.A(_05987_),
    .B(_07671_),
    .X(_07695_));
 sg13g2_o21ai_1 _26900_ (.B1(_07660_),
    .Y(_07696_),
    .A1(net122),
    .A2(_07695_));
 sg13g2_a22oi_1 _26901_ (.Y(_07697_),
    .B1(_07696_),
    .B2(\cpu.genblk1.mmu.r_valid_d[22] ),
    .A2(_07676_),
    .A1(_07642_));
 sg13g2_nor2_1 _26902_ (.A(net588),
    .B(_07697_),
    .Y(_01079_));
 sg13g2_nor2_2 _26903_ (.A(_07653_),
    .B(_05884_),
    .Y(_07698_));
 sg13g2_buf_1 _26904_ (.A(net162),
    .X(_07699_));
 sg13g2_o21ai_1 _26905_ (.B1(net121),
    .Y(_07700_),
    .A1(net120),
    .A2(_07698_));
 sg13g2_a22oi_1 _26906_ (.Y(_07701_),
    .B1(_07700_),
    .B2(\cpu.genblk1.mmu.r_valid_d[23] ),
    .A2(_07698_),
    .A1(net97));
 sg13g2_nor2_1 _26907_ (.A(net588),
    .B(_07701_),
    .Y(_01080_));
 sg13g2_nor2b_1 _26908_ (.A(_07655_),
    .B_N(_07671_),
    .Y(_07702_));
 sg13g2_o21ai_1 _26909_ (.B1(net121),
    .Y(_07703_),
    .A1(net120),
    .A2(_07702_));
 sg13g2_a22oi_1 _26910_ (.Y(_07704_),
    .B1(_07703_),
    .B2(\cpu.genblk1.mmu.r_valid_d[24] ),
    .A2(_07676_),
    .A1(_07652_));
 sg13g2_nor2_1 _26911_ (.A(net588),
    .B(_07704_),
    .Y(_01081_));
 sg13g2_nor2_1 _26912_ (.A(_05848_),
    .B(_07614_),
    .Y(_07705_));
 sg13g2_or2_1 _26913_ (.X(_07706_),
    .B(_07705_),
    .A(_07597_));
 sg13g2_buf_1 _26914_ (.A(_07706_),
    .X(_07707_));
 sg13g2_and2_1 _26915_ (.A(_07664_),
    .B(_07707_),
    .X(_07708_));
 sg13g2_buf_1 _26916_ (.A(_07708_),
    .X(_07709_));
 sg13g2_o21ai_1 _26917_ (.B1(net121),
    .Y(_07710_),
    .A1(net120),
    .A2(_07709_));
 sg13g2_a22oi_1 _26918_ (.Y(_07711_),
    .B1(_07710_),
    .B2(\cpu.genblk1.mmu.r_valid_d[25] ),
    .A2(_07709_),
    .A1(net97));
 sg13g2_nor2_1 _26919_ (.A(net588),
    .B(_07711_),
    .Y(_01082_));
 sg13g2_buf_1 _26920_ (.A(_07577_),
    .X(_07712_));
 sg13g2_nor2b_1 _26921_ (.A(net162),
    .B_N(_07707_),
    .Y(_07713_));
 sg13g2_o21ai_1 _26922_ (.B1(_07659_),
    .Y(_07714_),
    .A1(_05942_),
    .A2(net124));
 sg13g2_a22oi_1 _26923_ (.Y(_07715_),
    .B1(_07714_),
    .B2(\cpu.genblk1.mmu.r_valid_d[26] ),
    .A2(_07713_),
    .A1(_07612_));
 sg13g2_nor2_1 _26924_ (.A(net587),
    .B(_07715_),
    .Y(_01083_));
 sg13g2_o21ai_1 _26925_ (.B1(_07659_),
    .Y(_07716_),
    .A1(_05948_),
    .A2(net124));
 sg13g2_a22oi_1 _26926_ (.Y(_07717_),
    .B1(_07716_),
    .B2(\cpu.genblk1.mmu.r_valid_d[27] ),
    .A2(_07608_),
    .A1(_05948_));
 sg13g2_nor2_1 _26927_ (.A(net587),
    .B(_07717_),
    .Y(_01084_));
 sg13g2_nor2b_1 _26928_ (.A(_07632_),
    .B_N(_07707_),
    .Y(_07718_));
 sg13g2_o21ai_1 _26929_ (.B1(_07659_),
    .Y(_07719_),
    .A1(net120),
    .A2(_07718_));
 sg13g2_a22oi_1 _26930_ (.Y(_07720_),
    .B1(_07719_),
    .B2(\cpu.genblk1.mmu.r_valid_d[28] ),
    .A2(_07713_),
    .A1(_07627_));
 sg13g2_nor2_1 _26931_ (.A(net587),
    .B(_07720_),
    .Y(_01085_));
 sg13g2_and2_1 _26932_ (.A(_07636_),
    .B(_07707_),
    .X(_07721_));
 sg13g2_buf_1 _26933_ (.A(_07721_),
    .X(_07722_));
 sg13g2_o21ai_1 _26934_ (.B1(_07659_),
    .Y(_07723_),
    .A1(net120),
    .A2(_07722_));
 sg13g2_a22oi_1 _26935_ (.Y(_07724_),
    .B1(_07723_),
    .B2(\cpu.genblk1.mmu.r_valid_d[29] ),
    .A2(_07722_),
    .A1(net97));
 sg13g2_nor2_1 _26936_ (.A(net587),
    .B(_07724_),
    .Y(_01086_));
 sg13g2_nor3_1 _26937_ (.A(net979),
    .B(net746),
    .C(_07684_),
    .Y(_07725_));
 sg13g2_o21ai_1 _26938_ (.B1(_07605_),
    .Y(_07726_),
    .A1(net162),
    .A2(_07725_));
 sg13g2_and2_1 _26939_ (.A(_12161_),
    .B(_07725_),
    .X(_07727_));
 sg13g2_inv_1 _26940_ (.Y(_07728_),
    .A(net124));
 sg13g2_a22oi_1 _26941_ (.Y(_07729_),
    .B1(_07727_),
    .B2(_07728_),
    .A2(_07726_),
    .A1(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_nor2_1 _26942_ (.A(net587),
    .B(_07729_),
    .Y(_01087_));
 sg13g2_and2_1 _26943_ (.A(_05987_),
    .B(_07707_),
    .X(_07730_));
 sg13g2_o21ai_1 _26944_ (.B1(_07659_),
    .Y(_07731_),
    .A1(net120),
    .A2(_07730_));
 sg13g2_a22oi_1 _26945_ (.Y(_07732_),
    .B1(_07731_),
    .B2(\cpu.genblk1.mmu.r_valid_d[30] ),
    .A2(_07713_),
    .A1(_07642_));
 sg13g2_nor2_1 _26946_ (.A(net587),
    .B(_07732_),
    .Y(_01088_));
 sg13g2_and2_1 _26947_ (.A(_05819_),
    .B(_07707_),
    .X(_07733_));
 sg13g2_buf_1 _26948_ (.A(_07733_),
    .X(_07734_));
 sg13g2_o21ai_1 _26949_ (.B1(_07659_),
    .Y(_07735_),
    .A1(net120),
    .A2(_07734_));
 sg13g2_a22oi_1 _26950_ (.Y(_07736_),
    .B1(_07735_),
    .B2(\cpu.genblk1.mmu.r_valid_d[31] ),
    .A2(_07734_),
    .A1(net97));
 sg13g2_nor2_1 _26951_ (.A(net587),
    .B(_07736_),
    .Y(_01089_));
 sg13g2_nor2b_1 _26952_ (.A(_07684_),
    .B_N(_07629_),
    .Y(_07737_));
 sg13g2_o21ai_1 _26953_ (.B1(net123),
    .Y(_07738_),
    .A1(_07699_),
    .A2(_07737_));
 sg13g2_a22oi_1 _26954_ (.Y(_07739_),
    .B1(_07738_),
    .B2(\cpu.genblk1.mmu.r_valid_d[3] ),
    .A2(_07737_),
    .A1(_07608_));
 sg13g2_nor2_1 _26955_ (.A(_07712_),
    .B(_07739_),
    .Y(_01090_));
 sg13g2_nor2_1 _26956_ (.A(net162),
    .B(_07684_),
    .Y(_07740_));
 sg13g2_nor2_1 _26957_ (.A(_07632_),
    .B(_07684_),
    .Y(_07741_));
 sg13g2_o21ai_1 _26958_ (.B1(net123),
    .Y(_07742_),
    .A1(_07699_),
    .A2(_07741_));
 sg13g2_a22oi_1 _26959_ (.Y(_07743_),
    .B1(_07742_),
    .B2(\cpu.genblk1.mmu.r_valid_d[4] ),
    .A2(_07740_),
    .A1(_07627_));
 sg13g2_nor2_1 _26960_ (.A(net587),
    .B(_07743_),
    .Y(_01091_));
 sg13g2_o21ai_1 _26961_ (.B1(_07620_),
    .Y(_07744_),
    .A1(_05983_),
    .A2(_07619_));
 sg13g2_a22oi_1 _26962_ (.Y(_07745_),
    .B1(_07744_),
    .B2(\cpu.genblk1.mmu.r_valid_d[5] ),
    .A2(_07608_),
    .A1(_05983_));
 sg13g2_nor2_1 _26963_ (.A(_07712_),
    .B(_07745_),
    .Y(_01092_));
 sg13g2_buf_1 _26964_ (.A(_07577_),
    .X(_07746_));
 sg13g2_o21ai_1 _26965_ (.B1(_07605_),
    .Y(_07747_),
    .A1(_05989_),
    .A2(net124));
 sg13g2_a22oi_1 _26966_ (.Y(_07748_),
    .B1(_07747_),
    .B2(\cpu.genblk1.mmu.r_valid_d[6] ),
    .A2(_07740_),
    .A1(_07642_));
 sg13g2_nor2_1 _26967_ (.A(net586),
    .B(_07748_),
    .Y(_01093_));
 sg13g2_o21ai_1 _26968_ (.B1(_07605_),
    .Y(_07749_),
    .A1(_05994_),
    .A2(net124));
 sg13g2_a22oi_1 _26969_ (.Y(_07750_),
    .B1(_07749_),
    .B2(\cpu.genblk1.mmu.r_valid_d[7] ),
    .A2(_07608_),
    .A1(_05994_));
 sg13g2_nor2_1 _26970_ (.A(net586),
    .B(_07750_),
    .Y(_01094_));
 sg13g2_nor2_1 _26971_ (.A(_07655_),
    .B(_07684_),
    .Y(_07751_));
 sg13g2_o21ai_1 _26972_ (.B1(_07605_),
    .Y(_07752_),
    .A1(net120),
    .A2(_07751_));
 sg13g2_a22oi_1 _26973_ (.Y(_07753_),
    .B1(_07752_),
    .B2(\cpu.genblk1.mmu.r_valid_d[8] ),
    .A2(_07740_),
    .A1(_07652_));
 sg13g2_nor2_1 _26974_ (.A(net586),
    .B(_07753_),
    .Y(_01095_));
 sg13g2_and2_1 _26975_ (.A(_07617_),
    .B(_07664_),
    .X(_07754_));
 sg13g2_buf_1 _26976_ (.A(_07754_),
    .X(_07755_));
 sg13g2_o21ai_1 _26977_ (.B1(_07605_),
    .Y(_07756_),
    .A1(_07602_),
    .A2(_07755_));
 sg13g2_a22oi_1 _26978_ (.Y(_07757_),
    .B1(_07756_),
    .B2(\cpu.genblk1.mmu.r_valid_d[9] ),
    .A2(_07755_),
    .A1(_07608_));
 sg13g2_nor2_1 _26979_ (.A(_07746_),
    .B(_07757_),
    .Y(_01096_));
 sg13g2_inv_1 _26980_ (.Y(_07758_),
    .A(_00247_));
 sg13g2_o21ai_1 _26981_ (.B1(_07598_),
    .Y(_07759_),
    .A1(_10984_),
    .A2(_07758_));
 sg13g2_a21oi_1 _26982_ (.A1(_05793_),
    .A2(_07759_),
    .Y(_07760_),
    .B1(_08419_));
 sg13g2_nand2_1 _26983_ (.Y(_07761_),
    .A(_05793_),
    .B(_07760_));
 sg13g2_buf_1 _26984_ (.A(_07761_),
    .X(_07762_));
 sg13g2_nand3_1 _26985_ (.B(_10590_),
    .C(_05791_),
    .A(_03447_),
    .Y(_07763_));
 sg13g2_and2_1 _26986_ (.A(_07760_),
    .B(_07763_),
    .X(_07764_));
 sg13g2_buf_2 _26987_ (.A(_07764_),
    .X(_07765_));
 sg13g2_o21ai_1 _26988_ (.B1(_07765_),
    .Y(_07766_),
    .A1(_07597_),
    .A2(net161));
 sg13g2_nor2_1 _26989_ (.A(_10039_),
    .B(_07761_),
    .Y(_07767_));
 sg13g2_buf_2 _26990_ (.A(_07767_),
    .X(_07768_));
 sg13g2_buf_1 _26991_ (.A(_07768_),
    .X(_07769_));
 sg13g2_a22oi_1 _26992_ (.Y(_07770_),
    .B1(net96),
    .B2(_07597_),
    .A2(_07766_),
    .A1(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_nor2_1 _26993_ (.A(net586),
    .B(_07770_),
    .Y(_01097_));
 sg13g2_nor2b_1 _26994_ (.A(net161),
    .B_N(_07617_),
    .Y(_07771_));
 sg13g2_buf_1 _26995_ (.A(net161),
    .X(_07772_));
 sg13g2_buf_1 _26996_ (.A(_07765_),
    .X(_07773_));
 sg13g2_o21ai_1 _26997_ (.B1(net118),
    .Y(_07774_),
    .A1(_05851_),
    .A2(net119));
 sg13g2_a22oi_1 _26998_ (.Y(_07775_),
    .B1(_07774_),
    .B2(\cpu.genblk1.mmu.r_valid_i[10] ),
    .A2(_07771_),
    .A1(_07612_));
 sg13g2_nor2_1 _26999_ (.A(net586),
    .B(_07775_),
    .Y(_01098_));
 sg13g2_o21ai_1 _27000_ (.B1(_07773_),
    .Y(_07776_),
    .A1(_05857_),
    .A2(_07772_));
 sg13g2_a22oi_1 _27001_ (.Y(_07777_),
    .B1(_07776_),
    .B2(\cpu.genblk1.mmu.r_valid_i[11] ),
    .A2(_07769_),
    .A1(_05857_));
 sg13g2_nor2_1 _27002_ (.A(net586),
    .B(_07777_),
    .Y(_01099_));
 sg13g2_o21ai_1 _27003_ (.B1(_07773_),
    .Y(_07778_),
    .A1(_07633_),
    .A2(net119));
 sg13g2_a22oi_1 _27004_ (.Y(_07779_),
    .B1(_07778_),
    .B2(\cpu.genblk1.mmu.r_valid_i[12] ),
    .A2(_07771_),
    .A1(_07627_));
 sg13g2_nor2_1 _27005_ (.A(net586),
    .B(_07779_),
    .Y(_01100_));
 sg13g2_o21ai_1 _27006_ (.B1(net118),
    .Y(_07780_),
    .A1(_07638_),
    .A2(net119));
 sg13g2_a22oi_1 _27007_ (.Y(_07781_),
    .B1(_07780_),
    .B2(\cpu.genblk1.mmu.r_valid_i[13] ),
    .A2(net96),
    .A1(_07638_));
 sg13g2_nor2_1 _27008_ (.A(_07746_),
    .B(_07781_),
    .Y(_01101_));
 sg13g2_o21ai_1 _27009_ (.B1(net118),
    .Y(_07782_),
    .A1(_07643_),
    .A2(net119));
 sg13g2_a22oi_1 _27010_ (.Y(_07783_),
    .B1(_07782_),
    .B2(\cpu.genblk1.mmu.r_valid_i[14] ),
    .A2(_07771_),
    .A1(_07642_));
 sg13g2_nor2_1 _27011_ (.A(net586),
    .B(_07783_),
    .Y(_01102_));
 sg13g2_buf_1 _27012_ (.A(_07577_),
    .X(_07784_));
 sg13g2_o21ai_1 _27013_ (.B1(net118),
    .Y(_07785_),
    .A1(_07647_),
    .A2(_07772_));
 sg13g2_a22oi_1 _27014_ (.Y(_07786_),
    .B1(_07785_),
    .B2(\cpu.genblk1.mmu.r_valid_i[15] ),
    .A2(_07769_),
    .A1(_07647_));
 sg13g2_nor2_1 _27015_ (.A(_07784_),
    .B(_07786_),
    .Y(_01103_));
 sg13g2_a21oi_1 _27016_ (.A1(_03447_),
    .A2(_11221_),
    .Y(_07787_),
    .B1(_05793_));
 sg13g2_nor2b_1 _27017_ (.A(_07787_),
    .B_N(_07760_),
    .Y(_07788_));
 sg13g2_buf_2 _27018_ (.A(_07788_),
    .X(_07789_));
 sg13g2_buf_1 _27019_ (.A(_07789_),
    .X(_07790_));
 sg13g2_o21ai_1 _27020_ (.B1(net117),
    .Y(_07791_),
    .A1(_07656_),
    .A2(net119));
 sg13g2_a22oi_1 _27021_ (.Y(_07792_),
    .B1(_07791_),
    .B2(\cpu.genblk1.mmu.r_valid_i[16] ),
    .A2(_07771_),
    .A1(_07652_));
 sg13g2_nor2_1 _27022_ (.A(net585),
    .B(_07792_),
    .Y(_01104_));
 sg13g2_o21ai_1 _27023_ (.B1(_07790_),
    .Y(_07793_),
    .A1(_07673_),
    .A2(net119));
 sg13g2_a22oi_1 _27024_ (.Y(_07794_),
    .B1(_07793_),
    .B2(\cpu.genblk1.mmu.r_valid_i[17] ),
    .A2(net96),
    .A1(_07673_));
 sg13g2_nor2_1 _27025_ (.A(net585),
    .B(_07794_),
    .Y(_01105_));
 sg13g2_nor2b_1 _27026_ (.A(net161),
    .B_N(_07671_),
    .Y(_07795_));
 sg13g2_o21ai_1 _27027_ (.B1(net117),
    .Y(_07796_),
    .A1(_05897_),
    .A2(net119));
 sg13g2_a22oi_1 _27028_ (.Y(_07797_),
    .B1(_07796_),
    .B2(\cpu.genblk1.mmu.r_valid_i[18] ),
    .A2(_07795_),
    .A1(_07612_));
 sg13g2_nor2_1 _27029_ (.A(net585),
    .B(_07797_),
    .Y(_01106_));
 sg13g2_buf_1 _27030_ (.A(net161),
    .X(_07798_));
 sg13g2_o21ai_1 _27031_ (.B1(net117),
    .Y(_07799_),
    .A1(_05906_),
    .A2(net116));
 sg13g2_a22oi_1 _27032_ (.Y(_07800_),
    .B1(_07799_),
    .B2(\cpu.genblk1.mmu.r_valid_i[19] ),
    .A2(net96),
    .A1(_05906_));
 sg13g2_nor2_1 _27033_ (.A(net585),
    .B(_07800_),
    .Y(_01107_));
 sg13g2_o21ai_1 _27034_ (.B1(net118),
    .Y(_07801_),
    .A1(_07685_),
    .A2(_07798_));
 sg13g2_a22oi_1 _27035_ (.Y(_07802_),
    .B1(_07801_),
    .B2(\cpu.genblk1.mmu.r_valid_i[1] ),
    .A2(net96),
    .A1(_07685_));
 sg13g2_nor2_1 _27036_ (.A(_07784_),
    .B(_07802_),
    .Y(_01108_));
 sg13g2_o21ai_1 _27037_ (.B1(net117),
    .Y(_07803_),
    .A1(_07688_),
    .A2(net116));
 sg13g2_a22oi_1 _27038_ (.Y(_07804_),
    .B1(_07803_),
    .B2(\cpu.genblk1.mmu.r_valid_i[20] ),
    .A2(_07795_),
    .A1(_07627_));
 sg13g2_nor2_1 _27039_ (.A(net585),
    .B(_07804_),
    .Y(_01109_));
 sg13g2_o21ai_1 _27040_ (.B1(net117),
    .Y(_07805_),
    .A1(_07692_),
    .A2(_07798_));
 sg13g2_a22oi_1 _27041_ (.Y(_07806_),
    .B1(_07805_),
    .B2(\cpu.genblk1.mmu.r_valid_i[21] ),
    .A2(net96),
    .A1(_07692_));
 sg13g2_nor2_1 _27042_ (.A(net585),
    .B(_07806_),
    .Y(_01110_));
 sg13g2_o21ai_1 _27043_ (.B1(net117),
    .Y(_07807_),
    .A1(_07695_),
    .A2(net116));
 sg13g2_a22oi_1 _27044_ (.Y(_07808_),
    .B1(_07807_),
    .B2(\cpu.genblk1.mmu.r_valid_i[22] ),
    .A2(_07795_),
    .A1(_07642_));
 sg13g2_nor2_1 _27045_ (.A(net585),
    .B(_07808_),
    .Y(_01111_));
 sg13g2_o21ai_1 _27046_ (.B1(net117),
    .Y(_07809_),
    .A1(_07698_),
    .A2(net116));
 sg13g2_a22oi_1 _27047_ (.Y(_07810_),
    .B1(_07809_),
    .B2(\cpu.genblk1.mmu.r_valid_i[23] ),
    .A2(net96),
    .A1(_07698_));
 sg13g2_nor2_1 _27048_ (.A(net585),
    .B(_07810_),
    .Y(_01112_));
 sg13g2_buf_1 _27049_ (.A(_07577_),
    .X(_07811_));
 sg13g2_o21ai_1 _27050_ (.B1(net117),
    .Y(_07812_),
    .A1(_07702_),
    .A2(net116));
 sg13g2_a22oi_1 _27051_ (.Y(_07813_),
    .B1(_07812_),
    .B2(\cpu.genblk1.mmu.r_valid_i[24] ),
    .A2(_07795_),
    .A1(_07652_));
 sg13g2_nor2_1 _27052_ (.A(net584),
    .B(_07813_),
    .Y(_01113_));
 sg13g2_o21ai_1 _27053_ (.B1(_07790_),
    .Y(_07814_),
    .A1(_07709_),
    .A2(net116));
 sg13g2_a22oi_1 _27054_ (.Y(_07815_),
    .B1(_07814_),
    .B2(\cpu.genblk1.mmu.r_valid_i[25] ),
    .A2(net96),
    .A1(_07709_));
 sg13g2_nor2_1 _27055_ (.A(net584),
    .B(_07815_),
    .Y(_01114_));
 sg13g2_nor2b_1 _27056_ (.A(net161),
    .B_N(_07707_),
    .Y(_07816_));
 sg13g2_o21ai_1 _27057_ (.B1(_07789_),
    .Y(_07817_),
    .A1(_05942_),
    .A2(net116));
 sg13g2_a22oi_1 _27058_ (.Y(_07818_),
    .B1(_07817_),
    .B2(\cpu.genblk1.mmu.r_valid_i[26] ),
    .A2(_07816_),
    .A1(_07612_));
 sg13g2_nor2_1 _27059_ (.A(net584),
    .B(_07818_),
    .Y(_01115_));
 sg13g2_o21ai_1 _27060_ (.B1(_07789_),
    .Y(_07819_),
    .A1(_05948_),
    .A2(net116));
 sg13g2_a22oi_1 _27061_ (.Y(_07820_),
    .B1(_07819_),
    .B2(\cpu.genblk1.mmu.r_valid_i[27] ),
    .A2(_07768_),
    .A1(_05948_));
 sg13g2_nor2_1 _27062_ (.A(net584),
    .B(_07820_),
    .Y(_01116_));
 sg13g2_buf_1 _27063_ (.A(net161),
    .X(_07821_));
 sg13g2_o21ai_1 _27064_ (.B1(_07789_),
    .Y(_07822_),
    .A1(_07718_),
    .A2(net115));
 sg13g2_a22oi_1 _27065_ (.Y(_07823_),
    .B1(_07822_),
    .B2(\cpu.genblk1.mmu.r_valid_i[28] ),
    .A2(_07816_),
    .A1(_07627_));
 sg13g2_nor2_1 _27066_ (.A(net584),
    .B(_07823_),
    .Y(_01117_));
 sg13g2_o21ai_1 _27067_ (.B1(_07789_),
    .Y(_07824_),
    .A1(_07722_),
    .A2(net115));
 sg13g2_a22oi_1 _27068_ (.Y(_07825_),
    .B1(_07824_),
    .B2(\cpu.genblk1.mmu.r_valid_i[29] ),
    .A2(_07768_),
    .A1(_07722_));
 sg13g2_nor2_1 _27069_ (.A(net584),
    .B(_07825_),
    .Y(_01118_));
 sg13g2_inv_1 _27070_ (.Y(_07826_),
    .A(net119));
 sg13g2_o21ai_1 _27071_ (.B1(net118),
    .Y(_07827_),
    .A1(_07725_),
    .A2(net115));
 sg13g2_a22oi_1 _27072_ (.Y(_07828_),
    .B1(_07827_),
    .B2(\cpu.genblk1.mmu.r_valid_i[2] ),
    .A2(_07826_),
    .A1(_07727_));
 sg13g2_nor2_1 _27073_ (.A(_07811_),
    .B(_07828_),
    .Y(_01119_));
 sg13g2_o21ai_1 _27074_ (.B1(_07789_),
    .Y(_07829_),
    .A1(_07730_),
    .A2(net115));
 sg13g2_a22oi_1 _27075_ (.Y(_07830_),
    .B1(_07829_),
    .B2(\cpu.genblk1.mmu.r_valid_i[30] ),
    .A2(_07816_),
    .A1(_07642_));
 sg13g2_nor2_1 _27076_ (.A(net584),
    .B(_07830_),
    .Y(_01120_));
 sg13g2_o21ai_1 _27077_ (.B1(_07789_),
    .Y(_07831_),
    .A1(_07734_),
    .A2(net115));
 sg13g2_a22oi_1 _27078_ (.Y(_07832_),
    .B1(_07831_),
    .B2(\cpu.genblk1.mmu.r_valid_i[31] ),
    .A2(_07768_),
    .A1(_07734_));
 sg13g2_nor2_1 _27079_ (.A(net584),
    .B(_07832_),
    .Y(_01121_));
 sg13g2_o21ai_1 _27080_ (.B1(net118),
    .Y(_07833_),
    .A1(_07737_),
    .A2(net115));
 sg13g2_a22oi_1 _27081_ (.Y(_07834_),
    .B1(_07833_),
    .B2(\cpu.genblk1.mmu.r_valid_i[3] ),
    .A2(_07768_),
    .A1(_07737_));
 sg13g2_nor2_1 _27082_ (.A(_07811_),
    .B(_07834_),
    .Y(_01122_));
 sg13g2_buf_1 _27083_ (.A(_07577_),
    .X(_07835_));
 sg13g2_nor2_1 _27084_ (.A(_07684_),
    .B(net161),
    .Y(_07836_));
 sg13g2_o21ai_1 _27085_ (.B1(net118),
    .Y(_07837_),
    .A1(_07741_),
    .A2(net115));
 sg13g2_a22oi_1 _27086_ (.Y(_07838_),
    .B1(_07837_),
    .B2(\cpu.genblk1.mmu.r_valid_i[4] ),
    .A2(_07836_),
    .A1(_07627_));
 sg13g2_nor2_1 _27087_ (.A(net583),
    .B(_07838_),
    .Y(_01123_));
 sg13g2_o21ai_1 _27088_ (.B1(_07765_),
    .Y(_07839_),
    .A1(_05983_),
    .A2(net115));
 sg13g2_a22oi_1 _27089_ (.Y(_07840_),
    .B1(_07839_),
    .B2(\cpu.genblk1.mmu.r_valid_i[5] ),
    .A2(_07768_),
    .A1(_05983_));
 sg13g2_nor2_1 _27090_ (.A(net583),
    .B(_07840_),
    .Y(_01124_));
 sg13g2_o21ai_1 _27091_ (.B1(_07765_),
    .Y(_07841_),
    .A1(_05989_),
    .A2(_07821_));
 sg13g2_a22oi_1 _27092_ (.Y(_07842_),
    .B1(_07841_),
    .B2(\cpu.genblk1.mmu.r_valid_i[6] ),
    .A2(_07836_),
    .A1(_07642_));
 sg13g2_nor2_1 _27093_ (.A(net583),
    .B(_07842_),
    .Y(_01125_));
 sg13g2_o21ai_1 _27094_ (.B1(_07765_),
    .Y(_07843_),
    .A1(_05994_),
    .A2(_07821_));
 sg13g2_a22oi_1 _27095_ (.Y(_07844_),
    .B1(_07843_),
    .B2(\cpu.genblk1.mmu.r_valid_i[7] ),
    .A2(_07768_),
    .A1(_05994_));
 sg13g2_nor2_1 _27096_ (.A(net583),
    .B(_07844_),
    .Y(_01126_));
 sg13g2_o21ai_1 _27097_ (.B1(_07765_),
    .Y(_07845_),
    .A1(_07751_),
    .A2(_07762_));
 sg13g2_a22oi_1 _27098_ (.Y(_07846_),
    .B1(_07845_),
    .B2(\cpu.genblk1.mmu.r_valid_i[8] ),
    .A2(_07836_),
    .A1(_07652_));
 sg13g2_nor2_1 _27099_ (.A(_07835_),
    .B(_07846_),
    .Y(_01127_));
 sg13g2_o21ai_1 _27100_ (.B1(_07765_),
    .Y(_07847_),
    .A1(_07755_),
    .A2(_07762_));
 sg13g2_a22oi_1 _27101_ (.Y(_07848_),
    .B1(_07847_),
    .B2(\cpu.genblk1.mmu.r_valid_i[9] ),
    .A2(_07768_),
    .A1(_07755_));
 sg13g2_nor2_1 _27102_ (.A(_07835_),
    .B(_07848_),
    .Y(_01128_));
 sg13g2_buf_1 _27103_ (.A(_06307_),
    .X(_07849_));
 sg13g2_and2_1 _27104_ (.A(_04891_),
    .B(net160),
    .X(_07850_));
 sg13g2_buf_2 _27105_ (.A(_07850_),
    .X(_07851_));
 sg13g2_nand2_1 _27106_ (.Y(_07852_),
    .A(net960),
    .B(_07851_));
 sg13g2_nand2_1 _27107_ (.Y(_07853_),
    .A(_04891_),
    .B(_06307_));
 sg13g2_buf_2 _27108_ (.A(_07853_),
    .X(_07854_));
 sg13g2_nand2_1 _27109_ (.Y(_07855_),
    .A(\cpu.gpio.r_enable_in[0] ),
    .B(_07854_));
 sg13g2_a21oi_1 _27110_ (.A1(_07852_),
    .A2(_07855_),
    .Y(_01929_),
    .B1(net589));
 sg13g2_nand2_1 _27111_ (.Y(_07856_),
    .A(net1055),
    .B(_07851_));
 sg13g2_nand2_1 _27112_ (.Y(_07857_),
    .A(_09125_),
    .B(_07854_));
 sg13g2_a21oi_1 _27113_ (.A1(_07856_),
    .A2(_07857_),
    .Y(_01930_),
    .B1(net589));
 sg13g2_nand2_1 _27114_ (.Y(_07858_),
    .A(_09985_),
    .B(_07851_));
 sg13g2_nand2_1 _27115_ (.Y(_07859_),
    .A(_09136_),
    .B(_07854_));
 sg13g2_a21oi_1 _27116_ (.A1(_07858_),
    .A2(_07859_),
    .Y(_01931_),
    .B1(net589));
 sg13g2_nand2_1 _27117_ (.Y(_07860_),
    .A(net1058),
    .B(_07851_));
 sg13g2_nand2_1 _27118_ (.Y(_07861_),
    .A(_09144_),
    .B(_07854_));
 sg13g2_a21oi_1 _27119_ (.A1(_07860_),
    .A2(_07861_),
    .Y(_01932_),
    .B1(net589));
 sg13g2_nand2_1 _27120_ (.Y(_07862_),
    .A(net1057),
    .B(_07851_));
 sg13g2_nand2_1 _27121_ (.Y(_07863_),
    .A(_09146_),
    .B(_07854_));
 sg13g2_a21oi_1 _27122_ (.A1(_07862_),
    .A2(_07863_),
    .Y(_01933_),
    .B1(net589));
 sg13g2_nand2_1 _27123_ (.Y(_07864_),
    .A(net1054),
    .B(_07851_));
 sg13g2_nand2_1 _27124_ (.Y(_07865_),
    .A(_09127_),
    .B(_07854_));
 sg13g2_a21oi_1 _27125_ (.A1(_07864_),
    .A2(_07865_),
    .Y(_01934_),
    .B1(_07591_));
 sg13g2_nand2_1 _27126_ (.Y(_07866_),
    .A(net1053),
    .B(_07851_));
 sg13g2_nand2_1 _27127_ (.Y(_07867_),
    .A(_09150_),
    .B(_07854_));
 sg13g2_a21oi_1 _27128_ (.A1(_07866_),
    .A2(_07867_),
    .Y(_01935_),
    .B1(net589));
 sg13g2_nand2_1 _27129_ (.Y(_07868_),
    .A(net1056),
    .B(_07851_));
 sg13g2_nand2_1 _27130_ (.Y(_07869_),
    .A(_09138_),
    .B(_07854_));
 sg13g2_a21oi_1 _27131_ (.A1(_07868_),
    .A2(_07869_),
    .Y(_01936_),
    .B1(net589));
 sg13g2_nand3_1 _27132_ (.B(net410),
    .C(net160),
    .A(_10000_),
    .Y(_07870_));
 sg13g2_nand2_1 _27133_ (.Y(_07871_),
    .A(net410),
    .B(net160));
 sg13g2_nand2_1 _27134_ (.Y(_07872_),
    .A(\cpu.gpio.r_enable_io[4] ),
    .B(_07871_));
 sg13g2_a21oi_1 _27135_ (.A1(_07870_),
    .A2(_07872_),
    .Y(_01937_),
    .B1(net589));
 sg13g2_nand3_1 _27136_ (.B(net410),
    .C(net160),
    .A(net1054),
    .Y(_07873_));
 sg13g2_nand2_1 _27137_ (.Y(_07874_),
    .A(\cpu.gpio.r_enable_io[5] ),
    .B(_07871_));
 sg13g2_buf_1 _27138_ (.A(_09772_),
    .X(_07875_));
 sg13g2_a21oi_1 _27139_ (.A1(_07873_),
    .A2(_07874_),
    .Y(_01938_),
    .B1(net582));
 sg13g2_nand3_1 _27140_ (.B(net410),
    .C(net160),
    .A(_10010_),
    .Y(_07876_));
 sg13g2_nand2_1 _27141_ (.Y(_07877_),
    .A(_09130_),
    .B(_07871_));
 sg13g2_a21oi_1 _27142_ (.A1(_07876_),
    .A2(_07877_),
    .Y(_01939_),
    .B1(net582));
 sg13g2_nand3_1 _27143_ (.B(net410),
    .C(net160),
    .A(_10015_),
    .Y(_07878_));
 sg13g2_nand2_1 _27144_ (.Y(_07879_),
    .A(\cpu.gpio.r_enable_io[7] ),
    .B(_07871_));
 sg13g2_a21oi_1 _27145_ (.A1(_07878_),
    .A2(_07879_),
    .Y(_01940_),
    .B1(net582));
 sg13g2_nand3_1 _27146_ (.B(net601),
    .C(_06307_),
    .A(net869),
    .Y(_07880_));
 sg13g2_buf_2 _27147_ (.A(_07880_),
    .X(_07881_));
 sg13g2_mux2_1 _27148_ (.A0(_09999_),
    .A1(net7),
    .S(_07881_),
    .X(_07882_));
 sg13g2_and2_1 _27149_ (.A(net717),
    .B(_07882_),
    .X(_01941_));
 sg13g2_nand2_1 _27150_ (.Y(_07883_),
    .A(net8),
    .B(_07881_));
 sg13g2_o21ai_1 _27151_ (.B1(_07883_),
    .Y(_07884_),
    .A1(_12261_),
    .A2(_07881_));
 sg13g2_and2_1 _27152_ (.A(net717),
    .B(_07884_),
    .X(_01942_));
 sg13g2_nand2_1 _27153_ (.Y(_07885_),
    .A(net9),
    .B(_07881_));
 sg13g2_o21ai_1 _27154_ (.B1(_07885_),
    .Y(_07886_),
    .A1(_12265_),
    .A2(_07881_));
 sg13g2_and2_1 _27155_ (.A(net717),
    .B(_07886_),
    .X(_01943_));
 sg13g2_nand2_1 _27156_ (.Y(_07887_),
    .A(net10),
    .B(_07881_));
 sg13g2_o21ai_1 _27157_ (.B1(_07887_),
    .Y(_07888_),
    .A1(_12269_),
    .A2(_07881_));
 sg13g2_and2_1 _27158_ (.A(net717),
    .B(_07888_),
    .X(_01944_));
 sg13g2_nand2b_1 _27159_ (.Y(_07889_),
    .B(_06307_),
    .A_N(_05340_));
 sg13g2_buf_2 _27160_ (.A(_07889_),
    .X(_07890_));
 sg13g2_nor2_1 _27161_ (.A(net960),
    .B(_07890_),
    .Y(_07891_));
 sg13g2_nor2b_1 _27162_ (.A(_04853_),
    .B_N(_07890_),
    .Y(_07892_));
 sg13g2_o21ai_1 _27163_ (.B1(net696),
    .Y(_01990_),
    .A1(_07891_),
    .A2(_07892_));
 sg13g2_buf_1 _27164_ (.A(\cpu.gpio.r_src_o[6][1] ),
    .X(_07893_));
 sg13g2_nand2_1 _27165_ (.Y(_07894_),
    .A(_07893_),
    .B(_07890_));
 sg13g2_o21ai_1 _27166_ (.B1(_07894_),
    .Y(_07895_),
    .A1(net897),
    .A2(_07890_));
 sg13g2_and2_1 _27167_ (.A(net717),
    .B(_07895_),
    .X(_01991_));
 sg13g2_nand2_1 _27168_ (.Y(_07896_),
    .A(\cpu.gpio.r_src_o[6][2] ),
    .B(_07890_));
 sg13g2_o21ai_1 _27169_ (.B1(_07896_),
    .Y(_07897_),
    .A1(_12240_),
    .A2(_07890_));
 sg13g2_and2_1 _27170_ (.A(net717),
    .B(_07897_),
    .X(_01992_));
 sg13g2_mux2_1 _27171_ (.A0(net1144),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .S(_07890_),
    .X(_07898_));
 sg13g2_and2_1 _27172_ (.A(net680),
    .B(_07898_),
    .X(_01993_));
 sg13g2_nand3_1 _27173_ (.B(net670),
    .C(net160),
    .A(net960),
    .Y(_07899_));
 sg13g2_nand2_1 _27174_ (.Y(_07900_),
    .A(net670),
    .B(_07849_));
 sg13g2_nand2_1 _27175_ (.Y(_07901_),
    .A(_04841_),
    .B(_07900_));
 sg13g2_a21oi_1 _27176_ (.A1(_07899_),
    .A2(_07901_),
    .Y(_01998_),
    .B1(net582));
 sg13g2_nand3_1 _27177_ (.B(_04843_),
    .C(net160),
    .A(net1055),
    .Y(_07902_));
 sg13g2_nand2_1 _27178_ (.Y(_07903_),
    .A(\cpu.gpio.r_uart_rx_src[1] ),
    .B(_07900_));
 sg13g2_a21oi_1 _27179_ (.A1(_07902_),
    .A2(_07903_),
    .Y(_01999_),
    .B1(_07875_));
 sg13g2_nand3_1 _27180_ (.B(_04843_),
    .C(_07849_),
    .A(net1059),
    .Y(_07904_));
 sg13g2_nand2_1 _27181_ (.Y(_07905_),
    .A(\cpu.gpio.r_uart_rx_src[2] ),
    .B(_07900_));
 sg13g2_a21oi_1 _27182_ (.A1(_07904_),
    .A2(_07905_),
    .Y(_02000_),
    .B1(_07875_));
 sg13g2_and2_1 _27183_ (.A(\cpu.i_wstrobe_d ),
    .B(_00307_),
    .X(_02257_));
 sg13g2_nor2_1 _27184_ (.A(_06384_),
    .B(_06396_),
    .Y(_07906_));
 sg13g2_nor2_1 _27185_ (.A(_06410_),
    .B(_07906_),
    .Y(_02258_));
 sg13g2_xor2_1 _27186_ (.B(_06391_),
    .A(\cpu.icache.r_offset[2] ),
    .X(_07907_));
 sg13g2_nor2_1 _27187_ (.A(_06410_),
    .B(_07907_),
    .Y(_02259_));
 sg13g2_xnor2_1 _27188_ (.Y(_07908_),
    .A(\cpu.intr.r_clock_cmp[26] ),
    .B(_05142_));
 sg13g2_xnor2_1 _27189_ (.Y(_07909_),
    .A(\cpu.intr.r_clock_cmp[13] ),
    .B(_10105_));
 sg13g2_xnor2_1 _27190_ (.Y(_07910_),
    .A(\cpu.intr.r_clock_cmp[16] ),
    .B(_04919_));
 sg13g2_xnor2_1 _27191_ (.Y(_07911_),
    .A(\cpu.intr.r_clock_cmp[6] ),
    .B(_10065_));
 sg13g2_nand4_1 _27192_ (.B(_07909_),
    .C(_07910_),
    .A(_07908_),
    .Y(_07912_),
    .D(_07911_));
 sg13g2_xnor2_1 _27193_ (.Y(_07913_),
    .A(\cpu.intr.r_clock_cmp[22] ),
    .B(_05659_));
 sg13g2_xnor2_1 _27194_ (.Y(_07914_),
    .A(\cpu.intr.r_clock_cmp[19] ),
    .B(_05495_));
 sg13g2_xnor2_1 _27195_ (.Y(_07915_),
    .A(\cpu.intr.r_clock_cmp[29] ),
    .B(_05222_));
 sg13g2_xnor2_1 _27196_ (.Y(_07916_),
    .A(\cpu.intr.r_clock_cmp[4] ),
    .B(_10053_));
 sg13g2_nand4_1 _27197_ (.B(_07914_),
    .C(_07915_),
    .A(_07913_),
    .Y(_07917_),
    .D(_07916_));
 sg13g2_xnor2_1 _27198_ (.Y(_07918_),
    .A(\cpu.intr.r_clock_cmp[5] ),
    .B(_10059_));
 sg13g2_xnor2_1 _27199_ (.Y(_07919_),
    .A(\cpu.intr.r_clock_cmp[30] ),
    .B(_05272_));
 sg13g2_xnor2_1 _27200_ (.Y(_07920_),
    .A(\cpu.intr.r_clock_cmp[11] ),
    .B(_10093_));
 sg13g2_xnor2_1 _27201_ (.Y(_07921_),
    .A(\cpu.intr.r_clock_cmp[20] ),
    .B(_05542_));
 sg13g2_nand4_1 _27202_ (.B(_07919_),
    .C(_07920_),
    .A(_07918_),
    .Y(_07922_),
    .D(_07921_));
 sg13g2_xnor2_1 _27203_ (.Y(_07923_),
    .A(\cpu.intr.r_clock_cmp[21] ),
    .B(_05636_));
 sg13g2_xnor2_1 _27204_ (.Y(_07924_),
    .A(\cpu.intr.r_clock_cmp[10] ),
    .B(_10088_));
 sg13g2_xnor2_1 _27205_ (.Y(_07925_),
    .A(\cpu.intr.r_clock_cmp[17] ),
    .B(_05359_));
 sg13g2_xnor2_1 _27206_ (.Y(_07926_),
    .A(\cpu.intr.r_clock_cmp[15] ),
    .B(_10116_));
 sg13g2_nand4_1 _27207_ (.B(_07924_),
    .C(_07925_),
    .A(_07923_),
    .Y(_07927_),
    .D(_07926_));
 sg13g2_nor4_1 _27208_ (.A(_07912_),
    .B(_07917_),
    .C(_07922_),
    .D(_07927_),
    .Y(_07928_));
 sg13g2_xnor2_1 _27209_ (.Y(_07929_),
    .A(\cpu.intr.r_clock_cmp[27] ),
    .B(_05165_));
 sg13g2_xnor2_1 _27210_ (.Y(_07930_),
    .A(\cpu.intr.r_clock_cmp[31] ),
    .B(_05282_));
 sg13g2_xnor2_1 _27211_ (.Y(_07931_),
    .A(\cpu.intr.r_clock_cmp[8] ),
    .B(_10076_));
 sg13g2_xnor2_1 _27212_ (.Y(_07932_),
    .A(\cpu.intr.r_clock_cmp[9] ),
    .B(_10083_));
 sg13g2_nand4_1 _27213_ (.B(_07930_),
    .C(_07931_),
    .A(_07929_),
    .Y(_07933_),
    .D(_07932_));
 sg13g2_xnor2_1 _27214_ (.Y(_07934_),
    .A(\cpu.intr.r_clock_cmp[7] ),
    .B(_10072_));
 sg13g2_xnor2_1 _27215_ (.Y(_07935_),
    .A(\cpu.intr.r_clock_cmp[1] ),
    .B(_10037_));
 sg13g2_xnor2_1 _27216_ (.Y(_07936_),
    .A(\cpu.intr.r_clock_cmp[12] ),
    .B(_10100_));
 sg13g2_xnor2_1 _27217_ (.Y(_07937_),
    .A(\cpu.intr.r_clock_cmp[23] ),
    .B(_05067_));
 sg13g2_nand4_1 _27218_ (.B(_07935_),
    .C(_07936_),
    .A(_07934_),
    .Y(_07938_),
    .D(_07937_));
 sg13g2_xnor2_1 _27219_ (.Y(_07939_),
    .A(\cpu.intr.r_clock_cmp[28] ),
    .B(_05208_));
 sg13g2_xnor2_1 _27220_ (.Y(_07940_),
    .A(\cpu.intr.r_clock_cmp[18] ),
    .B(_05408_));
 sg13g2_xnor2_1 _27221_ (.Y(_07941_),
    .A(\cpu.intr.r_clock_cmp[14] ),
    .B(_10110_));
 sg13g2_xnor2_1 _27222_ (.Y(_07942_),
    .A(\cpu.intr.r_clock_cmp[3] ),
    .B(_10049_));
 sg13g2_nand4_1 _27223_ (.B(_07940_),
    .C(_07941_),
    .A(_07939_),
    .Y(_07943_),
    .D(_07942_));
 sg13g2_xnor2_1 _27224_ (.Y(_07944_),
    .A(\cpu.intr.r_clock_cmp[2] ),
    .B(_10045_));
 sg13g2_xnor2_1 _27225_ (.Y(_07945_),
    .A(\cpu.intr.r_clock_cmp[0] ),
    .B(_10036_));
 sg13g2_xnor2_1 _27226_ (.Y(_07946_),
    .A(\cpu.intr.r_clock_cmp[25] ),
    .B(_05740_));
 sg13g2_xnor2_1 _27227_ (.Y(_07947_),
    .A(\cpu.intr.r_clock_cmp[24] ),
    .B(_05727_));
 sg13g2_nand4_1 _27228_ (.B(_07945_),
    .C(_07946_),
    .A(_07944_),
    .Y(_07948_),
    .D(_07947_));
 sg13g2_nor4_1 _27229_ (.A(_07933_),
    .B(_07938_),
    .C(_07943_),
    .D(_07948_),
    .Y(_07949_));
 sg13g2_a22oi_1 _27230_ (.Y(_07950_),
    .B1(_07928_),
    .B2(_07949_),
    .A2(_07547_),
    .A1(net1055));
 sg13g2_nand3_1 _27231_ (.B(net234),
    .C(_04966_),
    .A(_09978_),
    .Y(_07951_));
 sg13g2_nand2_1 _27232_ (.Y(_07952_),
    .A(\cpu.intr.r_clock ),
    .B(_07951_));
 sg13g2_a21oi_1 _27233_ (.A1(_07950_),
    .A2(_07952_),
    .Y(_02420_),
    .B1(net582));
 sg13g2_and2_1 _27234_ (.A(net234),
    .B(net408),
    .X(_07953_));
 sg13g2_buf_1 _27235_ (.A(_07953_),
    .X(_07954_));
 sg13g2_nand2_1 _27236_ (.Y(_07955_),
    .A(net960),
    .B(_07954_));
 sg13g2_nand2_1 _27237_ (.Y(_07956_),
    .A(net234),
    .B(net408));
 sg13g2_buf_1 _27238_ (.A(_07956_),
    .X(_07957_));
 sg13g2_nand2_1 _27239_ (.Y(_07958_),
    .A(_09116_),
    .B(_07957_));
 sg13g2_a21oi_1 _27240_ (.A1(_07955_),
    .A2(_07958_),
    .Y(_02469_),
    .B1(net582));
 sg13g2_nand2_1 _27241_ (.Y(_07959_),
    .A(net1055),
    .B(_07954_));
 sg13g2_nand2_1 _27242_ (.Y(_07960_),
    .A(\cpu.intr.r_enable[1] ),
    .B(_07957_));
 sg13g2_a21oi_1 _27243_ (.A1(_07959_),
    .A2(_07960_),
    .Y(_02470_),
    .B1(net582));
 sg13g2_nand2_1 _27244_ (.Y(_07961_),
    .A(net1059),
    .B(_07954_));
 sg13g2_nand2_1 _27245_ (.Y(_07962_),
    .A(\cpu.intr.r_enable[2] ),
    .B(_07957_));
 sg13g2_a21oi_1 _27246_ (.A1(_07961_),
    .A2(_07962_),
    .Y(_02471_),
    .B1(net582));
 sg13g2_nand2_1 _27247_ (.Y(_07963_),
    .A(net1058),
    .B(_07954_));
 sg13g2_nand2_1 _27248_ (.Y(_07964_),
    .A(\cpu.intr.r_enable[3] ),
    .B(_07957_));
 sg13g2_buf_1 _27249_ (.A(_09772_),
    .X(_07965_));
 sg13g2_a21oi_1 _27250_ (.A1(_07963_),
    .A2(_07964_),
    .Y(_02472_),
    .B1(net581));
 sg13g2_nand2_1 _27251_ (.Y(_07966_),
    .A(_10000_),
    .B(_07954_));
 sg13g2_nand2_1 _27252_ (.Y(_07967_),
    .A(_09155_),
    .B(_07957_));
 sg13g2_a21oi_1 _27253_ (.A1(_07966_),
    .A2(_07967_),
    .Y(_02473_),
    .B1(net581));
 sg13g2_nand2_1 _27254_ (.Y(_07968_),
    .A(net1054),
    .B(_07954_));
 sg13g2_nand2_1 _27255_ (.Y(_07969_),
    .A(_09120_),
    .B(_07957_));
 sg13g2_a21oi_1 _27256_ (.A1(_07968_),
    .A2(_07969_),
    .Y(_02474_),
    .B1(net581));
 sg13g2_nand3_1 _27257_ (.B(net234),
    .C(_04966_),
    .A(net1059),
    .Y(_07970_));
 sg13g2_a22oi_1 _27258_ (.Y(_07971_),
    .B1(_07970_),
    .B2(_09112_),
    .A2(_07547_),
    .A1(net1059));
 sg13g2_a21oi_1 _27259_ (.A1(_09930_),
    .A2(_07971_),
    .Y(_02475_),
    .B1(net581));
 sg13g2_inv_1 _27260_ (.Y(_07972_),
    .A(_06772_));
 sg13g2_or4_1 _27261_ (.A(_09832_),
    .B(_09781_),
    .C(net1149),
    .D(_06770_),
    .X(_07973_));
 sg13g2_nor2_1 _27262_ (.A(_09779_),
    .B(_07973_),
    .Y(_07974_));
 sg13g2_nand2_1 _27263_ (.Y(_07975_),
    .A(_09760_),
    .B(_07974_));
 sg13g2_or4_1 _27264_ (.A(net1147),
    .B(_09809_),
    .C(_07972_),
    .D(_07975_),
    .X(_07976_));
 sg13g2_buf_1 _27265_ (.A(_07976_),
    .X(_07977_));
 sg13g2_o21ai_1 _27266_ (.B1(_09106_),
    .Y(_07978_),
    .A1(_06831_),
    .A2(_07977_));
 sg13g2_nor2b_1 _27267_ (.A(_09800_),
    .B_N(_09784_),
    .Y(_07979_));
 sg13g2_o21ai_1 _27268_ (.B1(net19),
    .Y(_07980_),
    .A1(_07977_),
    .A2(_07979_));
 sg13g2_nand2b_1 _27269_ (.Y(_02505_),
    .B(_07980_),
    .A_N(_07978_));
 sg13g2_nand3b_1 _27270_ (.B(_06784_),
    .C(_09762_),
    .Y(_07981_),
    .A_N(_09784_));
 sg13g2_a21o_1 _27271_ (.A2(_07981_),
    .A1(_06831_),
    .B1(_07977_),
    .X(_07982_));
 sg13g2_nand2_1 _27272_ (.Y(_07983_),
    .A(_09784_),
    .B(_06831_));
 sg13g2_nor2_1 _27273_ (.A(_09795_),
    .B(_07983_),
    .Y(_07984_));
 sg13g2_o21ai_1 _27274_ (.B1(net20),
    .Y(_07985_),
    .A1(_07977_),
    .A2(_07984_));
 sg13g2_nand3_1 _27275_ (.B(_07982_),
    .C(_07985_),
    .A(net663),
    .Y(_02506_));
 sg13g2_nor2b_1 _27276_ (.A(_09798_),
    .B_N(_09784_),
    .Y(_07986_));
 sg13g2_buf_1 _27277_ (.A(\cpu.gpio.genblk1[3].srcs_o[11] ),
    .X(_07987_));
 sg13g2_o21ai_1 _27278_ (.B1(_07987_),
    .Y(_07988_),
    .A1(_07977_),
    .A2(_07986_));
 sg13g2_nand2b_1 _27279_ (.Y(_02507_),
    .B(_07988_),
    .A_N(_07978_));
 sg13g2_nor4_1 _27280_ (.A(\cpu.qspi.r_state[17] ),
    .B(_09769_),
    .C(_09785_),
    .D(_06784_),
    .Y(_07989_));
 sg13g2_nand2_1 _27281_ (.Y(_07990_),
    .A(_06688_),
    .B(_07989_));
 sg13g2_nor4_1 _27282_ (.A(_09770_),
    .B(net1147),
    .C(_07973_),
    .D(_07990_),
    .Y(_07991_));
 sg13g2_a21oi_1 _27283_ (.A1(_12013_),
    .A2(_07991_),
    .Y(_07992_),
    .B1(_09762_));
 sg13g2_nor2_1 _27284_ (.A(net583),
    .B(_07992_),
    .Y(_02508_));
 sg13g2_nand2_1 _27285_ (.Y(_07993_),
    .A(net1056),
    .B(_06734_));
 sg13g2_nand2_1 _27286_ (.Y(_07994_),
    .A(\cpu.qspi.r_mask[0] ),
    .B(_06737_));
 sg13g2_a21oi_1 _27287_ (.A1(_07993_),
    .A2(_07994_),
    .Y(_02509_),
    .B1(_07965_));
 sg13g2_a21oi_1 _27288_ (.A1(net604),
    .A2(_04900_),
    .Y(_07995_),
    .B1(net1030));
 sg13g2_nand2_1 _27289_ (.Y(_07996_),
    .A(_06732_),
    .B(_07995_));
 sg13g2_o21ai_1 _27290_ (.B1(_09106_),
    .Y(_07997_),
    .A1(_07194_),
    .A2(_07996_));
 sg13g2_a21o_1 _27291_ (.A2(_06750_),
    .A1(\cpu.qspi.r_mask[1] ),
    .B1(_07997_),
    .X(_02510_));
 sg13g2_nor2_1 _27292_ (.A(_07194_),
    .B(_06762_),
    .Y(_07998_));
 sg13g2_a21oi_1 _27293_ (.A1(\cpu.qspi.r_mask[2] ),
    .A2(_06762_),
    .Y(_07999_),
    .B1(_07998_));
 sg13g2_nor2_1 _27294_ (.A(net583),
    .B(_07999_),
    .Y(_02511_));
 sg13g2_nand2_1 _27295_ (.Y(_08000_),
    .A(\cpu.qspi.r_quad[0] ),
    .B(_06737_));
 sg13g2_nand2_1 _27296_ (.Y(_08001_),
    .A(_10069_),
    .B(_06734_));
 sg13g2_nand3_1 _27297_ (.B(_08000_),
    .C(_08001_),
    .A(net663),
    .Y(_02512_));
 sg13g2_nor2_1 _27298_ (.A(_07190_),
    .B(_07996_),
    .Y(_08002_));
 sg13g2_a21oi_1 _27299_ (.A1(\cpu.qspi.r_quad[1] ),
    .A2(_06750_),
    .Y(_08003_),
    .B1(_08002_));
 sg13g2_nor2_1 _27300_ (.A(net583),
    .B(_08003_),
    .Y(_02513_));
 sg13g2_nand2_1 _27301_ (.Y(_08004_),
    .A(_07190_),
    .B(_06759_));
 sg13g2_o21ai_1 _27302_ (.B1(_08004_),
    .Y(_08005_),
    .A1(\cpu.qspi.r_quad[2] ),
    .A2(_06759_));
 sg13g2_nand2_1 _27303_ (.Y(_02514_),
    .A(net696),
    .B(_08005_));
 sg13g2_nand2b_1 _27304_ (.Y(_08006_),
    .B(_06732_),
    .A_N(_04866_));
 sg13g2_buf_1 _27305_ (.A(_08006_),
    .X(_08007_));
 sg13g2_nor2_1 _27306_ (.A(_06673_),
    .B(_08007_),
    .Y(_08008_));
 sg13g2_nor2b_1 _27307_ (.A(_09788_),
    .B_N(_08007_),
    .Y(_08009_));
 sg13g2_o21ai_1 _27308_ (.B1(net696),
    .Y(_02527_),
    .A1(_08008_),
    .A2(_08009_));
 sg13g2_nor2_1 _27309_ (.A(_10042_),
    .B(_08007_),
    .Y(_08010_));
 sg13g2_nor2b_1 _27310_ (.A(_09787_),
    .B_N(_08007_),
    .Y(_08011_));
 sg13g2_o21ai_1 _27311_ (.B1(net696),
    .Y(_02528_),
    .A1(_08010_),
    .A2(_08011_));
 sg13g2_nor2b_1 _27312_ (.A(_06829_),
    .B_N(_12018_),
    .Y(_08012_));
 sg13g2_or4_1 _27313_ (.A(_12015_),
    .B(_09769_),
    .C(net1148),
    .D(_09782_),
    .X(_08013_));
 sg13g2_nor3_2 _27314_ (.A(_07975_),
    .B(_08012_),
    .C(_08013_),
    .Y(_08014_));
 sg13g2_nand2b_1 _27315_ (.Y(_08015_),
    .B(net3),
    .A_N(_08014_));
 sg13g2_nor4_1 _27316_ (.A(_12018_),
    .B(_09770_),
    .C(_09761_),
    .D(_09807_),
    .Y(_08016_));
 sg13g2_nor3_1 _27317_ (.A(_12016_),
    .B(_06784_),
    .C(_08016_),
    .Y(_08017_));
 sg13g2_nand2b_1 _27318_ (.Y(_08018_),
    .B(_08014_),
    .A_N(_08017_));
 sg13g2_a21oi_1 _27319_ (.A1(_08015_),
    .A2(_08018_),
    .Y(_02529_),
    .B1(net581));
 sg13g2_nand2b_1 _27320_ (.Y(_08019_),
    .B(net6),
    .A_N(_08014_));
 sg13g2_nand2b_1 _27321_ (.Y(_08020_),
    .B(_08016_),
    .A_N(_06784_));
 sg13g2_o21ai_1 _27322_ (.B1(_12017_),
    .Y(_08021_),
    .A1(_09803_),
    .A2(_08020_));
 sg13g2_nand2_1 _27323_ (.Y(_08022_),
    .A(_08014_),
    .B(_08021_));
 sg13g2_a21oi_1 _27324_ (.A1(_08019_),
    .A2(_08022_),
    .Y(_02530_),
    .B1(_07965_));
 sg13g2_nor3_1 _27325_ (.A(net1151),
    .B(net1152),
    .C(_09265_),
    .Y(_08023_));
 sg13g2_nor3_1 _27326_ (.A(_09262_),
    .B(_09270_),
    .C(_08023_),
    .Y(_08024_));
 sg13g2_buf_1 _27327_ (.A(_08024_),
    .X(_08025_));
 sg13g2_nand3_1 _27328_ (.B(net1151),
    .C(_08025_),
    .A(_09204_),
    .Y(_08026_));
 sg13g2_o21ai_1 _27329_ (.B1(_08026_),
    .Y(_08027_),
    .A1(_09204_),
    .A2(_08025_));
 sg13g2_nand2_1 _27330_ (.Y(_02536_),
    .A(net696),
    .B(_08027_));
 sg13g2_nand2_1 _27331_ (.Y(_08028_),
    .A(_09204_),
    .B(_12048_));
 sg13g2_a21oi_1 _27332_ (.A1(_08025_),
    .A2(_08028_),
    .Y(_08029_),
    .B1(_09205_));
 sg13g2_inv_1 _27333_ (.Y(_08030_),
    .A(_09204_));
 sg13g2_and4_1 _27334_ (.A(_08030_),
    .B(_09205_),
    .C(_12048_),
    .D(_08025_),
    .X(_08031_));
 sg13g2_o21ai_1 _27335_ (.B1(net696),
    .Y(_02537_),
    .A1(_08029_),
    .A2(_08031_));
 sg13g2_nor2_1 _27336_ (.A(_09204_),
    .B(_09205_),
    .Y(_08032_));
 sg13g2_or2_1 _27337_ (.X(_08033_),
    .B(_08032_),
    .A(_00219_));
 sg13g2_a21oi_1 _27338_ (.A1(_08025_),
    .A2(_08033_),
    .Y(_08034_),
    .B1(\cpu.spi.r_bits[2] ));
 sg13g2_and4_1 _27339_ (.A(\cpu.spi.r_bits[2] ),
    .B(_12048_),
    .C(_08032_),
    .D(_08025_),
    .X(_08035_));
 sg13g2_o21ai_1 _27340_ (.B1(net696),
    .Y(_02538_),
    .A1(_08034_),
    .A2(_08035_));
 sg13g2_buf_1 _27341_ (.A(\cpu.gpio.genblk1[3].srcs_o[6] ),
    .X(_08036_));
 sg13g2_inv_1 _27342_ (.Y(_08037_),
    .A(net1094));
 sg13g2_nor2b_1 _27343_ (.A(_09199_),
    .B_N(_09185_),
    .Y(_08038_));
 sg13g2_or2_1 _27344_ (.X(_08039_),
    .B(_09263_),
    .A(\cpu.spi.r_state[1] ));
 sg13g2_buf_1 _27345_ (.A(_08039_),
    .X(_08040_));
 sg13g2_nand2_1 _27346_ (.Y(_08041_),
    .A(net353),
    .B(_08040_));
 sg13g2_nor3_1 _27347_ (.A(net1150),
    .B(_09239_),
    .C(_08040_),
    .Y(_08042_));
 sg13g2_a21oi_1 _27348_ (.A1(_12051_),
    .A2(_06971_),
    .Y(_08043_),
    .B1(_09249_));
 sg13g2_nor3_1 _27349_ (.A(_00271_),
    .B(_08042_),
    .C(_08043_),
    .Y(_08044_));
 sg13g2_a21oi_1 _27350_ (.A1(_00271_),
    .A2(_08041_),
    .Y(_08045_),
    .B1(_08044_));
 sg13g2_o21ai_1 _27351_ (.B1(_08045_),
    .Y(_08046_),
    .A1(_06964_),
    .A2(_08038_));
 sg13g2_nor3_1 _27352_ (.A(_12051_),
    .B(net1032),
    .C(_08046_),
    .Y(_08047_));
 sg13g2_inv_1 _27353_ (.Y(_08048_),
    .A(_08046_));
 sg13g2_a21oi_1 _27354_ (.A1(_08040_),
    .A2(_08048_),
    .Y(_08049_),
    .B1(net815));
 sg13g2_o21ai_1 _27355_ (.B1(_08049_),
    .Y(_02571_),
    .A1(_08037_),
    .A2(_08047_));
 sg13g2_buf_1 _27356_ (.A(\cpu.gpio.genblk1[3].srcs_o[7] ),
    .X(_08050_));
 sg13g2_inv_1 _27357_ (.Y(_08051_),
    .A(net1093));
 sg13g2_nor3_1 _27358_ (.A(net772),
    .B(_12068_),
    .C(_08046_),
    .Y(_08052_));
 sg13g2_o21ai_1 _27359_ (.B1(_08049_),
    .Y(_02572_),
    .A1(_08051_),
    .A2(_08052_));
 sg13g2_buf_1 _27360_ (.A(\cpu.gpio.genblk1[3].srcs_o[8] ),
    .X(_08053_));
 sg13g2_nand3_1 _27361_ (.B(_12068_),
    .C(_08048_),
    .A(_12065_),
    .Y(_08054_));
 sg13g2_nand2_1 _27362_ (.Y(_08055_),
    .A(_08053_),
    .B(_08054_));
 sg13g2_nand2_1 _27363_ (.Y(_02573_),
    .A(_08049_),
    .B(_08055_));
 sg13g2_a21oi_1 _27364_ (.A1(_09227_),
    .A2(_09239_),
    .Y(_08056_),
    .B1(_09251_));
 sg13g2_nor3_1 _27365_ (.A(_06964_),
    .B(_09185_),
    .C(_09199_),
    .Y(_08057_));
 sg13g2_nor3_1 _27366_ (.A(_09301_),
    .B(_08056_),
    .C(_08057_),
    .Y(_08058_));
 sg13g2_o21ai_1 _27367_ (.B1(_08058_),
    .Y(_08059_),
    .A1(_12102_),
    .A2(_09265_));
 sg13g2_a22oi_1 _27368_ (.Y(_08060_),
    .B1(_08059_),
    .B2(_09119_),
    .A2(_08058_),
    .A1(net1151));
 sg13g2_nor2_1 _27369_ (.A(net583),
    .B(_08060_),
    .Y(_02582_));
 sg13g2_nor3_1 _27370_ (.A(_09203_),
    .B(_09265_),
    .C(_08040_),
    .Y(_08061_));
 sg13g2_nor2b_1 _27371_ (.A(_08061_),
    .B_N(_08058_),
    .Y(_08062_));
 sg13g2_nor2_1 _27372_ (.A(_09263_),
    .B(_09262_),
    .Y(_08063_));
 sg13g2_a22oi_1 _27373_ (.Y(_08064_),
    .B1(_08062_),
    .B2(_08063_),
    .A2(_09250_),
    .A1(_04945_));
 sg13g2_nor2_1 _27374_ (.A(net1151),
    .B(_08064_),
    .Y(_08065_));
 sg13g2_nor2_1 _27375_ (.A(\cpu.spi.r_ready ),
    .B(_08062_),
    .Y(_08066_));
 sg13g2_o21ai_1 _27376_ (.B1(net663),
    .Y(_02597_),
    .A1(_08065_),
    .A2(_08066_));
 sg13g2_nor2_1 _27377_ (.A(_06964_),
    .B(_09183_),
    .Y(_08067_));
 sg13g2_nor3_1 _27378_ (.A(_09262_),
    .B(_08023_),
    .C(_08056_),
    .Y(_08068_));
 sg13g2_mux2_1 _27379_ (.A0(\cpu.spi.r_searching ),
    .A1(_08067_),
    .S(_08068_),
    .X(_08069_));
 sg13g2_and2_1 _27380_ (.A(net680),
    .B(_08069_),
    .X(_02598_));
 sg13g2_buf_1 _27381_ (.A(_07265_),
    .X(_08070_));
 sg13g2_and2_1 _27382_ (.A(net375),
    .B(_08070_),
    .X(_08071_));
 sg13g2_buf_2 _27383_ (.A(_08071_),
    .X(_08072_));
 sg13g2_nand2_1 _27384_ (.Y(_08073_),
    .A(net841),
    .B(_08072_));
 sg13g2_nand2_1 _27385_ (.Y(_08074_),
    .A(net375),
    .B(net159));
 sg13g2_buf_2 _27386_ (.A(_08074_),
    .X(_08075_));
 sg13g2_nand2_1 _27387_ (.Y(_08076_),
    .A(\cpu.uart.r_div_value[0] ),
    .B(_08075_));
 sg13g2_nand3_1 _27388_ (.B(_08073_),
    .C(_08076_),
    .A(net663),
    .Y(_02620_));
 sg13g2_nand2_2 _27389_ (.Y(_08077_),
    .A(net409),
    .B(net159));
 sg13g2_nor2_1 _27390_ (.A(_12240_),
    .B(_08077_),
    .Y(_08078_));
 sg13g2_a21oi_1 _27391_ (.A1(\cpu.uart.r_div_value[10] ),
    .A2(_08077_),
    .Y(_08079_),
    .B1(_08078_));
 sg13g2_nor2_1 _27392_ (.A(net637),
    .B(_08079_),
    .Y(_02621_));
 sg13g2_nand3_1 _27393_ (.B(net409),
    .C(net159),
    .A(net1058),
    .Y(_08080_));
 sg13g2_nand2_1 _27394_ (.Y(_08081_),
    .A(\cpu.uart.r_div_value[11] ),
    .B(_08077_));
 sg13g2_a21oi_1 _27395_ (.A1(_08080_),
    .A2(_08081_),
    .Y(_02622_),
    .B1(net581));
 sg13g2_nand2_1 _27396_ (.Y(_08082_),
    .A(net1055),
    .B(_08072_));
 sg13g2_nand2_1 _27397_ (.Y(_08083_),
    .A(\cpu.uart.r_div_value[1] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27398_ (.A1(_08082_),
    .A2(_08083_),
    .Y(_02623_),
    .B1(net581));
 sg13g2_nand2_1 _27399_ (.Y(_08084_),
    .A(net1059),
    .B(_08072_));
 sg13g2_nand2_1 _27400_ (.Y(_08085_),
    .A(\cpu.uart.r_div_value[2] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27401_ (.A1(_08084_),
    .A2(_08085_),
    .Y(_02624_),
    .B1(net581));
 sg13g2_nand2_1 _27402_ (.Y(_08086_),
    .A(net1058),
    .B(_08072_));
 sg13g2_nand2_1 _27403_ (.Y(_08087_),
    .A(\cpu.uart.r_div_value[3] ),
    .B(_08075_));
 sg13g2_buf_1 _27404_ (.A(_09772_),
    .X(_08088_));
 sg13g2_a21oi_1 _27405_ (.A1(_08086_),
    .A2(_08087_),
    .Y(_02625_),
    .B1(net580));
 sg13g2_nand2_1 _27406_ (.Y(_08089_),
    .A(net1057),
    .B(_08072_));
 sg13g2_nand2_1 _27407_ (.Y(_08090_),
    .A(\cpu.uart.r_div_value[4] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27408_ (.A1(_08089_),
    .A2(_08090_),
    .Y(_02626_),
    .B1(net580));
 sg13g2_nand2_1 _27409_ (.Y(_08091_),
    .A(net1054),
    .B(_08072_));
 sg13g2_nand2_1 _27410_ (.Y(_08092_),
    .A(\cpu.uart.r_div_value[5] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27411_ (.A1(_08091_),
    .A2(_08092_),
    .Y(_02627_),
    .B1(net580));
 sg13g2_nand2_1 _27412_ (.Y(_08093_),
    .A(net1053),
    .B(_08072_));
 sg13g2_nand2_1 _27413_ (.Y(_08094_),
    .A(\cpu.uart.r_div_value[6] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27414_ (.A1(_08093_),
    .A2(_08094_),
    .Y(_02628_),
    .B1(net580));
 sg13g2_nand2_1 _27415_ (.Y(_08095_),
    .A(net1056),
    .B(_08072_));
 sg13g2_nand2_1 _27416_ (.Y(_08096_),
    .A(\cpu.uart.r_div_value[7] ),
    .B(_08075_));
 sg13g2_a21oi_1 _27417_ (.A1(_08095_),
    .A2(_08096_),
    .Y(_02629_),
    .B1(_08088_));
 sg13g2_nand3_1 _27418_ (.B(net409),
    .C(net159),
    .A(net960),
    .Y(_08097_));
 sg13g2_nand2_1 _27419_ (.Y(_08098_),
    .A(\cpu.uart.r_div_value[8] ),
    .B(_08077_));
 sg13g2_a21oi_1 _27420_ (.A1(_08097_),
    .A2(_08098_),
    .Y(_02630_),
    .B1(net580));
 sg13g2_nand3_1 _27421_ (.B(net409),
    .C(net159),
    .A(net1055),
    .Y(_08099_));
 sg13g2_nand2_1 _27422_ (.Y(_08100_),
    .A(\cpu.uart.r_div_value[9] ),
    .B(_08077_));
 sg13g2_a21oi_1 _27423_ (.A1(_08099_),
    .A2(_08100_),
    .Y(_02631_),
    .B1(net580));
 sg13g2_nor2_1 _27424_ (.A(_00195_),
    .B(_09163_),
    .Y(_08101_));
 sg13g2_nand2_1 _27425_ (.Y(_08102_),
    .A(net992),
    .B(net877));
 sg13g2_nand2_1 _27426_ (.Y(_08103_),
    .A(_12085_),
    .B(_07263_));
 sg13g2_nor4_1 _27427_ (.A(net1161),
    .B(net1000),
    .C(_04859_),
    .D(_08103_),
    .Y(_08104_));
 sg13g2_nand4_1 _27428_ (.B(_09181_),
    .C(_08102_),
    .A(_08101_),
    .Y(_08105_),
    .D(_08104_));
 sg13g2_nand3_1 _27429_ (.B(net408),
    .C(_08070_),
    .A(_09978_),
    .Y(_08106_));
 sg13g2_nand4_1 _27430_ (.B(net818),
    .C(_08105_),
    .A(_09115_),
    .Y(_08107_),
    .D(_08106_));
 sg13g2_nand2b_1 _27431_ (.Y(_02655_),
    .B(_08107_),
    .A_N(net188));
 sg13g2_nand3_1 _27432_ (.B(net515),
    .C(net159),
    .A(net1055),
    .Y(_08108_));
 sg13g2_nand2_1 _27433_ (.Y(_08109_),
    .A(net515),
    .B(net159));
 sg13g2_nand2_1 _27434_ (.Y(_08110_),
    .A(\cpu.uart.r_r_invert ),
    .B(_08109_));
 sg13g2_a21oi_1 _27435_ (.A1(_08108_),
    .A2(_08110_),
    .Y(_02656_),
    .B1(net580));
 sg13g2_a21oi_1 _27436_ (.A1(_07254_),
    .A2(net349),
    .Y(_08111_),
    .B1(_07248_));
 sg13g2_a21oi_1 _27437_ (.A1(_07255_),
    .A2(net349),
    .Y(_08112_),
    .B1(_07323_));
 sg13g2_a221oi_1 _27438_ (.B2(_08111_),
    .C1(_08112_),
    .B1(_07253_),
    .A1(net956),
    .Y(_08113_),
    .A2(_07248_));
 sg13g2_a21oi_1 _27439_ (.A1(_07246_),
    .A2(_08113_),
    .Y(_08114_),
    .B1(_07331_));
 sg13g2_buf_2 _27440_ (.A(_08114_),
    .X(_08115_));
 sg13g2_o21ai_1 _27441_ (.B1(_08115_),
    .Y(_08116_),
    .A1(net956),
    .A2(_07323_));
 sg13g2_xnor2_1 _27442_ (.Y(_08117_),
    .A(_07255_),
    .B(_08116_));
 sg13g2_nor2_1 _27443_ (.A(net637),
    .B(_08117_),
    .Y(_02659_));
 sg13g2_o21ai_1 _27444_ (.B1(_08115_),
    .Y(_08118_),
    .A1(_07254_),
    .A2(net957));
 sg13g2_nand2_1 _27445_ (.Y(_08119_),
    .A(net1099),
    .B(_08118_));
 sg13g2_nand2b_1 _27446_ (.Y(_08120_),
    .B(net956),
    .A_N(net957));
 sg13g2_o21ai_1 _27447_ (.B1(_08120_),
    .Y(_08121_),
    .A1(net956),
    .A2(_07332_));
 sg13g2_nand3_1 _27448_ (.B(_08115_),
    .C(_08121_),
    .A(_07333_),
    .Y(_08122_));
 sg13g2_a21oi_1 _27449_ (.A1(_08119_),
    .A2(_08122_),
    .Y(_02660_),
    .B1(_08088_));
 sg13g2_nand2_1 _27450_ (.Y(_08123_),
    .A(_07254_),
    .B(_07250_));
 sg13g2_nor3_1 _27451_ (.A(_07252_),
    .B(net957),
    .C(_08123_),
    .Y(_08124_));
 sg13g2_o21ai_1 _27452_ (.B1(_08115_),
    .Y(_08125_),
    .A1(net957),
    .A2(_07340_));
 sg13g2_a22oi_1 _27453_ (.Y(_08126_),
    .B1(_08125_),
    .B2(net956),
    .A2(_08124_),
    .A1(_08115_));
 sg13g2_nor2_1 _27454_ (.A(net637),
    .B(_08126_),
    .Y(_02661_));
 sg13g2_a21oi_1 _27455_ (.A1(_07340_),
    .A2(_08115_),
    .Y(_08127_),
    .B1(net957));
 sg13g2_nor2b_1 _27456_ (.A(_07252_),
    .B_N(net1099),
    .Y(_08128_));
 sg13g2_a21oi_1 _27457_ (.A1(_08115_),
    .A2(_08128_),
    .Y(_08129_),
    .B1(_09772_));
 sg13g2_nor2b_1 _27458_ (.A(_08127_),
    .B_N(_08129_),
    .Y(_02662_));
 sg13g2_and2_1 _27459_ (.A(_09857_),
    .B(_07281_),
    .X(_08130_));
 sg13g2_buf_1 _27460_ (.A(_08130_),
    .X(_08131_));
 sg13g2_nor2_1 _27461_ (.A(_07269_),
    .B(_07275_),
    .Y(_08132_));
 sg13g2_o21ai_1 _27462_ (.B1(net668),
    .Y(_08133_),
    .A1(_00216_),
    .A2(net604));
 sg13g2_and2_1 _27463_ (.A(net669),
    .B(_08133_),
    .X(_08134_));
 sg13g2_a22oi_1 _27464_ (.Y(_08135_),
    .B1(_08132_),
    .B2(_08134_),
    .A2(_07350_),
    .A1(_07272_));
 sg13g2_a21o_1 _27465_ (.A2(net408),
    .A1(_09968_),
    .B1(net517),
    .X(_08136_));
 sg13g2_a21oi_1 _27466_ (.A1(_07265_),
    .A2(_08136_),
    .Y(_08137_),
    .B1(_07278_));
 sg13g2_nor3_1 _27467_ (.A(_07295_),
    .B(_08135_),
    .C(_08137_),
    .Y(_08138_));
 sg13g2_a21oi_1 _27468_ (.A1(_08131_),
    .A2(_08138_),
    .Y(_08139_),
    .B1(_09114_));
 sg13g2_nand3b_1 _27469_ (.B(_07367_),
    .C(_07272_),
    .Y(_08140_),
    .A_N(_07287_));
 sg13g2_a21oi_1 _27470_ (.A1(_08138_),
    .A2(_08140_),
    .Y(_08141_),
    .B1(_09772_));
 sg13g2_nor2b_1 _27471_ (.A(_08139_),
    .B_N(_08141_),
    .Y(_02664_));
 sg13g2_nand3_1 _27472_ (.B(net515),
    .C(net159),
    .A(net960),
    .Y(_08142_));
 sg13g2_nand2_1 _27473_ (.Y(_08143_),
    .A(_04969_),
    .B(_08109_));
 sg13g2_a21oi_1 _27474_ (.A1(_08142_),
    .A2(_08143_),
    .Y(_02665_),
    .B1(net580));
 sg13g2_o21ai_1 _27475_ (.B1(_07275_),
    .Y(_08144_),
    .A1(_07278_),
    .A2(_08131_));
 sg13g2_and2_1 _27476_ (.A(_07274_),
    .B(_07382_),
    .X(_08145_));
 sg13g2_a221oi_1 _27477_ (.B2(_07283_),
    .C1(_07377_),
    .B1(_08145_),
    .A1(_07267_),
    .Y(_08146_),
    .A2(_08144_));
 sg13g2_buf_2 _27478_ (.A(_08146_),
    .X(_08147_));
 sg13g2_nand2_1 _27479_ (.Y(_08148_),
    .A(_08131_),
    .B(_07373_));
 sg13g2_nand4_1 _27480_ (.B(_07361_),
    .C(_08147_),
    .A(net954),
    .Y(_08149_),
    .D(_08148_));
 sg13g2_o21ai_1 _27481_ (.B1(_08149_),
    .Y(_08150_),
    .A1(net954),
    .A2(_08147_));
 sg13g2_nor2_1 _27482_ (.A(net637),
    .B(_08150_),
    .Y(_02668_));
 sg13g2_o21ai_1 _27483_ (.B1(_08147_),
    .Y(_08151_),
    .A1(net954),
    .A2(_07382_));
 sg13g2_nand2_1 _27484_ (.Y(_08152_),
    .A(net955),
    .B(_08151_));
 sg13g2_nand4_1 _27485_ (.B(_07287_),
    .C(_07361_),
    .A(_07358_),
    .Y(_08153_),
    .D(_08147_));
 sg13g2_a21oi_1 _27486_ (.A1(_08152_),
    .A2(_08153_),
    .Y(_02669_),
    .B1(net714));
 sg13g2_inv_1 _27487_ (.Y(_08154_),
    .A(_08147_));
 sg13g2_nand2_1 _27488_ (.Y(_08155_),
    .A(_07388_),
    .B(_08147_));
 sg13g2_nand2_1 _27489_ (.Y(_08156_),
    .A(net953),
    .B(_07387_));
 sg13g2_a21oi_1 _27490_ (.A1(_08155_),
    .A2(_08156_),
    .Y(_08157_),
    .B1(net952));
 sg13g2_a221oi_1 _27491_ (.B2(net953),
    .C1(_08157_),
    .B1(_08154_),
    .A1(_07283_),
    .Y(_08158_),
    .A2(_07373_));
 sg13g2_nor2_1 _27492_ (.A(net637),
    .B(_08158_),
    .Y(_02670_));
 sg13g2_nand2b_1 _27493_ (.Y(_08159_),
    .B(net953),
    .A_N(net952));
 sg13g2_nand2_1 _27494_ (.Y(_08160_),
    .A(_07283_),
    .B(_07373_));
 sg13g2_o21ai_1 _27495_ (.B1(_08160_),
    .Y(_08161_),
    .A1(_07387_),
    .A2(_08159_));
 sg13g2_o21ai_1 _27496_ (.B1(_08147_),
    .Y(_08162_),
    .A1(net953),
    .A2(_07277_));
 sg13g2_a22oi_1 _27497_ (.Y(_08163_),
    .B1(_08162_),
    .B2(net952),
    .A2(_08161_),
    .A1(_08147_));
 sg13g2_nor2_1 _27498_ (.A(net637),
    .B(_08163_),
    .Y(_02671_));
 sg13g2_or2_1 _27499_ (.X(\cpu.ex.genblk3.c_supmode ),
    .B(_07556_),
    .A(_07553_));
 sg13g2_and2_1 _27500_ (.A(_09811_),
    .B(_07991_),
    .X(_08164_));
 sg13g2_a22oi_1 _27501_ (.Y(_08165_),
    .B1(_09778_),
    .B2(_08164_),
    .A2(net799),
    .A1(net1149));
 sg13g2_inv_1 _27502_ (.Y(\cpu.qspi.c_rstrobe_d ),
    .A(_08165_));
 sg13g2_nor4_1 _27503_ (.A(_09770_),
    .B(_09761_),
    .C(net799),
    .D(_07990_),
    .Y(_08166_));
 sg13g2_a21oi_2 _27504_ (.B1(_09809_),
    .Y(_08167_),
    .A2(_08166_),
    .A1(_07974_));
 sg13g2_nor2_1 _27505_ (.A(net840),
    .B(_08167_),
    .Y(\cpu.qspi.c_wstrobe_d ));
 sg13g2_nor2_1 _27506_ (.A(_08245_),
    .B(_08167_),
    .Y(\cpu.qspi.c_wstrobe_i ));
 sg13g2_mux4_1 _27507_ (.S0(_04841_),
    .A0(_09149_),
    .A1(_09126_),
    .A2(_09137_),
    .A3(_09145_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08168_));
 sg13g2_mux4_1 _27508_ (.S0(_04841_),
    .A0(_09147_),
    .A1(_09128_),
    .A2(_09151_),
    .A3(_09139_),
    .S1(\cpu.gpio.r_uart_rx_src[1] ),
    .X(_08169_));
 sg13g2_mux2_1 _27509_ (.A0(_08168_),
    .A1(_08169_),
    .S(\cpu.gpio.r_uart_rx_src[2] ),
    .X(\cpu.gpio.uart_rx ));
 sg13g2_mux4_1 _27510_ (.S0(_04872_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(net1093),
    .S1(_05341_),
    .X(_08170_));
 sg13g2_mux4_1 _27511_ (.S0(_04872_),
    .A0(\cpu.gpio.genblk2[4].srcs_io[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_05341_),
    .X(_08171_));
 sg13g2_nor2b_1 _27512_ (.A(_05421_),
    .B_N(_08171_),
    .Y(_08172_));
 sg13g2_a21oi_1 _27513_ (.A1(_05421_),
    .A2(_08170_),
    .Y(_08173_),
    .B1(_08172_));
 sg13g2_nand2b_1 _27514_ (.Y(_08174_),
    .B(net1092),
    .A_N(_04872_));
 sg13g2_nand3_1 _27515_ (.B(_05341_),
    .C(net1095),
    .A(_04872_),
    .Y(_08175_));
 sg13g2_o21ai_1 _27516_ (.B1(_08175_),
    .Y(_08176_),
    .A1(_05341_),
    .A2(_08174_));
 sg13g2_nand3_1 _27517_ (.B(_00185_),
    .C(_08176_),
    .A(_05482_),
    .Y(_08177_));
 sg13g2_o21ai_1 _27518_ (.B1(_08177_),
    .Y(net15),
    .A1(_05482_),
    .A2(_08173_));
 sg13g2_mux4_1 _27519_ (.S0(_05558_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(net1093),
    .S1(_05622_),
    .X(_08178_));
 sg13g2_mux4_1 _27520_ (.S0(_05558_),
    .A0(\cpu.gpio.genblk2[5].srcs_io[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_05622_),
    .X(_08179_));
 sg13g2_nor2b_1 _27521_ (.A(_05664_),
    .B_N(_08179_),
    .Y(_08180_));
 sg13g2_a21oi_1 _27522_ (.A1(_05664_),
    .A2(_08178_),
    .Y(_08181_),
    .B1(_08180_));
 sg13g2_nand2b_1 _27523_ (.Y(_08182_),
    .B(net1092),
    .A_N(_05558_));
 sg13g2_nand3_1 _27524_ (.B(_05622_),
    .C(net1095),
    .A(_05558_),
    .Y(_08183_));
 sg13g2_o21ai_1 _27525_ (.B1(_08183_),
    .Y(_08184_),
    .A1(_05622_),
    .A2(_08182_));
 sg13g2_nand3_1 _27526_ (.B(_00184_),
    .C(_08184_),
    .A(_05078_),
    .Y(_08185_));
 sg13g2_o21ai_1 _27527_ (.B1(_08185_),
    .Y(net16),
    .A1(_05078_),
    .A2(_08181_));
 sg13g2_mux4_1 _27528_ (.S0(_04865_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(net1093),
    .S1(_06345_),
    .X(_08186_));
 sg13g2_mux4_1 _27529_ (.S0(_04865_),
    .A0(\cpu.gpio.genblk2[6].srcs_io[0] ),
    .A1(_07349_),
    .A2(net1115),
    .A3(net1116),
    .S1(_06345_),
    .X(_08187_));
 sg13g2_nor2b_1 _27530_ (.A(\cpu.gpio.r_src_io[6][2] ),
    .B_N(_08187_),
    .Y(_08188_));
 sg13g2_a21oi_1 _27531_ (.A1(\cpu.gpio.r_src_io[6][2] ),
    .A2(_08186_),
    .Y(_08189_),
    .B1(_08188_));
 sg13g2_nand2b_1 _27532_ (.Y(_08190_),
    .B(net1092),
    .A_N(_04865_));
 sg13g2_nand3_1 _27533_ (.B(net1095),
    .C(_06345_),
    .A(_04865_),
    .Y(_08191_));
 sg13g2_o21ai_1 _27534_ (.B1(_08191_),
    .Y(_08192_),
    .A1(_06345_),
    .A2(_08190_));
 sg13g2_nand3_1 _27535_ (.B(\cpu.gpio.r_src_io[6][3] ),
    .C(_08192_),
    .A(_00098_),
    .Y(_08193_));
 sg13g2_o21ai_1 _27536_ (.B1(_08193_),
    .Y(net17),
    .A1(\cpu.gpio.r_src_io[6][3] ),
    .A2(_08189_));
 sg13g2_mux4_1 _27537_ (.S0(_05557_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(_08050_),
    .S1(_06348_),
    .X(_08194_));
 sg13g2_mux4_1 _27538_ (.S0(_05557_),
    .A0(\cpu.gpio.genblk2[7].srcs_io[0] ),
    .A1(_07349_),
    .A2(net1115),
    .A3(net1116),
    .S1(_06348_),
    .X(_08195_));
 sg13g2_nor2b_1 _27539_ (.A(\cpu.gpio.r_src_io[7][2] ),
    .B_N(_08195_),
    .Y(_08196_));
 sg13g2_a21oi_1 _27540_ (.A1(\cpu.gpio.r_src_io[7][2] ),
    .A2(_08194_),
    .Y(_08197_),
    .B1(_08196_));
 sg13g2_nand2b_1 _27541_ (.Y(_08198_),
    .B(net1092),
    .A_N(_05557_));
 sg13g2_nand3_1 _27542_ (.B(net1095),
    .C(_06348_),
    .A(_05557_),
    .Y(_08199_));
 sg13g2_o21ai_1 _27543_ (.B1(_08199_),
    .Y(_08200_),
    .A1(_06348_),
    .A2(_08198_));
 sg13g2_nand3_1 _27544_ (.B(\cpu.gpio.r_src_io[7][3] ),
    .C(_08200_),
    .A(_00139_),
    .Y(_08201_));
 sg13g2_o21ai_1 _27545_ (.B1(_08201_),
    .Y(net18),
    .A1(\cpu.gpio.r_src_io[7][3] ),
    .A2(_08197_));
 sg13g2_xor2_1 _27546_ (.B(clknet_leaf_75_clk),
    .A(\cpu.r_clk_invert ),
    .X(net21));
 sg13g2_mux4_1 _27547_ (.S0(_05567_),
    .A0(net1117),
    .A1(net1118),
    .A2(_08036_),
    .A3(_08050_),
    .S1(_06354_),
    .X(_08202_));
 sg13g2_mux4_1 _27548_ (.S0(_05567_),
    .A0(\cpu.gpio.genblk1[3].srcs_o[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_06354_),
    .X(_08203_));
 sg13g2_nor2b_1 _27549_ (.A(\cpu.gpio.r_src_o[3][2] ),
    .B_N(_08203_),
    .Y(_08204_));
 sg13g2_a21oi_1 _27550_ (.A1(\cpu.gpio.r_src_o[3][2] ),
    .A2(_08202_),
    .Y(_08205_),
    .B1(_08204_));
 sg13g2_nand2b_1 _27551_ (.Y(_08206_),
    .B(net1092),
    .A_N(_05567_));
 sg13g2_nand3_1 _27552_ (.B(net1095),
    .C(_06354_),
    .A(_05567_),
    .Y(_08207_));
 sg13g2_o21ai_1 _27553_ (.B1(_08207_),
    .Y(_08208_),
    .A1(_06354_),
    .A2(_08206_));
 sg13g2_nand3_1 _27554_ (.B(\cpu.gpio.r_src_o[3][3] ),
    .C(_08208_),
    .A(_00142_),
    .Y(_08209_));
 sg13g2_o21ai_1 _27555_ (.B1(_08209_),
    .Y(net22),
    .A1(\cpu.gpio.r_src_o[3][3] ),
    .A2(_08205_));
 sg13g2_mux4_1 _27556_ (.S0(_04858_),
    .A0(_12100_),
    .A1(net1118),
    .A2(_08036_),
    .A3(net1093),
    .S1(_06362_),
    .X(_08210_));
 sg13g2_mux4_1 _27557_ (.S0(_04858_),
    .A0(\cpu.gpio.genblk1[4].srcs_o[0] ),
    .A1(net1096),
    .A2(_12120_),
    .A3(_12104_),
    .S1(_06362_),
    .X(_08211_));
 sg13g2_nor2b_1 _27558_ (.A(\cpu.gpio.r_src_o[4][2] ),
    .B_N(_08211_),
    .Y(_08212_));
 sg13g2_a21oi_1 _27559_ (.A1(\cpu.gpio.r_src_o[4][2] ),
    .A2(_08210_),
    .Y(_08213_),
    .B1(_08212_));
 sg13g2_nand2b_1 _27560_ (.Y(_08214_),
    .B(net1092),
    .A_N(_04858_));
 sg13g2_nand3_1 _27561_ (.B(net1095),
    .C(_06362_),
    .A(_04858_),
    .Y(_08215_));
 sg13g2_o21ai_1 _27562_ (.B1(_08215_),
    .Y(_08216_),
    .A1(_06362_),
    .A2(_08214_));
 sg13g2_nand3_1 _27563_ (.B(\cpu.gpio.r_src_o[4][3] ),
    .C(_08216_),
    .A(_00100_),
    .Y(_08217_));
 sg13g2_o21ai_1 _27564_ (.B1(_08217_),
    .Y(net23),
    .A1(\cpu.gpio.r_src_o[4][3] ),
    .A2(_08213_));
 sg13g2_mux4_1 _27565_ (.S0(_05561_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(net1093),
    .S1(_06365_),
    .X(_08218_));
 sg13g2_mux4_1 _27566_ (.S0(_05561_),
    .A0(\cpu.gpio.genblk1[5].srcs_o[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_06365_),
    .X(_08219_));
 sg13g2_nor2b_1 _27567_ (.A(\cpu.gpio.r_src_o[5][2] ),
    .B_N(_08219_),
    .Y(_08220_));
 sg13g2_a21oi_1 _27568_ (.A1(\cpu.gpio.r_src_o[5][2] ),
    .A2(_08218_),
    .Y(_08221_),
    .B1(_08220_));
 sg13g2_nand2b_1 _27569_ (.Y(_08222_),
    .B(_08053_),
    .A_N(_05561_));
 sg13g2_nand3_1 _27570_ (.B(net1095),
    .C(_06365_),
    .A(_05561_),
    .Y(_08223_));
 sg13g2_o21ai_1 _27571_ (.B1(_08223_),
    .Y(_08224_),
    .A1(_06365_),
    .A2(_08222_));
 sg13g2_nand3_1 _27572_ (.B(\cpu.gpio.r_src_o[5][3] ),
    .C(_08224_),
    .A(_00141_),
    .Y(_08225_));
 sg13g2_o21ai_1 _27573_ (.B1(_08225_),
    .Y(net24),
    .A1(\cpu.gpio.r_src_o[5][3] ),
    .A2(_08221_));
 sg13g2_mux4_1 _27574_ (.S0(_04853_),
    .A0(net1117),
    .A1(net1118),
    .A2(net1094),
    .A3(net1093),
    .S1(_07893_),
    .X(_08226_));
 sg13g2_mux4_1 _27575_ (.S0(_04853_),
    .A0(\cpu.gpio.genblk1[6].srcs_o[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_07893_),
    .X(_08227_));
 sg13g2_nor2b_1 _27576_ (.A(\cpu.gpio.r_src_o[6][2] ),
    .B_N(_08227_),
    .Y(_08228_));
 sg13g2_a21oi_1 _27577_ (.A1(\cpu.gpio.r_src_o[6][2] ),
    .A2(_08226_),
    .Y(_08229_),
    .B1(_08228_));
 sg13g2_nand2b_1 _27578_ (.Y(_08230_),
    .B(net1092),
    .A_N(_04853_));
 sg13g2_nand3_1 _27579_ (.B(net1095),
    .C(_07893_),
    .A(_04853_),
    .Y(_08231_));
 sg13g2_o21ai_1 _27580_ (.B1(_08231_),
    .Y(_08232_),
    .A1(_07893_),
    .A2(_08230_));
 sg13g2_nand3_1 _27581_ (.B(\cpu.gpio.r_src_o[6][3] ),
    .C(_08232_),
    .A(_00099_),
    .Y(_08233_));
 sg13g2_o21ai_1 _27582_ (.B1(_08233_),
    .Y(net25),
    .A1(\cpu.gpio.r_src_o[6][3] ),
    .A2(_08229_));
 sg13g2_mux4_1 _27583_ (.S0(_05559_),
    .A0(net1117),
    .A1(_12094_),
    .A2(net1094),
    .A3(net1093),
    .S1(_06371_),
    .X(_08234_));
 sg13g2_mux4_1 _27584_ (.S0(_05559_),
    .A0(\cpu.gpio.genblk1[7].srcs_o[0] ),
    .A1(net1096),
    .A2(net1115),
    .A3(net1116),
    .S1(_06371_),
    .X(_08235_));
 sg13g2_nor2b_1 _27585_ (.A(\cpu.gpio.r_src_o[7][2] ),
    .B_N(_08235_),
    .Y(_08236_));
 sg13g2_a21oi_1 _27586_ (.A1(\cpu.gpio.r_src_o[7][2] ),
    .A2(_08234_),
    .Y(_08237_),
    .B1(_08236_));
 sg13g2_nand2b_1 _27587_ (.Y(_08238_),
    .B(net1092),
    .A_N(_05559_));
 sg13g2_nand3_1 _27588_ (.B(_07987_),
    .C(_06371_),
    .A(_05559_),
    .Y(_08239_));
 sg13g2_o21ai_1 _27589_ (.B1(_08239_),
    .Y(_08240_),
    .A1(_06371_),
    .A2(_08238_));
 sg13g2_nand3_1 _27590_ (.B(\cpu.gpio.r_src_o[7][3] ),
    .C(_08240_),
    .A(_00140_),
    .Y(_08241_));
 sg13g2_o21ai_1 _27591_ (.B1(_08241_),
    .Y(net26),
    .A1(\cpu.gpio.r_src_o[7][3] ),
    .A2(_08237_));
 sg13g2_dfrbp_1 _27592_ (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1167),
    .D(_00308_),
    .Q_N(_14919_),
    .Q(\cpu.intr.r_swi ));
 sg13g2_dfrbp_1 _27593_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1168),
    .D(_00309_),
    .Q_N(_14918_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[5] ));
 sg13g2_dfrbp_1 _27594_ (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1169),
    .D(_00310_),
    .Q_N(_14917_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[4] ));
 sg13g2_dfrbp_1 _27595_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1170),
    .D(_00311_),
    .Q_N(_14916_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[3] ));
 sg13g2_dfrbp_1 _27596_ (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1171),
    .D(_00312_),
    .Q_N(_14915_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[2] ));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_buf_1 _27598_ (.A(net6),
    .X(net4));
 sg13g2_buf_1 _27599_ (.A(net6),
    .X(net5));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1172),
    .D(_00313_),
    .Q_N(_14914_),
    .Q(\cpu.dcache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1173),
    .D(_00314_),
    .Q_N(_00095_),
    .Q(\cpu.dcache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1174),
    .D(_00315_),
    .Q_N(_00106_),
    .Q(\cpu.dcache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1175),
    .D(_00316_),
    .Q_N(_00117_),
    .Q(\cpu.dcache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1176),
    .D(_00317_),
    .Q_N(_00124_),
    .Q(\cpu.dcache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1177),
    .D(_00318_),
    .Q_N(_00136_),
    .Q(\cpu.dcache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1178),
    .D(_00319_),
    .Q_N(_00148_),
    .Q(\cpu.dcache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1179),
    .D(_00320_),
    .Q_N(_14913_),
    .Q(\cpu.dcache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1180),
    .D(_00321_),
    .Q_N(_00296_),
    .Q(\cpu.dcache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1181),
    .D(_00322_),
    .Q_N(_00093_),
    .Q(\cpu.dcache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1182),
    .D(_00323_),
    .Q_N(_00104_),
    .Q(\cpu.dcache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1183),
    .D(_00324_),
    .Q_N(_14912_),
    .Q(\cpu.dcache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1184),
    .D(_00325_),
    .Q_N(_00115_),
    .Q(\cpu.dcache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1185),
    .D(_00326_),
    .Q_N(_00122_),
    .Q(\cpu.dcache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1186),
    .D(_00327_),
    .Q_N(_00134_),
    .Q(\cpu.dcache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1187),
    .D(_00328_),
    .Q_N(_00146_),
    .Q(\cpu.dcache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1188),
    .D(_00329_),
    .Q_N(_00292_),
    .Q(\cpu.dcache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1189),
    .D(_00330_),
    .Q_N(_00297_),
    .Q(\cpu.dcache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1190),
    .D(_00331_),
    .Q_N(_00094_),
    .Q(\cpu.dcache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1191),
    .D(_00332_),
    .Q_N(_00105_),
    .Q(\cpu.dcache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1192),
    .D(_00333_),
    .Q_N(_00116_),
    .Q(\cpu.dcache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1193),
    .D(_00334_),
    .Q_N(_00123_),
    .Q(\cpu.dcache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1194),
    .D(_00335_),
    .Q_N(_14911_),
    .Q(\cpu.dcache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1195),
    .D(_00336_),
    .Q_N(_00135_),
    .Q(\cpu.dcache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1196),
    .D(_00337_),
    .Q_N(_00147_),
    .Q(\cpu.dcache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1197),
    .D(_00338_),
    .Q_N(_14910_),
    .Q(\cpu.dcache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1198),
    .D(_00339_),
    .Q_N(_00114_),
    .Q(\cpu.dcache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1199),
    .D(_00340_),
    .Q_N(_00121_),
    .Q(\cpu.dcache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1200),
    .D(_00341_),
    .Q_N(_00133_),
    .Q(\cpu.dcache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1201),
    .D(_00342_),
    .Q_N(_00145_),
    .Q(\cpu.dcache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1202),
    .D(_00343_),
    .Q_N(_00293_),
    .Q(\cpu.dcache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1203),
    .D(_00344_),
    .Q_N(_00298_),
    .Q(\cpu.dcache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1204),
    .D(_00345_),
    .Q_N(_14909_),
    .Q(\cpu.dcache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1205),
    .D(_00346_),
    .Q_N(_14908_),
    .Q(\cpu.dcache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1206),
    .D(_00347_),
    .Q_N(_14907_),
    .Q(\cpu.dcache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1207),
    .D(_00348_),
    .Q_N(_14906_),
    .Q(\cpu.dcache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1208),
    .D(_00349_),
    .Q_N(_14905_),
    .Q(\cpu.dcache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1209),
    .D(_00350_),
    .Q_N(_14904_),
    .Q(\cpu.dcache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1210),
    .D(_00351_),
    .Q_N(_14903_),
    .Q(\cpu.dcache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1211),
    .D(_00352_),
    .Q_N(_14902_),
    .Q(\cpu.dcache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1212),
    .D(_00353_),
    .Q_N(_14901_),
    .Q(\cpu.dcache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1213),
    .D(_00354_),
    .Q_N(_14900_),
    .Q(\cpu.dcache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1214),
    .D(_00355_),
    .Q_N(_14899_),
    .Q(\cpu.dcache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1215),
    .D(_00356_),
    .Q_N(_14898_),
    .Q(\cpu.dcache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1216),
    .D(_00357_),
    .Q_N(_14897_),
    .Q(\cpu.dcache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1217),
    .D(_00358_),
    .Q_N(_14896_),
    .Q(\cpu.dcache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1218),
    .D(_00359_),
    .Q_N(_14895_),
    .Q(\cpu.dcache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1219),
    .D(_00360_),
    .Q_N(_14894_),
    .Q(\cpu.dcache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1220),
    .D(_00361_),
    .Q_N(_14893_),
    .Q(\cpu.dcache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1221),
    .D(_00362_),
    .Q_N(_14892_),
    .Q(\cpu.dcache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1222),
    .D(_00363_),
    .Q_N(_14891_),
    .Q(\cpu.dcache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1223),
    .D(_00364_),
    .Q_N(_14890_),
    .Q(\cpu.dcache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1224),
    .D(_00365_),
    .Q_N(_14889_),
    .Q(\cpu.dcache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1225),
    .D(_00366_),
    .Q_N(_14888_),
    .Q(\cpu.dcache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1226),
    .D(_00367_),
    .Q_N(_14887_),
    .Q(\cpu.dcache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1227),
    .D(_00368_),
    .Q_N(_14886_),
    .Q(\cpu.dcache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1228),
    .D(_00369_),
    .Q_N(_14885_),
    .Q(\cpu.dcache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1229),
    .D(_00370_),
    .Q_N(_14884_),
    .Q(\cpu.dcache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1230),
    .D(_00371_),
    .Q_N(_14883_),
    .Q(\cpu.dcache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1231),
    .D(_00372_),
    .Q_N(_14882_),
    .Q(\cpu.dcache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1232),
    .D(_00373_),
    .Q_N(_14881_),
    .Q(\cpu.dcache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1233),
    .D(_00374_),
    .Q_N(_14880_),
    .Q(\cpu.dcache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1234),
    .D(_00375_),
    .Q_N(_14879_),
    .Q(\cpu.dcache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1235),
    .D(_00376_),
    .Q_N(_14878_),
    .Q(\cpu.dcache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1236),
    .D(_00377_),
    .Q_N(_14877_),
    .Q(\cpu.dcache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1237),
    .D(_00378_),
    .Q_N(_14876_),
    .Q(\cpu.dcache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1238),
    .D(_00379_),
    .Q_N(_14875_),
    .Q(\cpu.dcache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1239),
    .D(_00380_),
    .Q_N(_14874_),
    .Q(\cpu.dcache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1240),
    .D(_00381_),
    .Q_N(_14873_),
    .Q(\cpu.dcache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1241),
    .D(_00382_),
    .Q_N(_14872_),
    .Q(\cpu.dcache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1242),
    .D(_00383_),
    .Q_N(_14871_),
    .Q(\cpu.dcache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1243),
    .D(_00384_),
    .Q_N(_14870_),
    .Q(\cpu.dcache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1244),
    .D(_00385_),
    .Q_N(_14869_),
    .Q(\cpu.dcache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1245),
    .D(_00386_),
    .Q_N(_14868_),
    .Q(\cpu.dcache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1246),
    .D(_00387_),
    .Q_N(_14867_),
    .Q(\cpu.dcache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1247),
    .D(_00388_),
    .Q_N(_14866_),
    .Q(\cpu.dcache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1248),
    .D(_00389_),
    .Q_N(_14865_),
    .Q(\cpu.dcache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1249),
    .D(_00390_),
    .Q_N(_14864_),
    .Q(\cpu.dcache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1250),
    .D(_00391_),
    .Q_N(_14863_),
    .Q(\cpu.dcache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1251),
    .D(_00392_),
    .Q_N(_14862_),
    .Q(\cpu.dcache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1252),
    .D(_00393_),
    .Q_N(_14861_),
    .Q(\cpu.dcache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1253),
    .D(_00394_),
    .Q_N(_14860_),
    .Q(\cpu.dcache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1254),
    .D(_00395_),
    .Q_N(_14859_),
    .Q(\cpu.dcache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1255),
    .D(_00396_),
    .Q_N(_14858_),
    .Q(\cpu.dcache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1256),
    .D(_00397_),
    .Q_N(_14857_),
    .Q(\cpu.dcache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1257),
    .D(_00398_),
    .Q_N(_14856_),
    .Q(\cpu.dcache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1258),
    .D(_00399_),
    .Q_N(_14855_),
    .Q(\cpu.dcache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1259),
    .D(_00400_),
    .Q_N(_14854_),
    .Q(\cpu.dcache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1260),
    .D(_00401_),
    .Q_N(_14853_),
    .Q(\cpu.dcache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1261),
    .D(_00402_),
    .Q_N(_14852_),
    .Q(\cpu.dcache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1262),
    .D(_00403_),
    .Q_N(_14851_),
    .Q(\cpu.dcache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1263),
    .D(_00404_),
    .Q_N(_14850_),
    .Q(\cpu.dcache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1264),
    .D(_00405_),
    .Q_N(_14849_),
    .Q(\cpu.dcache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1265),
    .D(_00406_),
    .Q_N(_14848_),
    .Q(\cpu.dcache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1266),
    .D(_00407_),
    .Q_N(_14847_),
    .Q(\cpu.dcache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1267),
    .D(_00408_),
    .Q_N(_14846_),
    .Q(\cpu.dcache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1268),
    .D(_00409_),
    .Q_N(_14845_),
    .Q(\cpu.dcache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1269),
    .D(_00410_),
    .Q_N(_14844_),
    .Q(\cpu.dcache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1270),
    .D(_00411_),
    .Q_N(_14843_),
    .Q(\cpu.dcache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1271),
    .D(_00412_),
    .Q_N(_14842_),
    .Q(\cpu.dcache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1272),
    .D(_00413_),
    .Q_N(_14841_),
    .Q(\cpu.dcache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1273),
    .D(_00414_),
    .Q_N(_14840_),
    .Q(\cpu.dcache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1274),
    .D(_00415_),
    .Q_N(_14839_),
    .Q(\cpu.dcache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1275),
    .D(_00416_),
    .Q_N(_14838_),
    .Q(\cpu.dcache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1276),
    .D(_00417_),
    .Q_N(_14837_),
    .Q(\cpu.dcache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1277),
    .D(_00418_),
    .Q_N(_14836_),
    .Q(\cpu.dcache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1278),
    .D(_00419_),
    .Q_N(_14835_),
    .Q(\cpu.dcache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1279),
    .D(_00420_),
    .Q_N(_14834_),
    .Q(\cpu.dcache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1280),
    .D(_00421_),
    .Q_N(_14833_),
    .Q(\cpu.dcache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1281),
    .D(_00422_),
    .Q_N(_14832_),
    .Q(\cpu.dcache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1282),
    .D(_00423_),
    .Q_N(_14831_),
    .Q(\cpu.dcache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1283),
    .D(_00424_),
    .Q_N(_14830_),
    .Q(\cpu.dcache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1284),
    .D(_00425_),
    .Q_N(_14829_),
    .Q(\cpu.dcache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1285),
    .D(_00426_),
    .Q_N(_14828_),
    .Q(\cpu.dcache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1286),
    .D(_00427_),
    .Q_N(_14827_),
    .Q(\cpu.dcache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1287),
    .D(_00428_),
    .Q_N(_14826_),
    .Q(\cpu.dcache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1288),
    .D(_00429_),
    .Q_N(_14825_),
    .Q(\cpu.dcache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1289),
    .D(_00430_),
    .Q_N(_14824_),
    .Q(\cpu.dcache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1290),
    .D(_00431_),
    .Q_N(_14823_),
    .Q(\cpu.dcache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1291),
    .D(_00432_),
    .Q_N(_14822_),
    .Q(\cpu.dcache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1292),
    .D(_00433_),
    .Q_N(_14821_),
    .Q(\cpu.dcache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1293),
    .D(_00434_),
    .Q_N(_14820_),
    .Q(\cpu.dcache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1294),
    .D(_00435_),
    .Q_N(_14819_),
    .Q(\cpu.dcache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1295),
    .D(_00436_),
    .Q_N(_14818_),
    .Q(\cpu.dcache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1296),
    .D(_00437_),
    .Q_N(_14817_),
    .Q(\cpu.dcache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1297),
    .D(_00438_),
    .Q_N(_14816_),
    .Q(\cpu.dcache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1298),
    .D(_00439_),
    .Q_N(_14815_),
    .Q(\cpu.dcache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1299),
    .D(_00440_),
    .Q_N(_14814_),
    .Q(\cpu.dcache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1300),
    .D(_00441_),
    .Q_N(_14813_),
    .Q(\cpu.dcache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1301),
    .D(_00442_),
    .Q_N(_14812_),
    .Q(\cpu.dcache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1302),
    .D(_00443_),
    .Q_N(_14811_),
    .Q(\cpu.dcache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1303),
    .D(_00444_),
    .Q_N(_14810_),
    .Q(\cpu.dcache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1304),
    .D(_00445_),
    .Q_N(_14809_),
    .Q(\cpu.dcache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1305),
    .D(_00446_),
    .Q_N(_14808_),
    .Q(\cpu.dcache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1306),
    .D(_00447_),
    .Q_N(_14807_),
    .Q(\cpu.dcache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1307),
    .D(_00448_),
    .Q_N(_14806_),
    .Q(\cpu.dcache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1308),
    .D(_00449_),
    .Q_N(_14805_),
    .Q(\cpu.dcache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1309),
    .D(_00450_),
    .Q_N(_14804_),
    .Q(\cpu.dcache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1310),
    .D(_00451_),
    .Q_N(_14803_),
    .Q(\cpu.dcache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1311),
    .D(_00452_),
    .Q_N(_14802_),
    .Q(\cpu.dcache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1312),
    .D(_00453_),
    .Q_N(_14801_),
    .Q(\cpu.dcache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1313),
    .D(_00454_),
    .Q_N(_14800_),
    .Q(\cpu.dcache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1314),
    .D(_00455_),
    .Q_N(_14799_),
    .Q(\cpu.dcache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1315),
    .D(_00456_),
    .Q_N(_14798_),
    .Q(\cpu.dcache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1316),
    .D(_00457_),
    .Q_N(_14797_),
    .Q(\cpu.dcache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1317),
    .D(_00458_),
    .Q_N(_14796_),
    .Q(\cpu.dcache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1318),
    .D(_00459_),
    .Q_N(_14795_),
    .Q(\cpu.dcache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1319),
    .D(_00460_),
    .Q_N(_14794_),
    .Q(\cpu.dcache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1320),
    .D(_00461_),
    .Q_N(_14793_),
    .Q(\cpu.dcache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1321),
    .D(_00462_),
    .Q_N(_14792_),
    .Q(\cpu.dcache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1322),
    .D(_00463_),
    .Q_N(_14791_),
    .Q(\cpu.dcache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1323),
    .D(_00464_),
    .Q_N(_14790_),
    .Q(\cpu.dcache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1324),
    .D(_00465_),
    .Q_N(_14789_),
    .Q(\cpu.dcache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1325),
    .D(_00466_),
    .Q_N(_14788_),
    .Q(\cpu.dcache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1326),
    .D(_00467_),
    .Q_N(_14787_),
    .Q(\cpu.dcache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1327),
    .D(_00468_),
    .Q_N(_14786_),
    .Q(\cpu.dcache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1328),
    .D(_00469_),
    .Q_N(_14785_),
    .Q(\cpu.dcache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1329),
    .D(_00470_),
    .Q_N(_14784_),
    .Q(\cpu.dcache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1330),
    .D(_00471_),
    .Q_N(_14783_),
    .Q(\cpu.dcache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1331),
    .D(_00472_),
    .Q_N(_14782_),
    .Q(\cpu.dcache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1332),
    .D(_00473_),
    .Q_N(_14781_),
    .Q(\cpu.dcache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1333),
    .D(_00474_),
    .Q_N(_14780_),
    .Q(\cpu.dcache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1334),
    .D(_00475_),
    .Q_N(_14779_),
    .Q(\cpu.dcache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1335),
    .D(_00476_),
    .Q_N(_14778_),
    .Q(\cpu.dcache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1336),
    .D(_00477_),
    .Q_N(_14777_),
    .Q(\cpu.dcache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1337),
    .D(_00478_),
    .Q_N(_14776_),
    .Q(\cpu.dcache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1338),
    .D(_00479_),
    .Q_N(_14775_),
    .Q(\cpu.dcache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1339),
    .D(_00480_),
    .Q_N(_14774_),
    .Q(\cpu.dcache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1340),
    .D(_00481_),
    .Q_N(_14773_),
    .Q(\cpu.dcache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1341),
    .D(_00482_),
    .Q_N(_14772_),
    .Q(\cpu.dcache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1342),
    .D(_00483_),
    .Q_N(_14771_),
    .Q(\cpu.dcache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1343),
    .D(_00484_),
    .Q_N(_14770_),
    .Q(\cpu.dcache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1344),
    .D(_00485_),
    .Q_N(_14769_),
    .Q(\cpu.dcache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1345),
    .D(_00486_),
    .Q_N(_14768_),
    .Q(\cpu.dcache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1346),
    .D(_00487_),
    .Q_N(_14767_),
    .Q(\cpu.dcache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1347),
    .D(_00488_),
    .Q_N(_14766_),
    .Q(\cpu.dcache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1348),
    .D(_00489_),
    .Q_N(_14765_),
    .Q(\cpu.dcache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1349),
    .D(_00490_),
    .Q_N(_14764_),
    .Q(\cpu.dcache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1350),
    .D(_00491_),
    .Q_N(_14763_),
    .Q(\cpu.dcache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1351),
    .D(_00492_),
    .Q_N(_14762_),
    .Q(\cpu.dcache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1352),
    .D(_00493_),
    .Q_N(_14761_),
    .Q(\cpu.dcache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1353),
    .D(_00494_),
    .Q_N(_14760_),
    .Q(\cpu.dcache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1354),
    .D(_00495_),
    .Q_N(_14759_),
    .Q(\cpu.dcache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1355),
    .D(_00496_),
    .Q_N(_14758_),
    .Q(\cpu.dcache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1356),
    .D(_00497_),
    .Q_N(_14757_),
    .Q(\cpu.dcache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1357),
    .D(_00498_),
    .Q_N(_14756_),
    .Q(\cpu.dcache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1358),
    .D(_00499_),
    .Q_N(_14755_),
    .Q(\cpu.dcache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1359),
    .D(_00500_),
    .Q_N(_14754_),
    .Q(\cpu.dcache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net1360),
    .D(_00501_),
    .Q_N(_14753_),
    .Q(\cpu.dcache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net1361),
    .D(_00502_),
    .Q_N(_14752_),
    .Q(\cpu.dcache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1362),
    .D(_00503_),
    .Q_N(_14751_),
    .Q(\cpu.dcache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1363),
    .D(_00504_),
    .Q_N(_14750_),
    .Q(\cpu.dcache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1364),
    .D(_00505_),
    .Q_N(_14749_),
    .Q(\cpu.dcache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1365),
    .D(_00506_),
    .Q_N(_14748_),
    .Q(\cpu.dcache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1366),
    .D(_00507_),
    .Q_N(_14747_),
    .Q(\cpu.dcache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1367),
    .D(_00508_),
    .Q_N(_14746_),
    .Q(\cpu.dcache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1368),
    .D(_00509_),
    .Q_N(_14745_),
    .Q(\cpu.dcache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1369),
    .D(_00510_),
    .Q_N(_14744_),
    .Q(\cpu.dcache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1370),
    .D(_00511_),
    .Q_N(_14743_),
    .Q(\cpu.dcache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1371),
    .D(_00512_),
    .Q_N(_14742_),
    .Q(\cpu.dcache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1372),
    .D(_00513_),
    .Q_N(_14741_),
    .Q(\cpu.dcache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1373),
    .D(_00514_),
    .Q_N(_14740_),
    .Q(\cpu.dcache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1374),
    .D(_00515_),
    .Q_N(_14739_),
    .Q(\cpu.dcache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1375),
    .D(_00516_),
    .Q_N(_14738_),
    .Q(\cpu.dcache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1376),
    .D(_00517_),
    .Q_N(_14737_),
    .Q(\cpu.dcache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1377),
    .D(_00518_),
    .Q_N(_14736_),
    .Q(\cpu.dcache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1378),
    .D(_00519_),
    .Q_N(_14735_),
    .Q(\cpu.dcache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1379),
    .D(_00520_),
    .Q_N(_14734_),
    .Q(\cpu.dcache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1380),
    .D(_00521_),
    .Q_N(_14733_),
    .Q(\cpu.dcache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1381),
    .D(_00522_),
    .Q_N(_14732_),
    .Q(\cpu.dcache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1382),
    .D(_00523_),
    .Q_N(_14731_),
    .Q(\cpu.dcache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1383),
    .D(_00524_),
    .Q_N(_14730_),
    .Q(\cpu.dcache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1384),
    .D(_00525_),
    .Q_N(_14729_),
    .Q(\cpu.dcache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1385),
    .D(_00526_),
    .Q_N(_14728_),
    .Q(\cpu.dcache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1386),
    .D(_00527_),
    .Q_N(_14727_),
    .Q(\cpu.dcache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1387),
    .D(_00528_),
    .Q_N(_14726_),
    .Q(\cpu.dcache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1388),
    .D(_00529_),
    .Q_N(_14725_),
    .Q(\cpu.dcache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1389),
    .D(_00530_),
    .Q_N(_14724_),
    .Q(\cpu.dcache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1390),
    .D(_00531_),
    .Q_N(_14723_),
    .Q(\cpu.dcache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1391),
    .D(_00532_),
    .Q_N(_14722_),
    .Q(\cpu.dcache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1392),
    .D(_00533_),
    .Q_N(_14721_),
    .Q(\cpu.dcache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1393),
    .D(_00534_),
    .Q_N(_14720_),
    .Q(\cpu.dcache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1394),
    .D(_00535_),
    .Q_N(_14719_),
    .Q(\cpu.dcache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1395),
    .D(_00536_),
    .Q_N(_14718_),
    .Q(\cpu.dcache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1396),
    .D(_00537_),
    .Q_N(_14717_),
    .Q(\cpu.dcache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1397),
    .D(_00538_),
    .Q_N(_14716_),
    .Q(\cpu.dcache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1398),
    .D(_00539_),
    .Q_N(_14715_),
    .Q(\cpu.dcache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1399),
    .D(_00540_),
    .Q_N(_14714_),
    .Q(\cpu.dcache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1400),
    .D(_00541_),
    .Q_N(_14713_),
    .Q(\cpu.dcache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1401),
    .D(_00542_),
    .Q_N(_14712_),
    .Q(\cpu.dcache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1402),
    .D(_00543_),
    .Q_N(_14711_),
    .Q(\cpu.dcache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1403),
    .D(_00544_),
    .Q_N(_14710_),
    .Q(\cpu.dcache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1404),
    .D(_00545_),
    .Q_N(_14709_),
    .Q(\cpu.dcache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1405),
    .D(_00546_),
    .Q_N(_14708_),
    .Q(\cpu.dcache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1406),
    .D(_00547_),
    .Q_N(_14707_),
    .Q(\cpu.dcache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1407),
    .D(_00548_),
    .Q_N(_14706_),
    .Q(\cpu.dcache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1408),
    .D(_00549_),
    .Q_N(_14705_),
    .Q(\cpu.dcache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1409),
    .D(_00550_),
    .Q_N(_14704_),
    .Q(\cpu.dcache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1410),
    .D(_00551_),
    .Q_N(_14703_),
    .Q(\cpu.dcache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1411),
    .D(_00552_),
    .Q_N(_14702_),
    .Q(\cpu.dcache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1412),
    .D(_00553_),
    .Q_N(_14701_),
    .Q(\cpu.dcache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1413),
    .D(_00554_),
    .Q_N(_14700_),
    .Q(\cpu.dcache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1414),
    .D(_00555_),
    .Q_N(_14699_),
    .Q(\cpu.dcache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1415),
    .D(_00556_),
    .Q_N(_14698_),
    .Q(\cpu.dcache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1416),
    .D(_00557_),
    .Q_N(_14697_),
    .Q(\cpu.dcache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1417),
    .D(_00558_),
    .Q_N(_14696_),
    .Q(\cpu.dcache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1418),
    .D(_00559_),
    .Q_N(_14695_),
    .Q(\cpu.dcache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1419),
    .D(_00560_),
    .Q_N(_14694_),
    .Q(\cpu.dcache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1420),
    .D(_00561_),
    .Q_N(_14693_),
    .Q(\cpu.dcache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1421),
    .D(_00562_),
    .Q_N(_14692_),
    .Q(\cpu.dcache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1422),
    .D(_00563_),
    .Q_N(_14691_),
    .Q(\cpu.dcache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1423),
    .D(_00564_),
    .Q_N(_14690_),
    .Q(\cpu.dcache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1424),
    .D(_00565_),
    .Q_N(_14689_),
    .Q(\cpu.dcache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1425),
    .D(_00566_),
    .Q_N(_14688_),
    .Q(\cpu.dcache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1426),
    .D(_00567_),
    .Q_N(_14687_),
    .Q(\cpu.dcache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1427),
    .D(_00568_),
    .Q_N(_14686_),
    .Q(\cpu.dcache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1428),
    .D(_00569_),
    .Q_N(_14685_),
    .Q(\cpu.dcache.r_dirty[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1429),
    .D(_00570_),
    .Q_N(_14684_),
    .Q(\cpu.dcache.r_dirty[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1430),
    .D(_00571_),
    .Q_N(_14683_),
    .Q(\cpu.dcache.r_dirty[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1431),
    .D(_00572_),
    .Q_N(_14682_),
    .Q(\cpu.dcache.r_dirty[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1432),
    .D(_00573_),
    .Q_N(_14681_),
    .Q(\cpu.dcache.r_dirty[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1433),
    .D(_00574_),
    .Q_N(_14680_),
    .Q(\cpu.dcache.r_dirty[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1434),
    .D(_00575_),
    .Q_N(_14679_),
    .Q(\cpu.dcache.r_dirty[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1435),
    .D(_00576_),
    .Q_N(_14678_),
    .Q(\cpu.dcache.r_dirty[7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1436),
    .D(_00577_),
    .Q_N(_00306_),
    .Q(\cpu.dcache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1437),
    .D(_00578_),
    .Q_N(_14677_),
    .Q(\cpu.dcache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1438),
    .D(_00579_),
    .Q_N(_00269_),
    .Q(\cpu.dcache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1439),
    .D(_00580_),
    .Q_N(_00222_),
    .Q(\cpu.dcache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1440),
    .D(_00581_),
    .Q_N(_00238_),
    .Q(\cpu.dcache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1441),
    .D(_00582_),
    .Q_N(_00239_),
    .Q(\cpu.dcache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1442),
    .D(_00583_),
    .Q_N(_00240_),
    .Q(\cpu.dcache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1443),
    .D(_00584_),
    .Q_N(_00241_),
    .Q(\cpu.dcache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1444),
    .D(_00585_),
    .Q_N(_00242_),
    .Q(\cpu.dcache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1445),
    .D(_00586_),
    .Q_N(_14676_),
    .Q(\cpu.dcache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1446),
    .D(_00587_),
    .Q_N(_14675_),
    .Q(\cpu.dcache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1447),
    .D(_00588_),
    .Q_N(_14674_),
    .Q(\cpu.dcache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1448),
    .D(_00589_),
    .Q_N(_00243_),
    .Q(\cpu.dcache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1449),
    .D(_00590_),
    .Q_N(_00224_),
    .Q(\cpu.dcache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1450),
    .D(_00591_),
    .Q_N(_00226_),
    .Q(\cpu.dcache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1451),
    .D(_00592_),
    .Q_N(_00228_),
    .Q(\cpu.dcache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1452),
    .D(_00593_),
    .Q_N(_00230_),
    .Q(\cpu.dcache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1453),
    .D(_00594_),
    .Q_N(_00232_),
    .Q(\cpu.dcache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1454),
    .D(_00595_),
    .Q_N(_00234_),
    .Q(\cpu.dcache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1455),
    .D(_00596_),
    .Q_N(_00235_),
    .Q(\cpu.dcache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1456),
    .D(_00597_),
    .Q_N(_00236_),
    .Q(\cpu.dcache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1457),
    .D(_00598_),
    .Q_N(_00237_),
    .Q(\cpu.dcache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1458),
    .D(_00599_),
    .Q_N(_14673_),
    .Q(\cpu.dcache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1459),
    .D(_00600_),
    .Q_N(_14672_),
    .Q(\cpu.dcache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1460),
    .D(_00601_),
    .Q_N(_14671_),
    .Q(\cpu.dcache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1461),
    .D(_00602_),
    .Q_N(_14670_),
    .Q(\cpu.dcache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1462),
    .D(_00603_),
    .Q_N(_14669_),
    .Q(\cpu.dcache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1463),
    .D(_00604_),
    .Q_N(_14668_),
    .Q(\cpu.dcache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1464),
    .D(_00605_),
    .Q_N(_14667_),
    .Q(\cpu.dcache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1465),
    .D(_00606_),
    .Q_N(_14666_),
    .Q(\cpu.dcache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1466),
    .D(_00607_),
    .Q_N(_14665_),
    .Q(\cpu.dcache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1467),
    .D(_00608_),
    .Q_N(_14664_),
    .Q(\cpu.dcache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1468),
    .D(_00609_),
    .Q_N(_14663_),
    .Q(\cpu.dcache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1469),
    .D(_00610_),
    .Q_N(_14662_),
    .Q(\cpu.dcache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1470),
    .D(_00611_),
    .Q_N(_14661_),
    .Q(\cpu.dcache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1471),
    .D(_00612_),
    .Q_N(_14660_),
    .Q(\cpu.dcache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1472),
    .D(_00613_),
    .Q_N(_14659_),
    .Q(\cpu.dcache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1473),
    .D(_00614_),
    .Q_N(_14658_),
    .Q(\cpu.dcache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1474),
    .D(_00615_),
    .Q_N(_14657_),
    .Q(\cpu.dcache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1475),
    .D(_00616_),
    .Q_N(_14656_),
    .Q(\cpu.dcache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1476),
    .D(_00617_),
    .Q_N(_14655_),
    .Q(\cpu.dcache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1477),
    .D(_00618_),
    .Q_N(_14654_),
    .Q(\cpu.dcache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1478),
    .D(_00619_),
    .Q_N(_14653_),
    .Q(\cpu.dcache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1479),
    .D(_00620_),
    .Q_N(_14652_),
    .Q(\cpu.dcache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1480),
    .D(_00621_),
    .Q_N(_14651_),
    .Q(\cpu.dcache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1481),
    .D(_00622_),
    .Q_N(_14650_),
    .Q(\cpu.dcache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1482),
    .D(_00623_),
    .Q_N(_14649_),
    .Q(\cpu.dcache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1483),
    .D(_00624_),
    .Q_N(_14648_),
    .Q(\cpu.dcache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1484),
    .D(_00625_),
    .Q_N(_14647_),
    .Q(\cpu.dcache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1485),
    .D(_00626_),
    .Q_N(_14646_),
    .Q(\cpu.dcache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1486),
    .D(_00627_),
    .Q_N(_14645_),
    .Q(\cpu.dcache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1487),
    .D(_00628_),
    .Q_N(_14644_),
    .Q(\cpu.dcache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1488),
    .D(_00629_),
    .Q_N(_14643_),
    .Q(\cpu.dcache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1489),
    .D(_00630_),
    .Q_N(_14642_),
    .Q(\cpu.dcache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1490),
    .D(_00631_),
    .Q_N(_14641_),
    .Q(\cpu.dcache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1491),
    .D(_00632_),
    .Q_N(_14640_),
    .Q(\cpu.dcache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1492),
    .D(_00633_),
    .Q_N(_14639_),
    .Q(\cpu.dcache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1493),
    .D(_00634_),
    .Q_N(_14638_),
    .Q(\cpu.dcache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1494),
    .D(_00635_),
    .Q_N(_14637_),
    .Q(\cpu.dcache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1495),
    .D(_00636_),
    .Q_N(_14636_),
    .Q(\cpu.dcache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1496),
    .D(_00637_),
    .Q_N(_14635_),
    .Q(\cpu.dcache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1497),
    .D(_00638_),
    .Q_N(_14634_),
    .Q(\cpu.dcache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1498),
    .D(_00639_),
    .Q_N(_14633_),
    .Q(\cpu.dcache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1499),
    .D(_00640_),
    .Q_N(_14632_),
    .Q(\cpu.dcache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1500),
    .D(_00641_),
    .Q_N(_14631_),
    .Q(\cpu.dcache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1501),
    .D(_00642_),
    .Q_N(_14630_),
    .Q(\cpu.dcache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1502),
    .D(_00643_),
    .Q_N(_14629_),
    .Q(\cpu.dcache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1503),
    .D(_00644_),
    .Q_N(_14628_),
    .Q(\cpu.dcache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1504),
    .D(_00645_),
    .Q_N(_14627_),
    .Q(\cpu.dcache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1505),
    .D(_00646_),
    .Q_N(_14626_),
    .Q(\cpu.dcache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1506),
    .D(_00647_),
    .Q_N(_14625_),
    .Q(\cpu.dcache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1507),
    .D(_00648_),
    .Q_N(_14624_),
    .Q(\cpu.dcache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1508),
    .D(_00649_),
    .Q_N(_14623_),
    .Q(\cpu.dcache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1509),
    .D(_00650_),
    .Q_N(_14622_),
    .Q(\cpu.dcache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1510),
    .D(_00651_),
    .Q_N(_14621_),
    .Q(\cpu.dcache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1511),
    .D(_00652_),
    .Q_N(_14620_),
    .Q(\cpu.dcache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1512),
    .D(_00653_),
    .Q_N(_14619_),
    .Q(\cpu.dcache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1513),
    .D(_00654_),
    .Q_N(_14618_),
    .Q(\cpu.dcache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1514),
    .D(_00655_),
    .Q_N(_14617_),
    .Q(\cpu.dcache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1515),
    .D(_00656_),
    .Q_N(_14616_),
    .Q(\cpu.dcache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1516),
    .D(_00657_),
    .Q_N(_14615_),
    .Q(\cpu.dcache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1517),
    .D(_00658_),
    .Q_N(_14614_),
    .Q(\cpu.dcache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1518),
    .D(_00659_),
    .Q_N(_14613_),
    .Q(\cpu.dcache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1519),
    .D(_00660_),
    .Q_N(_14612_),
    .Q(\cpu.dcache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1520),
    .D(_00661_),
    .Q_N(_14611_),
    .Q(\cpu.dcache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1521),
    .D(_00662_),
    .Q_N(_14610_),
    .Q(\cpu.dcache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1522),
    .D(_00663_),
    .Q_N(_14609_),
    .Q(\cpu.dcache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1523),
    .D(_00664_),
    .Q_N(_14608_),
    .Q(\cpu.dcache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1524),
    .D(_00665_),
    .Q_N(_14607_),
    .Q(\cpu.dcache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1525),
    .D(_00666_),
    .Q_N(_14606_),
    .Q(\cpu.dcache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1526),
    .D(_00667_),
    .Q_N(_14605_),
    .Q(\cpu.dcache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1527),
    .D(_00668_),
    .Q_N(_14604_),
    .Q(\cpu.dcache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1528),
    .D(_00669_),
    .Q_N(_14603_),
    .Q(\cpu.dcache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1529),
    .D(_00670_),
    .Q_N(_14602_),
    .Q(\cpu.dcache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1530),
    .D(_00671_),
    .Q_N(_14601_),
    .Q(\cpu.dcache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1531),
    .D(_00672_),
    .Q_N(_14600_),
    .Q(\cpu.dcache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1532),
    .D(_00673_),
    .Q_N(_14599_),
    .Q(\cpu.dcache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1533),
    .D(_00674_),
    .Q_N(_14598_),
    .Q(\cpu.dcache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1534),
    .D(_00675_),
    .Q_N(_14597_),
    .Q(\cpu.dcache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1535),
    .D(_00676_),
    .Q_N(_14596_),
    .Q(\cpu.dcache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1536),
    .D(_00677_),
    .Q_N(_14595_),
    .Q(\cpu.dcache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1537),
    .D(_00678_),
    .Q_N(_14594_),
    .Q(\cpu.dcache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1538),
    .D(_00679_),
    .Q_N(_14593_),
    .Q(\cpu.dcache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1539),
    .D(_00680_),
    .Q_N(_14592_),
    .Q(\cpu.dcache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1540),
    .D(_00681_),
    .Q_N(_14591_),
    .Q(\cpu.dcache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1541),
    .D(_00682_),
    .Q_N(_14590_),
    .Q(\cpu.dcache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1542),
    .D(_00683_),
    .Q_N(_14589_),
    .Q(\cpu.dcache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1543),
    .D(_00684_),
    .Q_N(_14588_),
    .Q(\cpu.dcache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1544),
    .D(_00685_),
    .Q_N(_14587_),
    .Q(\cpu.dcache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1545),
    .D(_00686_),
    .Q_N(_14586_),
    .Q(\cpu.dcache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1546),
    .D(_00687_),
    .Q_N(_14585_),
    .Q(\cpu.dcache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1547),
    .D(_00688_),
    .Q_N(_14584_),
    .Q(\cpu.dcache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1548),
    .D(_00689_),
    .Q_N(_14583_),
    .Q(\cpu.dcache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1549),
    .D(_00690_),
    .Q_N(_14582_),
    .Q(\cpu.dcache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1550),
    .D(_00691_),
    .Q_N(_14581_),
    .Q(\cpu.dcache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1551),
    .D(_00692_),
    .Q_N(_14580_),
    .Q(\cpu.dcache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1552),
    .D(_00693_),
    .Q_N(_14579_),
    .Q(\cpu.dcache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1553),
    .D(_00694_),
    .Q_N(_14578_),
    .Q(\cpu.dcache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1554),
    .D(_00695_),
    .Q_N(_14577_),
    .Q(\cpu.dcache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1555),
    .D(_00696_),
    .Q_N(_14576_),
    .Q(\cpu.dcache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1556),
    .D(_00697_),
    .Q_N(_14575_),
    .Q(\cpu.dcache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1557),
    .D(_00698_),
    .Q_N(_14574_),
    .Q(\cpu.dcache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1558),
    .D(_00699_),
    .Q_N(_14573_),
    .Q(\cpu.dcache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1559),
    .D(_00700_),
    .Q_N(_14572_),
    .Q(\cpu.dcache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1560),
    .D(_00701_),
    .Q_N(_14571_),
    .Q(\cpu.dcache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1561),
    .D(_00702_),
    .Q_N(_14570_),
    .Q(\cpu.dcache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1562),
    .D(_00703_),
    .Q_N(_14569_),
    .Q(\cpu.dcache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1563),
    .D(_00704_),
    .Q_N(_14568_),
    .Q(\cpu.dcache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1564),
    .D(_00705_),
    .Q_N(_14567_),
    .Q(\cpu.dcache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1565),
    .D(_00706_),
    .Q_N(_14566_),
    .Q(\cpu.dcache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1566),
    .D(_00707_),
    .Q_N(_14565_),
    .Q(\cpu.dcache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1567),
    .D(_00708_),
    .Q_N(_14564_),
    .Q(\cpu.dcache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1568),
    .D(_00709_),
    .Q_N(_14563_),
    .Q(\cpu.dcache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1569),
    .D(_00710_),
    .Q_N(_14562_),
    .Q(\cpu.dcache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1570),
    .D(_00711_),
    .Q_N(_14561_),
    .Q(\cpu.dcache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1571),
    .D(_00712_),
    .Q_N(_14560_),
    .Q(\cpu.dcache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1572),
    .D(_00713_),
    .Q_N(_14559_),
    .Q(\cpu.dcache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1573),
    .D(_00714_),
    .Q_N(_14558_),
    .Q(\cpu.dcache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1574),
    .D(_00715_),
    .Q_N(_14557_),
    .Q(\cpu.dcache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1575),
    .D(_00716_),
    .Q_N(_14556_),
    .Q(\cpu.dcache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1576),
    .D(_00717_),
    .Q_N(_14555_),
    .Q(\cpu.dcache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1577),
    .D(_00718_),
    .Q_N(_14554_),
    .Q(\cpu.dcache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1578),
    .D(_00719_),
    .Q_N(_14553_),
    .Q(\cpu.dcache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1579),
    .D(_00720_),
    .Q_N(_14552_),
    .Q(\cpu.dcache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1580),
    .D(_00721_),
    .Q_N(_14551_),
    .Q(\cpu.dcache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1581),
    .D(_00722_),
    .Q_N(_14550_),
    .Q(\cpu.dcache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1582),
    .D(_00723_),
    .Q_N(_14549_),
    .Q(\cpu.dcache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1583),
    .D(_00724_),
    .Q_N(_14548_),
    .Q(\cpu.dcache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1584),
    .D(_00725_),
    .Q_N(_14547_),
    .Q(\cpu.dcache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1585),
    .D(_00726_),
    .Q_N(_14546_),
    .Q(\cpu.dcache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1586),
    .D(_00727_),
    .Q_N(_14545_),
    .Q(\cpu.dcache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1587),
    .D(_00728_),
    .Q_N(_14544_),
    .Q(\cpu.dcache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1588),
    .D(_00729_),
    .Q_N(_14543_),
    .Q(\cpu.dcache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1589),
    .D(_00730_),
    .Q_N(_14542_),
    .Q(\cpu.dcache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1590),
    .D(_00731_),
    .Q_N(_14541_),
    .Q(\cpu.dcache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1591),
    .D(_00732_),
    .Q_N(_14540_),
    .Q(\cpu.dcache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1592),
    .D(_00733_),
    .Q_N(_14539_),
    .Q(\cpu.dcache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1593),
    .D(_00734_),
    .Q_N(_14538_),
    .Q(\cpu.dcache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1594),
    .D(_00735_),
    .Q_N(_14537_),
    .Q(\cpu.dcache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1595),
    .D(_00736_),
    .Q_N(_14536_),
    .Q(\cpu.dcache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1596),
    .D(_00737_),
    .Q_N(_14535_),
    .Q(\cpu.dcache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1597),
    .D(_00738_),
    .Q_N(_14534_),
    .Q(\cpu.dcache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.dcache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1598),
    .D(_00739_),
    .Q_N(_14533_),
    .Q(\cpu.dcache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_br$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1599),
    .D(_00740_),
    .Q_N(_14532_),
    .Q(\cpu.br ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[0]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1600),
    .D(_00741_),
    .Q_N(_14531_),
    .Q(\cpu.cond[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[1]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1601),
    .D(_00742_),
    .Q_N(_14530_),
    .Q(\cpu.cond[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_cond[2]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1602),
    .D(_00743_),
    .Q_N(_00266_),
    .Q(\cpu.cond[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_div$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1603),
    .D(_00744_),
    .Q_N(_14529_),
    .Q(\cpu.dec.div ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_all$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1604),
    .D(_00745_),
    .Q_N(_14528_),
    .Q(\cpu.dec.do_flush_all ));
 sg13g2_dfrbp_1 \cpu.dec.r_flush_write$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1605),
    .D(_00746_),
    .Q_N(_14527_),
    .Q(\cpu.dec.do_flush_write ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[0]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1606),
    .D(_00747_),
    .Q_N(_14526_),
    .Q(\cpu.dec.imm[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[10]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1607),
    .D(_00748_),
    .Q_N(_14525_),
    .Q(\cpu.dec.imm[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[11]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1608),
    .D(_00749_),
    .Q_N(_14524_),
    .Q(\cpu.dec.imm[11] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[12]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1609),
    .D(_00750_),
    .Q_N(_14523_),
    .Q(\cpu.dec.imm[12] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[13]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1610),
    .D(_00751_),
    .Q_N(_14522_),
    .Q(\cpu.dec.imm[13] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[14]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1611),
    .D(_00752_),
    .Q_N(_14521_),
    .Q(\cpu.dec.imm[14] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[15]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1612),
    .D(_00753_),
    .Q_N(_14520_),
    .Q(\cpu.dec.imm[15] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[1]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1613),
    .D(_00754_),
    .Q_N(_14519_),
    .Q(\cpu.dec.imm[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1614),
    .D(_00755_),
    .Q_N(_14518_),
    .Q(\cpu.dec.imm[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1615),
    .D(_00756_),
    .Q_N(_14517_),
    .Q(\cpu.dec.imm[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[4]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1616),
    .D(_00757_),
    .Q_N(_14516_),
    .Q(\cpu.dec.imm[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[5]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1617),
    .D(_00758_),
    .Q_N(_14515_),
    .Q(\cpu.dec.imm[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[6]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1618),
    .D(_00759_),
    .Q_N(_14514_),
    .Q(\cpu.dec.imm[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[7]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1619),
    .D(_00760_),
    .Q_N(_14513_),
    .Q(\cpu.dec.imm[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[8]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1620),
    .D(_00761_),
    .Q_N(_14512_),
    .Q(\cpu.dec.imm[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_imm[9]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1621),
    .D(_00762_),
    .Q_N(_14511_),
    .Q(\cpu.dec.imm[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_inv_mmu$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1622),
    .D(_00763_),
    .Q_N(_14510_),
    .Q(\cpu.dec.do_inv_mmu ));
 sg13g2_dfrbp_1 \cpu.dec.r_io$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1623),
    .D(_00764_),
    .Q_N(_14509_),
    .Q(\cpu.dec.io ));
 sg13g2_dfrbp_1 \cpu.dec.r_jmp$_SDFFCE_PP0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1624),
    .D(_00765_),
    .Q_N(_00250_),
    .Q(\cpu.dec.jmp ));
 sg13g2_dfrbp_1 \cpu.dec.r_load$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1625),
    .D(_00766_),
    .Q_N(_14508_),
    .Q(\cpu.dec.load ));
 sg13g2_dfrbp_1 \cpu.dec.r_mult$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1626),
    .D(_00767_),
    .Q_N(_14507_),
    .Q(\cpu.dec.mult ));
 sg13g2_dfrbp_1 \cpu.dec.r_needs_rs2$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1627),
    .D(_00768_),
    .Q_N(_14920_),
    .Q(\cpu.dec.needs_rs2 ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[10]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1628),
    .D(_00011_),
    .Q_N(_14921_),
    .Q(\cpu.dec.r_op[10] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[1]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1629),
    .D(_00012_),
    .Q_N(_14922_),
    .Q(\cpu.dec.r_op[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[2]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1630),
    .D(_00013_),
    .Q_N(_14923_),
    .Q(\cpu.dec.r_op[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[3]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1631),
    .D(_00014_),
    .Q_N(_14924_),
    .Q(\cpu.dec.r_op[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[4]$_DFF_P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1632),
    .D(_00015_),
    .Q_N(_14925_),
    .Q(\cpu.dec.r_op[4] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[5]$_DFF_P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1633),
    .D(_00016_),
    .Q_N(_14926_),
    .Q(\cpu.dec.r_op[5] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[6]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1634),
    .D(_00017_),
    .Q_N(_14927_),
    .Q(\cpu.dec.r_op[6] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[7]$_DFF_P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1635),
    .D(_00018_),
    .Q_N(_14928_),
    .Q(\cpu.dec.r_op[7] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[8]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1636),
    .D(_00019_),
    .Q_N(_14929_),
    .Q(\cpu.dec.r_op[8] ));
 sg13g2_dfrbp_1 \cpu.dec.r_op[9]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1637),
    .D(_00020_),
    .Q_N(_14506_),
    .Q(\cpu.dec.r_op[9] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[0]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1638),
    .D(_00769_),
    .Q_N(_14505_),
    .Q(\cpu.dec.r_rd[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[1]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1639),
    .D(_00770_),
    .Q_N(_14504_),
    .Q(\cpu.dec.r_rd[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1640),
    .D(_00771_),
    .Q_N(_14503_),
    .Q(\cpu.dec.r_rd[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rd[3]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1641),
    .D(_00772_),
    .Q_N(_14930_),
    .Q(\cpu.dec.r_rd[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_ready$_DFF_P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1642),
    .D(_00052_),
    .Q_N(_14502_),
    .Q(\cpu.dec.iready ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[0]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1643),
    .D(_00773_),
    .Q_N(_14501_),
    .Q(\cpu.dec.r_rs1[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[1]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1644),
    .D(_00774_),
    .Q_N(_14500_),
    .Q(\cpu.dec.r_rs1[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1645),
    .D(_00775_),
    .Q_N(_14499_),
    .Q(\cpu.dec.r_rs1[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs1[3]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1646),
    .D(_00776_),
    .Q_N(_14498_),
    .Q(\cpu.dec.r_rs1[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[0]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1647),
    .D(_00777_),
    .Q_N(_14497_),
    .Q(\cpu.dec.r_rs2[0] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[1]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1648),
    .D(_00778_),
    .Q_N(_14496_),
    .Q(\cpu.dec.r_rs2[1] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1649),
    .D(_00779_),
    .Q_N(_14495_),
    .Q(\cpu.dec.r_rs2[2] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2[3]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1650),
    .D(_00780_),
    .Q_N(_14494_),
    .Q(\cpu.dec.r_rs2[3] ));
 sg13g2_dfrbp_1 \cpu.dec.r_rs2_pc$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1651),
    .D(_00781_),
    .Q_N(_14493_),
    .Q(\cpu.dec.r_rs2_pc ));
 sg13g2_dfrbp_1 \cpu.dec.r_set_cc$_SDFFCE_PP0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1652),
    .D(_00782_),
    .Q_N(_14492_),
    .Q(\cpu.dec.r_set_cc ));
 sg13g2_dfrbp_1 \cpu.dec.r_store$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1653),
    .D(_00783_),
    .Q_N(_00291_),
    .Q(\cpu.dec.r_store ));
 sg13g2_dfrbp_1 \cpu.dec.r_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1654),
    .D(_00784_),
    .Q_N(_14491_),
    .Q(\cpu.dec.r_swapsp ));
 sg13g2_dfrbp_1 \cpu.dec.r_sys_call$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1655),
    .D(_00785_),
    .Q_N(_00267_),
    .Q(\cpu.dec.r_sys_call ));
 sg13g2_dfrbp_1 \cpu.dec.r_trap$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1656),
    .D(_00786_),
    .Q_N(_14490_),
    .Q(\cpu.dec.r_trap ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1657),
    .D(_00787_),
    .Q_N(_14489_),
    .Q(\cpu.ex.genblk3.r_mmu_d_proxy ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1658),
    .D(_00788_),
    .Q_N(_00190_),
    .Q(\cpu.ex.genblk3.r_mmu_enable ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1659),
    .D(_00789_),
    .Q_N(_14931_),
    .Q(\cpu.ex.genblk3.r_prev_supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_supmode$_DFF_P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1660),
    .D(\cpu.ex.genblk3.c_supmode ),
    .Q_N(_00191_),
    .Q(\cpu.dec.supmode ));
 sg13g2_dfrbp_1 \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1661),
    .D(_00790_),
    .Q_N(_14488_),
    .Q(\cpu.dec.user_io ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[0]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1662),
    .D(_00791_),
    .Q_N(_14487_),
    .Q(\cpu.ex.r_10[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[10]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1663),
    .D(_00792_),
    .Q_N(_14486_),
    .Q(\cpu.ex.r_10[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[11]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1664),
    .D(_00793_),
    .Q_N(_14485_),
    .Q(\cpu.ex.r_10[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1665),
    .D(_00794_),
    .Q_N(_14484_),
    .Q(\cpu.ex.r_10[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1666),
    .D(_00795_),
    .Q_N(_14483_),
    .Q(\cpu.ex.r_10[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[14]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1667),
    .D(_00796_),
    .Q_N(_14482_),
    .Q(\cpu.ex.r_10[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1668),
    .D(_00797_),
    .Q_N(_14481_),
    .Q(\cpu.ex.r_10[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[1]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1669),
    .D(_00798_),
    .Q_N(_14480_),
    .Q(\cpu.ex.r_10[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[2]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1670),
    .D(_00799_),
    .Q_N(_14479_),
    .Q(\cpu.ex.r_10[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[3]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1671),
    .D(_00800_),
    .Q_N(_14478_),
    .Q(\cpu.ex.r_10[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[4]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1672),
    .D(_00801_),
    .Q_N(_14477_),
    .Q(\cpu.ex.r_10[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[5]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1673),
    .D(_00802_),
    .Q_N(_14476_),
    .Q(\cpu.ex.r_10[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[6]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1674),
    .D(_00803_),
    .Q_N(_14475_),
    .Q(\cpu.ex.r_10[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[7]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1675),
    .D(_00804_),
    .Q_N(_14474_),
    .Q(\cpu.ex.r_10[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[8]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1676),
    .D(_00805_),
    .Q_N(_14473_),
    .Q(\cpu.ex.r_10[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_10[9]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1677),
    .D(_00806_),
    .Q_N(_14472_),
    .Q(\cpu.ex.r_10[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1678),
    .D(_00807_),
    .Q_N(_14471_),
    .Q(\cpu.ex.r_11[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[10]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1679),
    .D(_00808_),
    .Q_N(_14470_),
    .Q(\cpu.ex.r_11[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[11]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1680),
    .D(_00809_),
    .Q_N(_14469_),
    .Q(\cpu.ex.r_11[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1681),
    .D(_00810_),
    .Q_N(_14468_),
    .Q(\cpu.ex.r_11[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[13]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1682),
    .D(_00811_),
    .Q_N(_14467_),
    .Q(\cpu.ex.r_11[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[14]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1683),
    .D(_00812_),
    .Q_N(_14466_),
    .Q(\cpu.ex.r_11[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[15]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1684),
    .D(_00813_),
    .Q_N(_14465_),
    .Q(\cpu.ex.r_11[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1685),
    .D(_00814_),
    .Q_N(_14464_),
    .Q(\cpu.ex.r_11[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[2]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1686),
    .D(_00815_),
    .Q_N(_14463_),
    .Q(\cpu.ex.r_11[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1687),
    .D(_00816_),
    .Q_N(_14462_),
    .Q(\cpu.ex.r_11[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[4]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1688),
    .D(_00817_),
    .Q_N(_14461_),
    .Q(\cpu.ex.r_11[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1689),
    .D(_00818_),
    .Q_N(_14460_),
    .Q(\cpu.ex.r_11[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[6]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1690),
    .D(_00819_),
    .Q_N(_14459_),
    .Q(\cpu.ex.r_11[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[7]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1691),
    .D(_00820_),
    .Q_N(_14458_),
    .Q(\cpu.ex.r_11[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1692),
    .D(_00821_),
    .Q_N(_14457_),
    .Q(\cpu.ex.r_11[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_11[9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1693),
    .D(_00822_),
    .Q_N(_14456_),
    .Q(\cpu.ex.r_11[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1694),
    .D(_00823_),
    .Q_N(_14455_),
    .Q(\cpu.ex.r_12[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1695),
    .D(_00824_),
    .Q_N(_14454_),
    .Q(\cpu.ex.r_12[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1696),
    .D(_00825_),
    .Q_N(_14453_),
    .Q(\cpu.ex.r_12[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1697),
    .D(_00826_),
    .Q_N(_14452_),
    .Q(\cpu.ex.r_12[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1698),
    .D(_00827_),
    .Q_N(_14451_),
    .Q(\cpu.ex.r_12[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1699),
    .D(_00828_),
    .Q_N(_14450_),
    .Q(\cpu.ex.r_12[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[15]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1700),
    .D(_00829_),
    .Q_N(_14449_),
    .Q(\cpu.ex.r_12[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[1]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1701),
    .D(_00830_),
    .Q_N(_14448_),
    .Q(\cpu.ex.r_12[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1702),
    .D(_00831_),
    .Q_N(_14447_),
    .Q(\cpu.ex.r_12[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1703),
    .D(_00832_),
    .Q_N(_14446_),
    .Q(\cpu.ex.r_12[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[4]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1704),
    .D(_00833_),
    .Q_N(_14445_),
    .Q(\cpu.ex.r_12[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[5]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1705),
    .D(_00834_),
    .Q_N(_14444_),
    .Q(\cpu.ex.r_12[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[6]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1706),
    .D(_00835_),
    .Q_N(_14443_),
    .Q(\cpu.ex.r_12[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1707),
    .D(_00836_),
    .Q_N(_14442_),
    .Q(\cpu.ex.r_12[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[8]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1708),
    .D(_00837_),
    .Q_N(_14441_),
    .Q(\cpu.ex.r_12[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_12[9]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1709),
    .D(_00838_),
    .Q_N(_14440_),
    .Q(\cpu.ex.r_12[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[0]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1710),
    .D(_00839_),
    .Q_N(_14439_),
    .Q(\cpu.ex.r_13[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1711),
    .D(_00840_),
    .Q_N(_14438_),
    .Q(\cpu.ex.r_13[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[11]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1712),
    .D(_00841_),
    .Q_N(_14437_),
    .Q(\cpu.ex.r_13[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1713),
    .D(_00842_),
    .Q_N(_14436_),
    .Q(\cpu.ex.r_13[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1714),
    .D(_00843_),
    .Q_N(_14435_),
    .Q(\cpu.ex.r_13[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[14]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1715),
    .D(_00844_),
    .Q_N(_14434_),
    .Q(\cpu.ex.r_13[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[15]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1716),
    .D(_00845_),
    .Q_N(_14433_),
    .Q(\cpu.ex.r_13[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1717),
    .D(_00846_),
    .Q_N(_14432_),
    .Q(\cpu.ex.r_13[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1718),
    .D(_00847_),
    .Q_N(_14431_),
    .Q(\cpu.ex.r_13[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[3]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1719),
    .D(_00848_),
    .Q_N(_14430_),
    .Q(\cpu.ex.r_13[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[4]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1720),
    .D(_00849_),
    .Q_N(_14429_),
    .Q(\cpu.ex.r_13[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1721),
    .D(_00850_),
    .Q_N(_14428_),
    .Q(\cpu.ex.r_13[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[6]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1722),
    .D(_00851_),
    .Q_N(_14427_),
    .Q(\cpu.ex.r_13[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[7]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1723),
    .D(_00852_),
    .Q_N(_14426_),
    .Q(\cpu.ex.r_13[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[8]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1724),
    .D(_00853_),
    .Q_N(_14425_),
    .Q(\cpu.ex.r_13[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_13[9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1725),
    .D(_00854_),
    .Q_N(_14424_),
    .Q(\cpu.ex.r_13[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[0]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1726),
    .D(_00855_),
    .Q_N(_14423_),
    .Q(\cpu.ex.r_14[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[10]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1727),
    .D(_00856_),
    .Q_N(_14422_),
    .Q(\cpu.ex.r_14[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[11]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1728),
    .D(_00857_),
    .Q_N(_14421_),
    .Q(\cpu.ex.r_14[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[12]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1729),
    .D(_00858_),
    .Q_N(_14420_),
    .Q(\cpu.ex.r_14[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[13]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1730),
    .D(_00859_),
    .Q_N(_14419_),
    .Q(\cpu.ex.r_14[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[14]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1731),
    .D(_00860_),
    .Q_N(_14418_),
    .Q(\cpu.ex.r_14[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1732),
    .D(_00861_),
    .Q_N(_14417_),
    .Q(\cpu.ex.r_14[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[1]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1733),
    .D(_00862_),
    .Q_N(_14416_),
    .Q(\cpu.ex.r_14[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1734),
    .D(_00863_),
    .Q_N(_14415_),
    .Q(\cpu.ex.r_14[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1735),
    .D(_00864_),
    .Q_N(_14414_),
    .Q(\cpu.ex.r_14[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1736),
    .D(_00865_),
    .Q_N(_14413_),
    .Q(\cpu.ex.r_14[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[5]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1737),
    .D(_00866_),
    .Q_N(_14412_),
    .Q(\cpu.ex.r_14[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[6]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1738),
    .D(_00867_),
    .Q_N(_14411_),
    .Q(\cpu.ex.r_14[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[7]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1739),
    .D(_00868_),
    .Q_N(_14410_),
    .Q(\cpu.ex.r_14[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[8]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1740),
    .D(_00869_),
    .Q_N(_14409_),
    .Q(\cpu.ex.r_14[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_14[9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1741),
    .D(_00870_),
    .Q_N(_14408_),
    .Q(\cpu.ex.r_14[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1742),
    .D(_00871_),
    .Q_N(_14407_),
    .Q(\cpu.ex.r_15[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[10]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1743),
    .D(_00872_),
    .Q_N(_00260_),
    .Q(\cpu.ex.r_15[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1744),
    .D(_00873_),
    .Q_N(_00261_),
    .Q(\cpu.ex.r_15[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[12]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1745),
    .D(_00874_),
    .Q_N(_00262_),
    .Q(\cpu.ex.r_15[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[13]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1746),
    .D(_00875_),
    .Q_N(_00263_),
    .Q(\cpu.ex.r_15[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[14]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1747),
    .D(_00876_),
    .Q_N(_00264_),
    .Q(\cpu.ex.r_15[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[15]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1748),
    .D(_00877_),
    .Q_N(_00265_),
    .Q(\cpu.ex.r_15[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[1]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1749),
    .D(_00878_),
    .Q_N(_00251_),
    .Q(\cpu.ex.r_15[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[2]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1750),
    .D(_00879_),
    .Q_N(_00252_),
    .Q(\cpu.ex.r_15[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1751),
    .D(_00880_),
    .Q_N(_00253_),
    .Q(\cpu.ex.r_15[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[4]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1752),
    .D(_00881_),
    .Q_N(_00254_),
    .Q(\cpu.ex.r_15[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1753),
    .D(_00882_),
    .Q_N(_00255_),
    .Q(\cpu.ex.r_15[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[6]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1754),
    .D(_00883_),
    .Q_N(_00256_),
    .Q(\cpu.ex.r_15[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[7]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1755),
    .D(_00884_),
    .Q_N(_00257_),
    .Q(\cpu.ex.r_15[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1756),
    .D(_00885_),
    .Q_N(_00258_),
    .Q(\cpu.ex.r_15[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_15[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1757),
    .D(_00886_),
    .Q_N(_00259_),
    .Q(\cpu.ex.r_15[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1758),
    .D(_00887_),
    .Q_N(_14406_),
    .Q(\cpu.ex.r_8[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1759),
    .D(_00888_),
    .Q_N(_14405_),
    .Q(\cpu.ex.r_8[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[11]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1760),
    .D(_00889_),
    .Q_N(_14404_),
    .Q(\cpu.ex.r_8[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[12]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1761),
    .D(_00890_),
    .Q_N(_14403_),
    .Q(\cpu.ex.r_8[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[13]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1762),
    .D(_00891_),
    .Q_N(_14402_),
    .Q(\cpu.ex.r_8[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[14]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1763),
    .D(_00892_),
    .Q_N(_14401_),
    .Q(\cpu.ex.r_8[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[15]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1764),
    .D(_00893_),
    .Q_N(_14400_),
    .Q(\cpu.ex.r_8[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1765),
    .D(_00894_),
    .Q_N(_14399_),
    .Q(\cpu.ex.r_8[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[2]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1766),
    .D(_00895_),
    .Q_N(_14398_),
    .Q(\cpu.ex.r_8[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1767),
    .D(_00896_),
    .Q_N(_14397_),
    .Q(\cpu.ex.r_8[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[4]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1768),
    .D(_00897_),
    .Q_N(_14396_),
    .Q(\cpu.ex.r_8[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1769),
    .D(_00898_),
    .Q_N(_14395_),
    .Q(\cpu.ex.r_8[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[6]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1770),
    .D(_00899_),
    .Q_N(_14394_),
    .Q(\cpu.ex.r_8[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[7]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1771),
    .D(_00900_),
    .Q_N(_14393_),
    .Q(\cpu.ex.r_8[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[8]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1772),
    .D(_00901_),
    .Q_N(_14392_),
    .Q(\cpu.ex.r_8[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_8[9]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1773),
    .D(_00902_),
    .Q_N(_14391_),
    .Q(\cpu.ex.r_8[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[0]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1774),
    .D(_00903_),
    .Q_N(_14390_),
    .Q(\cpu.ex.r_9[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[10]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1775),
    .D(_00904_),
    .Q_N(_14389_),
    .Q(\cpu.ex.r_9[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[11]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1776),
    .D(_00905_),
    .Q_N(_14388_),
    .Q(\cpu.ex.r_9[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[12]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1777),
    .D(_00906_),
    .Q_N(_14387_),
    .Q(\cpu.ex.r_9[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[13]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1778),
    .D(_00907_),
    .Q_N(_14386_),
    .Q(\cpu.ex.r_9[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[14]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1779),
    .D(_00908_),
    .Q_N(_14385_),
    .Q(\cpu.ex.r_9[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[15]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1780),
    .D(_00909_),
    .Q_N(_14384_),
    .Q(\cpu.ex.r_9[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[1]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1781),
    .D(_00910_),
    .Q_N(_14383_),
    .Q(\cpu.ex.r_9[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[2]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1782),
    .D(_00911_),
    .Q_N(_14382_),
    .Q(\cpu.ex.r_9[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[3]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1783),
    .D(_00912_),
    .Q_N(_14381_),
    .Q(\cpu.ex.r_9[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[4]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1784),
    .D(_00913_),
    .Q_N(_14380_),
    .Q(\cpu.ex.r_9[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[5]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1785),
    .D(_00914_),
    .Q_N(_14379_),
    .Q(\cpu.ex.r_9[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[6]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1786),
    .D(_00915_),
    .Q_N(_14378_),
    .Q(\cpu.ex.r_9[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[7]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1787),
    .D(_00916_),
    .Q_N(_14377_),
    .Q(\cpu.ex.r_9[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[8]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1788),
    .D(_00917_),
    .Q_N(_14376_),
    .Q(\cpu.ex.r_9[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_9[9]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1789),
    .D(_00918_),
    .Q_N(_14932_),
    .Q(\cpu.ex.r_9[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_branch_stall$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1790),
    .D(_00053_),
    .Q_N(_14375_),
    .Q(\cpu.ex.r_branch_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_d_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net1791),
    .D(_00919_),
    .Q_N(_14933_),
    .Q(\cpu.d_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_div_running$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1792),
    .D(\cpu.ex.c_div_running ),
    .Q_N(_14374_),
    .Q(\cpu.ex.r_div_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1793),
    .D(_00920_),
    .Q_N(_14373_),
    .Q(\cpu.ex.r_epc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[10]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1794),
    .D(_00921_),
    .Q_N(_14372_),
    .Q(\cpu.ex.r_epc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1795),
    .D(_00922_),
    .Q_N(_14371_),
    .Q(\cpu.ex.r_epc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1796),
    .D(_00923_),
    .Q_N(_14370_),
    .Q(\cpu.ex.r_epc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1797),
    .D(_00924_),
    .Q_N(_14369_),
    .Q(\cpu.ex.r_epc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[14]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1798),
    .D(_00925_),
    .Q_N(_14368_),
    .Q(\cpu.ex.r_epc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[1]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1799),
    .D(_00926_),
    .Q_N(_14367_),
    .Q(\cpu.ex.r_epc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1800),
    .D(_00927_),
    .Q_N(_14366_),
    .Q(\cpu.ex.r_epc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[3]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1801),
    .D(_00928_),
    .Q_N(_14365_),
    .Q(\cpu.ex.r_epc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[4]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1802),
    .D(_00929_),
    .Q_N(_14364_),
    .Q(\cpu.ex.r_epc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1803),
    .D(_00930_),
    .Q_N(_14363_),
    .Q(\cpu.ex.r_epc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[6]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1804),
    .D(_00931_),
    .Q_N(_14362_),
    .Q(\cpu.ex.r_epc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[7]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1805),
    .D(_00932_),
    .Q_N(_14361_),
    .Q(\cpu.ex.r_epc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[8]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1806),
    .D(_00933_),
    .Q_N(_14360_),
    .Q(\cpu.ex.r_epc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_epc[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1807),
    .D(_00934_),
    .Q_N(_14359_),
    .Q(\cpu.ex.r_epc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_fetch$_SDFF_PN1_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1808),
    .D(_00935_),
    .Q_N(_00187_),
    .Q(\cpu.ex.ifetch ));
 sg13g2_dfrbp_1 \cpu.ex.r_flush_write$_SDFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1809),
    .D(_00936_),
    .Q_N(_14358_),
    .Q(\cpu.dcache.flush_write ));
 sg13g2_dfrbp_1 \cpu.ex.r_i_flush_all$_SDFF_PP0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1810),
    .D(_00937_),
    .Q_N(_14357_),
    .Q(\cpu.ex.i_flush_all ));
 sg13g2_dfrbp_1 \cpu.ex.r_ie$_SDFFE_PP0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1811),
    .D(_00938_),
    .Q_N(_14356_),
    .Q(\cpu.ex.r_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_io_access$_SDFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1812),
    .D(_00939_),
    .Q_N(_00195_),
    .Q(\cpu.ex.io_access ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[0]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1813),
    .D(_00940_),
    .Q_N(_14355_),
    .Q(\cpu.ex.r_lr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[10]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net1814),
    .D(_00941_),
    .Q_N(_14354_),
    .Q(\cpu.ex.r_lr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[11]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1815),
    .D(_00942_),
    .Q_N(_14353_),
    .Q(\cpu.ex.r_lr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[12]$_DFFE_PP_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1816),
    .D(_00943_),
    .Q_N(_14352_),
    .Q(\cpu.ex.r_lr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[13]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1817),
    .D(_00944_),
    .Q_N(_14351_),
    .Q(\cpu.ex.r_lr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[14]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1818),
    .D(_00945_),
    .Q_N(_14350_),
    .Q(\cpu.ex.r_lr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[1]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1819),
    .D(_00946_),
    .Q_N(_14349_),
    .Q(\cpu.ex.r_lr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[2]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1820),
    .D(_00947_),
    .Q_N(_14348_),
    .Q(\cpu.ex.r_lr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[3]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1821),
    .D(_00948_),
    .Q_N(_14347_),
    .Q(\cpu.ex.r_lr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[4]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1822),
    .D(_00949_),
    .Q_N(_14346_),
    .Q(\cpu.ex.r_lr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[5]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1823),
    .D(_00950_),
    .Q_N(_14345_),
    .Q(\cpu.ex.r_lr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[6]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1824),
    .D(_00951_),
    .Q_N(_14344_),
    .Q(\cpu.ex.r_lr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[7]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1825),
    .D(_00952_),
    .Q_N(_14343_),
    .Q(\cpu.ex.r_lr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[8]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1826),
    .D(_00953_),
    .Q_N(_14342_),
    .Q(\cpu.ex.r_lr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_lr[9]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1827),
    .D(_00954_),
    .Q_N(_14934_),
    .Q(\cpu.ex.r_lr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[0]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1828),
    .D(\cpu.ex.c_mult[0] ),
    .Q_N(_00091_),
    .Q(\cpu.ex.r_mult[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[10]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1829),
    .D(\cpu.ex.c_mult[10] ),
    .Q_N(_00159_),
    .Q(\cpu.ex.r_mult[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[11]$_DFF_P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1830),
    .D(\cpu.ex.c_mult[11] ),
    .Q_N(_00160_),
    .Q(\cpu.ex.r_mult[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[12]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1831),
    .D(\cpu.ex.c_mult[12] ),
    .Q_N(_00161_),
    .Q(\cpu.ex.r_mult[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[13]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1832),
    .D(\cpu.ex.c_mult[13] ),
    .Q_N(_00162_),
    .Q(\cpu.ex.r_mult[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[14]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1833),
    .D(\cpu.ex.c_mult[14] ),
    .Q_N(_00163_),
    .Q(\cpu.ex.r_mult[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[15]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1834),
    .D(\cpu.ex.c_mult[15] ),
    .Q_N(_14341_),
    .Q(\cpu.ex.r_mult[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[16]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1835),
    .D(_00955_),
    .Q_N(_14340_),
    .Q(\cpu.ex.r_mult[16] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[17]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1836),
    .D(_00956_),
    .Q_N(_14339_),
    .Q(\cpu.ex.r_mult[17] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[18]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1837),
    .D(_00957_),
    .Q_N(_14338_),
    .Q(\cpu.ex.r_mult[18] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[19]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1838),
    .D(_00958_),
    .Q_N(_14935_),
    .Q(\cpu.ex.r_mult[19] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[1]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1839),
    .D(\cpu.ex.c_mult[1] ),
    .Q_N(_00092_),
    .Q(\cpu.ex.r_mult[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[20]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1840),
    .D(_00959_),
    .Q_N(_14337_),
    .Q(\cpu.ex.r_mult[20] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[21]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1841),
    .D(_00960_),
    .Q_N(_14336_),
    .Q(\cpu.ex.r_mult[21] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[22]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1842),
    .D(_00961_),
    .Q_N(_14335_),
    .Q(\cpu.ex.r_mult[22] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[23]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1843),
    .D(_00962_),
    .Q_N(_14334_),
    .Q(\cpu.ex.r_mult[23] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[24]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1844),
    .D(_00963_),
    .Q_N(_14333_),
    .Q(\cpu.ex.r_mult[24] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[25]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1845),
    .D(_00964_),
    .Q_N(_14332_),
    .Q(\cpu.ex.r_mult[25] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[26]$_DFFE_PP_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1846),
    .D(_00965_),
    .Q_N(_14331_),
    .Q(\cpu.ex.r_mult[26] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[27]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1847),
    .D(_00966_),
    .Q_N(_14330_),
    .Q(\cpu.ex.r_mult[27] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[28]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1848),
    .D(_00967_),
    .Q_N(_14329_),
    .Q(\cpu.ex.r_mult[28] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[29]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1849),
    .D(_00968_),
    .Q_N(_14936_),
    .Q(\cpu.ex.r_mult[29] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[2]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1850),
    .D(\cpu.ex.c_mult[2] ),
    .Q_N(_00103_),
    .Q(\cpu.ex.r_mult[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[30]$_DFFE_PP_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1851),
    .D(_00969_),
    .Q_N(_14328_),
    .Q(\cpu.ex.r_mult[30] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[31]$_DFFE_PP_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1852),
    .D(_00970_),
    .Q_N(_14937_),
    .Q(\cpu.ex.r_mult[31] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[3]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1853),
    .D(\cpu.ex.c_mult[3] ),
    .Q_N(_00113_),
    .Q(\cpu.ex.r_mult[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[4]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1854),
    .D(\cpu.ex.c_mult[4] ),
    .Q_N(_00120_),
    .Q(\cpu.ex.r_mult[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[5]$_DFF_P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1855),
    .D(\cpu.ex.c_mult[5] ),
    .Q_N(_00132_),
    .Q(\cpu.ex.r_mult[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[6]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1856),
    .D(\cpu.ex.c_mult[6] ),
    .Q_N(_00144_),
    .Q(\cpu.ex.r_mult[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[7]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1857),
    .D(\cpu.ex.c_mult[7] ),
    .Q_N(_00156_),
    .Q(\cpu.ex.r_mult[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[8]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1858),
    .D(\cpu.ex.c_mult[8] ),
    .Q_N(_00157_),
    .Q(\cpu.ex.r_mult[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult[9]$_DFF_P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1859),
    .D(\cpu.ex.c_mult[9] ),
    .Q_N(_00158_),
    .Q(\cpu.ex.r_mult[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[0]$_DFF_P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1860),
    .D(\cpu.ex.c_mult_off[0] ),
    .Q_N(_14938_),
    .Q(\cpu.ex.r_mult_off[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[1]$_DFF_P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1861),
    .D(\cpu.ex.c_mult_off[1] ),
    .Q_N(_14939_),
    .Q(\cpu.ex.r_mult_off[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[2]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1862),
    .D(\cpu.ex.c_mult_off[2] ),
    .Q_N(_14940_),
    .Q(\cpu.ex.r_mult_off[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_off[3]$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1863),
    .D(\cpu.ex.c_mult_off[3] ),
    .Q_N(_14941_),
    .Q(\cpu.ex.r_mult_off[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_mult_running$_DFF_P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1864),
    .D(\cpu.ex.c_mult_running ),
    .Q_N(_00197_),
    .Q(\cpu.ex.r_mult_running ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1865),
    .D(_00971_),
    .Q_N(_00198_),
    .Q(\cpu.ex.pc[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[10]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1866),
    .D(_00972_),
    .Q_N(_00285_),
    .Q(\cpu.ex.pc[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[11]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1867),
    .D(_00973_),
    .Q_N(_00284_),
    .Q(\cpu.ex.pc[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[12]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1868),
    .D(_00974_),
    .Q_N(_00194_),
    .Q(\cpu.ex.pc[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[13]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1869),
    .D(_00975_),
    .Q_N(_00193_),
    .Q(\cpu.ex.pc[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[14]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1870),
    .D(_00976_),
    .Q_N(_00192_),
    .Q(\cpu.ex.pc[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1871),
    .D(_00977_),
    .Q_N(_00283_),
    .Q(\cpu.ex.pc[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1872),
    .D(_00978_),
    .Q_N(_00189_),
    .Q(\cpu.ex.pc[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1873),
    .D(_00979_),
    .Q_N(_00188_),
    .Q(\cpu.ex.pc[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1874),
    .D(_00980_),
    .Q_N(_00290_),
    .Q(\cpu.ex.pc[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1875),
    .D(_00981_),
    .Q_N(_00289_),
    .Q(\cpu.ex.pc[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1876),
    .D(_00982_),
    .Q_N(_00288_),
    .Q(\cpu.ex.pc[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1877),
    .D(_00983_),
    .Q_N(_00282_),
    .Q(\cpu.ex.pc[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[8]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1878),
    .D(_00984_),
    .Q_N(_00287_),
    .Q(\cpu.ex.pc[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_pc[9]$_DFFE_PP_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1879),
    .D(_00985_),
    .Q_N(_00286_),
    .Q(\cpu.ex.pc[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_prev_ie$_SDFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1880),
    .D(_00986_),
    .Q_N(_14327_),
    .Q(\cpu.ex.r_prev_ie ));
 sg13g2_dfrbp_1 \cpu.ex.r_read_stall$_SDFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1881),
    .D(_00987_),
    .Q_N(_00196_),
    .Q(\cpu.ex.r_read_stall ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[0]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1882),
    .D(_00988_),
    .Q_N(_14326_),
    .Q(\cpu.ex.r_sp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[10]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1883),
    .D(_00989_),
    .Q_N(_14325_),
    .Q(\cpu.ex.r_sp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[11]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1884),
    .D(_00990_),
    .Q_N(_14324_),
    .Q(\cpu.ex.r_sp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[12]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1885),
    .D(_00991_),
    .Q_N(_14323_),
    .Q(\cpu.ex.r_sp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[13]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1886),
    .D(_00992_),
    .Q_N(_14322_),
    .Q(\cpu.ex.r_sp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[14]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1887),
    .D(_00993_),
    .Q_N(_14321_),
    .Q(\cpu.ex.r_sp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[1]$_DFFE_PP_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1888),
    .D(_00994_),
    .Q_N(_14320_),
    .Q(\cpu.ex.r_sp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[2]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1889),
    .D(_00995_),
    .Q_N(_14319_),
    .Q(\cpu.ex.r_sp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[3]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1890),
    .D(_00996_),
    .Q_N(_14318_),
    .Q(\cpu.ex.r_sp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[4]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1891),
    .D(_00997_),
    .Q_N(_14317_),
    .Q(\cpu.ex.r_sp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[5]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1892),
    .D(_00998_),
    .Q_N(_14316_),
    .Q(\cpu.ex.r_sp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[6]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1893),
    .D(_00999_),
    .Q_N(_14315_),
    .Q(\cpu.ex.r_sp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[7]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1894),
    .D(_01000_),
    .Q_N(_14314_),
    .Q(\cpu.ex.r_sp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1895),
    .D(_01001_),
    .Q_N(_14313_),
    .Q(\cpu.ex.r_sp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_sp[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1896),
    .D(_01002_),
    .Q_N(_14312_),
    .Q(\cpu.ex.r_sp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1897),
    .D(_01003_),
    .Q_N(_14311_),
    .Q(\cpu.ex.r_stmp[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1898),
    .D(_01004_),
    .Q_N(_14310_),
    .Q(\cpu.ex.r_stmp[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1899),
    .D(_01005_),
    .Q_N(_14309_),
    .Q(\cpu.ex.r_stmp[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1900),
    .D(_01006_),
    .Q_N(_14308_),
    .Q(\cpu.ex.r_stmp[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1901),
    .D(_01007_),
    .Q_N(_14307_),
    .Q(\cpu.ex.r_stmp[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1902),
    .D(_01008_),
    .Q_N(_14306_),
    .Q(\cpu.ex.r_stmp[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1903),
    .D(_01009_),
    .Q_N(_14305_),
    .Q(\cpu.ex.r_stmp[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1904),
    .D(_01010_),
    .Q_N(_14304_),
    .Q(\cpu.ex.r_stmp[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1905),
    .D(_01011_),
    .Q_N(_14303_),
    .Q(\cpu.ex.r_stmp[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1906),
    .D(_01012_),
    .Q_N(_14302_),
    .Q(\cpu.ex.r_stmp[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1907),
    .D(_01013_),
    .Q_N(_14301_),
    .Q(\cpu.ex.r_stmp[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1908),
    .D(_01014_),
    .Q_N(_14300_),
    .Q(\cpu.ex.r_stmp[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1909),
    .D(_01015_),
    .Q_N(_14299_),
    .Q(\cpu.ex.r_stmp[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1910),
    .D(_01016_),
    .Q_N(_14298_),
    .Q(\cpu.ex.r_stmp[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1911),
    .D(_01017_),
    .Q_N(_14297_),
    .Q(\cpu.ex.r_stmp[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_stmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1912),
    .D(_01018_),
    .Q_N(_14296_),
    .Q(\cpu.ex.r_stmp[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[0]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1913),
    .D(_01019_),
    .Q_N(_00249_),
    .Q(\cpu.ex.mmu_reg_data[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[10]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1914),
    .D(_01020_),
    .Q_N(_00231_),
    .Q(\cpu.addr[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[11]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1915),
    .D(_01021_),
    .Q_N(_00233_),
    .Q(\cpu.addr[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[12]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1916),
    .D(_01022_),
    .Q_N(_14295_),
    .Q(\cpu.addr[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[13]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1917),
    .D(_01023_),
    .Q_N(_14294_),
    .Q(\cpu.addr[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[14]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1918),
    .D(_01024_),
    .Q_N(_14293_),
    .Q(\cpu.addr[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[15]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1919),
    .D(_01025_),
    .Q_N(_14292_),
    .Q(\cpu.addr[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[1]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1920),
    .D(_01026_),
    .Q_N(_00268_),
    .Q(\cpu.addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[2]$_DFFE_PP_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1921),
    .D(_01027_),
    .Q_N(_14291_),
    .Q(\cpu.addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[3]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1922),
    .D(_01028_),
    .Q_N(_00215_),
    .Q(\cpu.addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[4]$_DFFE_PP_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1923),
    .D(_01029_),
    .Q_N(_00220_),
    .Q(\cpu.addr[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[5]$_DFFE_PP_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1924),
    .D(_01030_),
    .Q_N(_00221_),
    .Q(\cpu.addr[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[6]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1925),
    .D(_01031_),
    .Q_N(_00223_),
    .Q(\cpu.addr[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[7]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1926),
    .D(_01032_),
    .Q_N(_00225_),
    .Q(\cpu.addr[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[8]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1927),
    .D(_01033_),
    .Q_N(_00227_),
    .Q(\cpu.addr[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb[9]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1928),
    .D(_01034_),
    .Q_N(_00229_),
    .Q(\cpu.addr[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1929),
    .D(_01035_),
    .Q_N(_14290_),
    .Q(\cpu.ex.r_wb_addr[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1930),
    .D(_01036_),
    .Q_N(_14289_),
    .Q(\cpu.ex.r_wb_addr[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1931),
    .D(_01037_),
    .Q_N(_14288_),
    .Q(\cpu.ex.r_wb_addr[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1932),
    .D(_01038_),
    .Q_N(_14287_),
    .Q(\cpu.ex.r_wb_addr[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_swapsp$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1933),
    .D(_01039_),
    .Q_N(_14942_),
    .Q(\cpu.ex.r_wb_swapsp ));
 sg13g2_dfrbp_1 \cpu.ex.r_wb_valid$_DFF_P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1934),
    .D(_00054_),
    .Q_N(_00248_),
    .Q(\cpu.ex.r_wb_valid ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1935),
    .D(_01040_),
    .Q_N(_00216_),
    .Q(\cpu.dcache.wdata[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[10]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1936),
    .D(_01041_),
    .Q_N(_14286_),
    .Q(\cpu.dcache.wdata[10] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[11]$_DFFE_PP_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1937),
    .D(_01042_),
    .Q_N(_14285_),
    .Q(\cpu.dcache.wdata[11] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[12]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1938),
    .D(_01043_),
    .Q_N(_14284_),
    .Q(\cpu.dcache.wdata[12] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[13]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1939),
    .D(_01044_),
    .Q_N(_14283_),
    .Q(\cpu.dcache.wdata[13] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1940),
    .D(_01045_),
    .Q_N(_14282_),
    .Q(\cpu.dcache.wdata[14] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[15]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1941),
    .D(_01046_),
    .Q_N(_14281_),
    .Q(\cpu.dcache.wdata[15] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[1]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1942),
    .D(_01047_),
    .Q_N(_00176_),
    .Q(\cpu.dcache.wdata[1] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[2]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1943),
    .D(_01048_),
    .Q_N(_00177_),
    .Q(\cpu.dcache.wdata[2] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1944),
    .D(_01049_),
    .Q_N(_00280_),
    .Q(\cpu.dcache.wdata[3] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1945),
    .D(_01050_),
    .Q_N(_00178_),
    .Q(\cpu.dcache.wdata[4] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1946),
    .D(_01051_),
    .Q_N(_00179_),
    .Q(\cpu.dcache.wdata[5] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[6]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1947),
    .D(_01052_),
    .Q_N(_00180_),
    .Q(\cpu.dcache.wdata[6] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[7]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1948),
    .D(_01053_),
    .Q_N(_00274_),
    .Q(\cpu.dcache.wdata[7] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[8]$_DFFE_PP_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1949),
    .D(_01054_),
    .Q_N(_14280_),
    .Q(\cpu.dcache.wdata[8] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wdata[9]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1950),
    .D(_01055_),
    .Q_N(_14279_),
    .Q(\cpu.dcache.wdata[9] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1951),
    .D(_01056_),
    .Q_N(_14278_),
    .Q(\cpu.ex.r_wmask[0] ));
 sg13g2_dfrbp_1 \cpu.ex.r_wmask[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1952),
    .D(_01057_),
    .Q_N(_14277_),
    .Q(\cpu.ex.r_wmask[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1953),
    .D(_01058_),
    .Q_N(_00281_),
    .Q(\cpu.ex.mmu_read[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1954),
    .D(_01059_),
    .Q_N(_14276_),
    .Q(\cpu.ex.mmu_read[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1955),
    .D(_01060_),
    .Q_N(_00186_),
    .Q(\cpu.ex.mmu_read[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1956),
    .D(_01061_),
    .Q_N(_14275_),
    .Q(\cpu.ex.mmu_read[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1957),
    .D(_01062_),
    .Q_N(_00247_),
    .Q(\cpu.ex.mmu_read[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1958),
    .D(_01063_),
    .Q_N(_14274_),
    .Q(\cpu.ex.mmu_read[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1959),
    .D(_01064_),
    .Q_N(_14273_),
    .Q(\cpu.ex.mmu_read[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1960),
    .D(_01065_),
    .Q_N(_14272_),
    .Q(\cpu.genblk1.mmu.r_valid_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1961),
    .D(_01066_),
    .Q_N(_14271_),
    .Q(\cpu.genblk1.mmu.r_valid_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1962),
    .D(_01067_),
    .Q_N(_14270_),
    .Q(\cpu.genblk1.mmu.r_valid_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1963),
    .D(_01068_),
    .Q_N(_14269_),
    .Q(\cpu.genblk1.mmu.r_valid_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1964),
    .D(_01069_),
    .Q_N(_14268_),
    .Q(\cpu.genblk1.mmu.r_valid_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1965),
    .D(_01070_),
    .Q_N(_14267_),
    .Q(\cpu.genblk1.mmu.r_valid_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1966),
    .D(_01071_),
    .Q_N(_14266_),
    .Q(\cpu.genblk1.mmu.r_valid_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1967),
    .D(_01072_),
    .Q_N(_14265_),
    .Q(\cpu.genblk1.mmu.r_valid_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1968),
    .D(_01073_),
    .Q_N(_14264_),
    .Q(\cpu.genblk1.mmu.r_valid_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1969),
    .D(_01074_),
    .Q_N(_14263_),
    .Q(\cpu.genblk1.mmu.r_valid_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1970),
    .D(_01075_),
    .Q_N(_14262_),
    .Q(\cpu.genblk1.mmu.r_valid_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1971),
    .D(_01076_),
    .Q_N(_14261_),
    .Q(\cpu.genblk1.mmu.r_valid_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1972),
    .D(_01077_),
    .Q_N(_14260_),
    .Q(\cpu.genblk1.mmu.r_valid_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1973),
    .D(_01078_),
    .Q_N(_14259_),
    .Q(\cpu.genblk1.mmu.r_valid_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1974),
    .D(_01079_),
    .Q_N(_14258_),
    .Q(\cpu.genblk1.mmu.r_valid_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1975),
    .D(_01080_),
    .Q_N(_14257_),
    .Q(\cpu.genblk1.mmu.r_valid_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1976),
    .D(_01081_),
    .Q_N(_14256_),
    .Q(\cpu.genblk1.mmu.r_valid_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1977),
    .D(_01082_),
    .Q_N(_14255_),
    .Q(\cpu.genblk1.mmu.r_valid_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1978),
    .D(_01083_),
    .Q_N(_14254_),
    .Q(\cpu.genblk1.mmu.r_valid_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1979),
    .D(_01084_),
    .Q_N(_14253_),
    .Q(\cpu.genblk1.mmu.r_valid_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1980),
    .D(_01085_),
    .Q_N(_14252_),
    .Q(\cpu.genblk1.mmu.r_valid_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1981),
    .D(_01086_),
    .Q_N(_14251_),
    .Q(\cpu.genblk1.mmu.r_valid_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1982),
    .D(_01087_),
    .Q_N(_14250_),
    .Q(\cpu.genblk1.mmu.r_valid_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1983),
    .D(_01088_),
    .Q_N(_14249_),
    .Q(\cpu.genblk1.mmu.r_valid_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1984),
    .D(_01089_),
    .Q_N(_14248_),
    .Q(\cpu.genblk1.mmu.r_valid_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1985),
    .D(_01090_),
    .Q_N(_14247_),
    .Q(\cpu.genblk1.mmu.r_valid_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1986),
    .D(_01091_),
    .Q_N(_14246_),
    .Q(\cpu.genblk1.mmu.r_valid_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1987),
    .D(_01092_),
    .Q_N(_14245_),
    .Q(\cpu.genblk1.mmu.r_valid_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1988),
    .D(_01093_),
    .Q_N(_14244_),
    .Q(\cpu.genblk1.mmu.r_valid_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1989),
    .D(_01094_),
    .Q_N(_14243_),
    .Q(\cpu.genblk1.mmu.r_valid_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1990),
    .D(_01095_),
    .Q_N(_14242_),
    .Q(\cpu.genblk1.mmu.r_valid_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1991),
    .D(_01096_),
    .Q_N(_14241_),
    .Q(\cpu.genblk1.mmu.r_valid_d[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1992),
    .D(_01097_),
    .Q_N(_14240_),
    .Q(\cpu.genblk1.mmu.r_valid_i[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1993),
    .D(_01098_),
    .Q_N(_14239_),
    .Q(\cpu.genblk1.mmu.r_valid_i[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1994),
    .D(_01099_),
    .Q_N(_14238_),
    .Q(\cpu.genblk1.mmu.r_valid_i[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1995),
    .D(_01100_),
    .Q_N(_14237_),
    .Q(\cpu.genblk1.mmu.r_valid_i[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1996),
    .D(_01101_),
    .Q_N(_14236_),
    .Q(\cpu.genblk1.mmu.r_valid_i[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1997),
    .D(_01102_),
    .Q_N(_14235_),
    .Q(\cpu.genblk1.mmu.r_valid_i[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1998),
    .D(_01103_),
    .Q_N(_14234_),
    .Q(\cpu.genblk1.mmu.r_valid_i[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1999),
    .D(_01104_),
    .Q_N(_14233_),
    .Q(\cpu.genblk1.mmu.r_valid_i[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2000),
    .D(_01105_),
    .Q_N(_14232_),
    .Q(\cpu.genblk1.mmu.r_valid_i[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2001),
    .D(_01106_),
    .Q_N(_14231_),
    .Q(\cpu.genblk1.mmu.r_valid_i[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2002),
    .D(_01107_),
    .Q_N(_14230_),
    .Q(\cpu.genblk1.mmu.r_valid_i[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2003),
    .D(_01108_),
    .Q_N(_14229_),
    .Q(\cpu.genblk1.mmu.r_valid_i[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net2004),
    .D(_01109_),
    .Q_N(_14228_),
    .Q(\cpu.genblk1.mmu.r_valid_i[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2005),
    .D(_01110_),
    .Q_N(_14227_),
    .Q(\cpu.genblk1.mmu.r_valid_i[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2006),
    .D(_01111_),
    .Q_N(_14226_),
    .Q(\cpu.genblk1.mmu.r_valid_i[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2007),
    .D(_01112_),
    .Q_N(_14225_),
    .Q(\cpu.genblk1.mmu.r_valid_i[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2008),
    .D(_01113_),
    .Q_N(_14224_),
    .Q(\cpu.genblk1.mmu.r_valid_i[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net2009),
    .D(_01114_),
    .Q_N(_14223_),
    .Q(\cpu.genblk1.mmu.r_valid_i[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2010),
    .D(_01115_),
    .Q_N(_14222_),
    .Q(\cpu.genblk1.mmu.r_valid_i[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2011),
    .D(_01116_),
    .Q_N(_14221_),
    .Q(\cpu.genblk1.mmu.r_valid_i[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2012),
    .D(_01117_),
    .Q_N(_14220_),
    .Q(\cpu.genblk1.mmu.r_valid_i[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2013),
    .D(_01118_),
    .Q_N(_14219_),
    .Q(\cpu.genblk1.mmu.r_valid_i[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2014),
    .D(_01119_),
    .Q_N(_14218_),
    .Q(\cpu.genblk1.mmu.r_valid_i[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net2015),
    .D(_01120_),
    .Q_N(_14217_),
    .Q(\cpu.genblk1.mmu.r_valid_i[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net2016),
    .D(_01121_),
    .Q_N(_14216_),
    .Q(\cpu.genblk1.mmu.r_valid_i[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net2017),
    .D(_01122_),
    .Q_N(_14215_),
    .Q(\cpu.genblk1.mmu.r_valid_i[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2018),
    .D(_01123_),
    .Q_N(_14214_),
    .Q(\cpu.genblk1.mmu.r_valid_i[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net2019),
    .D(_01124_),
    .Q_N(_14213_),
    .Q(\cpu.genblk1.mmu.r_valid_i[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2020),
    .D(_01125_),
    .Q_N(_14212_),
    .Q(\cpu.genblk1.mmu.r_valid_i[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net2021),
    .D(_01126_),
    .Q_N(_14211_),
    .Q(\cpu.genblk1.mmu.r_valid_i[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2022),
    .D(_01127_),
    .Q_N(_14210_),
    .Q(\cpu.genblk1.mmu.r_valid_i[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2023),
    .D(_01128_),
    .Q_N(_14209_),
    .Q(\cpu.genblk1.mmu.r_valid_i[9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2024),
    .D(_01129_),
    .Q_N(_14208_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2025),
    .D(_01130_),
    .Q_N(_14207_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2026),
    .D(_01131_),
    .Q_N(_14206_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2027),
    .D(_01132_),
    .Q_N(_14205_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2028),
    .D(_01133_),
    .Q_N(_14204_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2029),
    .D(_01134_),
    .Q_N(_14203_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2030),
    .D(_01135_),
    .Q_N(_14202_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2031),
    .D(_01136_),
    .Q_N(_14201_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2032),
    .D(_01137_),
    .Q_N(_14200_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2033),
    .D(_01138_),
    .Q_N(_14199_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2034),
    .D(_01139_),
    .Q_N(_14198_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2035),
    .D(_01140_),
    .Q_N(_14197_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2036),
    .D(_01141_),
    .Q_N(_14196_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2037),
    .D(_01142_),
    .Q_N(_14195_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2038),
    .D(_01143_),
    .Q_N(_14194_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2039),
    .D(_01144_),
    .Q_N(_14193_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2040),
    .D(_01145_),
    .Q_N(_14192_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2041),
    .D(_01146_),
    .Q_N(_14191_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2042),
    .D(_01147_),
    .Q_N(_14190_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2043),
    .D(_01148_),
    .Q_N(_14189_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2044),
    .D(_01149_),
    .Q_N(_14188_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2045),
    .D(_01150_),
    .Q_N(_14187_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2046),
    .D(_01151_),
    .Q_N(_14186_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2047),
    .D(_01152_),
    .Q_N(_14185_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2048),
    .D(_01153_),
    .Q_N(_14184_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2049),
    .D(_01154_),
    .Q_N(_14183_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2050),
    .D(_01155_),
    .Q_N(_14182_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2051),
    .D(_01156_),
    .Q_N(_14181_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2052),
    .D(_01157_),
    .Q_N(_14180_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2053),
    .D(_01158_),
    .Q_N(_14179_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2054),
    .D(_01159_),
    .Q_N(_14178_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2055),
    .D(_01160_),
    .Q_N(_14177_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2056),
    .D(_01161_),
    .Q_N(_14176_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2057),
    .D(_01162_),
    .Q_N(_14175_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2058),
    .D(_01163_),
    .Q_N(_14174_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2059),
    .D(_01164_),
    .Q_N(_14173_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2060),
    .D(_01165_),
    .Q_N(_14172_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2061),
    .D(_01166_),
    .Q_N(_14171_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2062),
    .D(_01167_),
    .Q_N(_14170_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2063),
    .D(_01168_),
    .Q_N(_14169_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2064),
    .D(_01169_),
    .Q_N(_14168_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2065),
    .D(_01170_),
    .Q_N(_14167_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2066),
    .D(_01171_),
    .Q_N(_14166_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2067),
    .D(_01172_),
    .Q_N(_14165_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2068),
    .D(_01173_),
    .Q_N(_14164_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2069),
    .D(_01174_),
    .Q_N(_14163_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2070),
    .D(_01175_),
    .Q_N(_14162_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2071),
    .D(_01176_),
    .Q_N(_14161_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2072),
    .D(_01177_),
    .Q_N(_14160_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2073),
    .D(_01178_),
    .Q_N(_14159_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2074),
    .D(_01179_),
    .Q_N(_14158_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2075),
    .D(_01180_),
    .Q_N(_14157_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2076),
    .D(_01181_),
    .Q_N(_14156_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2077),
    .D(_01182_),
    .Q_N(_14155_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2078),
    .D(_01183_),
    .Q_N(_14154_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2079),
    .D(_01184_),
    .Q_N(_14153_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2080),
    .D(_01185_),
    .Q_N(_14152_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2081),
    .D(_01186_),
    .Q_N(_14151_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2082),
    .D(_01187_),
    .Q_N(_14150_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2083),
    .D(_01188_),
    .Q_N(_14149_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2084),
    .D(_01189_),
    .Q_N(_14148_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2085),
    .D(_01190_),
    .Q_N(_14147_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2086),
    .D(_01191_),
    .Q_N(_14146_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2087),
    .D(_01192_),
    .Q_N(_14145_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2088),
    .D(_01193_),
    .Q_N(_14144_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2089),
    .D(_01194_),
    .Q_N(_14143_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2090),
    .D(_01195_),
    .Q_N(_14142_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2091),
    .D(_01196_),
    .Q_N(_14141_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2092),
    .D(_01197_),
    .Q_N(_14140_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2093),
    .D(_01198_),
    .Q_N(_14139_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2094),
    .D(_01199_),
    .Q_N(_14138_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2095),
    .D(_01200_),
    .Q_N(_14137_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2096),
    .D(_01201_),
    .Q_N(_14136_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2097),
    .D(_01202_),
    .Q_N(_14135_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2098),
    .D(_01203_),
    .Q_N(_14134_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2099),
    .D(_01204_),
    .Q_N(_14133_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2100),
    .D(_01205_),
    .Q_N(_14132_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2101),
    .D(_01206_),
    .Q_N(_14131_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2102),
    .D(_01207_),
    .Q_N(_14130_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2103),
    .D(_01208_),
    .Q_N(_14129_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2104),
    .D(_01209_),
    .Q_N(_14128_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2105),
    .D(_01210_),
    .Q_N(_14127_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2106),
    .D(_01211_),
    .Q_N(_14126_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2107),
    .D(_01212_),
    .Q_N(_14125_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2108),
    .D(_01213_),
    .Q_N(_14124_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2109),
    .D(_01214_),
    .Q_N(_14123_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2110),
    .D(_01215_),
    .Q_N(_14122_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2111),
    .D(_01216_),
    .Q_N(_14121_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2112),
    .D(_01217_),
    .Q_N(_14120_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2113),
    .D(_01218_),
    .Q_N(_14119_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2114),
    .D(_01219_),
    .Q_N(_14118_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2115),
    .D(_01220_),
    .Q_N(_14117_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2116),
    .D(_01221_),
    .Q_N(_14116_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2117),
    .D(_01222_),
    .Q_N(_14115_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2118),
    .D(_01223_),
    .Q_N(_14114_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2119),
    .D(_01224_),
    .Q_N(_14113_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2120),
    .D(_01225_),
    .Q_N(_14112_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2121),
    .D(_01226_),
    .Q_N(_14111_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2122),
    .D(_01227_),
    .Q_N(_14110_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2123),
    .D(_01228_),
    .Q_N(_14109_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2124),
    .D(_01229_),
    .Q_N(_14108_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2125),
    .D(_01230_),
    .Q_N(_14107_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2126),
    .D(_01231_),
    .Q_N(_14106_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2127),
    .D(_01232_),
    .Q_N(_14105_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2128),
    .D(_01233_),
    .Q_N(_14104_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2129),
    .D(_01234_),
    .Q_N(_14103_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2130),
    .D(_01235_),
    .Q_N(_14102_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2131),
    .D(_01236_),
    .Q_N(_14101_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2132),
    .D(_01237_),
    .Q_N(_14100_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2133),
    .D(_01238_),
    .Q_N(_14099_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2134),
    .D(_01239_),
    .Q_N(_14098_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2135),
    .D(_01240_),
    .Q_N(_14097_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2136),
    .D(_01241_),
    .Q_N(_14096_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2137),
    .D(_01242_),
    .Q_N(_14095_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2138),
    .D(_01243_),
    .Q_N(_14094_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2139),
    .D(_01244_),
    .Q_N(_14093_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2140),
    .D(_01245_),
    .Q_N(_14092_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2141),
    .D(_01246_),
    .Q_N(_14091_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2142),
    .D(_01247_),
    .Q_N(_14090_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2143),
    .D(_01248_),
    .Q_N(_14089_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2144),
    .D(_01249_),
    .Q_N(_14088_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2145),
    .D(_01250_),
    .Q_N(_14087_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2146),
    .D(_01251_),
    .Q_N(_14086_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2147),
    .D(_01252_),
    .Q_N(_14085_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2148),
    .D(_01253_),
    .Q_N(_14084_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2149),
    .D(_01254_),
    .Q_N(_14083_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2150),
    .D(_01255_),
    .Q_N(_14082_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2151),
    .D(_01256_),
    .Q_N(_14081_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2152),
    .D(_01257_),
    .Q_N(_14080_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2153),
    .D(_01258_),
    .Q_N(_14079_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2154),
    .D(_01259_),
    .Q_N(_14078_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2155),
    .D(_01260_),
    .Q_N(_14077_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2156),
    .D(_01261_),
    .Q_N(_14076_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2157),
    .D(_01262_),
    .Q_N(_14075_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2158),
    .D(_01263_),
    .Q_N(_14074_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2159),
    .D(_01264_),
    .Q_N(_14073_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2160),
    .D(_01265_),
    .Q_N(_14072_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2161),
    .D(_01266_),
    .Q_N(_14071_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2162),
    .D(_01267_),
    .Q_N(_14070_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2163),
    .D(_01268_),
    .Q_N(_14069_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2164),
    .D(_01269_),
    .Q_N(_14068_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2165),
    .D(_01270_),
    .Q_N(_14067_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2166),
    .D(_01271_),
    .Q_N(_14066_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2167),
    .D(_01272_),
    .Q_N(_14065_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2168),
    .D(_01273_),
    .Q_N(_14064_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2169),
    .D(_01274_),
    .Q_N(_14063_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2170),
    .D(_01275_),
    .Q_N(_14062_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2171),
    .D(_01276_),
    .Q_N(_14061_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2172),
    .D(_01277_),
    .Q_N(_14060_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2173),
    .D(_01278_),
    .Q_N(_14059_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2174),
    .D(_01279_),
    .Q_N(_14058_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2175),
    .D(_01280_),
    .Q_N(_14057_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2176),
    .D(_01281_),
    .Q_N(_14056_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2177),
    .D(_01282_),
    .Q_N(_14055_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2178),
    .D(_01283_),
    .Q_N(_14054_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2179),
    .D(_01284_),
    .Q_N(_14053_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2180),
    .D(_01285_),
    .Q_N(_14052_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2181),
    .D(_01286_),
    .Q_N(_14051_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2182),
    .D(_01287_),
    .Q_N(_14050_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2183),
    .D(_01288_),
    .Q_N(_14049_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2184),
    .D(_01289_),
    .Q_N(_14048_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2185),
    .D(_01290_),
    .Q_N(_14047_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2186),
    .D(_01291_),
    .Q_N(_14046_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2187),
    .D(_01292_),
    .Q_N(_14045_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2188),
    .D(_01293_),
    .Q_N(_14044_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2189),
    .D(_01294_),
    .Q_N(_14043_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2190),
    .D(_01295_),
    .Q_N(_14042_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2191),
    .D(_01296_),
    .Q_N(_14041_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2192),
    .D(_01297_),
    .Q_N(_14040_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2193),
    .D(_01298_),
    .Q_N(_14039_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2194),
    .D(_01299_),
    .Q_N(_14038_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2195),
    .D(_01300_),
    .Q_N(_14037_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2196),
    .D(_01301_),
    .Q_N(_14036_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2197),
    .D(_01302_),
    .Q_N(_14035_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2198),
    .D(_01303_),
    .Q_N(_14034_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2199),
    .D(_01304_),
    .Q_N(_14033_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2200),
    .D(_01305_),
    .Q_N(_14032_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2201),
    .D(_01306_),
    .Q_N(_14031_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2202),
    .D(_01307_),
    .Q_N(_14030_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2203),
    .D(_01308_),
    .Q_N(_14029_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2204),
    .D(_01309_),
    .Q_N(_14028_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2205),
    .D(_01310_),
    .Q_N(_14027_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2206),
    .D(_01311_),
    .Q_N(_14026_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net2207),
    .D(_01312_),
    .Q_N(_14025_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2208),
    .D(_01313_),
    .Q_N(_14024_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2209),
    .D(_01314_),
    .Q_N(_14023_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2210),
    .D(_01315_),
    .Q_N(_14022_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2211),
    .D(_01316_),
    .Q_N(_14021_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2212),
    .D(_01317_),
    .Q_N(_14020_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net2213),
    .D(_01318_),
    .Q_N(_14019_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2214),
    .D(_01319_),
    .Q_N(_14018_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2215),
    .D(_01320_),
    .Q_N(_14017_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2216),
    .D(_01321_),
    .Q_N(_14016_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2217),
    .D(_01322_),
    .Q_N(_14015_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net2218),
    .D(_01323_),
    .Q_N(_14014_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2219),
    .D(_01324_),
    .Q_N(_14013_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2220),
    .D(_01325_),
    .Q_N(_14012_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net2221),
    .D(_01326_),
    .Q_N(_14011_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2222),
    .D(_01327_),
    .Q_N(_14010_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2223),
    .D(_01328_),
    .Q_N(_14009_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2224),
    .D(_01329_),
    .Q_N(_14008_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2225),
    .D(_01330_),
    .Q_N(_14007_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2226),
    .D(_01331_),
    .Q_N(_14006_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2227),
    .D(_01332_),
    .Q_N(_14005_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2228),
    .D(_01333_),
    .Q_N(_14004_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2229),
    .D(_01334_),
    .Q_N(_14003_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net2230),
    .D(_01335_),
    .Q_N(_14002_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2231),
    .D(_01336_),
    .Q_N(_14001_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2232),
    .D(_01337_),
    .Q_N(_14000_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2233),
    .D(_01338_),
    .Q_N(_13999_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net2234),
    .D(_01339_),
    .Q_N(_13998_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2235),
    .D(_01340_),
    .Q_N(_13997_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2236),
    .D(_01341_),
    .Q_N(_13996_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2237),
    .D(_01342_),
    .Q_N(_13995_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2238),
    .D(_01343_),
    .Q_N(_13994_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net2239),
    .D(_01344_),
    .Q_N(_13993_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2240),
    .D(_01345_),
    .Q_N(_13992_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net2241),
    .D(_01346_),
    .Q_N(_13991_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2242),
    .D(_01347_),
    .Q_N(_13990_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2243),
    .D(_01348_),
    .Q_N(_13989_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2244),
    .D(_01349_),
    .Q_N(_13988_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2245),
    .D(_01350_),
    .Q_N(_13987_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2246),
    .D(_01351_),
    .Q_N(_13986_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2247),
    .D(_01352_),
    .Q_N(_13985_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2248),
    .D(_01353_),
    .Q_N(_13984_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2249),
    .D(_01354_),
    .Q_N(_13983_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2250),
    .D(_01355_),
    .Q_N(_13982_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2251),
    .D(_01356_),
    .Q_N(_13981_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2252),
    .D(_01357_),
    .Q_N(_13980_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2253),
    .D(_01358_),
    .Q_N(_13979_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2254),
    .D(_01359_),
    .Q_N(_13978_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2255),
    .D(_01360_),
    .Q_N(_13977_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2256),
    .D(_01361_),
    .Q_N(_13976_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2257),
    .D(_01362_),
    .Q_N(_13975_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net2258),
    .D(_01363_),
    .Q_N(_13974_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2259),
    .D(_01364_),
    .Q_N(_13973_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2260),
    .D(_01365_),
    .Q_N(_13972_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net2261),
    .D(_01366_),
    .Q_N(_13971_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2262),
    .D(_01367_),
    .Q_N(_13970_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2263),
    .D(_01368_),
    .Q_N(_13969_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2264),
    .D(_01369_),
    .Q_N(_13968_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2265),
    .D(_01370_),
    .Q_N(_13967_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2266),
    .D(_01371_),
    .Q_N(_13966_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2267),
    .D(_01372_),
    .Q_N(_13965_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2268),
    .D(_01373_),
    .Q_N(_13964_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2269),
    .D(_01374_),
    .Q_N(_13963_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2270),
    .D(_01375_),
    .Q_N(_13962_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2271),
    .D(_01376_),
    .Q_N(_13961_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2272),
    .D(_01377_),
    .Q_N(_13960_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2273),
    .D(_01378_),
    .Q_N(_13959_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2274),
    .D(_01379_),
    .Q_N(_13958_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2275),
    .D(_01380_),
    .Q_N(_13957_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2276),
    .D(_01381_),
    .Q_N(_13956_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2277),
    .D(_01382_),
    .Q_N(_13955_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2278),
    .D(_01383_),
    .Q_N(_13954_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2279),
    .D(_01384_),
    .Q_N(_13953_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2280),
    .D(_01385_),
    .Q_N(_13952_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2281),
    .D(_01386_),
    .Q_N(_13951_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2282),
    .D(_01387_),
    .Q_N(_13950_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2283),
    .D(_01388_),
    .Q_N(_13949_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2284),
    .D(_01389_),
    .Q_N(_13948_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2285),
    .D(_01390_),
    .Q_N(_13947_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2286),
    .D(_01391_),
    .Q_N(_13946_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2287),
    .D(_01392_),
    .Q_N(_13945_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2288),
    .D(_01393_),
    .Q_N(_13944_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2289),
    .D(_01394_),
    .Q_N(_13943_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2290),
    .D(_01395_),
    .Q_N(_13942_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2291),
    .D(_01396_),
    .Q_N(_13941_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2292),
    .D(_01397_),
    .Q_N(_13940_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2293),
    .D(_01398_),
    .Q_N(_13939_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2294),
    .D(_01399_),
    .Q_N(_13938_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2295),
    .D(_01400_),
    .Q_N(_13937_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2296),
    .D(_01401_),
    .Q_N(_13936_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2297),
    .D(_01402_),
    .Q_N(_13935_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2298),
    .D(_01403_),
    .Q_N(_13934_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2299),
    .D(_01404_),
    .Q_N(_13933_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2300),
    .D(_01405_),
    .Q_N(_13932_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2301),
    .D(_01406_),
    .Q_N(_13931_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2302),
    .D(_01407_),
    .Q_N(_13930_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2303),
    .D(_01408_),
    .Q_N(_13929_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net2304),
    .D(_01409_),
    .Q_N(_13928_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2305),
    .D(_01410_),
    .Q_N(_13927_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net2306),
    .D(_01411_),
    .Q_N(_13926_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2307),
    .D(_01412_),
    .Q_N(_13925_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2308),
    .D(_01413_),
    .Q_N(_13924_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2309),
    .D(_01414_),
    .Q_N(_13923_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2310),
    .D(_01415_),
    .Q_N(_13922_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2311),
    .D(_01416_),
    .Q_N(_13921_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net2312),
    .D(_01417_),
    .Q_N(_13920_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net2313),
    .D(_01418_),
    .Q_N(_13919_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net2314),
    .D(_01419_),
    .Q_N(_13918_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2315),
    .D(_01420_),
    .Q_N(_13917_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2316),
    .D(_01421_),
    .Q_N(_13916_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net2317),
    .D(_01422_),
    .Q_N(_13915_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2318),
    .D(_01423_),
    .Q_N(_13914_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net2319),
    .D(_01424_),
    .Q_N(_13913_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2320),
    .D(_01425_),
    .Q_N(_13912_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net2321),
    .D(_01426_),
    .Q_N(_13911_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net2322),
    .D(_01427_),
    .Q_N(_13910_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2323),
    .D(_01428_),
    .Q_N(_13909_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2324),
    .D(_01429_),
    .Q_N(_13908_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2325),
    .D(_01430_),
    .Q_N(_13907_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2326),
    .D(_01431_),
    .Q_N(_13906_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2327),
    .D(_01432_),
    .Q_N(_13905_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net2328),
    .D(_01433_),
    .Q_N(_13904_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2329),
    .D(_01434_),
    .Q_N(_13903_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2330),
    .D(_01435_),
    .Q_N(_13902_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2331),
    .D(_01436_),
    .Q_N(_13901_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net2332),
    .D(_01437_),
    .Q_N(_13900_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2333),
    .D(_01438_),
    .Q_N(_13899_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2334),
    .D(_01439_),
    .Q_N(_13898_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2335),
    .D(_01440_),
    .Q_N(_13897_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2336),
    .D(_01441_),
    .Q_N(_13896_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2337),
    .D(_01442_),
    .Q_N(_13895_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net2338),
    .D(_01443_),
    .Q_N(_13894_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2339),
    .D(_01444_),
    .Q_N(_13893_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2340),
    .D(_01445_),
    .Q_N(_13892_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net2341),
    .D(_01446_),
    .Q_N(_13891_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2342),
    .D(_01447_),
    .Q_N(_13890_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2343),
    .D(_01448_),
    .Q_N(_13889_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2344),
    .D(_01449_),
    .Q_N(_13888_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net2345),
    .D(_01450_),
    .Q_N(_13887_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2346),
    .D(_01451_),
    .Q_N(_13886_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2347),
    .D(_01452_),
    .Q_N(_13885_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2348),
    .D(_01453_),
    .Q_N(_13884_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net2349),
    .D(_01454_),
    .Q_N(_13883_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2350),
    .D(_01455_),
    .Q_N(_13882_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2351),
    .D(_01456_),
    .Q_N(_13881_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2352),
    .D(_01457_),
    .Q_N(_13880_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2353),
    .D(_01458_),
    .Q_N(_13879_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2354),
    .D(_01459_),
    .Q_N(_13878_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2355),
    .D(_01460_),
    .Q_N(_13877_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2356),
    .D(_01461_),
    .Q_N(_13876_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2357),
    .D(_01462_),
    .Q_N(_13875_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2358),
    .D(_01463_),
    .Q_N(_13874_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2359),
    .D(_01464_),
    .Q_N(_13873_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2360),
    .D(_01465_),
    .Q_N(_13872_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2361),
    .D(_01466_),
    .Q_N(_13871_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2362),
    .D(_01467_),
    .Q_N(_13870_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2363),
    .D(_01468_),
    .Q_N(_13869_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2364),
    .D(_01469_),
    .Q_N(_13868_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net2365),
    .D(_01470_),
    .Q_N(_13867_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2366),
    .D(_01471_),
    .Q_N(_13866_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2367),
    .D(_01472_),
    .Q_N(_13865_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2368),
    .D(_01473_),
    .Q_N(_13864_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net2369),
    .D(_01474_),
    .Q_N(_13863_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2370),
    .D(_01475_),
    .Q_N(_13862_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2371),
    .D(_01476_),
    .Q_N(_13861_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2372),
    .D(_01477_),
    .Q_N(_13860_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net2373),
    .D(_01478_),
    .Q_N(_13859_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2374),
    .D(_01479_),
    .Q_N(_13858_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net2375),
    .D(_01480_),
    .Q_N(_13857_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2376),
    .D(_01481_),
    .Q_N(_13856_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net2377),
    .D(_01482_),
    .Q_N(_13855_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net2378),
    .D(_01483_),
    .Q_N(_13854_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2379),
    .D(_01484_),
    .Q_N(_13853_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2380),
    .D(_01485_),
    .Q_N(_13852_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2381),
    .D(_01486_),
    .Q_N(_13851_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2382),
    .D(_01487_),
    .Q_N(_13850_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net2383),
    .D(_01488_),
    .Q_N(_13849_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2384),
    .D(_01489_),
    .Q_N(_13848_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2385),
    .D(_01490_),
    .Q_N(_13847_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net2386),
    .D(_01491_),
    .Q_N(_13846_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2387),
    .D(_01492_),
    .Q_N(_13845_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2388),
    .D(_01493_),
    .Q_N(_13844_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2389),
    .D(_01494_),
    .Q_N(_13843_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2390),
    .D(_01495_),
    .Q_N(_13842_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2391),
    .D(_01496_),
    .Q_N(_13841_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2392),
    .D(_01497_),
    .Q_N(_13840_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2393),
    .D(_01498_),
    .Q_N(_13839_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2394),
    .D(_01499_),
    .Q_N(_13838_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net2395),
    .D(_01500_),
    .Q_N(_13837_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net2396),
    .D(_01501_),
    .Q_N(_13836_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net2397),
    .D(_01502_),
    .Q_N(_13835_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net2398),
    .D(_01503_),
    .Q_N(_13834_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net2399),
    .D(_01504_),
    .Q_N(_13833_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2400),
    .D(_01505_),
    .Q_N(_13832_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net2401),
    .D(_01506_),
    .Q_N(_13831_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net2402),
    .D(_01507_),
    .Q_N(_13830_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2403),
    .D(_01508_),
    .Q_N(_13829_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net2404),
    .D(_01509_),
    .Q_N(_13828_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net2405),
    .D(_01510_),
    .Q_N(_13827_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2406),
    .D(_01511_),
    .Q_N(_13826_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net2407),
    .D(_01512_),
    .Q_N(_13825_),
    .Q(\cpu.genblk1.mmu.r_vtop_d[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2408),
    .D(_01513_),
    .Q_N(_13824_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2409),
    .D(_01514_),
    .Q_N(_13823_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2410),
    .D(_01515_),
    .Q_N(_13822_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2411),
    .D(_01516_),
    .Q_N(_13821_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2412),
    .D(_01517_),
    .Q_N(_13820_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2413),
    .D(_01518_),
    .Q_N(_13819_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2414),
    .D(_01519_),
    .Q_N(_13818_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2415),
    .D(_01520_),
    .Q_N(_13817_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2416),
    .D(_01521_),
    .Q_N(_13816_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net2417),
    .D(_01522_),
    .Q_N(_13815_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2418),
    .D(_01523_),
    .Q_N(_13814_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2419),
    .D(_01524_),
    .Q_N(_13813_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[0][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2420),
    .D(_01525_),
    .Q_N(_13812_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2421),
    .D(_01526_),
    .Q_N(_13811_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2422),
    .D(_01527_),
    .Q_N(_13810_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2423),
    .D(_01528_),
    .Q_N(_13809_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2424),
    .D(_01529_),
    .Q_N(_13808_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2425),
    .D(_01530_),
    .Q_N(_13807_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2426),
    .D(_01531_),
    .Q_N(_13806_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2427),
    .D(_01532_),
    .Q_N(_13805_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2428),
    .D(_01533_),
    .Q_N(_13804_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2429),
    .D(_01534_),
    .Q_N(_13803_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2430),
    .D(_01535_),
    .Q_N(_13802_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2431),
    .D(_01536_),
    .Q_N(_13801_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[10][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2432),
    .D(_01537_),
    .Q_N(_13800_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2433),
    .D(_01538_),
    .Q_N(_13799_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2434),
    .D(_01539_),
    .Q_N(_13798_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net2435),
    .D(_01540_),
    .Q_N(_13797_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2436),
    .D(_01541_),
    .Q_N(_13796_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2437),
    .D(_01542_),
    .Q_N(_13795_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2438),
    .D(_01543_),
    .Q_N(_13794_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2439),
    .D(_01544_),
    .Q_N(_13793_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2440),
    .D(_01545_),
    .Q_N(_13792_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2441),
    .D(_01546_),
    .Q_N(_13791_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2442),
    .D(_01547_),
    .Q_N(_13790_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2443),
    .D(_01548_),
    .Q_N(_13789_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[11][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2444),
    .D(_01549_),
    .Q_N(_13788_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2445),
    .D(_01550_),
    .Q_N(_13787_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2446),
    .D(_01551_),
    .Q_N(_13786_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2447),
    .D(_01552_),
    .Q_N(_13785_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2448),
    .D(_01553_),
    .Q_N(_13784_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2449),
    .D(_01554_),
    .Q_N(_13783_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2450),
    .D(_01555_),
    .Q_N(_13782_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2451),
    .D(_01556_),
    .Q_N(_13781_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2452),
    .D(_01557_),
    .Q_N(_13780_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2453),
    .D(_01558_),
    .Q_N(_13779_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2454),
    .D(_01559_),
    .Q_N(_13778_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2455),
    .D(_01560_),
    .Q_N(_13777_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[12][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2456),
    .D(_01561_),
    .Q_N(_13776_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2457),
    .D(_01562_),
    .Q_N(_13775_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2458),
    .D(_01563_),
    .Q_N(_13774_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2459),
    .D(_01564_),
    .Q_N(_13773_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2460),
    .D(_01565_),
    .Q_N(_13772_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2461),
    .D(_01566_),
    .Q_N(_13771_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2462),
    .D(_01567_),
    .Q_N(_13770_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2463),
    .D(_01568_),
    .Q_N(_13769_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2464),
    .D(_01569_),
    .Q_N(_13768_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2465),
    .D(_01570_),
    .Q_N(_13767_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2466),
    .D(_01571_),
    .Q_N(_13766_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2467),
    .D(_01572_),
    .Q_N(_13765_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[13][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2468),
    .D(_01573_),
    .Q_N(_13764_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2469),
    .D(_01574_),
    .Q_N(_13763_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2470),
    .D(_01575_),
    .Q_N(_13762_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2471),
    .D(_01576_),
    .Q_N(_13761_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2472),
    .D(_01577_),
    .Q_N(_13760_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2473),
    .D(_01578_),
    .Q_N(_13759_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2474),
    .D(_01579_),
    .Q_N(_13758_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2475),
    .D(_01580_),
    .Q_N(_13757_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2476),
    .D(_01581_),
    .Q_N(_13756_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2477),
    .D(_01582_),
    .Q_N(_13755_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2478),
    .D(_01583_),
    .Q_N(_13754_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2479),
    .D(_01584_),
    .Q_N(_13753_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[14][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2480),
    .D(_01585_),
    .Q_N(_13752_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2481),
    .D(_01586_),
    .Q_N(_13751_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2482),
    .D(_01587_),
    .Q_N(_13750_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2483),
    .D(_01588_),
    .Q_N(_13749_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2484),
    .D(_01589_),
    .Q_N(_13748_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2485),
    .D(_01590_),
    .Q_N(_13747_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2486),
    .D(_01591_),
    .Q_N(_13746_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2487),
    .D(_01592_),
    .Q_N(_13745_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2488),
    .D(_01593_),
    .Q_N(_13744_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net2489),
    .D(_01594_),
    .Q_N(_13743_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2490),
    .D(_01595_),
    .Q_N(_13742_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2491),
    .D(_01596_),
    .Q_N(_13741_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[15][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2492),
    .D(_01597_),
    .Q_N(_13740_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2493),
    .D(_01598_),
    .Q_N(_13739_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2494),
    .D(_01599_),
    .Q_N(_13738_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2495),
    .D(_01600_),
    .Q_N(_13737_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2496),
    .D(_01601_),
    .Q_N(_13736_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2497),
    .D(_01602_),
    .Q_N(_13735_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2498),
    .D(_01603_),
    .Q_N(_13734_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2499),
    .D(_01604_),
    .Q_N(_13733_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2500),
    .D(_01605_),
    .Q_N(_13732_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net2501),
    .D(_01606_),
    .Q_N(_13731_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2502),
    .D(_01607_),
    .Q_N(_13730_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2503),
    .D(_01608_),
    .Q_N(_13729_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[16][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2504),
    .D(_01609_),
    .Q_N(_13728_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net2505),
    .D(_01610_),
    .Q_N(_13727_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2506),
    .D(_01611_),
    .Q_N(_13726_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2507),
    .D(_01612_),
    .Q_N(_13725_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2508),
    .D(_01613_),
    .Q_N(_13724_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2509),
    .D(_01614_),
    .Q_N(_13723_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2510),
    .D(_01615_),
    .Q_N(_13722_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2511),
    .D(_01616_),
    .Q_N(_13721_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net2512),
    .D(_01617_),
    .Q_N(_13720_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2513),
    .D(_01618_),
    .Q_N(_13719_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2514),
    .D(_01619_),
    .Q_N(_13718_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2515),
    .D(_01620_),
    .Q_N(_13717_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[17][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2516),
    .D(_01621_),
    .Q_N(_13716_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2517),
    .D(_01622_),
    .Q_N(_13715_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2518),
    .D(_01623_),
    .Q_N(_13714_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2519),
    .D(_01624_),
    .Q_N(_13713_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2520),
    .D(_01625_),
    .Q_N(_13712_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2521),
    .D(_01626_),
    .Q_N(_13711_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2522),
    .D(_01627_),
    .Q_N(_13710_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2523),
    .D(_01628_),
    .Q_N(_13709_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2524),
    .D(_01629_),
    .Q_N(_13708_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2525),
    .D(_01630_),
    .Q_N(_13707_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2526),
    .D(_01631_),
    .Q_N(_13706_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2527),
    .D(_01632_),
    .Q_N(_13705_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[18][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2528),
    .D(_01633_),
    .Q_N(_13704_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2529),
    .D(_01634_),
    .Q_N(_13703_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2530),
    .D(_01635_),
    .Q_N(_13702_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2531),
    .D(_01636_),
    .Q_N(_13701_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2532),
    .D(_01637_),
    .Q_N(_13700_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2533),
    .D(_01638_),
    .Q_N(_13699_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2534),
    .D(_01639_),
    .Q_N(_13698_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2535),
    .D(_01640_),
    .Q_N(_13697_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2536),
    .D(_01641_),
    .Q_N(_13696_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2537),
    .D(_01642_),
    .Q_N(_13695_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2538),
    .D(_01643_),
    .Q_N(_13694_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2539),
    .D(_01644_),
    .Q_N(_13693_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[19][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2540),
    .D(_01645_),
    .Q_N(_13692_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2541),
    .D(_01646_),
    .Q_N(_13691_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2542),
    .D(_01647_),
    .Q_N(_13690_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2543),
    .D(_01648_),
    .Q_N(_13689_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net2544),
    .D(_01649_),
    .Q_N(_13688_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2545),
    .D(_01650_),
    .Q_N(_13687_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2546),
    .D(_01651_),
    .Q_N(_13686_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2547),
    .D(_01652_),
    .Q_N(_13685_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2548),
    .D(_01653_),
    .Q_N(_13684_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2549),
    .D(_01654_),
    .Q_N(_13683_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2550),
    .D(_01655_),
    .Q_N(_13682_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2551),
    .D(_01656_),
    .Q_N(_13681_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[1][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2552),
    .D(_01657_),
    .Q_N(_13680_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2553),
    .D(_01658_),
    .Q_N(_13679_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2554),
    .D(_01659_),
    .Q_N(_13678_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2555),
    .D(_01660_),
    .Q_N(_13677_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2556),
    .D(_01661_),
    .Q_N(_13676_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2557),
    .D(_01662_),
    .Q_N(_13675_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2558),
    .D(_01663_),
    .Q_N(_13674_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2559),
    .D(_01664_),
    .Q_N(_13673_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2560),
    .D(_01665_),
    .Q_N(_13672_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net2561),
    .D(_01666_),
    .Q_N(_13671_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2562),
    .D(_01667_),
    .Q_N(_13670_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2563),
    .D(_01668_),
    .Q_N(_13669_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[20][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2564),
    .D(_01669_),
    .Q_N(_13668_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net2565),
    .D(_01670_),
    .Q_N(_13667_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2566),
    .D(_01671_),
    .Q_N(_13666_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2567),
    .D(_01672_),
    .Q_N(_13665_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2568),
    .D(_01673_),
    .Q_N(_13664_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2569),
    .D(_01674_),
    .Q_N(_13663_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2570),
    .D(_01675_),
    .Q_N(_13662_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2571),
    .D(_01676_),
    .Q_N(_13661_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2572),
    .D(_01677_),
    .Q_N(_13660_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2573),
    .D(_01678_),
    .Q_N(_13659_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2574),
    .D(_01679_),
    .Q_N(_13658_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2575),
    .D(_01680_),
    .Q_N(_13657_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[21][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2576),
    .D(_01681_),
    .Q_N(_13656_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2577),
    .D(_01682_),
    .Q_N(_13655_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2578),
    .D(_01683_),
    .Q_N(_13654_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2579),
    .D(_01684_),
    .Q_N(_13653_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2580),
    .D(_01685_),
    .Q_N(_13652_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2581),
    .D(_01686_),
    .Q_N(_13651_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2582),
    .D(_01687_),
    .Q_N(_13650_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2583),
    .D(_01688_),
    .Q_N(_13649_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2584),
    .D(_01689_),
    .Q_N(_13648_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2585),
    .D(_01690_),
    .Q_N(_13647_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2586),
    .D(_01691_),
    .Q_N(_13646_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2587),
    .D(_01692_),
    .Q_N(_13645_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[22][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2588),
    .D(_01693_),
    .Q_N(_13644_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2589),
    .D(_01694_),
    .Q_N(_13643_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2590),
    .D(_01695_),
    .Q_N(_13642_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net2591),
    .D(_01696_),
    .Q_N(_13641_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net2592),
    .D(_01697_),
    .Q_N(_13640_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net2593),
    .D(_01698_),
    .Q_N(_13639_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2594),
    .D(_01699_),
    .Q_N(_13638_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net2595),
    .D(_01700_),
    .Q_N(_13637_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2596),
    .D(_01701_),
    .Q_N(_13636_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net2597),
    .D(_01702_),
    .Q_N(_13635_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2598),
    .D(_01703_),
    .Q_N(_13634_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2599),
    .D(_01704_),
    .Q_N(_13633_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[23][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2600),
    .D(_01705_),
    .Q_N(_13632_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2601),
    .D(_01706_),
    .Q_N(_13631_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2602),
    .D(_01707_),
    .Q_N(_13630_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2603),
    .D(_01708_),
    .Q_N(_13629_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2604),
    .D(_01709_),
    .Q_N(_13628_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2605),
    .D(_01710_),
    .Q_N(_13627_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2606),
    .D(_01711_),
    .Q_N(_13626_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2607),
    .D(_01712_),
    .Q_N(_13625_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net2608),
    .D(_01713_),
    .Q_N(_13624_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2609),
    .D(_01714_),
    .Q_N(_13623_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2610),
    .D(_01715_),
    .Q_N(_13622_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2611),
    .D(_01716_),
    .Q_N(_13621_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[24][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2612),
    .D(_01717_),
    .Q_N(_13620_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net2613),
    .D(_01718_),
    .Q_N(_13619_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2614),
    .D(_01719_),
    .Q_N(_13618_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2615),
    .D(_01720_),
    .Q_N(_13617_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2616),
    .D(_01721_),
    .Q_N(_13616_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2617),
    .D(_01722_),
    .Q_N(_13615_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2618),
    .D(_01723_),
    .Q_N(_13614_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2619),
    .D(_01724_),
    .Q_N(_13613_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2620),
    .D(_01725_),
    .Q_N(_13612_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2621),
    .D(_01726_),
    .Q_N(_13611_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2622),
    .D(_01727_),
    .Q_N(_13610_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2623),
    .D(_01728_),
    .Q_N(_13609_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[25][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2624),
    .D(_01729_),
    .Q_N(_13608_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net2625),
    .D(_01730_),
    .Q_N(_13607_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2626),
    .D(_01731_),
    .Q_N(_13606_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2627),
    .D(_01732_),
    .Q_N(_13605_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2628),
    .D(_01733_),
    .Q_N(_13604_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2629),
    .D(_01734_),
    .Q_N(_13603_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2630),
    .D(_01735_),
    .Q_N(_13602_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2631),
    .D(_01736_),
    .Q_N(_13601_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2632),
    .D(_01737_),
    .Q_N(_13600_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2633),
    .D(_01738_),
    .Q_N(_13599_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net2634),
    .D(_01739_),
    .Q_N(_13598_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2635),
    .D(_01740_),
    .Q_N(_13597_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[26][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2636),
    .D(_01741_),
    .Q_N(_13596_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2637),
    .D(_01742_),
    .Q_N(_13595_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2638),
    .D(_01743_),
    .Q_N(_13594_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net2639),
    .D(_01744_),
    .Q_N(_13593_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net2640),
    .D(_01745_),
    .Q_N(_13592_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2641),
    .D(_01746_),
    .Q_N(_13591_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net2642),
    .D(_01747_),
    .Q_N(_13590_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2643),
    .D(_01748_),
    .Q_N(_13589_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net2644),
    .D(_01749_),
    .Q_N(_13588_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2645),
    .D(_01750_),
    .Q_N(_13587_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net2646),
    .D(_01751_),
    .Q_N(_13586_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2647),
    .D(_01752_),
    .Q_N(_13585_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[27][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2648),
    .D(_01753_),
    .Q_N(_13584_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2649),
    .D(_01754_),
    .Q_N(_13583_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2650),
    .D(_01755_),
    .Q_N(_13582_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2651),
    .D(_01756_),
    .Q_N(_13581_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2652),
    .D(_01757_),
    .Q_N(_13580_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2653),
    .D(_01758_),
    .Q_N(_13579_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2654),
    .D(_01759_),
    .Q_N(_13578_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2655),
    .D(_01760_),
    .Q_N(_13577_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2656),
    .D(_01761_),
    .Q_N(_13576_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net2657),
    .D(_01762_),
    .Q_N(_13575_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2658),
    .D(_01763_),
    .Q_N(_13574_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net2659),
    .D(_01764_),
    .Q_N(_13573_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[28][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2660),
    .D(_01765_),
    .Q_N(_13572_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2661),
    .D(_01766_),
    .Q_N(_13571_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2662),
    .D(_01767_),
    .Q_N(_13570_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2663),
    .D(_01768_),
    .Q_N(_13569_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2664),
    .D(_01769_),
    .Q_N(_13568_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2665),
    .D(_01770_),
    .Q_N(_13567_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2666),
    .D(_01771_),
    .Q_N(_13566_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2667),
    .D(_01772_),
    .Q_N(_13565_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net2668),
    .D(_01773_),
    .Q_N(_13564_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2669),
    .D(_01774_),
    .Q_N(_13563_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2670),
    .D(_01775_),
    .Q_N(_13562_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2671),
    .D(_01776_),
    .Q_N(_13561_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[29][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2672),
    .D(_01777_),
    .Q_N(_13560_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2673),
    .D(_01778_),
    .Q_N(_13559_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2674),
    .D(_01779_),
    .Q_N(_13558_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2675),
    .D(_01780_),
    .Q_N(_13557_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2676),
    .D(_01781_),
    .Q_N(_13556_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2677),
    .D(_01782_),
    .Q_N(_13555_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2678),
    .D(_01783_),
    .Q_N(_13554_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2679),
    .D(_01784_),
    .Q_N(_13553_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2680),
    .D(_01785_),
    .Q_N(_13552_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2681),
    .D(_01786_),
    .Q_N(_13551_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2682),
    .D(_01787_),
    .Q_N(_13550_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2683),
    .D(_01788_),
    .Q_N(_13549_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[2][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2684),
    .D(_01789_),
    .Q_N(_13548_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net2685),
    .D(_01790_),
    .Q_N(_13547_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2686),
    .D(_01791_),
    .Q_N(_13546_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2687),
    .D(_01792_),
    .Q_N(_13545_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2688),
    .D(_01793_),
    .Q_N(_13544_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2689),
    .D(_01794_),
    .Q_N(_13543_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2690),
    .D(_01795_),
    .Q_N(_13542_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2691),
    .D(_01796_),
    .Q_N(_13541_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2692),
    .D(_01797_),
    .Q_N(_13540_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2693),
    .D(_01798_),
    .Q_N(_13539_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2694),
    .D(_01799_),
    .Q_N(_13538_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2695),
    .D(_01800_),
    .Q_N(_13537_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[30][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net2696),
    .D(_01801_),
    .Q_N(_13536_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net2697),
    .D(_01802_),
    .Q_N(_13535_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net2698),
    .D(_01803_),
    .Q_N(_13534_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net2699),
    .D(_01804_),
    .Q_N(_13533_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net2700),
    .D(_01805_),
    .Q_N(_13532_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net2701),
    .D(_01806_),
    .Q_N(_13531_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2702),
    .D(_01807_),
    .Q_N(_13530_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net2703),
    .D(_01808_),
    .Q_N(_13529_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net2704),
    .D(_01809_),
    .Q_N(_13528_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2705),
    .D(_01810_),
    .Q_N(_13527_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2706),
    .D(_01811_),
    .Q_N(_13526_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net2707),
    .D(_01812_),
    .Q_N(_13525_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[31][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2708),
    .D(_01813_),
    .Q_N(_13524_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2709),
    .D(_01814_),
    .Q_N(_13523_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net2710),
    .D(_01815_),
    .Q_N(_13522_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2711),
    .D(_01816_),
    .Q_N(_13521_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net2712),
    .D(_01817_),
    .Q_N(_13520_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net2713),
    .D(_01818_),
    .Q_N(_13519_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2714),
    .D(_01819_),
    .Q_N(_13518_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net2715),
    .D(_01820_),
    .Q_N(_13517_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net2716),
    .D(_01821_),
    .Q_N(_13516_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net2717),
    .D(_01822_),
    .Q_N(_13515_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net2718),
    .D(_01823_),
    .Q_N(_13514_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2719),
    .D(_01824_),
    .Q_N(_13513_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[3][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net2720),
    .D(_01825_),
    .Q_N(_13512_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2721),
    .D(_01826_),
    .Q_N(_13511_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2722),
    .D(_01827_),
    .Q_N(_13510_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_42_clk),
    .RESET_B(net2723),
    .D(_01828_),
    .Q_N(_13509_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2724),
    .D(_01829_),
    .Q_N(_13508_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2725),
    .D(_01830_),
    .Q_N(_13507_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2726),
    .D(_01831_),
    .Q_N(_13506_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2727),
    .D(_01832_),
    .Q_N(_13505_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2728),
    .D(_01833_),
    .Q_N(_13504_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2729),
    .D(_01834_),
    .Q_N(_13503_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2730),
    .D(_01835_),
    .Q_N(_13502_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2731),
    .D(_01836_),
    .Q_N(_13501_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[4][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2732),
    .D(_01837_),
    .Q_N(_13500_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2733),
    .D(_01838_),
    .Q_N(_13499_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2734),
    .D(_01839_),
    .Q_N(_13498_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2735),
    .D(_01840_),
    .Q_N(_13497_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2736),
    .D(_01841_),
    .Q_N(_13496_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2737),
    .D(_01842_),
    .Q_N(_13495_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2738),
    .D(_01843_),
    .Q_N(_13494_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2739),
    .D(_01844_),
    .Q_N(_13493_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2740),
    .D(_01845_),
    .Q_N(_13492_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2741),
    .D(_01846_),
    .Q_N(_13491_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net2742),
    .D(_01847_),
    .Q_N(_13490_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2743),
    .D(_01848_),
    .Q_N(_13489_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[5][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2744),
    .D(_01849_),
    .Q_N(_13488_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net2745),
    .D(_01850_),
    .Q_N(_13487_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2746),
    .D(_01851_),
    .Q_N(_13486_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2747),
    .D(_01852_),
    .Q_N(_13485_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2748),
    .D(_01853_),
    .Q_N(_13484_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2749),
    .D(_01854_),
    .Q_N(_13483_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2750),
    .D(_01855_),
    .Q_N(_13482_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2751),
    .D(_01856_),
    .Q_N(_13481_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2752),
    .D(_01857_),
    .Q_N(_13480_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2753),
    .D(_01858_),
    .Q_N(_13479_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2754),
    .D(_01859_),
    .Q_N(_13478_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2755),
    .D(_01860_),
    .Q_N(_13477_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[6][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2756),
    .D(_01861_),
    .Q_N(_13476_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2757),
    .D(_01862_),
    .Q_N(_13475_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2758),
    .D(_01863_),
    .Q_N(_13474_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2759),
    .D(_01864_),
    .Q_N(_13473_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2760),
    .D(_01865_),
    .Q_N(_13472_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net2761),
    .D(_01866_),
    .Q_N(_13471_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2762),
    .D(_01867_),
    .Q_N(_13470_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_41_clk),
    .RESET_B(net2763),
    .D(_01868_),
    .Q_N(_13469_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net2764),
    .D(_01869_),
    .Q_N(_13468_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net2765),
    .D(_01870_),
    .Q_N(_13467_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2766),
    .D(_01871_),
    .Q_N(_13466_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net2767),
    .D(_01872_),
    .Q_N(_13465_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[7][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2768),
    .D(_01873_),
    .Q_N(_13464_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2769),
    .D(_01874_),
    .Q_N(_13463_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_39_clk),
    .RESET_B(net2770),
    .D(_01875_),
    .Q_N(_13462_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2771),
    .D(_01876_),
    .Q_N(_13461_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2772),
    .D(_01877_),
    .Q_N(_13460_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2773),
    .D(_01878_),
    .Q_N(_13459_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2774),
    .D(_01879_),
    .Q_N(_13458_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net2775),
    .D(_01880_),
    .Q_N(_13457_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2776),
    .D(_01881_),
    .Q_N(_13456_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2777),
    .D(_01882_),
    .Q_N(_13455_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net2778),
    .D(_01883_),
    .Q_N(_13454_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net2779),
    .D(_01884_),
    .Q_N(_13453_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[8][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net2780),
    .D(_01885_),
    .Q_N(_13452_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2781),
    .D(_01886_),
    .Q_N(_13451_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2782),
    .D(_01887_),
    .Q_N(_13450_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net2783),
    .D(_01888_),
    .Q_N(_13449_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net2784),
    .D(_01889_),
    .Q_N(_13448_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net2785),
    .D(_01890_),
    .Q_N(_13447_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net2786),
    .D(_01891_),
    .Q_N(_13446_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net2787),
    .D(_01892_),
    .Q_N(_13445_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net2788),
    .D(_01893_),
    .Q_N(_13444_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net2789),
    .D(_01894_),
    .Q_N(_13443_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net2790),
    .D(_01895_),
    .Q_N(_13442_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net2791),
    .D(_01896_),
    .Q_N(_13441_),
    .Q(\cpu.genblk1.mmu.r_vtop_i[9][9] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2792),
    .D(_01897_),
    .Q_N(_13440_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[0] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2793),
    .D(_01898_),
    .Q_N(_13439_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[10] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2794),
    .D(_01899_),
    .Q_N(_13438_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[11] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2795),
    .D(_01900_),
    .Q_N(_13437_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[12] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2796),
    .D(_01901_),
    .Q_N(_13436_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[13] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2797),
    .D(_01902_),
    .Q_N(_13435_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[14] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2798),
    .D(_01903_),
    .Q_N(_13434_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[15] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2799),
    .D(_01904_),
    .Q_N(_13433_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[16] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2800),
    .D(_01905_),
    .Q_N(_13432_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[17] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2801),
    .D(_01906_),
    .Q_N(_13431_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[18] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2802),
    .D(_01907_),
    .Q_N(_13430_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[19] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2803),
    .D(_01908_),
    .Q_N(_13429_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[1] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2804),
    .D(_01909_),
    .Q_N(_13428_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[20] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net2805),
    .D(_01910_),
    .Q_N(_13427_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[21] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2806),
    .D(_01911_),
    .Q_N(_13426_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[22] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net2807),
    .D(_01912_),
    .Q_N(_13425_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[23] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2808),
    .D(_01913_),
    .Q_N(_13424_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[24] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2809),
    .D(_01914_),
    .Q_N(_13423_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[25] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2810),
    .D(_01915_),
    .Q_N(_13422_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[26] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net2811),
    .D(_01916_),
    .Q_N(_13421_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[27] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net2812),
    .D(_01917_),
    .Q_N(_13420_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[28] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net2813),
    .D(_01918_),
    .Q_N(_13419_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[29] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net2814),
    .D(_01919_),
    .Q_N(_13418_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[2] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2815),
    .D(_01920_),
    .Q_N(_13417_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[30] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net2816),
    .D(_01921_),
    .Q_N(_13416_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[31] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2817),
    .D(_01922_),
    .Q_N(_13415_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[3] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2818),
    .D(_01923_),
    .Q_N(_13414_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[4] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net2819),
    .D(_01924_),
    .Q_N(_13413_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[5] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net2820),
    .D(_01925_),
    .Q_N(_13412_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[6] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net2821),
    .D(_01926_),
    .Q_N(_13411_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[7] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net2822),
    .D(_01927_),
    .Q_N(_13410_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[8] ));
 sg13g2_dfrbp_1 \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net2823),
    .D(_01928_),
    .Q_N(_13409_),
    .Q(\cpu.genblk1.mmu.r_writeable_d[9] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2824),
    .D(_01929_),
    .Q_N(_13408_),
    .Q(\cpu.gpio.r_enable_in[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2825),
    .D(_01930_),
    .Q_N(_13407_),
    .Q(\cpu.gpio.r_enable_in[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2826),
    .D(_01931_),
    .Q_N(_13406_),
    .Q(\cpu.gpio.r_enable_in[2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2827),
    .D(_01932_),
    .Q_N(_13405_),
    .Q(\cpu.gpio.r_enable_in[3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2828),
    .D(_01933_),
    .Q_N(_13404_),
    .Q(\cpu.gpio.r_enable_in[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net2829),
    .D(_01934_),
    .Q_N(_13403_),
    .Q(\cpu.gpio.r_enable_in[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2830),
    .D(_01935_),
    .Q_N(_13402_),
    .Q(\cpu.gpio.r_enable_in[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net2831),
    .D(_01936_),
    .Q_N(_13401_),
    .Q(\cpu.gpio.r_enable_in[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2832),
    .D(_01937_),
    .Q_N(_13400_),
    .Q(\cpu.gpio.r_enable_io[4] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2833),
    .D(_01938_),
    .Q_N(_13399_),
    .Q(\cpu.gpio.r_enable_io[5] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2834),
    .D(_01939_),
    .Q_N(_13398_),
    .Q(\cpu.gpio.r_enable_io[6] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2835),
    .D(_01940_),
    .Q_N(_13397_),
    .Q(\cpu.gpio.r_enable_io[7] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2836),
    .D(_01941_),
    .Q_N(_13396_),
    .Q(net7));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2837),
    .D(_01942_),
    .Q_N(_13395_),
    .Q(net8));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2838),
    .D(_01943_),
    .Q_N(_13394_),
    .Q(net9));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2839),
    .D(_01944_),
    .Q_N(_13393_),
    .Q(net10));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2840),
    .D(_01945_),
    .Q_N(_13392_),
    .Q(\cpu.gpio.genblk2[4].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2841),
    .D(_01946_),
    .Q_N(_13391_),
    .Q(\cpu.gpio.genblk2[5].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2842),
    .D(_01947_),
    .Q_N(_13390_),
    .Q(\cpu.gpio.genblk2[6].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_io[3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2843),
    .D(_01948_),
    .Q_N(_13389_),
    .Q(\cpu.gpio.genblk2[7].srcs_io[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[0]$_DFFE_PP_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2844),
    .D(_01949_),
    .Q_N(_13388_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[1]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2845),
    .D(_01950_),
    .Q_N(_13387_),
    .Q(\cpu.gpio.genblk1[4].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[2]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2846),
    .D(_01951_),
    .Q_N(_13386_),
    .Q(\cpu.gpio.genblk1[5].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[3]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net2847),
    .D(_01952_),
    .Q_N(_13385_),
    .Q(\cpu.gpio.genblk1[6].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_gpio_o[4]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2848),
    .D(_01953_),
    .Q_N(_13384_),
    .Q(\cpu.gpio.genblk1[7].srcs_o[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2849),
    .D(_01954_),
    .Q_N(_13383_),
    .Q(\cpu.gpio.r_spi_miso_src[0][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2850),
    .D(_01955_),
    .Q_N(_00305_),
    .Q(\cpu.gpio.r_spi_miso_src[0][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2851),
    .D(_01956_),
    .Q_N(_00102_),
    .Q(\cpu.gpio.r_spi_miso_src[0][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net2852),
    .D(_01957_),
    .Q_N(_00112_),
    .Q(\cpu.gpio.r_spi_miso_src[0][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2853),
    .D(_01958_),
    .Q_N(_13382_),
    .Q(\cpu.gpio.r_spi_miso_src[1][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2854),
    .D(_01959_),
    .Q_N(_00131_),
    .Q(\cpu.gpio.r_spi_miso_src[1][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2855),
    .D(_01960_),
    .Q_N(_00143_),
    .Q(\cpu.gpio.r_spi_miso_src[1][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net2856),
    .D(_01961_),
    .Q_N(_00155_),
    .Q(\cpu.gpio.r_spi_miso_src[1][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2857),
    .D(_01962_),
    .Q_N(_13381_),
    .Q(\cpu.gpio.r_src_io[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2858),
    .D(_01963_),
    .Q_N(_13380_),
    .Q(\cpu.gpio.r_src_io[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2859),
    .D(_01964_),
    .Q_N(_00185_),
    .Q(\cpu.gpio.r_src_io[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2860),
    .D(_01965_),
    .Q_N(_13379_),
    .Q(\cpu.gpio.r_src_io[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2861),
    .D(_01966_),
    .Q_N(_13378_),
    .Q(\cpu.gpio.r_src_io[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2862),
    .D(_01967_),
    .Q_N(_13377_),
    .Q(\cpu.gpio.r_src_io[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2863),
    .D(_01968_),
    .Q_N(_00184_),
    .Q(\cpu.gpio.r_src_io[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net2864),
    .D(_01969_),
    .Q_N(_13376_),
    .Q(\cpu.gpio.r_src_io[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2865),
    .D(_01970_),
    .Q_N(_13375_),
    .Q(\cpu.gpio.r_src_io[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2866),
    .D(_01971_),
    .Q_N(_00301_),
    .Q(\cpu.gpio.r_src_io[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2867),
    .D(_01972_),
    .Q_N(_00098_),
    .Q(\cpu.gpio.r_src_io[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2868),
    .D(_01973_),
    .Q_N(_00109_),
    .Q(\cpu.gpio.r_src_io[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2869),
    .D(_01974_),
    .Q_N(_13374_),
    .Q(\cpu.gpio.r_src_io[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2870),
    .D(_01975_),
    .Q_N(_00127_),
    .Q(\cpu.gpio.r_src_io[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net2871),
    .D(_01976_),
    .Q_N(_00139_),
    .Q(\cpu.gpio.r_src_io[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_io[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2872),
    .D(_01977_),
    .Q_N(_00151_),
    .Q(\cpu.gpio.r_src_io[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2873),
    .D(_01978_),
    .Q_N(_13373_),
    .Q(\cpu.gpio.r_src_o[3][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2874),
    .D(_01979_),
    .Q_N(_00130_),
    .Q(\cpu.gpio.r_src_o[3][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2875),
    .D(_01980_),
    .Q_N(_00142_),
    .Q(\cpu.gpio.r_src_o[3][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2876),
    .D(_01981_),
    .Q_N(_00154_),
    .Q(\cpu.gpio.r_src_o[3][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2877),
    .D(_01982_),
    .Q_N(_13372_),
    .Q(\cpu.gpio.r_src_o[4][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2878),
    .D(_01983_),
    .Q_N(_00303_),
    .Q(\cpu.gpio.r_src_o[4][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2879),
    .D(_01984_),
    .Q_N(_00100_),
    .Q(\cpu.gpio.r_src_o[4][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2880),
    .D(_01985_),
    .Q_N(_00111_),
    .Q(\cpu.gpio.r_src_o[4][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2881),
    .D(_01986_),
    .Q_N(_13371_),
    .Q(\cpu.gpio.r_src_o[5][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2882),
    .D(_01987_),
    .Q_N(_00129_),
    .Q(\cpu.gpio.r_src_o[5][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net2883),
    .D(_01988_),
    .Q_N(_00141_),
    .Q(\cpu.gpio.r_src_o[5][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2884),
    .D(_01989_),
    .Q_N(_00153_),
    .Q(\cpu.gpio.r_src_o[5][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2885),
    .D(_01990_),
    .Q_N(_13370_),
    .Q(\cpu.gpio.r_src_o[6][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2886),
    .D(_01991_),
    .Q_N(_00302_),
    .Q(\cpu.gpio.r_src_o[6][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net2887),
    .D(_01992_),
    .Q_N(_00099_),
    .Q(\cpu.gpio.r_src_o[6][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net2888),
    .D(_01993_),
    .Q_N(_00110_),
    .Q(\cpu.gpio.r_src_o[6][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2889),
    .D(_01994_),
    .Q_N(_13369_),
    .Q(\cpu.gpio.r_src_o[7][0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net2890),
    .D(_01995_),
    .Q_N(_00128_),
    .Q(\cpu.gpio.r_src_o[7][1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2891),
    .D(_01996_),
    .Q_N(_00140_),
    .Q(\cpu.gpio.r_src_o[7][2] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_src_o[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net2892),
    .D(_01997_),
    .Q_N(_00152_),
    .Q(\cpu.gpio.r_src_o[7][3] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2893),
    .D(_01998_),
    .Q_N(_13368_),
    .Q(\cpu.gpio.r_uart_rx_src[0] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2894),
    .D(_01999_),
    .Q_N(_00304_),
    .Q(\cpu.gpio.r_uart_rx_src[1] ));
 sg13g2_dfrbp_1 \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net2895),
    .D(_02000_),
    .Q_N(_00101_),
    .Q(\cpu.gpio.r_uart_rx_src[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2896),
    .D(_02001_),
    .Q_N(_13367_),
    .Q(\cpu.icache.r_data[0][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2897),
    .D(_02002_),
    .Q_N(_00199_),
    .Q(\cpu.icache.r_data[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2898),
    .D(_02003_),
    .Q_N(_00201_),
    .Q(\cpu.icache.r_data[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2899),
    .D(_02004_),
    .Q_N(_00211_),
    .Q(\cpu.icache.r_data[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2900),
    .D(_02005_),
    .Q_N(_13366_),
    .Q(\cpu.icache.r_data[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2901),
    .D(_02006_),
    .Q_N(_00203_),
    .Q(\cpu.icache.r_data[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2902),
    .D(_02007_),
    .Q_N(_00205_),
    .Q(\cpu.icache.r_data[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2903),
    .D(_02008_),
    .Q_N(_13365_),
    .Q(\cpu.icache.r_data[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2904),
    .D(_02009_),
    .Q_N(_13364_),
    .Q(\cpu.icache.r_data[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2905),
    .D(_02010_),
    .Q_N(_00171_),
    .Q(\cpu.icache.r_data[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][19]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2906),
    .D(_02011_),
    .Q_N(_00173_),
    .Q(\cpu.icache.r_data[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2907),
    .D(_02012_),
    .Q_N(_13363_),
    .Q(\cpu.icache.r_data[0][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][20]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2908),
    .D(_02013_),
    .Q_N(_00175_),
    .Q(\cpu.icache.r_data[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][21]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2909),
    .D(_02014_),
    .Q_N(_00208_),
    .Q(\cpu.icache.r_data[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][22]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2910),
    .D(_02015_),
    .Q_N(_00210_),
    .Q(\cpu.icache.r_data[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][23]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2911),
    .D(_02016_),
    .Q_N(_00165_),
    .Q(\cpu.icache.r_data[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][24]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2912),
    .D(_02017_),
    .Q_N(_00167_),
    .Q(\cpu.icache.r_data[0][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2913),
    .D(_02018_),
    .Q_N(_00169_),
    .Q(\cpu.icache.r_data[0][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][26]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2914),
    .D(_02019_),
    .Q_N(_00200_),
    .Q(\cpu.icache.r_data[0][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][27]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net2915),
    .D(_02020_),
    .Q_N(_00202_),
    .Q(\cpu.icache.r_data[0][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][28]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2916),
    .D(_02021_),
    .Q_N(_00212_),
    .Q(\cpu.icache.r_data[0][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][29]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2917),
    .D(_02022_),
    .Q_N(_13362_),
    .Q(\cpu.icache.r_data[0][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2918),
    .D(_02023_),
    .Q_N(_00170_),
    .Q(\cpu.icache.r_data[0][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2919),
    .D(_02024_),
    .Q_N(_00204_),
    .Q(\cpu.icache.r_data[0][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][31]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2920),
    .D(_02025_),
    .Q_N(_00206_),
    .Q(\cpu.icache.r_data[0][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net2921),
    .D(_02026_),
    .Q_N(_00172_),
    .Q(\cpu.icache.r_data[0][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2922),
    .D(_02027_),
    .Q_N(_00174_),
    .Q(\cpu.icache.r_data[0][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2923),
    .D(_02028_),
    .Q_N(_00207_),
    .Q(\cpu.icache.r_data[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2924),
    .D(_02029_),
    .Q_N(_00209_),
    .Q(\cpu.icache.r_data[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2925),
    .D(_02030_),
    .Q_N(_00164_),
    .Q(\cpu.icache.r_data[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net2926),
    .D(_02031_),
    .Q_N(_00166_),
    .Q(\cpu.icache.r_data[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2927),
    .D(_02032_),
    .Q_N(_00168_),
    .Q(\cpu.icache.r_data[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net2928),
    .D(_02033_),
    .Q_N(_13361_),
    .Q(\cpu.icache.r_data[1][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2929),
    .D(_02034_),
    .Q_N(_13360_),
    .Q(\cpu.icache.r_data[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2930),
    .D(_02035_),
    .Q_N(_13359_),
    .Q(\cpu.icache.r_data[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2931),
    .D(_02036_),
    .Q_N(_13358_),
    .Q(\cpu.icache.r_data[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2932),
    .D(_02037_),
    .Q_N(_13357_),
    .Q(\cpu.icache.r_data[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net2933),
    .D(_02038_),
    .Q_N(_13356_),
    .Q(\cpu.icache.r_data[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2934),
    .D(_02039_),
    .Q_N(_13355_),
    .Q(\cpu.icache.r_data[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2935),
    .D(_02040_),
    .Q_N(_13354_),
    .Q(\cpu.icache.r_data[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2936),
    .D(_02041_),
    .Q_N(_13353_),
    .Q(\cpu.icache.r_data[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2937),
    .D(_02042_),
    .Q_N(_13352_),
    .Q(\cpu.icache.r_data[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][19]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net2938),
    .D(_02043_),
    .Q_N(_13351_),
    .Q(\cpu.icache.r_data[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2939),
    .D(_02044_),
    .Q_N(_13350_),
    .Q(\cpu.icache.r_data[1][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net2940),
    .D(_02045_),
    .Q_N(_13349_),
    .Q(\cpu.icache.r_data[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][21]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2941),
    .D(_02046_),
    .Q_N(_13348_),
    .Q(\cpu.icache.r_data[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][22]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2942),
    .D(_02047_),
    .Q_N(_13347_),
    .Q(\cpu.icache.r_data[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][23]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2943),
    .D(_02048_),
    .Q_N(_13346_),
    .Q(\cpu.icache.r_data[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][24]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2944),
    .D(_02049_),
    .Q_N(_13345_),
    .Q(\cpu.icache.r_data[1][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][25]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net2945),
    .D(_02050_),
    .Q_N(_13344_),
    .Q(\cpu.icache.r_data[1][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2946),
    .D(_02051_),
    .Q_N(_13343_),
    .Q(\cpu.icache.r_data[1][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][27]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2947),
    .D(_02052_),
    .Q_N(_13342_),
    .Q(\cpu.icache.r_data[1][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][28]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2948),
    .D(_02053_),
    .Q_N(_13341_),
    .Q(\cpu.icache.r_data[1][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][29]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2949),
    .D(_02054_),
    .Q_N(_13340_),
    .Q(\cpu.icache.r_data[1][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2950),
    .D(_02055_),
    .Q_N(_13339_),
    .Q(\cpu.icache.r_data[1][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net2951),
    .D(_02056_),
    .Q_N(_13338_),
    .Q(\cpu.icache.r_data[1][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][31]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2952),
    .D(_02057_),
    .Q_N(_13337_),
    .Q(\cpu.icache.r_data[1][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2953),
    .D(_02058_),
    .Q_N(_13336_),
    .Q(\cpu.icache.r_data[1][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2954),
    .D(_02059_),
    .Q_N(_13335_),
    .Q(\cpu.icache.r_data[1][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2955),
    .D(_02060_),
    .Q_N(_13334_),
    .Q(\cpu.icache.r_data[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2956),
    .D(_02061_),
    .Q_N(_13333_),
    .Q(\cpu.icache.r_data[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2957),
    .D(_02062_),
    .Q_N(_13332_),
    .Q(\cpu.icache.r_data[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2958),
    .D(_02063_),
    .Q_N(_13331_),
    .Q(\cpu.icache.r_data[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net2959),
    .D(_02064_),
    .Q_N(_13330_),
    .Q(\cpu.icache.r_data[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2960),
    .D(_02065_),
    .Q_N(_13329_),
    .Q(\cpu.icache.r_data[2][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2961),
    .D(_02066_),
    .Q_N(_13328_),
    .Q(\cpu.icache.r_data[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2962),
    .D(_02067_),
    .Q_N(_13327_),
    .Q(\cpu.icache.r_data[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2963),
    .D(_02068_),
    .Q_N(_13326_),
    .Q(\cpu.icache.r_data[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net2964),
    .D(_02069_),
    .Q_N(_13325_),
    .Q(\cpu.icache.r_data[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2965),
    .D(_02070_),
    .Q_N(_13324_),
    .Q(\cpu.icache.r_data[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net2966),
    .D(_02071_),
    .Q_N(_13323_),
    .Q(\cpu.icache.r_data[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net2967),
    .D(_02072_),
    .Q_N(_13322_),
    .Q(\cpu.icache.r_data[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2968),
    .D(_02073_),
    .Q_N(_13321_),
    .Q(\cpu.icache.r_data[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2969),
    .D(_02074_),
    .Q_N(_13320_),
    .Q(\cpu.icache.r_data[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][19]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net2970),
    .D(_02075_),
    .Q_N(_13319_),
    .Q(\cpu.icache.r_data[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2971),
    .D(_02076_),
    .Q_N(_13318_),
    .Q(\cpu.icache.r_data[2][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][20]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2972),
    .D(_02077_),
    .Q_N(_13317_),
    .Q(\cpu.icache.r_data[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][21]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2973),
    .D(_02078_),
    .Q_N(_13316_),
    .Q(\cpu.icache.r_data[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][22]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net2974),
    .D(_02079_),
    .Q_N(_13315_),
    .Q(\cpu.icache.r_data[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][23]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net2975),
    .D(_02080_),
    .Q_N(_13314_),
    .Q(\cpu.icache.r_data[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][24]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2976),
    .D(_02081_),
    .Q_N(_13313_),
    .Q(\cpu.icache.r_data[2][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][25]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2977),
    .D(_02082_),
    .Q_N(_13312_),
    .Q(\cpu.icache.r_data[2][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][26]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2978),
    .D(_02083_),
    .Q_N(_13311_),
    .Q(\cpu.icache.r_data[2][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][27]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net2979),
    .D(_02084_),
    .Q_N(_13310_),
    .Q(\cpu.icache.r_data[2][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][28]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net2980),
    .D(_02085_),
    .Q_N(_13309_),
    .Q(\cpu.icache.r_data[2][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][29]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net2981),
    .D(_02086_),
    .Q_N(_13308_),
    .Q(\cpu.icache.r_data[2][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net2982),
    .D(_02087_),
    .Q_N(_13307_),
    .Q(\cpu.icache.r_data[2][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][30]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2983),
    .D(_02088_),
    .Q_N(_13306_),
    .Q(\cpu.icache.r_data[2][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][31]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2984),
    .D(_02089_),
    .Q_N(_13305_),
    .Q(\cpu.icache.r_data[2][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2985),
    .D(_02090_),
    .Q_N(_13304_),
    .Q(\cpu.icache.r_data[2][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2986),
    .D(_02091_),
    .Q_N(_13303_),
    .Q(\cpu.icache.r_data[2][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2987),
    .D(_02092_),
    .Q_N(_13302_),
    .Q(\cpu.icache.r_data[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net2988),
    .D(_02093_),
    .Q_N(_13301_),
    .Q(\cpu.icache.r_data[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net2989),
    .D(_02094_),
    .Q_N(_13300_),
    .Q(\cpu.icache.r_data[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2990),
    .D(_02095_),
    .Q_N(_13299_),
    .Q(\cpu.icache.r_data[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net2991),
    .D(_02096_),
    .Q_N(_13298_),
    .Q(\cpu.icache.r_data[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net2992),
    .D(_02097_),
    .Q_N(_13297_),
    .Q(\cpu.icache.r_data[3][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net2993),
    .D(_02098_),
    .Q_N(_13296_),
    .Q(\cpu.icache.r_data[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net2994),
    .D(_02099_),
    .Q_N(_13295_),
    .Q(\cpu.icache.r_data[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2995),
    .D(_02100_),
    .Q_N(_13294_),
    .Q(\cpu.icache.r_data[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2996),
    .D(_02101_),
    .Q_N(_13293_),
    .Q(\cpu.icache.r_data[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net2997),
    .D(_02102_),
    .Q_N(_13292_),
    .Q(\cpu.icache.r_data[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2998),
    .D(_02103_),
    .Q_N(_13291_),
    .Q(\cpu.icache.r_data[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net2999),
    .D(_02104_),
    .Q_N(_13290_),
    .Q(\cpu.icache.r_data[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3000),
    .D(_02105_),
    .Q_N(_13289_),
    .Q(\cpu.icache.r_data[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3001),
    .D(_02106_),
    .Q_N(_13288_),
    .Q(\cpu.icache.r_data[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][19]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3002),
    .D(_02107_),
    .Q_N(_13287_),
    .Q(\cpu.icache.r_data[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net3003),
    .D(_02108_),
    .Q_N(_13286_),
    .Q(\cpu.icache.r_data[3][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][20]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3004),
    .D(_02109_),
    .Q_N(_13285_),
    .Q(\cpu.icache.r_data[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][21]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3005),
    .D(_02110_),
    .Q_N(_13284_),
    .Q(\cpu.icache.r_data[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][22]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3006),
    .D(_02111_),
    .Q_N(_13283_),
    .Q(\cpu.icache.r_data[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][23]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3007),
    .D(_02112_),
    .Q_N(_13282_),
    .Q(\cpu.icache.r_data[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][24]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3008),
    .D(_02113_),
    .Q_N(_13281_),
    .Q(\cpu.icache.r_data[3][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3009),
    .D(_02114_),
    .Q_N(_13280_),
    .Q(\cpu.icache.r_data[3][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][26]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3010),
    .D(_02115_),
    .Q_N(_13279_),
    .Q(\cpu.icache.r_data[3][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][27]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3011),
    .D(_02116_),
    .Q_N(_13278_),
    .Q(\cpu.icache.r_data[3][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][28]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3012),
    .D(_02117_),
    .Q_N(_13277_),
    .Q(\cpu.icache.r_data[3][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3013),
    .D(_02118_),
    .Q_N(_13276_),
    .Q(\cpu.icache.r_data[3][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3014),
    .D(_02119_),
    .Q_N(_13275_),
    .Q(\cpu.icache.r_data[3][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][30]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3015),
    .D(_02120_),
    .Q_N(_13274_),
    .Q(\cpu.icache.r_data[3][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][31]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3016),
    .D(_02121_),
    .Q_N(_13273_),
    .Q(\cpu.icache.r_data[3][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net3017),
    .D(_02122_),
    .Q_N(_13272_),
    .Q(\cpu.icache.r_data[3][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3018),
    .D(_02123_),
    .Q_N(_13271_),
    .Q(\cpu.icache.r_data[3][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3019),
    .D(_02124_),
    .Q_N(_13270_),
    .Q(\cpu.icache.r_data[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net3020),
    .D(_02125_),
    .Q_N(_13269_),
    .Q(\cpu.icache.r_data[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3021),
    .D(_02126_),
    .Q_N(_13268_),
    .Q(\cpu.icache.r_data[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3022),
    .D(_02127_),
    .Q_N(_13267_),
    .Q(\cpu.icache.r_data[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3023),
    .D(_02128_),
    .Q_N(_13266_),
    .Q(\cpu.icache.r_data[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3024),
    .D(_02129_),
    .Q_N(_13265_),
    .Q(\cpu.icache.r_data[4][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3025),
    .D(_02130_),
    .Q_N(_13264_),
    .Q(\cpu.icache.r_data[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3026),
    .D(_02131_),
    .Q_N(_13263_),
    .Q(\cpu.icache.r_data[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3027),
    .D(_02132_),
    .Q_N(_13262_),
    .Q(\cpu.icache.r_data[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3028),
    .D(_02133_),
    .Q_N(_13261_),
    .Q(\cpu.icache.r_data[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3029),
    .D(_02134_),
    .Q_N(_13260_),
    .Q(\cpu.icache.r_data[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3030),
    .D(_02135_),
    .Q_N(_13259_),
    .Q(\cpu.icache.r_data[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3031),
    .D(_02136_),
    .Q_N(_13258_),
    .Q(\cpu.icache.r_data[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3032),
    .D(_02137_),
    .Q_N(_13257_),
    .Q(\cpu.icache.r_data[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3033),
    .D(_02138_),
    .Q_N(_13256_),
    .Q(\cpu.icache.r_data[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][19]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net3034),
    .D(_02139_),
    .Q_N(_13255_),
    .Q(\cpu.icache.r_data[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3035),
    .D(_02140_),
    .Q_N(_13254_),
    .Q(\cpu.icache.r_data[4][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][20]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3036),
    .D(_02141_),
    .Q_N(_13253_),
    .Q(\cpu.icache.r_data[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][21]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3037),
    .D(_02142_),
    .Q_N(_13252_),
    .Q(\cpu.icache.r_data[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][22]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3038),
    .D(_02143_),
    .Q_N(_13251_),
    .Q(\cpu.icache.r_data[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][23]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3039),
    .D(_02144_),
    .Q_N(_13250_),
    .Q(\cpu.icache.r_data[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][24]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3040),
    .D(_02145_),
    .Q_N(_13249_),
    .Q(\cpu.icache.r_data[4][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][25]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3041),
    .D(_02146_),
    .Q_N(_13248_),
    .Q(\cpu.icache.r_data[4][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][26]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3042),
    .D(_02147_),
    .Q_N(_13247_),
    .Q(\cpu.icache.r_data[4][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][27]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3043),
    .D(_02148_),
    .Q_N(_13246_),
    .Q(\cpu.icache.r_data[4][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3044),
    .D(_02149_),
    .Q_N(_13245_),
    .Q(\cpu.icache.r_data[4][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][29]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3045),
    .D(_02150_),
    .Q_N(_13244_),
    .Q(\cpu.icache.r_data[4][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3046),
    .D(_02151_),
    .Q_N(_13243_),
    .Q(\cpu.icache.r_data[4][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3047),
    .D(_02152_),
    .Q_N(_13242_),
    .Q(\cpu.icache.r_data[4][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][31]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3048),
    .D(_02153_),
    .Q_N(_13241_),
    .Q(\cpu.icache.r_data[4][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3049),
    .D(_02154_),
    .Q_N(_13240_),
    .Q(\cpu.icache.r_data[4][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3050),
    .D(_02155_),
    .Q_N(_13239_),
    .Q(\cpu.icache.r_data[4][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3051),
    .D(_02156_),
    .Q_N(_13238_),
    .Q(\cpu.icache.r_data[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3052),
    .D(_02157_),
    .Q_N(_13237_),
    .Q(\cpu.icache.r_data[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3053),
    .D(_02158_),
    .Q_N(_13236_),
    .Q(\cpu.icache.r_data[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3054),
    .D(_02159_),
    .Q_N(_13235_),
    .Q(\cpu.icache.r_data[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3055),
    .D(_02160_),
    .Q_N(_13234_),
    .Q(\cpu.icache.r_data[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3056),
    .D(_02161_),
    .Q_N(_13233_),
    .Q(\cpu.icache.r_data[5][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3057),
    .D(_02162_),
    .Q_N(_13232_),
    .Q(\cpu.icache.r_data[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3058),
    .D(_02163_),
    .Q_N(_13231_),
    .Q(\cpu.icache.r_data[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3059),
    .D(_02164_),
    .Q_N(_13230_),
    .Q(\cpu.icache.r_data[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3060),
    .D(_02165_),
    .Q_N(_13229_),
    .Q(\cpu.icache.r_data[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3061),
    .D(_02166_),
    .Q_N(_13228_),
    .Q(\cpu.icache.r_data[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3062),
    .D(_02167_),
    .Q_N(_13227_),
    .Q(\cpu.icache.r_data[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3063),
    .D(_02168_),
    .Q_N(_13226_),
    .Q(\cpu.icache.r_data[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3064),
    .D(_02169_),
    .Q_N(_13225_),
    .Q(\cpu.icache.r_data[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3065),
    .D(_02170_),
    .Q_N(_13224_),
    .Q(\cpu.icache.r_data[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][19]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3066),
    .D(_02171_),
    .Q_N(_13223_),
    .Q(\cpu.icache.r_data[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3067),
    .D(_02172_),
    .Q_N(_13222_),
    .Q(\cpu.icache.r_data[5][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3068),
    .D(_02173_),
    .Q_N(_13221_),
    .Q(\cpu.icache.r_data[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][21]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3069),
    .D(_02174_),
    .Q_N(_13220_),
    .Q(\cpu.icache.r_data[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][22]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3070),
    .D(_02175_),
    .Q_N(_13219_),
    .Q(\cpu.icache.r_data[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][23]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3071),
    .D(_02176_),
    .Q_N(_13218_),
    .Q(\cpu.icache.r_data[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][24]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3072),
    .D(_02177_),
    .Q_N(_13217_),
    .Q(\cpu.icache.r_data[5][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][25]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3073),
    .D(_02178_),
    .Q_N(_13216_),
    .Q(\cpu.icache.r_data[5][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3074),
    .D(_02179_),
    .Q_N(_13215_),
    .Q(\cpu.icache.r_data[5][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][27]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3075),
    .D(_02180_),
    .Q_N(_13214_),
    .Q(\cpu.icache.r_data[5][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][28]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net3076),
    .D(_02181_),
    .Q_N(_13213_),
    .Q(\cpu.icache.r_data[5][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3077),
    .D(_02182_),
    .Q_N(_13212_),
    .Q(\cpu.icache.r_data[5][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3078),
    .D(_02183_),
    .Q_N(_13211_),
    .Q(\cpu.icache.r_data[5][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][30]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3079),
    .D(_02184_),
    .Q_N(_13210_),
    .Q(\cpu.icache.r_data[5][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][31]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3080),
    .D(_02185_),
    .Q_N(_13209_),
    .Q(\cpu.icache.r_data[5][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3081),
    .D(_02186_),
    .Q_N(_13208_),
    .Q(\cpu.icache.r_data[5][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3082),
    .D(_02187_),
    .Q_N(_13207_),
    .Q(\cpu.icache.r_data[5][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3083),
    .D(_02188_),
    .Q_N(_13206_),
    .Q(\cpu.icache.r_data[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3084),
    .D(_02189_),
    .Q_N(_13205_),
    .Q(\cpu.icache.r_data[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3085),
    .D(_02190_),
    .Q_N(_13204_),
    .Q(\cpu.icache.r_data[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net3086),
    .D(_02191_),
    .Q_N(_13203_),
    .Q(\cpu.icache.r_data[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3087),
    .D(_02192_),
    .Q_N(_13202_),
    .Q(\cpu.icache.r_data[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3088),
    .D(_02193_),
    .Q_N(_13201_),
    .Q(\cpu.icache.r_data[6][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3089),
    .D(_02194_),
    .Q_N(_13200_),
    .Q(\cpu.icache.r_data[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3090),
    .D(_02195_),
    .Q_N(_13199_),
    .Q(\cpu.icache.r_data[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3091),
    .D(_02196_),
    .Q_N(_13198_),
    .Q(\cpu.icache.r_data[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3092),
    .D(_02197_),
    .Q_N(_13197_),
    .Q(\cpu.icache.r_data[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3093),
    .D(_02198_),
    .Q_N(_13196_),
    .Q(\cpu.icache.r_data[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3094),
    .D(_02199_),
    .Q_N(_13195_),
    .Q(\cpu.icache.r_data[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3095),
    .D(_02200_),
    .Q_N(_13194_),
    .Q(\cpu.icache.r_data[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3096),
    .D(_02201_),
    .Q_N(_13193_),
    .Q(\cpu.icache.r_data[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3097),
    .D(_02202_),
    .Q_N(_13192_),
    .Q(\cpu.icache.r_data[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][19]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3098),
    .D(_02203_),
    .Q_N(_13191_),
    .Q(\cpu.icache.r_data[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3099),
    .D(_02204_),
    .Q_N(_13190_),
    .Q(\cpu.icache.r_data[6][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][20]$_DFFE_PP_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net3100),
    .D(_02205_),
    .Q_N(_13189_),
    .Q(\cpu.icache.r_data[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][21]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net3101),
    .D(_02206_),
    .Q_N(_13188_),
    .Q(\cpu.icache.r_data[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][22]$_DFFE_PP_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net3102),
    .D(_02207_),
    .Q_N(_13187_),
    .Q(\cpu.icache.r_data[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][23]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3103),
    .D(_02208_),
    .Q_N(_13186_),
    .Q(\cpu.icache.r_data[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][24]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3104),
    .D(_02209_),
    .Q_N(_13185_),
    .Q(\cpu.icache.r_data[6][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][25]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3105),
    .D(_02210_),
    .Q_N(_13184_),
    .Q(\cpu.icache.r_data[6][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][26]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3106),
    .D(_02211_),
    .Q_N(_13183_),
    .Q(\cpu.icache.r_data[6][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][27]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3107),
    .D(_02212_),
    .Q_N(_13182_),
    .Q(\cpu.icache.r_data[6][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3108),
    .D(_02213_),
    .Q_N(_13181_),
    .Q(\cpu.icache.r_data[6][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3109),
    .D(_02214_),
    .Q_N(_13180_),
    .Q(\cpu.icache.r_data[6][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net3110),
    .D(_02215_),
    .Q_N(_13179_),
    .Q(\cpu.icache.r_data[6][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][30]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3111),
    .D(_02216_),
    .Q_N(_13178_),
    .Q(\cpu.icache.r_data[6][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][31]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3112),
    .D(_02217_),
    .Q_N(_13177_),
    .Q(\cpu.icache.r_data[6][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3113),
    .D(_02218_),
    .Q_N(_13176_),
    .Q(\cpu.icache.r_data[6][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3114),
    .D(_02219_),
    .Q_N(_13175_),
    .Q(\cpu.icache.r_data[6][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3115),
    .D(_02220_),
    .Q_N(_13174_),
    .Q(\cpu.icache.r_data[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3116),
    .D(_02221_),
    .Q_N(_13173_),
    .Q(\cpu.icache.r_data[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net3117),
    .D(_02222_),
    .Q_N(_13172_),
    .Q(\cpu.icache.r_data[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3118),
    .D(_02223_),
    .Q_N(_13171_),
    .Q(\cpu.icache.r_data[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net3119),
    .D(_02224_),
    .Q_N(_13170_),
    .Q(\cpu.icache.r_data[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net3120),
    .D(_02225_),
    .Q_N(_13169_),
    .Q(\cpu.icache.r_data[7][0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net3121),
    .D(_02226_),
    .Q_N(_13168_),
    .Q(\cpu.icache.r_data[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3122),
    .D(_02227_),
    .Q_N(_13167_),
    .Q(\cpu.icache.r_data[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3123),
    .D(_02228_),
    .Q_N(_13166_),
    .Q(\cpu.icache.r_data[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3124),
    .D(_02229_),
    .Q_N(_13165_),
    .Q(\cpu.icache.r_data[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3125),
    .D(_02230_),
    .Q_N(_13164_),
    .Q(\cpu.icache.r_data[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net3126),
    .D(_02231_),
    .Q_N(_13163_),
    .Q(\cpu.icache.r_data[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net3127),
    .D(_02232_),
    .Q_N(_13162_),
    .Q(\cpu.icache.r_data[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net3128),
    .D(_02233_),
    .Q_N(_13161_),
    .Q(\cpu.icache.r_data[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3129),
    .D(_02234_),
    .Q_N(_13160_),
    .Q(\cpu.icache.r_data[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][19]$_DFFE_PP_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net3130),
    .D(_02235_),
    .Q_N(_13159_),
    .Q(\cpu.icache.r_data[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3131),
    .D(_02236_),
    .Q_N(_13158_),
    .Q(\cpu.icache.r_data[7][1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][20]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3132),
    .D(_02237_),
    .Q_N(_13157_),
    .Q(\cpu.icache.r_data[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][21]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net3133),
    .D(_02238_),
    .Q_N(_13156_),
    .Q(\cpu.icache.r_data[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][22]$_DFFE_PP_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net3134),
    .D(_02239_),
    .Q_N(_13155_),
    .Q(\cpu.icache.r_data[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][23]$_DFFE_PP_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net3135),
    .D(_02240_),
    .Q_N(_13154_),
    .Q(\cpu.icache.r_data[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][24]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3136),
    .D(_02241_),
    .Q_N(_13153_),
    .Q(\cpu.icache.r_data[7][24] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][25]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3137),
    .D(_02242_),
    .Q_N(_13152_),
    .Q(\cpu.icache.r_data[7][25] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][26]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3138),
    .D(_02243_),
    .Q_N(_13151_),
    .Q(\cpu.icache.r_data[7][26] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][27]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3139),
    .D(_02244_),
    .Q_N(_13150_),
    .Q(\cpu.icache.r_data[7][27] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][28]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net3140),
    .D(_02245_),
    .Q_N(_13149_),
    .Q(\cpu.icache.r_data[7][28] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][29]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3141),
    .D(_02246_),
    .Q_N(_13148_),
    .Q(\cpu.icache.r_data[7][29] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3142),
    .D(_02247_),
    .Q_N(_13147_),
    .Q(\cpu.icache.r_data[7][2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][30]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3143),
    .D(_02248_),
    .Q_N(_13146_),
    .Q(\cpu.icache.r_data[7][30] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][31]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3144),
    .D(_02249_),
    .Q_N(_13145_),
    .Q(\cpu.icache.r_data[7][31] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net3145),
    .D(_02250_),
    .Q_N(_13144_),
    .Q(\cpu.icache.r_data[7][3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net3146),
    .D(_02251_),
    .Q_N(_13143_),
    .Q(\cpu.icache.r_data[7][4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3147),
    .D(_02252_),
    .Q_N(_13142_),
    .Q(\cpu.icache.r_data[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net3148),
    .D(_02253_),
    .Q_N(_13141_),
    .Q(\cpu.icache.r_data[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net3149),
    .D(_02254_),
    .Q_N(_13140_),
    .Q(\cpu.icache.r_data[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3150),
    .D(_02255_),
    .Q_N(_13139_),
    .Q(\cpu.icache.r_data[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_data[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3151),
    .D(_02256_),
    .Q_N(_13138_),
    .Q(\cpu.icache.r_data[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[0]$_SDFF_PN0_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3152),
    .D(_02257_),
    .Q_N(_00307_),
    .Q(\cpu.icache.r_offset[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[1]$_SDFF_PN0_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3153),
    .D(_02258_),
    .Q_N(_13137_),
    .Q(\cpu.icache.r_offset[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_offset[2]$_SDFF_PN0_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3154),
    .D(_02259_),
    .Q_N(_00246_),
    .Q(\cpu.icache.r_offset[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3155),
    .D(_02260_),
    .Q_N(_13136_),
    .Q(\cpu.icache.r_tag[0][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3156),
    .D(_02261_),
    .Q_N(_13135_),
    .Q(\cpu.icache.r_tag[0][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3157),
    .D(_02262_),
    .Q_N(_13134_),
    .Q(\cpu.icache.r_tag[0][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][12]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3158),
    .D(_02263_),
    .Q_N(_13133_),
    .Q(\cpu.icache.r_tag[0][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3159),
    .D(_02264_),
    .Q_N(_13132_),
    .Q(\cpu.icache.r_tag[0][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3160),
    .D(_02265_),
    .Q_N(_13131_),
    .Q(\cpu.icache.r_tag[0][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][15]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3161),
    .D(_02266_),
    .Q_N(_13130_),
    .Q(\cpu.icache.r_tag[0][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][16]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3162),
    .D(_02267_),
    .Q_N(_13129_),
    .Q(\cpu.icache.r_tag[0][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][17]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net3163),
    .D(_02268_),
    .Q_N(_13128_),
    .Q(\cpu.icache.r_tag[0][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][18]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3164),
    .D(_02269_),
    .Q_N(_13127_),
    .Q(\cpu.icache.r_tag[0][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3165),
    .D(_02270_),
    .Q_N(_13126_),
    .Q(\cpu.icache.r_tag[0][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3166),
    .D(_02271_),
    .Q_N(_13125_),
    .Q(\cpu.icache.r_tag[0][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net3167),
    .D(_02272_),
    .Q_N(_13124_),
    .Q(\cpu.icache.r_tag[0][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3168),
    .D(_02273_),
    .Q_N(_13123_),
    .Q(\cpu.icache.r_tag[0][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3169),
    .D(_02274_),
    .Q_N(_13122_),
    .Q(\cpu.icache.r_tag[0][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3170),
    .D(_02275_),
    .Q_N(_13121_),
    .Q(\cpu.icache.r_tag[0][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3171),
    .D(_02276_),
    .Q_N(_13120_),
    .Q(\cpu.icache.r_tag[0][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3172),
    .D(_02277_),
    .Q_N(_13119_),
    .Q(\cpu.icache.r_tag[0][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3173),
    .D(_02278_),
    .Q_N(_13118_),
    .Q(\cpu.icache.r_tag[0][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3174),
    .D(_02279_),
    .Q_N(_13117_),
    .Q(\cpu.icache.r_tag[1][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3175),
    .D(_02280_),
    .Q_N(_13116_),
    .Q(\cpu.icache.r_tag[1][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3176),
    .D(_02281_),
    .Q_N(_13115_),
    .Q(\cpu.icache.r_tag[1][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][12]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3177),
    .D(_02282_),
    .Q_N(_13114_),
    .Q(\cpu.icache.r_tag[1][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3178),
    .D(_02283_),
    .Q_N(_13113_),
    .Q(\cpu.icache.r_tag[1][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3179),
    .D(_02284_),
    .Q_N(_13112_),
    .Q(\cpu.icache.r_tag[1][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3180),
    .D(_02285_),
    .Q_N(_13111_),
    .Q(\cpu.icache.r_tag[1][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][16]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3181),
    .D(_02286_),
    .Q_N(_13110_),
    .Q(\cpu.icache.r_tag[1][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][17]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3182),
    .D(_02287_),
    .Q_N(_13109_),
    .Q(\cpu.icache.r_tag[1][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][18]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3183),
    .D(_02288_),
    .Q_N(_13108_),
    .Q(\cpu.icache.r_tag[1][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3184),
    .D(_02289_),
    .Q_N(_13107_),
    .Q(\cpu.icache.r_tag[1][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3185),
    .D(_02290_),
    .Q_N(_13106_),
    .Q(\cpu.icache.r_tag[1][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3186),
    .D(_02291_),
    .Q_N(_13105_),
    .Q(\cpu.icache.r_tag[1][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3187),
    .D(_02292_),
    .Q_N(_13104_),
    .Q(\cpu.icache.r_tag[1][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3188),
    .D(_02293_),
    .Q_N(_13103_),
    .Q(\cpu.icache.r_tag[1][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3189),
    .D(_02294_),
    .Q_N(_13102_),
    .Q(\cpu.icache.r_tag[1][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3190),
    .D(_02295_),
    .Q_N(_13101_),
    .Q(\cpu.icache.r_tag[1][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3191),
    .D(_02296_),
    .Q_N(_13100_),
    .Q(\cpu.icache.r_tag[1][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3192),
    .D(_02297_),
    .Q_N(_13099_),
    .Q(\cpu.icache.r_tag[1][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3193),
    .D(_02298_),
    .Q_N(_13098_),
    .Q(\cpu.icache.r_tag[2][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3194),
    .D(_02299_),
    .Q_N(_13097_),
    .Q(\cpu.icache.r_tag[2][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3195),
    .D(_02300_),
    .Q_N(_13096_),
    .Q(\cpu.icache.r_tag[2][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][12]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3196),
    .D(_02301_),
    .Q_N(_13095_),
    .Q(\cpu.icache.r_tag[2][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][13]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3197),
    .D(_02302_),
    .Q_N(_13094_),
    .Q(\cpu.icache.r_tag[2][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][14]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3198),
    .D(_02303_),
    .Q_N(_13093_),
    .Q(\cpu.icache.r_tag[2][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][15]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3199),
    .D(_02304_),
    .Q_N(_13092_),
    .Q(\cpu.icache.r_tag[2][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][16]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3200),
    .D(_02305_),
    .Q_N(_13091_),
    .Q(\cpu.icache.r_tag[2][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][17]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3201),
    .D(_02306_),
    .Q_N(_13090_),
    .Q(\cpu.icache.r_tag[2][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][18]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3202),
    .D(_02307_),
    .Q_N(_13089_),
    .Q(\cpu.icache.r_tag[2][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3203),
    .D(_02308_),
    .Q_N(_13088_),
    .Q(\cpu.icache.r_tag[2][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3204),
    .D(_02309_),
    .Q_N(_13087_),
    .Q(\cpu.icache.r_tag[2][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3205),
    .D(_02310_),
    .Q_N(_13086_),
    .Q(\cpu.icache.r_tag[2][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3206),
    .D(_02311_),
    .Q_N(_13085_),
    .Q(\cpu.icache.r_tag[2][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3207),
    .D(_02312_),
    .Q_N(_13084_),
    .Q(\cpu.icache.r_tag[2][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3208),
    .D(_02313_),
    .Q_N(_13083_),
    .Q(\cpu.icache.r_tag[2][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net3209),
    .D(_02314_),
    .Q_N(_13082_),
    .Q(\cpu.icache.r_tag[2][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3210),
    .D(_02315_),
    .Q_N(_13081_),
    .Q(\cpu.icache.r_tag[2][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3211),
    .D(_02316_),
    .Q_N(_13080_),
    .Q(\cpu.icache.r_tag[2][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3212),
    .D(_02317_),
    .Q_N(_13079_),
    .Q(\cpu.icache.r_tag[3][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3213),
    .D(_02318_),
    .Q_N(_13078_),
    .Q(\cpu.icache.r_tag[3][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3214),
    .D(_02319_),
    .Q_N(_13077_),
    .Q(\cpu.icache.r_tag[3][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][12]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3215),
    .D(_02320_),
    .Q_N(_13076_),
    .Q(\cpu.icache.r_tag[3][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3216),
    .D(_02321_),
    .Q_N(_13075_),
    .Q(\cpu.icache.r_tag[3][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3217),
    .D(_02322_),
    .Q_N(_13074_),
    .Q(\cpu.icache.r_tag[3][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3218),
    .D(_02323_),
    .Q_N(_13073_),
    .Q(\cpu.icache.r_tag[3][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][16]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3219),
    .D(_02324_),
    .Q_N(_13072_),
    .Q(\cpu.icache.r_tag[3][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][17]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3220),
    .D(_02325_),
    .Q_N(_13071_),
    .Q(\cpu.icache.r_tag[3][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][18]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net3221),
    .D(_02326_),
    .Q_N(_13070_),
    .Q(\cpu.icache.r_tag[3][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3222),
    .D(_02327_),
    .Q_N(_13069_),
    .Q(\cpu.icache.r_tag[3][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3223),
    .D(_02328_),
    .Q_N(_13068_),
    .Q(\cpu.icache.r_tag[3][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3224),
    .D(_02329_),
    .Q_N(_13067_),
    .Q(\cpu.icache.r_tag[3][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3225),
    .D(_02330_),
    .Q_N(_13066_),
    .Q(\cpu.icache.r_tag[3][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3226),
    .D(_02331_),
    .Q_N(_13065_),
    .Q(\cpu.icache.r_tag[3][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3227),
    .D(_02332_),
    .Q_N(_13064_),
    .Q(\cpu.icache.r_tag[3][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3228),
    .D(_02333_),
    .Q_N(_13063_),
    .Q(\cpu.icache.r_tag[3][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3229),
    .D(_02334_),
    .Q_N(_13062_),
    .Q(\cpu.icache.r_tag[3][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3230),
    .D(_02335_),
    .Q_N(_13061_),
    .Q(\cpu.icache.r_tag[3][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3231),
    .D(_02336_),
    .Q_N(_13060_),
    .Q(\cpu.icache.r_tag[4][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3232),
    .D(_02337_),
    .Q_N(_13059_),
    .Q(\cpu.icache.r_tag[4][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3233),
    .D(_02338_),
    .Q_N(_13058_),
    .Q(\cpu.icache.r_tag[4][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][12]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3234),
    .D(_02339_),
    .Q_N(_13057_),
    .Q(\cpu.icache.r_tag[4][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3235),
    .D(_02340_),
    .Q_N(_13056_),
    .Q(\cpu.icache.r_tag[4][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3236),
    .D(_02341_),
    .Q_N(_13055_),
    .Q(\cpu.icache.r_tag[4][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3237),
    .D(_02342_),
    .Q_N(_13054_),
    .Q(\cpu.icache.r_tag[4][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][16]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3238),
    .D(_02343_),
    .Q_N(_13053_),
    .Q(\cpu.icache.r_tag[4][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][17]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3239),
    .D(_02344_),
    .Q_N(_13052_),
    .Q(\cpu.icache.r_tag[4][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][18]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3240),
    .D(_02345_),
    .Q_N(_13051_),
    .Q(\cpu.icache.r_tag[4][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3241),
    .D(_02346_),
    .Q_N(_13050_),
    .Q(\cpu.icache.r_tag[4][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3242),
    .D(_02347_),
    .Q_N(_13049_),
    .Q(\cpu.icache.r_tag[4][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3243),
    .D(_02348_),
    .Q_N(_13048_),
    .Q(\cpu.icache.r_tag[4][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3244),
    .D(_02349_),
    .Q_N(_13047_),
    .Q(\cpu.icache.r_tag[4][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3245),
    .D(_02350_),
    .Q_N(_13046_),
    .Q(\cpu.icache.r_tag[4][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3246),
    .D(_02351_),
    .Q_N(_13045_),
    .Q(\cpu.icache.r_tag[4][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3247),
    .D(_02352_),
    .Q_N(_13044_),
    .Q(\cpu.icache.r_tag[4][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3248),
    .D(_02353_),
    .Q_N(_13043_),
    .Q(\cpu.icache.r_tag[4][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3249),
    .D(_02354_),
    .Q_N(_13042_),
    .Q(\cpu.icache.r_tag[4][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3250),
    .D(_02355_),
    .Q_N(_13041_),
    .Q(\cpu.icache.r_tag[5][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3251),
    .D(_02356_),
    .Q_N(_13040_),
    .Q(\cpu.icache.r_tag[5][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3252),
    .D(_02357_),
    .Q_N(_13039_),
    .Q(\cpu.icache.r_tag[5][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][12]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3253),
    .D(_02358_),
    .Q_N(_13038_),
    .Q(\cpu.icache.r_tag[5][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][13]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net3254),
    .D(_02359_),
    .Q_N(_13037_),
    .Q(\cpu.icache.r_tag[5][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][14]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3255),
    .D(_02360_),
    .Q_N(_13036_),
    .Q(\cpu.icache.r_tag[5][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3256),
    .D(_02361_),
    .Q_N(_13035_),
    .Q(\cpu.icache.r_tag[5][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][16]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3257),
    .D(_02362_),
    .Q_N(_13034_),
    .Q(\cpu.icache.r_tag[5][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][17]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net3258),
    .D(_02363_),
    .Q_N(_13033_),
    .Q(\cpu.icache.r_tag[5][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][18]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3259),
    .D(_02364_),
    .Q_N(_13032_),
    .Q(\cpu.icache.r_tag[5][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3260),
    .D(_02365_),
    .Q_N(_13031_),
    .Q(\cpu.icache.r_tag[5][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3261),
    .D(_02366_),
    .Q_N(_13030_),
    .Q(\cpu.icache.r_tag[5][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3262),
    .D(_02367_),
    .Q_N(_13029_),
    .Q(\cpu.icache.r_tag[5][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3263),
    .D(_02368_),
    .Q_N(_13028_),
    .Q(\cpu.icache.r_tag[5][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net3264),
    .D(_02369_),
    .Q_N(_13027_),
    .Q(\cpu.icache.r_tag[5][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net3265),
    .D(_02370_),
    .Q_N(_13026_),
    .Q(\cpu.icache.r_tag[5][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3266),
    .D(_02371_),
    .Q_N(_13025_),
    .Q(\cpu.icache.r_tag[5][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3267),
    .D(_02372_),
    .Q_N(_13024_),
    .Q(\cpu.icache.r_tag[5][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3268),
    .D(_02373_),
    .Q_N(_13023_),
    .Q(\cpu.icache.r_tag[5][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3269),
    .D(_02374_),
    .Q_N(_13022_),
    .Q(\cpu.icache.r_tag[6][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3270),
    .D(_02375_),
    .Q_N(_13021_),
    .Q(\cpu.icache.r_tag[6][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3271),
    .D(_02376_),
    .Q_N(_13020_),
    .Q(\cpu.icache.r_tag[6][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][12]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net3272),
    .D(_02377_),
    .Q_N(_13019_),
    .Q(\cpu.icache.r_tag[6][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][13]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3273),
    .D(_02378_),
    .Q_N(_13018_),
    .Q(\cpu.icache.r_tag[6][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3274),
    .D(_02379_),
    .Q_N(_13017_),
    .Q(\cpu.icache.r_tag[6][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3275),
    .D(_02380_),
    .Q_N(_13016_),
    .Q(\cpu.icache.r_tag[6][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][16]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net3276),
    .D(_02381_),
    .Q_N(_13015_),
    .Q(\cpu.icache.r_tag[6][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][17]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3277),
    .D(_02382_),
    .Q_N(_13014_),
    .Q(\cpu.icache.r_tag[6][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][18]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3278),
    .D(_02383_),
    .Q_N(_13013_),
    .Q(\cpu.icache.r_tag[6][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net3279),
    .D(_02384_),
    .Q_N(_13012_),
    .Q(\cpu.icache.r_tag[6][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3280),
    .D(_02385_),
    .Q_N(_13011_),
    .Q(\cpu.icache.r_tag[6][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net3281),
    .D(_02386_),
    .Q_N(_13010_),
    .Q(\cpu.icache.r_tag[6][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3282),
    .D(_02387_),
    .Q_N(_13009_),
    .Q(\cpu.icache.r_tag[6][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net3283),
    .D(_02388_),
    .Q_N(_13008_),
    .Q(\cpu.icache.r_tag[6][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net3284),
    .D(_02389_),
    .Q_N(_13007_),
    .Q(\cpu.icache.r_tag[6][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3285),
    .D(_02390_),
    .Q_N(_13006_),
    .Q(\cpu.icache.r_tag[6][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3286),
    .D(_02391_),
    .Q_N(_13005_),
    .Q(\cpu.icache.r_tag[6][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net3287),
    .D(_02392_),
    .Q_N(_13004_),
    .Q(\cpu.icache.r_tag[6][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3288),
    .D(_02393_),
    .Q_N(_13003_),
    .Q(\cpu.icache.r_tag[7][5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3289),
    .D(_02394_),
    .Q_N(_13002_),
    .Q(\cpu.icache.r_tag[7][15] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3290),
    .D(_02395_),
    .Q_N(_13001_),
    .Q(\cpu.icache.r_tag[7][16] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][12]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3291),
    .D(_02396_),
    .Q_N(_13000_),
    .Q(\cpu.icache.r_tag[7][17] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][13]$_DFFE_PP_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net3292),
    .D(_02397_),
    .Q_N(_12999_),
    .Q(\cpu.icache.r_tag[7][18] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net3293),
    .D(_02398_),
    .Q_N(_12998_),
    .Q(\cpu.icache.r_tag[7][19] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][15]$_DFFE_PP_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net3294),
    .D(_02399_),
    .Q_N(_12997_),
    .Q(\cpu.icache.r_tag[7][20] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][16]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3295),
    .D(_02400_),
    .Q_N(_12996_),
    .Q(\cpu.icache.r_tag[7][21] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][17]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net3296),
    .D(_02401_),
    .Q_N(_12995_),
    .Q(\cpu.icache.r_tag[7][22] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][18]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3297),
    .D(_02402_),
    .Q_N(_12994_),
    .Q(\cpu.icache.r_tag[7][23] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3298),
    .D(_02403_),
    .Q_N(_12993_),
    .Q(\cpu.icache.r_tag[7][6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3299),
    .D(_02404_),
    .Q_N(_12992_),
    .Q(\cpu.icache.r_tag[7][7] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net3300),
    .D(_02405_),
    .Q_N(_12991_),
    .Q(\cpu.icache.r_tag[7][8] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3301),
    .D(_02406_),
    .Q_N(_12990_),
    .Q(\cpu.icache.r_tag[7][9] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net3302),
    .D(_02407_),
    .Q_N(_12989_),
    .Q(\cpu.icache.r_tag[7][10] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3303),
    .D(_02408_),
    .Q_N(_12988_),
    .Q(\cpu.icache.r_tag[7][11] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net3304),
    .D(_02409_),
    .Q_N(_12987_),
    .Q(\cpu.icache.r_tag[7][12] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net3305),
    .D(_02410_),
    .Q_N(_12986_),
    .Q(\cpu.icache.r_tag[7][13] ));
 sg13g2_dfrbp_1 \cpu.icache.r_tag[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net3306),
    .D(_02411_),
    .Q_N(_12985_),
    .Q(\cpu.icache.r_tag[7][14] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[0]$_SDFFE_PP0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3307),
    .D(_02412_),
    .Q_N(_12984_),
    .Q(\cpu.icache.r_valid[0] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[1]$_SDFFE_PP0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3308),
    .D(_02413_),
    .Q_N(_12983_),
    .Q(\cpu.icache.r_valid[1] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[2]$_SDFFE_PP0P_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net3309),
    .D(_02414_),
    .Q_N(_12982_),
    .Q(\cpu.icache.r_valid[2] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[3]$_SDFFE_PP0P_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net3310),
    .D(_02415_),
    .Q_N(_12981_),
    .Q(\cpu.icache.r_valid[3] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net3311),
    .D(_02416_),
    .Q_N(_12980_),
    .Q(\cpu.icache.r_valid[4] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3312),
    .D(_02417_),
    .Q_N(_12979_),
    .Q(\cpu.icache.r_valid[5] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3313),
    .D(_02418_),
    .Q_N(_12978_),
    .Q(\cpu.icache.r_valid[6] ));
 sg13g2_dfrbp_1 \cpu.icache.r_valid[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net3314),
    .D(_02419_),
    .Q_N(_12977_),
    .Q(\cpu.icache.r_valid[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3315),
    .D(_02420_),
    .Q_N(_12976_),
    .Q(\cpu.intr.r_clock ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[0]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3316),
    .D(_02421_),
    .Q_N(_12975_),
    .Q(\cpu.intr.r_clock_cmp[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[10]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3317),
    .D(_02422_),
    .Q_N(_12974_),
    .Q(\cpu.intr.r_clock_cmp[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[11]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3318),
    .D(_02423_),
    .Q_N(_12973_),
    .Q(\cpu.intr.r_clock_cmp[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[12]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3319),
    .D(_02424_),
    .Q_N(_12972_),
    .Q(\cpu.intr.r_clock_cmp[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[13]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3320),
    .D(_02425_),
    .Q_N(_12971_),
    .Q(\cpu.intr.r_clock_cmp[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[14]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3321),
    .D(_02426_),
    .Q_N(_12970_),
    .Q(\cpu.intr.r_clock_cmp[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[15]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3322),
    .D(_02427_),
    .Q_N(_12969_),
    .Q(\cpu.intr.r_clock_cmp[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[16]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3323),
    .D(_02428_),
    .Q_N(_12968_),
    .Q(\cpu.intr.r_clock_cmp[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[17]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3324),
    .D(_02429_),
    .Q_N(_12967_),
    .Q(\cpu.intr.r_clock_cmp[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[18]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3325),
    .D(_02430_),
    .Q_N(_12966_),
    .Q(\cpu.intr.r_clock_cmp[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[19]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3326),
    .D(_02431_),
    .Q_N(_12965_),
    .Q(\cpu.intr.r_clock_cmp[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[1]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3327),
    .D(_02432_),
    .Q_N(_12964_),
    .Q(\cpu.intr.r_clock_cmp[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[20]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3328),
    .D(_02433_),
    .Q_N(_12963_),
    .Q(\cpu.intr.r_clock_cmp[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[21]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3329),
    .D(_02434_),
    .Q_N(_12962_),
    .Q(\cpu.intr.r_clock_cmp[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[22]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3330),
    .D(_02435_),
    .Q_N(_12961_),
    .Q(\cpu.intr.r_clock_cmp[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[23]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3331),
    .D(_02436_),
    .Q_N(_12960_),
    .Q(\cpu.intr.r_clock_cmp[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[24]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3332),
    .D(_02437_),
    .Q_N(_12959_),
    .Q(\cpu.intr.r_clock_cmp[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[25]$_DFFE_PP_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3333),
    .D(_02438_),
    .Q_N(_12958_),
    .Q(\cpu.intr.r_clock_cmp[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[26]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3334),
    .D(_02439_),
    .Q_N(_12957_),
    .Q(\cpu.intr.r_clock_cmp[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[27]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3335),
    .D(_02440_),
    .Q_N(_12956_),
    .Q(\cpu.intr.r_clock_cmp[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[28]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3336),
    .D(_02441_),
    .Q_N(_12955_),
    .Q(\cpu.intr.r_clock_cmp[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[29]$_DFFE_PP_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net3337),
    .D(_02442_),
    .Q_N(_12954_),
    .Q(\cpu.intr.r_clock_cmp[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[2]$_DFFE_PP_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3338),
    .D(_02443_),
    .Q_N(_12953_),
    .Q(\cpu.intr.r_clock_cmp[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[30]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3339),
    .D(_02444_),
    .Q_N(_12952_),
    .Q(\cpu.intr.r_clock_cmp[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[31]$_DFFE_PP_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3340),
    .D(_02445_),
    .Q_N(_12951_),
    .Q(\cpu.intr.r_clock_cmp[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[3]$_DFFE_PP_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3341),
    .D(_02446_),
    .Q_N(_12950_),
    .Q(\cpu.intr.r_clock_cmp[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[4]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3342),
    .D(_02447_),
    .Q_N(_12949_),
    .Q(\cpu.intr.r_clock_cmp[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[5]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3343),
    .D(_02448_),
    .Q_N(_12948_),
    .Q(\cpu.intr.r_clock_cmp[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[6]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3344),
    .D(_02449_),
    .Q_N(_12947_),
    .Q(\cpu.intr.r_clock_cmp[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[7]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3345),
    .D(_02450_),
    .Q_N(_12946_),
    .Q(\cpu.intr.r_clock_cmp[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[8]$_DFFE_PP_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net3346),
    .D(_02451_),
    .Q_N(_12945_),
    .Q(\cpu.intr.r_clock_cmp[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_cmp[9]$_DFFE_PP_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3347),
    .D(_02452_),
    .Q_N(_14943_),
    .Q(\cpu.intr.r_clock_cmp[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[0]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3348),
    .D(_00036_),
    .Q_N(_00279_),
    .Q(\cpu.intr.r_clock_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[10]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3349),
    .D(_00037_),
    .Q_N(_14944_),
    .Q(\cpu.intr.r_clock_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[11]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3350),
    .D(_00038_),
    .Q_N(_14945_),
    .Q(\cpu.intr.r_clock_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[12]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3351),
    .D(_00039_),
    .Q_N(_14946_),
    .Q(\cpu.intr.r_clock_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[13]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3352),
    .D(_00040_),
    .Q_N(_14947_),
    .Q(\cpu.intr.r_clock_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[14]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3353),
    .D(_00041_),
    .Q_N(_14948_),
    .Q(\cpu.intr.r_clock_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[15]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3354),
    .D(_00042_),
    .Q_N(_12944_),
    .Q(\cpu.intr.r_clock_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[16]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3355),
    .D(_02453_),
    .Q_N(_12943_),
    .Q(\cpu.intr.r_clock_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[17]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3356),
    .D(_02454_),
    .Q_N(_12942_),
    .Q(\cpu.intr.r_clock_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[18]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3357),
    .D(_02455_),
    .Q_N(_12941_),
    .Q(\cpu.intr.r_clock_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[19]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3358),
    .D(_02456_),
    .Q_N(_14949_),
    .Q(\cpu.intr.r_clock_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[1]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3359),
    .D(_00043_),
    .Q_N(_12940_),
    .Q(\cpu.intr.r_clock_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[20]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3360),
    .D(_02457_),
    .Q_N(_12939_),
    .Q(\cpu.intr.r_clock_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[21]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3361),
    .D(_02458_),
    .Q_N(_12938_),
    .Q(\cpu.intr.r_clock_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[22]$_DFFE_PN_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3362),
    .D(_02459_),
    .Q_N(_12937_),
    .Q(\cpu.intr.r_clock_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[23]$_DFFE_PN_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3363),
    .D(_02460_),
    .Q_N(_12936_),
    .Q(\cpu.intr.r_clock_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[24]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3364),
    .D(_02461_),
    .Q_N(_12935_),
    .Q(\cpu.intr.r_clock_count[24] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[25]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3365),
    .D(_02462_),
    .Q_N(_12934_),
    .Q(\cpu.intr.r_clock_count[25] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[26]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3366),
    .D(_02463_),
    .Q_N(_12933_),
    .Q(\cpu.intr.r_clock_count[26] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[27]$_DFFE_PN_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3367),
    .D(_02464_),
    .Q_N(_12932_),
    .Q(\cpu.intr.r_clock_count[27] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[28]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3368),
    .D(_02465_),
    .Q_N(_12931_),
    .Q(\cpu.intr.r_clock_count[28] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[29]$_DFFE_PN_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3369),
    .D(_02466_),
    .Q_N(_14950_),
    .Q(\cpu.intr.r_clock_count[29] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[2]$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3370),
    .D(_00044_),
    .Q_N(_12930_),
    .Q(\cpu.intr.r_clock_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[30]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3371),
    .D(_02467_),
    .Q_N(_12929_),
    .Q(\cpu.intr.r_clock_count[30] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[31]$_DFFE_PN_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3372),
    .D(_02468_),
    .Q_N(_14951_),
    .Q(\cpu.intr.r_clock_count[31] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[3]$_DFF_P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net3373),
    .D(_00045_),
    .Q_N(_14952_),
    .Q(\cpu.intr.r_clock_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[4]$_DFF_P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net3374),
    .D(_00046_),
    .Q_N(_14953_),
    .Q(\cpu.intr.r_clock_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[5]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3375),
    .D(_00047_),
    .Q_N(_14954_),
    .Q(\cpu.intr.r_clock_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[6]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3376),
    .D(_00048_),
    .Q_N(_14955_),
    .Q(\cpu.intr.r_clock_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[7]$_DFF_P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net3377),
    .D(_00049_),
    .Q_N(_14956_),
    .Q(\cpu.intr.r_clock_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[8]$_DFF_P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net3378),
    .D(_00050_),
    .Q_N(_14957_),
    .Q(\cpu.intr.r_clock_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_clock_count[9]$_DFF_P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net3379),
    .D(_00051_),
    .Q_N(_12928_),
    .Q(\cpu.intr.r_clock_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3380),
    .D(_02469_),
    .Q_N(_12927_),
    .Q(\cpu.intr.r_enable[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3381),
    .D(_02470_),
    .Q_N(_12926_),
    .Q(\cpu.intr.r_enable[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3382),
    .D(_02471_),
    .Q_N(_12925_),
    .Q(\cpu.intr.r_enable[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3383),
    .D(_02472_),
    .Q_N(_12924_),
    .Q(\cpu.intr.r_enable[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3384),
    .D(_02473_),
    .Q_N(_12923_),
    .Q(\cpu.intr.r_enable[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_enable[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net3385),
    .D(_02474_),
    .Q_N(_12922_),
    .Q(\cpu.intr.r_enable[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3386),
    .D(_02475_),
    .Q_N(_14958_),
    .Q(\cpu.intr.r_timer ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[0]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3387),
    .D(_00055_),
    .Q_N(_00278_),
    .Q(\cpu.intr.r_timer_count[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[10]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3388),
    .D(_00056_),
    .Q_N(_14959_),
    .Q(\cpu.intr.r_timer_count[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[11]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3389),
    .D(_00057_),
    .Q_N(_14960_),
    .Q(\cpu.intr.r_timer_count[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[12]$_DFF_P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3390),
    .D(_00058_),
    .Q_N(_14961_),
    .Q(\cpu.intr.r_timer_count[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[13]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3391),
    .D(_00059_),
    .Q_N(_14962_),
    .Q(\cpu.intr.r_timer_count[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[14]$_DFF_P_  (.CLK(clknet_leaf_51_clk),
    .RESET_B(net3392),
    .D(_00060_),
    .Q_N(_14963_),
    .Q(\cpu.intr.r_timer_count[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[15]$_DFF_P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3393),
    .D(_00061_),
    .Q_N(_14964_),
    .Q(\cpu.intr.r_timer_count[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[16]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3394),
    .D(_00062_),
    .Q_N(_14965_),
    .Q(\cpu.intr.r_timer_count[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[17]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3395),
    .D(_00063_),
    .Q_N(_14966_),
    .Q(\cpu.intr.r_timer_count[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[18]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3396),
    .D(_00064_),
    .Q_N(_14967_),
    .Q(\cpu.intr.r_timer_count[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[19]$_DFF_P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3397),
    .D(_00065_),
    .Q_N(_14968_),
    .Q(\cpu.intr.r_timer_count[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[1]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3398),
    .D(_00066_),
    .Q_N(_14969_),
    .Q(\cpu.intr.r_timer_count[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[20]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3399),
    .D(_00067_),
    .Q_N(_14970_),
    .Q(\cpu.intr.r_timer_count[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[21]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3400),
    .D(_00068_),
    .Q_N(_14971_),
    .Q(\cpu.intr.r_timer_count[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[22]$_DFF_P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3401),
    .D(_00069_),
    .Q_N(_14972_),
    .Q(\cpu.intr.r_timer_count[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[23]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3402),
    .D(_00070_),
    .Q_N(_14973_),
    .Q(\cpu.intr.r_timer_count[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[2]$_DFF_P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3403),
    .D(_00071_),
    .Q_N(_14974_),
    .Q(\cpu.intr.r_timer_count[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[3]$_DFF_P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3404),
    .D(_00072_),
    .Q_N(_14975_),
    .Q(\cpu.intr.r_timer_count[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[4]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3405),
    .D(_00073_),
    .Q_N(_14976_),
    .Q(\cpu.intr.r_timer_count[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[5]$_DFF_P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3406),
    .D(_00074_),
    .Q_N(_14977_),
    .Q(\cpu.intr.r_timer_count[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[6]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3407),
    .D(_00075_),
    .Q_N(_14978_),
    .Q(\cpu.intr.r_timer_count[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[7]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3408),
    .D(_00076_),
    .Q_N(_14979_),
    .Q(\cpu.intr.r_timer_count[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[8]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3409),
    .D(_00077_),
    .Q_N(_14980_),
    .Q(\cpu.intr.r_timer_count[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_count[9]$_DFF_P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3410),
    .D(_00078_),
    .Q_N(_12921_),
    .Q(\cpu.intr.r_timer_count[9] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3411),
    .D(_02476_),
    .Q_N(_12920_),
    .Q(\cpu.intr.r_timer_reload[0] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[10]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3412),
    .D(_02477_),
    .Q_N(_12919_),
    .Q(\cpu.intr.r_timer_reload[10] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[11]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3413),
    .D(_02478_),
    .Q_N(_12918_),
    .Q(\cpu.intr.r_timer_reload[11] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[12]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3414),
    .D(_02479_),
    .Q_N(_12917_),
    .Q(\cpu.intr.r_timer_reload[12] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[13]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3415),
    .D(_02480_),
    .Q_N(_12916_),
    .Q(\cpu.intr.r_timer_reload[13] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[14]$_DFFE_PP_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net3416),
    .D(_02481_),
    .Q_N(_12915_),
    .Q(\cpu.intr.r_timer_reload[14] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[15]$_DFFE_PP_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net3417),
    .D(_02482_),
    .Q_N(_12914_),
    .Q(\cpu.intr.r_timer_reload[15] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[16]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3418),
    .D(_02483_),
    .Q_N(_12913_),
    .Q(\cpu.intr.r_timer_reload[16] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[17]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3419),
    .D(_02484_),
    .Q_N(_12912_),
    .Q(\cpu.intr.r_timer_reload[17] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[18]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3420),
    .D(_02485_),
    .Q_N(_12911_),
    .Q(\cpu.intr.r_timer_reload[18] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[19]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3421),
    .D(_02486_),
    .Q_N(_12910_),
    .Q(\cpu.intr.r_timer_reload[19] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[1]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3422),
    .D(_02487_),
    .Q_N(_12909_),
    .Q(\cpu.intr.r_timer_reload[1] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[20]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3423),
    .D(_02488_),
    .Q_N(_12908_),
    .Q(\cpu.intr.r_timer_reload[20] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[21]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3424),
    .D(_02489_),
    .Q_N(_12907_),
    .Q(\cpu.intr.r_timer_reload[21] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[22]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net3425),
    .D(_02490_),
    .Q_N(_12906_),
    .Q(\cpu.intr.r_timer_reload[22] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[23]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3426),
    .D(_02491_),
    .Q_N(_12905_),
    .Q(\cpu.intr.r_timer_reload[23] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[2]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3427),
    .D(_02492_),
    .Q_N(_12904_),
    .Q(\cpu.intr.r_timer_reload[2] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[3]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3428),
    .D(_02493_),
    .Q_N(_12903_),
    .Q(\cpu.intr.r_timer_reload[3] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[4]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3429),
    .D(_02494_),
    .Q_N(_12902_),
    .Q(\cpu.intr.r_timer_reload[4] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[5]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3430),
    .D(_02495_),
    .Q_N(_12901_),
    .Q(\cpu.intr.r_timer_reload[5] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[6]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net3431),
    .D(_02496_),
    .Q_N(_12900_),
    .Q(\cpu.intr.r_timer_reload[6] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[7]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net3432),
    .D(_02497_),
    .Q_N(_12899_),
    .Q(\cpu.intr.r_timer_reload[7] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[8]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3433),
    .D(_02498_),
    .Q_N(_12898_),
    .Q(\cpu.intr.r_timer_reload[8] ));
 sg13g2_dfrbp_1 \cpu.intr.r_timer_reload[9]$_DFFE_PP_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net3434),
    .D(_02499_),
    .Q_N(_12897_),
    .Q(\cpu.intr.r_timer_reload[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3435),
    .D(_02500_),
    .Q_N(_00181_),
    .Q(\cpu.qspi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3436),
    .D(_02501_),
    .Q_N(_12896_),
    .Q(\cpu.qspi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3437),
    .D(_02502_),
    .Q_N(_00182_),
    .Q(\cpu.qspi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3438),
    .D(_02503_),
    .Q_N(_12895_),
    .Q(\cpu.qspi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3439),
    .D(_02504_),
    .Q_N(_00244_),
    .Q(\cpu.qspi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3440),
    .D(_02505_),
    .Q_N(_12894_),
    .Q(net19));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3441),
    .D(_02506_),
    .Q_N(_12893_),
    .Q(net20));
 sg13g2_dfrbp_1 \cpu.qspi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3442),
    .D(_02507_),
    .Q_N(_12892_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_ind$_SDFFE_PN0N_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net3443),
    .D(_02508_),
    .Q_N(_12891_),
    .Q(\cpu.qspi.r_ind ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3444),
    .D(_02509_),
    .Q_N(_12890_),
    .Q(\cpu.qspi.r_mask[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3445),
    .D(_02510_),
    .Q_N(_12889_),
    .Q(\cpu.qspi.r_mask[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_mask[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3446),
    .D(_02511_),
    .Q_N(_12888_),
    .Q(\cpu.qspi.r_mask[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3447),
    .D(_02512_),
    .Q_N(_12887_),
    .Q(\cpu.qspi.r_quad[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net3448),
    .D(_02513_),
    .Q_N(_12886_),
    .Q(\cpu.qspi.r_quad[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_quad[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3449),
    .D(_02514_),
    .Q_N(_12885_),
    .Q(\cpu.qspi.r_quad[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3450),
    .D(_02515_),
    .Q_N(_12884_),
    .Q(\cpu.qspi.r_read_delay[0][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3451),
    .D(_02516_),
    .Q_N(_12883_),
    .Q(\cpu.qspi.r_read_delay[0][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3452),
    .D(_02517_),
    .Q_N(_12882_),
    .Q(\cpu.qspi.r_read_delay[0][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3453),
    .D(_02518_),
    .Q_N(_12881_),
    .Q(\cpu.qspi.r_read_delay[0][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net3454),
    .D(_02519_),
    .Q_N(_12880_),
    .Q(\cpu.qspi.r_read_delay[1][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3455),
    .D(_02520_),
    .Q_N(_12879_),
    .Q(\cpu.qspi.r_read_delay[1][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3456),
    .D(_02521_),
    .Q_N(_12878_),
    .Q(\cpu.qspi.r_read_delay[1][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3457),
    .D(_02522_),
    .Q_N(_12877_),
    .Q(\cpu.qspi.r_read_delay[1][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3458),
    .D(_02523_),
    .Q_N(_12876_),
    .Q(\cpu.qspi.r_read_delay[2][0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3459),
    .D(_02524_),
    .Q_N(_12875_),
    .Q(\cpu.qspi.r_read_delay[2][1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3460),
    .D(_02525_),
    .Q_N(_12874_),
    .Q(\cpu.qspi.r_read_delay[2][2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3461),
    .D(_02526_),
    .Q_N(_12873_),
    .Q(\cpu.qspi.r_read_delay[2][3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3462),
    .D(_02527_),
    .Q_N(_12872_),
    .Q(\cpu.qspi.r_rom_mode[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net3463),
    .D(_02528_),
    .Q_N(_14981_),
    .Q(\cpu.qspi.r_rom_mode[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_rstrobe_d$_DFF_P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net3464),
    .D(\cpu.qspi.c_rstrobe_d ),
    .Q_N(_14982_),
    .Q(\cpu.d_rstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3465),
    .D(_00021_),
    .Q_N(_00270_),
    .Q(\cpu.qspi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[10]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3466),
    .D(_00008_),
    .Q_N(_14983_),
    .Q(\cpu.qspi.r_state[10] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[11]$_DFF_P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3467),
    .D(_00022_),
    .Q_N(_14984_),
    .Q(\cpu.qspi.r_state[11] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[12]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3468),
    .D(_00023_),
    .Q_N(_14985_),
    .Q(\cpu.qspi.r_state[12] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[13]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3469),
    .D(_00009_),
    .Q_N(_14986_),
    .Q(\cpu.qspi.r_state[13] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[14]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3470),
    .D(_00024_),
    .Q_N(_14987_),
    .Q(\cpu.qspi.r_state[14] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[15]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3471),
    .D(_00010_),
    .Q_N(_14988_),
    .Q(\cpu.qspi.r_state[15] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[16]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3472),
    .D(_00025_),
    .Q_N(_14989_),
    .Q(\cpu.qspi.r_state[16] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[17]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3473),
    .D(_00026_),
    .Q_N(_14990_),
    .Q(\cpu.qspi.r_state[17] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3474),
    .D(_00001_),
    .Q_N(_14991_),
    .Q(\cpu.qspi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3475),
    .D(_00027_),
    .Q_N(_14992_),
    .Q(\cpu.qspi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net3476),
    .D(_00002_),
    .Q_N(_14993_),
    .Q(\cpu.qspi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3477),
    .D(_00028_),
    .Q_N(_14994_),
    .Q(\cpu.qspi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net3478),
    .D(_00003_),
    .Q_N(_14995_),
    .Q(\cpu.qspi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3479),
    .D(_00004_),
    .Q_N(_14996_),
    .Q(\cpu.qspi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[7]$_DFF_P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net3480),
    .D(_00005_),
    .Q_N(_14997_),
    .Q(\cpu.qspi.r_state[7] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[8]$_DFF_P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net3481),
    .D(_00006_),
    .Q_N(_00183_),
    .Q(\cpu.qspi.r_state[8] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_state[9]$_DFF_P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net3482),
    .D(_00007_),
    .Q_N(_12871_),
    .Q(\cpu.qspi.r_state[9] ));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3483),
    .D(_02529_),
    .Q_N(_12870_),
    .Q(net3));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net3484),
    .D(_02530_),
    .Q_N(_12869_),
    .Q(net6));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3485),
    .D(_02531_),
    .Q_N(_12868_),
    .Q(net11));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3486),
    .D(_02532_),
    .Q_N(_12867_),
    .Q(net12));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3487),
    .D(_02533_),
    .Q_N(_12866_),
    .Q(net13));
 sg13g2_dfrbp_1 \cpu.qspi.r_uio_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net3488),
    .D(_02534_),
    .Q_N(_14998_),
    .Q(net14));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_d$_DFF_P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net3489),
    .D(\cpu.qspi.c_wstrobe_d ),
    .Q_N(_14999_),
    .Q(\cpu.d_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.qspi.r_wstrobe_i$_DFF_P_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net3490),
    .D(\cpu.qspi.c_wstrobe_i ),
    .Q_N(_00245_),
    .Q(\cpu.i_wstrobe_d ));
 sg13g2_dfrbp_1 \cpu.r_clk_invert$_DFFE_PN_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net3491),
    .D(_02535_),
    .Q_N(_12865_),
    .Q(\cpu.r_clk_invert ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3492),
    .D(_02536_),
    .Q_N(_12864_),
    .Q(\cpu.spi.r_bits[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3493),
    .D(_02537_),
    .Q_N(_12863_),
    .Q(\cpu.spi.r_bits[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_bits[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3494),
    .D(_02538_),
    .Q_N(_12862_),
    .Q(\cpu.spi.r_bits[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3495),
    .D(_02539_),
    .Q_N(_00295_),
    .Q(\cpu.spi.r_clk_count[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3496),
    .D(_02540_),
    .Q_N(_00300_),
    .Q(\cpu.spi.r_clk_count[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3497),
    .D(_02541_),
    .Q_N(_00097_),
    .Q(\cpu.spi.r_clk_count[0][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3498),
    .D(_02542_),
    .Q_N(_00108_),
    .Q(\cpu.spi.r_clk_count[0][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3499),
    .D(_02543_),
    .Q_N(_00119_),
    .Q(\cpu.spi.r_clk_count[0][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3500),
    .D(_02544_),
    .Q_N(_00126_),
    .Q(\cpu.spi.r_clk_count[0][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3501),
    .D(_02545_),
    .Q_N(_00138_),
    .Q(\cpu.spi.r_clk_count[0][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3502),
    .D(_02546_),
    .Q_N(_00150_),
    .Q(\cpu.spi.r_clk_count[0][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3503),
    .D(_02547_),
    .Q_N(_00294_),
    .Q(\cpu.spi.r_clk_count[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3504),
    .D(_02548_),
    .Q_N(_00299_),
    .Q(\cpu.spi.r_clk_count[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3505),
    .D(_02549_),
    .Q_N(_00096_),
    .Q(\cpu.spi.r_clk_count[1][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3506),
    .D(_02550_),
    .Q_N(_00107_),
    .Q(\cpu.spi.r_clk_count[1][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3507),
    .D(_02551_),
    .Q_N(_00118_),
    .Q(\cpu.spi.r_clk_count[1][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3508),
    .D(_02552_),
    .Q_N(_00125_),
    .Q(\cpu.spi.r_clk_count[1][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3509),
    .D(_02553_),
    .Q_N(_00137_),
    .Q(\cpu.spi.r_clk_count[1][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3510),
    .D(_02554_),
    .Q_N(_00149_),
    .Q(\cpu.spi.r_clk_count[1][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3511),
    .D(_02555_),
    .Q_N(_12861_),
    .Q(\cpu.spi.r_clk_count[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3512),
    .D(_02556_),
    .Q_N(_12860_),
    .Q(\cpu.spi.r_clk_count[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3513),
    .D(_02557_),
    .Q_N(_12859_),
    .Q(\cpu.spi.r_clk_count[2][2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3514),
    .D(_02558_),
    .Q_N(_12858_),
    .Q(\cpu.spi.r_clk_count[2][3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3515),
    .D(_02559_),
    .Q_N(_12857_),
    .Q(\cpu.spi.r_clk_count[2][4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3516),
    .D(_02560_),
    .Q_N(_12856_),
    .Q(\cpu.spi.r_clk_count[2][5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3517),
    .D(_02561_),
    .Q_N(_12855_),
    .Q(\cpu.spi.r_clk_count[2][6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_clk_count[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3518),
    .D(_02562_),
    .Q_N(_12854_),
    .Q(\cpu.spi.r_clk_count[2][7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3519),
    .D(_02563_),
    .Q_N(_12853_),
    .Q(\cpu.spi.r_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3520),
    .D(_02564_),
    .Q_N(_12852_),
    .Q(\cpu.spi.r_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3521),
    .D(_02565_),
    .Q_N(_12851_),
    .Q(\cpu.spi.r_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3522),
    .D(_02566_),
    .Q_N(_12850_),
    .Q(\cpu.spi.r_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3523),
    .D(_02567_),
    .Q_N(_12849_),
    .Q(\cpu.spi.r_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net3524),
    .D(_02568_),
    .Q_N(_12848_),
    .Q(\cpu.spi.r_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3525),
    .D(_02569_),
    .Q_N(_12847_),
    .Q(\cpu.spi.r_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net3526),
    .D(_02570_),
    .Q_N(_12846_),
    .Q(\cpu.spi.r_count[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3527),
    .D(_02571_),
    .Q_N(_12845_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[1]$_SDFFE_PN1P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3528),
    .D(_02572_),
    .Q_N(_12844_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_cs[2]$_SDFFE_PN1P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3529),
    .D(_02573_),
    .Q_N(_12843_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[8] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net3530),
    .D(_02574_),
    .Q_N(_12842_),
    .Q(\cpu.spi.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3531),
    .D(_02575_),
    .Q_N(_12841_),
    .Q(\cpu.spi.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net3532),
    .D(_02576_),
    .Q_N(_12840_),
    .Q(\cpu.spi.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3533),
    .D(_02577_),
    .Q_N(_12839_),
    .Q(\cpu.spi.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net3534),
    .D(_02578_),
    .Q_N(_12838_),
    .Q(\cpu.spi.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3535),
    .D(_02579_),
    .Q_N(_12837_),
    .Q(\cpu.spi.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3536),
    .D(_02580_),
    .Q_N(_12836_),
    .Q(\cpu.spi.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net3537),
    .D(_02581_),
    .Q_N(_00214_),
    .Q(\cpu.spi.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_interrupt$_SDFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3538),
    .D(_02582_),
    .Q_N(_12835_),
    .Q(\cpu.intr.spi_intr ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3539),
    .D(_02583_),
    .Q_N(_00217_),
    .Q(\cpu.spi.r_mode[0][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3540),
    .D(_02584_),
    .Q_N(_12834_),
    .Q(\cpu.spi.r_mode[0][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3541),
    .D(_02585_),
    .Q_N(_12833_),
    .Q(\cpu.spi.r_mode[1][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net3542),
    .D(_02586_),
    .Q_N(_12832_),
    .Q(\cpu.spi.r_mode[1][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3543),
    .D(_02587_),
    .Q_N(_12831_),
    .Q(\cpu.spi.r_mode[2][0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_mode[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3544),
    .D(_02588_),
    .Q_N(_12830_),
    .Q(\cpu.spi.r_mode[2][1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3545),
    .D(_02589_),
    .Q_N(_12829_),
    .Q(\cpu.spi.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3546),
    .D(_02590_),
    .Q_N(_12828_),
    .Q(\cpu.spi.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3547),
    .D(_02591_),
    .Q_N(_12827_),
    .Q(\cpu.spi.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3548),
    .D(_02592_),
    .Q_N(_12826_),
    .Q(\cpu.spi.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3549),
    .D(_02593_),
    .Q_N(_12825_),
    .Q(\cpu.spi.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3550),
    .D(_02594_),
    .Q_N(_12824_),
    .Q(\cpu.spi.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3551),
    .D(_02595_),
    .Q_N(_12823_),
    .Q(\cpu.spi.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3552),
    .D(_02596_),
    .Q_N(_12822_),
    .Q(\cpu.spi.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_ready$_SDFFE_PN1P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3553),
    .D(_02597_),
    .Q_N(_12821_),
    .Q(\cpu.spi.r_ready ));
 sg13g2_dfrbp_1 \cpu.spi.r_searching$_SDFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3554),
    .D(_02598_),
    .Q_N(_00213_),
    .Q(\cpu.spi.r_searching ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[0]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3555),
    .D(_02599_),
    .Q_N(_12820_),
    .Q(\cpu.spi.r_sel[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_sel[1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3556),
    .D(_02600_),
    .Q_N(_12819_),
    .Q(\cpu.spi.r_sel[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[0]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3557),
    .D(_02601_),
    .Q_N(_00275_),
    .Q(\cpu.spi.r_src[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[1]$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net3558),
    .D(_02602_),
    .Q_N(_00276_),
    .Q(\cpu.spi.r_src[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_src[2]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net3559),
    .D(_02603_),
    .Q_N(_15000_),
    .Q(\cpu.spi.r_src[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[0]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3560),
    .D(_00029_),
    .Q_N(_15001_),
    .Q(\cpu.spi.r_state[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[1]$_DFF_P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net3561),
    .D(_00030_),
    .Q_N(_00218_),
    .Q(\cpu.spi.r_state[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[2]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3562),
    .D(_00031_),
    .Q_N(_15002_),
    .Q(\cpu.spi.r_state[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[3]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3563),
    .D(_00032_),
    .Q_N(_15003_),
    .Q(\cpu.spi.r_state[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[4]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3564),
    .D(_00033_),
    .Q_N(_00271_),
    .Q(\cpu.spi.r_state[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[5]$_DFF_P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3565),
    .D(_00034_),
    .Q_N(_15004_),
    .Q(\cpu.spi.r_state[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_state[6]$_DFF_P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net3566),
    .D(_00035_),
    .Q_N(_00219_),
    .Q(\cpu.spi.r_state[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[0]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3567),
    .D(_02604_),
    .Q_N(_12818_),
    .Q(\cpu.spi.r_timeout[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[1]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net3568),
    .D(_02605_),
    .Q_N(_12817_),
    .Q(\cpu.spi.r_timeout[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[2]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3569),
    .D(_02606_),
    .Q_N(_12816_),
    .Q(\cpu.spi.r_timeout[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[3]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3570),
    .D(_02607_),
    .Q_N(_12815_),
    .Q(\cpu.spi.r_timeout[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[4]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3571),
    .D(_02608_),
    .Q_N(_12814_),
    .Q(\cpu.spi.r_timeout[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[5]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3572),
    .D(_02609_),
    .Q_N(_12813_),
    .Q(\cpu.spi.r_timeout[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[6]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net3573),
    .D(_02610_),
    .Q_N(_12812_),
    .Q(\cpu.spi.r_timeout[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout[7]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net3574),
    .D(_02611_),
    .Q_N(_12811_),
    .Q(\cpu.spi.r_timeout[7] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[0]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3575),
    .D(_02612_),
    .Q_N(_00277_),
    .Q(\cpu.spi.r_timeout_count[0] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[1]$_DFFE_PP_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net3576),
    .D(_02613_),
    .Q_N(_12810_),
    .Q(\cpu.spi.r_timeout_count[1] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[2]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3577),
    .D(_02614_),
    .Q_N(_12809_),
    .Q(\cpu.spi.r_timeout_count[2] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[3]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3578),
    .D(_02615_),
    .Q_N(_12808_),
    .Q(\cpu.spi.r_timeout_count[3] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[4]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3579),
    .D(_02616_),
    .Q_N(_12807_),
    .Q(\cpu.spi.r_timeout_count[4] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[5]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3580),
    .D(_02617_),
    .Q_N(_12806_),
    .Q(\cpu.spi.r_timeout_count[5] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[6]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3581),
    .D(_02618_),
    .Q_N(_12805_),
    .Q(\cpu.spi.r_timeout_count[6] ));
 sg13g2_dfrbp_1 \cpu.spi.r_timeout_count[7]$_DFFE_PP_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net3582),
    .D(_02619_),
    .Q_N(_15005_),
    .Q(\cpu.spi.r_timeout_count[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[0]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3583),
    .D(_00079_),
    .Q_N(_00272_),
    .Q(\cpu.uart.r_div[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[10]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3584),
    .D(_00080_),
    .Q_N(_15006_),
    .Q(\cpu.uart.r_div[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[11]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3585),
    .D(_00081_),
    .Q_N(_15007_),
    .Q(\cpu.uart.r_div[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[1]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3586),
    .D(_00082_),
    .Q_N(_15008_),
    .Q(\cpu.uart.r_div[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[2]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3587),
    .D(_00083_),
    .Q_N(_15009_),
    .Q(\cpu.uart.r_div[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[3]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3588),
    .D(_00084_),
    .Q_N(_15010_),
    .Q(\cpu.uart.r_div[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[4]$_DFF_P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3589),
    .D(_00085_),
    .Q_N(_15011_),
    .Q(\cpu.uart.r_div[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[5]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3590),
    .D(_00086_),
    .Q_N(_15012_),
    .Q(\cpu.uart.r_div[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[6]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3591),
    .D(_00087_),
    .Q_N(_15013_),
    .Q(\cpu.uart.r_div[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[7]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3592),
    .D(_00088_),
    .Q_N(_15014_),
    .Q(\cpu.uart.r_div[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[8]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3593),
    .D(_00089_),
    .Q_N(_15015_),
    .Q(\cpu.uart.r_div[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div[9]$_DFF_P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3594),
    .D(_00090_),
    .Q_N(_12804_),
    .Q(\cpu.uart.r_div[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[0]$_SDFFE_PN1P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3595),
    .D(_02620_),
    .Q_N(_12803_),
    .Q(\cpu.uart.r_div_value[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[10]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3596),
    .D(_02621_),
    .Q_N(_12802_),
    .Q(\cpu.uart.r_div_value[10] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[11]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3597),
    .D(_02622_),
    .Q_N(_12801_),
    .Q(\cpu.uart.r_div_value[11] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3598),
    .D(_02623_),
    .Q_N(_12800_),
    .Q(\cpu.uart.r_div_value[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3599),
    .D(_02624_),
    .Q_N(_12799_),
    .Q(\cpu.uart.r_div_value[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3600),
    .D(_02625_),
    .Q_N(_12798_),
    .Q(\cpu.uart.r_div_value[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[4]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3601),
    .D(_02626_),
    .Q_N(_12797_),
    .Q(\cpu.uart.r_div_value[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[5]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3602),
    .D(_02627_),
    .Q_N(_12796_),
    .Q(\cpu.uart.r_div_value[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[6]$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3603),
    .D(_02628_),
    .Q_N(_12795_),
    .Q(\cpu.uart.r_div_value[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[7]$_SDFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3604),
    .D(_02629_),
    .Q_N(_12794_),
    .Q(\cpu.uart.r_div_value[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[8]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3605),
    .D(_02630_),
    .Q_N(_12793_),
    .Q(\cpu.uart.r_div_value[8] ));
 sg13g2_dfrbp_1 \cpu.uart.r_div_value[9]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3606),
    .D(_02631_),
    .Q_N(_12792_),
    .Q(\cpu.uart.r_div_value[9] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[0]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3607),
    .D(_02632_),
    .Q_N(_12791_),
    .Q(\cpu.uart.r_ib[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3608),
    .D(_02633_),
    .Q_N(_12790_),
    .Q(\cpu.uart.r_ib[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3609),
    .D(_02634_),
    .Q_N(_12789_),
    .Q(\cpu.uart.r_ib[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3610),
    .D(_02635_),
    .Q_N(_12788_),
    .Q(\cpu.uart.r_ib[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3611),
    .D(_02636_),
    .Q_N(_12787_),
    .Q(\cpu.uart.r_ib[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[5]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3612),
    .D(_02637_),
    .Q_N(_12786_),
    .Q(\cpu.uart.r_ib[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_ib[6]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3613),
    .D(_02638_),
    .Q_N(_12785_),
    .Q(\cpu.uart.r_ib[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[0]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3614),
    .D(_02639_),
    .Q_N(_12784_),
    .Q(\cpu.uart.r_in[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[1]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3615),
    .D(_02640_),
    .Q_N(_12783_),
    .Q(\cpu.uart.r_in[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[2]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3616),
    .D(_02641_),
    .Q_N(_12782_),
    .Q(\cpu.uart.r_in[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[3]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net3617),
    .D(_02642_),
    .Q_N(_12781_),
    .Q(\cpu.uart.r_in[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[4]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net3618),
    .D(_02643_),
    .Q_N(_12780_),
    .Q(\cpu.uart.r_in[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[5]$_DFFE_PP_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net3619),
    .D(_02644_),
    .Q_N(_12779_),
    .Q(\cpu.uart.r_in[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[6]$_DFFE_PP_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net3620),
    .D(_02645_),
    .Q_N(_12778_),
    .Q(\cpu.uart.r_in[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_in[7]$_DFFE_PP_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net3621),
    .D(_02646_),
    .Q_N(_12777_),
    .Q(\cpu.uart.r_in[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[0]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3622),
    .D(_02647_),
    .Q_N(_12776_),
    .Q(\cpu.uart.r_out[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[1]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3623),
    .D(_02648_),
    .Q_N(_12775_),
    .Q(\cpu.uart.r_out[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[2]$_DFFE_PP_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net3624),
    .D(_02649_),
    .Q_N(_12774_),
    .Q(\cpu.uart.r_out[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[3]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3625),
    .D(_02650_),
    .Q_N(_12773_),
    .Q(\cpu.uart.r_out[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[4]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3626),
    .D(_02651_),
    .Q_N(_12772_),
    .Q(\cpu.uart.r_out[4] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[5]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3627),
    .D(_02652_),
    .Q_N(_12771_),
    .Q(\cpu.uart.r_out[5] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[6]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3628),
    .D(_02653_),
    .Q_N(_12770_),
    .Q(\cpu.uart.r_out[6] ));
 sg13g2_dfrbp_1 \cpu.uart.r_out[7]$_DFFE_PP_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net3629),
    .D(_02654_),
    .Q_N(_15016_),
    .Q(\cpu.uart.r_out[7] ));
 sg13g2_dfrbp_1 \cpu.uart.r_r$_DFF_P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net3630),
    .D(\cpu.gpio.uart_rx ),
    .Q_N(_12769_),
    .Q(\cpu.uart.r_r ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net3631),
    .D(_02655_),
    .Q_N(_12768_),
    .Q(\cpu.uart.r_r_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_r_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3632),
    .D(_02656_),
    .Q_N(_12767_),
    .Q(\cpu.uart.r_r_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3633),
    .D(_02657_),
    .Q_N(_12766_),
    .Q(\cpu.uart.r_rcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net3634),
    .D(_02658_),
    .Q_N(_12765_),
    .Q(\cpu.uart.r_rcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3635),
    .D(_02659_),
    .Q_N(_12764_),
    .Q(\cpu.uart.r_rstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net3636),
    .D(_02660_),
    .Q_N(_12763_),
    .Q(\cpu.uart.r_rstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3637),
    .D(_02661_),
    .Q_N(_12762_),
    .Q(\cpu.uart.r_rstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_rstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net3638),
    .D(_02662_),
    .Q_N(_12761_),
    .Q(\cpu.uart.r_rstate[3] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x$_DFFE_PP_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3639),
    .D(_02663_),
    .Q_N(_12760_),
    .Q(\cpu.gpio.genblk1[3].srcs_o[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_int$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3640),
    .D(_02664_),
    .Q_N(_12759_),
    .Q(\cpu.uart.r_x_int ));
 sg13g2_dfrbp_1 \cpu.uart.r_x_invert$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3641),
    .D(_02665_),
    .Q_N(_00273_),
    .Q(\cpu.uart.r_x_invert ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[0]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3642),
    .D(_02666_),
    .Q_N(_12758_),
    .Q(\cpu.uart.r_xcnt[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xcnt[1]$_DFFE_PP_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3643),
    .D(_02667_),
    .Q_N(_12757_),
    .Q(\cpu.uart.r_xcnt[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[0]$_SDFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net3644),
    .D(_02668_),
    .Q_N(_12756_),
    .Q(\cpu.uart.r_xstate[0] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[1]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3645),
    .D(_02669_),
    .Q_N(_12755_),
    .Q(\cpu.uart.r_xstate[1] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[2]$_SDFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net3646),
    .D(_02670_),
    .Q_N(_12754_),
    .Q(\cpu.uart.r_xstate[2] ));
 sg13g2_dfrbp_1 \cpu.uart.r_xstate[3]$_SDFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net3647),
    .D(_02671_),
    .Q_N(_15017_),
    .Q(\cpu.uart.r_xstate[3] ));
 sg13g2_dfrbp_1 \r_reset$_DFF_P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net3648),
    .D(_00000_),
    .Q_N(_12753_),
    .Q(r_reset));
 sg13g2_buf_1 input1 (.A(ena),
    .X(net1));
 sg13g2_buf_1 input2 (.A(rst_n),
    .X(net2));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_oe[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_oe[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_oe[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_oe[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_oe[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_oe[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uio_oe[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_oe[7]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[0]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[1]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[2]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[3]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[4]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[5]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[6]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uio_out[7]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[0]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[1]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[2]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[3]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[4]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[5]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[6]));
 sg13g2_buf_1 output26 (.A(net26),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout27 (.A(_03699_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_06693_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_03698_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_03816_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_04088_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_03696_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_02964_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_02936_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_02915_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_02908_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_02859_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02832_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02812_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_02805_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_02754_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_02722_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_02702_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_02695_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_12706_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_12682_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_12675_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_12623_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_12596_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_12576_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_12569_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_12516_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_12487_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_12467_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_12460_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_12407_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_12378_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_12355_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_12345_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_12228_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_12165_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_12144_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_09946_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_09935_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_09933_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_07294_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_06989_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_05025_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_05024_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_04230_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_03977_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_12737_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_12286_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_11426_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_07212_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_07168_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_06360_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_06343_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_06334_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_06322_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04080_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_11676_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_07409_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_07401_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_06943_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_04139_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_04043_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_03268_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_03111_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_11644_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_11439_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_09820_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_09095_),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(_09094_));
 sg13g2_buf_2 fanout95 (.A(_08861_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_07769_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_07609_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_06952_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_05725_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_05448_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_04262_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_04111_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04042_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_04029_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_04013_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_04010_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_03397_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_03296_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_11604_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_11438_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_09245_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_09101_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_09056_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_08860_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_07821_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_07798_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_07790_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_07773_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_07772_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_07699_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_07660_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_07628_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_07620_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_07619_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_06809_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_06777_),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(_06683_));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(_06677_));
 sg13g2_buf_2 fanout129 (.A(_05454_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_05219_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_05023_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_04838_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_04295_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_04269_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_04266_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_04244_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_04134_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_04033_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_04012_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_04009_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_04004_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_03994_),
    .X(net142));
 sg13g2_buf_2 fanout143 (.A(_03262_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_03147_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_03145_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_12042_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_11955_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_11612_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_11602_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_11331_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_10070_),
    .X(net151));
 sg13g2_buf_2 fanout152 (.A(_10035_),
    .X(net152));
 sg13g2_buf_2 fanout153 (.A(_10024_),
    .X(net153));
 sg13g2_buf_2 fanout154 (.A(_09842_),
    .X(net154));
 sg13g2_buf_2 fanout155 (.A(_09838_),
    .X(net155));
 sg13g2_buf_2 fanout156 (.A(_09825_),
    .X(net156));
 sg13g2_buf_2 fanout157 (.A(_09244_),
    .X(net157));
 sg13g2_buf_2 fanout158 (.A(_09011_),
    .X(net158));
 sg13g2_buf_2 fanout159 (.A(_08070_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_07849_),
    .X(net160));
 sg13g2_buf_2 fanout161 (.A(_07762_),
    .X(net161));
 sg13g2_buf_2 fanout162 (.A(_07602_),
    .X(net162));
 sg13g2_buf_4 fanout163 (.X(net163),
    .A(_06680_));
 sg13g2_buf_2 fanout164 (.A(_04834_),
    .X(net164));
 sg13g2_buf_2 fanout165 (.A(_04291_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_04265_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_04260_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_04022_),
    .X(net168));
 sg13g2_buf_2 fanout169 (.A(_04014_),
    .X(net169));
 sg13g2_buf_2 fanout170 (.A(_03996_),
    .X(net170));
 sg13g2_buf_2 fanout171 (.A(_03995_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_03733_),
    .X(net172));
 sg13g2_buf_2 fanout173 (.A(_03114_),
    .X(net173));
 sg13g2_buf_2 fanout174 (.A(_03108_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_11632_),
    .X(net175));
 sg13g2_buf_2 fanout176 (.A(_11611_),
    .X(net176));
 sg13g2_buf_2 fanout177 (.A(_11468_),
    .X(net177));
 sg13g2_buf_2 fanout178 (.A(_11460_),
    .X(net178));
 sg13g2_buf_2 fanout179 (.A(_11389_),
    .X(net179));
 sg13g2_buf_2 fanout180 (.A(_11361_),
    .X(net180));
 sg13g2_buf_2 fanout181 (.A(_11296_),
    .X(net181));
 sg13g2_buf_2 fanout182 (.A(_10043_),
    .X(net182));
 sg13g2_buf_2 fanout183 (.A(_10034_),
    .X(net183));
 sg13g2_buf_2 fanout184 (.A(_09973_),
    .X(net184));
 sg13g2_buf_2 fanout185 (.A(_09972_),
    .X(net185));
 sg13g2_buf_2 fanout186 (.A(_09826_),
    .X(net186));
 sg13g2_buf_2 fanout187 (.A(_09096_),
    .X(net187));
 sg13g2_buf_2 fanout188 (.A(_07262_),
    .X(net188));
 sg13g2_buf_2 fanout189 (.A(_04129_),
    .X(net189));
 sg13g2_buf_2 fanout190 (.A(_04090_),
    .X(net190));
 sg13g2_buf_2 fanout191 (.A(_04020_),
    .X(net191));
 sg13g2_buf_2 fanout192 (.A(_03787_),
    .X(net192));
 sg13g2_buf_2 fanout193 (.A(_03732_),
    .X(net193));
 sg13g2_buf_2 fanout194 (.A(_03306_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_03137_),
    .X(net195));
 sg13g2_buf_2 fanout196 (.A(_03132_),
    .X(net196));
 sg13g2_buf_2 fanout197 (.A(_03128_),
    .X(net197));
 sg13g2_buf_2 fanout198 (.A(_03123_),
    .X(net198));
 sg13g2_buf_2 fanout199 (.A(_11684_),
    .X(net199));
 sg13g2_buf_2 fanout200 (.A(_11645_),
    .X(net200));
 sg13g2_buf_2 fanout201 (.A(_11594_),
    .X(net201));
 sg13g2_buf_2 fanout202 (.A(_11517_),
    .X(net202));
 sg13g2_buf_2 fanout203 (.A(_11510_),
    .X(net203));
 sg13g2_buf_2 fanout204 (.A(_11467_),
    .X(net204));
 sg13g2_buf_2 fanout205 (.A(_11418_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_11328_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_11321_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_11256_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_09827_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_09009_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_05157_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_04261_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_04053_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_03985_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_03735_),
    .X(net215));
 sg13g2_buf_2 fanout216 (.A(_03254_),
    .X(net216));
 sg13g2_buf_2 fanout217 (.A(_03230_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_03136_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_03131_),
    .X(net219));
 sg13g2_buf_2 fanout220 (.A(_03127_),
    .X(net220));
 sg13g2_buf_2 fanout221 (.A(_03122_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_03112_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_11776_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_11722_),
    .X(net224));
 sg13g2_buf_2 fanout225 (.A(_11694_),
    .X(net225));
 sg13g2_buf_2 fanout226 (.A(_11663_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_11475_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_11419_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_11247_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_11245_),
    .X(net230));
 sg13g2_buf_2 fanout231 (.A(_11226_),
    .X(net231));
 sg13g2_buf_2 fanout232 (.A(_10520_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_10365_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_10021_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_09861_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_09075_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_06255_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_06207_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_06129_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_06039_),
    .X(net240));
 sg13g2_buf_2 fanout241 (.A(_06013_),
    .X(net241));
 sg13g2_buf_2 fanout242 (.A(_04286_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_04025_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_04006_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_04001_),
    .X(net245));
 sg13g2_buf_2 fanout246 (.A(_03979_),
    .X(net246));
 sg13g2_buf_2 fanout247 (.A(_03972_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_03734_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_03356_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_03135_),
    .X(net250));
 sg13g2_buf_2 fanout251 (.A(_03116_),
    .X(net251));
 sg13g2_buf_2 fanout252 (.A(_11749_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_11704_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_11662_),
    .X(net254));
 sg13g2_buf_2 fanout255 (.A(_11580_),
    .X(net255));
 sg13g2_buf_2 fanout256 (.A(_11551_),
    .X(net256));
 sg13g2_buf_2 fanout257 (.A(_11502_),
    .X(net257));
 sg13g2_buf_2 fanout258 (.A(_11436_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_11416_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_10447_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_10444_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_09860_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_08969_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_06287_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_06279_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_06271_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_06263_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_06247_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_06239_));
 sg13g2_buf_4 fanout270 (.X(net270),
    .A(_06231_));
 sg13g2_buf_2 fanout271 (.A(_06223_),
    .X(net271));
 sg13g2_buf_4 fanout272 (.X(net272),
    .A(_06198_));
 sg13g2_buf_4 fanout273 (.X(net273),
    .A(_06186_));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_06162_));
 sg13g2_buf_2 fanout275 (.A(_06153_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_06145_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_06112_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_06104_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_06083_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_06067_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_06058_),
    .X(net281));
 sg13g2_buf_2 fanout282 (.A(_06030_),
    .X(net282));
 sg13g2_buf_2 fanout283 (.A(_06022_),
    .X(net283));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_06003_));
 sg13g2_buf_4 fanout285 (.X(net285),
    .A(_05964_));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_05939_));
 sg13g2_buf_4 fanout287 (.X(net287),
    .A(_05922_));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_05913_));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_05893_));
 sg13g2_buf_4 fanout290 (.X(net290),
    .A(_05872_));
 sg13g2_buf_2 fanout291 (.A(_05155_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_04476_),
    .X(net292));
 sg13g2_buf_2 fanout293 (.A(_03303_),
    .X(net293));
 sg13g2_buf_2 fanout294 (.A(_03125_),
    .X(net294));
 sg13g2_buf_4 fanout295 (.X(net295),
    .A(_03107_));
 sg13g2_buf_4 fanout296 (.X(net296),
    .A(_03106_));
 sg13g2_buf_4 fanout297 (.X(net297),
    .A(_03091_));
 sg13g2_buf_2 fanout298 (.A(_03090_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_11590_),
    .X(net299));
 sg13g2_buf_2 fanout300 (.A(_11537_),
    .X(net300));
 sg13g2_buf_2 fanout301 (.A(_10729_),
    .X(net301));
 sg13g2_buf_2 fanout302 (.A(_10596_),
    .X(net302));
 sg13g2_buf_2 fanout303 (.A(_10517_),
    .X(net303));
 sg13g2_buf_2 fanout304 (.A(_09089_),
    .X(net304));
 sg13g2_buf_2 fanout305 (.A(_06581_),
    .X(net305));
 sg13g2_buf_2 fanout306 (.A(_06567_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_06565_),
    .X(net307));
 sg13g2_buf_2 fanout308 (.A(_06564_),
    .X(net308));
 sg13g2_buf_2 fanout309 (.A(_06548_),
    .X(net309));
 sg13g2_buf_2 fanout310 (.A(_06546_),
    .X(net310));
 sg13g2_buf_2 fanout311 (.A(_06545_),
    .X(net311));
 sg13g2_buf_2 fanout312 (.A(_06477_),
    .X(net312));
 sg13g2_buf_2 fanout313 (.A(_06295_),
    .X(net313));
 sg13g2_buf_4 fanout314 (.X(net314),
    .A(_06215_));
 sg13g2_buf_2 fanout315 (.A(_06177_),
    .X(net315));
 sg13g2_buf_2 fanout316 (.A(_06137_),
    .X(net316));
 sg13g2_buf_2 fanout317 (.A(_06120_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_06092_),
    .X(net318));
 sg13g2_buf_2 fanout319 (.A(_06049_),
    .X(net319));
 sg13g2_buf_4 fanout320 (.X(net320),
    .A(_06000_));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_05997_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05992_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_05986_));
 sg13g2_buf_4 fanout324 (.X(net324),
    .A(_05977_));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_05974_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05971_));
 sg13g2_buf_4 fanout327 (.X(net327),
    .A(_05968_));
 sg13g2_buf_4 fanout328 (.X(net328),
    .A(_05951_));
 sg13g2_buf_4 fanout329 (.X(net329),
    .A(_05945_));
 sg13g2_buf_4 fanout330 (.X(net330),
    .A(_05935_));
 sg13g2_buf_4 fanout331 (.X(net331),
    .A(_05928_));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_05925_));
 sg13g2_buf_4 fanout333 (.X(net333),
    .A(_05909_));
 sg13g2_buf_4 fanout334 (.X(net334),
    .A(_05900_));
 sg13g2_buf_4 fanout335 (.X(net335),
    .A(_05888_));
 sg13g2_buf_4 fanout336 (.X(net336),
    .A(_05881_));
 sg13g2_buf_4 fanout337 (.X(net337),
    .A(_05876_));
 sg13g2_buf_4 fanout338 (.X(net338),
    .A(_05860_));
 sg13g2_buf_4 fanout339 (.X(net339),
    .A(_05854_));
 sg13g2_buf_2 fanout340 (.A(_05141_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_05139_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_03170_),
    .X(net342));
 sg13g2_buf_4 fanout343 (.X(net343),
    .A(_03089_));
 sg13g2_buf_4 fanout344 (.X(net344),
    .A(_03088_));
 sg13g2_buf_2 fanout345 (.A(_02966_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_12734_),
    .X(net346));
 sg13g2_buf_2 fanout347 (.A(_11014_),
    .X(net347));
 sg13g2_buf_2 fanout348 (.A(_10130_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_09858_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_09745_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_09441_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_09250_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_09240_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_09074_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_09050_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_09032_),
    .X(net356));
 sg13g2_buf_2 fanout357 (.A(_08907_),
    .X(net357));
 sg13g2_buf_2 fanout358 (.A(_08417_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_06640_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_06638_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_06637_),
    .X(net361));
 sg13g2_buf_2 fanout362 (.A(_06621_),
    .X(net362));
 sg13g2_buf_2 fanout363 (.A(_06619_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_06618_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_06582_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_06525_),
    .X(net366));
 sg13g2_buf_2 fanout367 (.A(_06476_),
    .X(net367));
 sg13g2_buf_2 fanout368 (.A(_06414_),
    .X(net368));
 sg13g2_buf_4 fanout369 (.X(net369),
    .A(_05981_));
 sg13g2_buf_4 fanout370 (.X(net370),
    .A(_05960_));
 sg13g2_buf_4 fanout371 (.X(net371),
    .A(_05919_));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(_05866_));
 sg13g2_buf_4 fanout373 (.X(net373),
    .A(_05841_));
 sg13g2_buf_2 fanout374 (.A(_05144_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_04931_),
    .X(net375));
 sg13g2_buf_2 fanout376 (.A(_04918_),
    .X(net376));
 sg13g2_buf_2 fanout377 (.A(_03731_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_03623_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_03052_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_03043_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_02905_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_12625_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_12313_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_12309_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_11785_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_10129_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_09635_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_09479_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_09412_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_09387_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_09331_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_08712_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_08692_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_08670_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_08646_),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(_08619_),
    .X(net396));
 sg13g2_buf_2 fanout397 (.A(_08591_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_08563_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_08511_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_08447_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_06602_),
    .X(net401));
 sg13g2_buf_2 fanout402 (.A(_06600_),
    .X(net402));
 sg13g2_buf_2 fanout403 (.A(_06599_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_06526_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_06413_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_06064_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_06019_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_05334_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_04966_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_04941_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_04930_),
    .X(net411));
 sg13g2_buf_2 fanout412 (.A(_04923_),
    .X(net412));
 sg13g2_buf_2 fanout413 (.A(_04871_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_04778_),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(_04775_),
    .X(net415));
 sg13g2_buf_2 fanout416 (.A(_03779_),
    .X(net416));
 sg13g2_buf_2 fanout417 (.A(_03726_),
    .X(net417));
 sg13g2_buf_2 fanout418 (.A(_03622_),
    .X(net418));
 sg13g2_buf_4 fanout419 (.X(net419),
    .A(_03053_));
 sg13g2_buf_2 fanout420 (.A(_03048_),
    .X(net420));
 sg13g2_buf_2 fanout421 (.A(_03042_),
    .X(net421));
 sg13g2_buf_2 fanout422 (.A(_03038_),
    .X(net422));
 sg13g2_buf_2 fanout423 (.A(_03033_),
    .X(net423));
 sg13g2_buf_2 fanout424 (.A(_03029_),
    .X(net424));
 sg13g2_buf_2 fanout425 (.A(_03025_),
    .X(net425));
 sg13g2_buf_2 fanout426 (.A(_12566_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_12302_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_12295_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_12294_),
    .X(net429));
 sg13g2_buf_2 fanout430 (.A(_12291_),
    .X(net430));
 sg13g2_buf_2 fanout431 (.A(_12282_),
    .X(net431));
 sg13g2_buf_2 fanout432 (.A(_12277_),
    .X(net432));
 sg13g2_buf_2 fanout433 (.A(_12181_),
    .X(net433));
 sg13g2_buf_2 fanout434 (.A(_11721_),
    .X(net434));
 sg13g2_buf_2 fanout435 (.A(_11660_),
    .X(net435));
 sg13g2_buf_2 fanout436 (.A(_11653_),
    .X(net436));
 sg13g2_buf_2 fanout437 (.A(_10631_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_10608_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_10606_),
    .X(net439));
 sg13g2_buf_2 fanout440 (.A(_10273_),
    .X(net440));
 sg13g2_buf_2 fanout441 (.A(_10019_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_09727_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_09700_),
    .X(net443));
 sg13g2_buf_2 fanout444 (.A(_09680_),
    .X(net444));
 sg13g2_buf_2 fanout445 (.A(_09658_),
    .X(net445));
 sg13g2_buf_2 fanout446 (.A(_09539_),
    .X(net446));
 sg13g2_buf_2 fanout447 (.A(_08757_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_08733_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_06969_),
    .X(net449));
 sg13g2_buf_2 fanout450 (.A(_06659_),
    .X(net450));
 sg13g2_buf_2 fanout451 (.A(_06657_),
    .X(net451));
 sg13g2_buf_2 fanout452 (.A(_06656_),
    .X(net452));
 sg13g2_buf_2 fanout453 (.A(_06303_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_06302_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_06301_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_06195_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_06194_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_06101_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_06100_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_05882_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_05873_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_05845_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_05125_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_03673_),
    .X(net464));
 sg13g2_buf_2 fanout465 (.A(_03672_),
    .X(net465));
 sg13g2_buf_2 fanout466 (.A(_03655_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_03643_),
    .X(net467));
 sg13g2_buf_1 fanout468 (.A(_03629_),
    .X(net468));
 sg13g2_buf_2 fanout469 (.A(_03621_),
    .X(net469));
 sg13g2_buf_2 fanout470 (.A(_03619_),
    .X(net470));
 sg13g2_buf_1 fanout471 (.A(_03614_),
    .X(net471));
 sg13g2_buf_4 fanout472 (.X(net472),
    .A(_03213_));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_03100_));
 sg13g2_buf_4 fanout474 (.X(net474),
    .A(_03097_));
 sg13g2_buf_4 fanout475 (.X(net475),
    .A(_03085_));
 sg13g2_buf_4 fanout476 (.X(net476),
    .A(_03076_));
 sg13g2_buf_4 fanout477 (.X(net477),
    .A(_03074_));
 sg13g2_buf_2 fanout478 (.A(_03047_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_03041_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_03037_),
    .X(net480));
 sg13g2_buf_2 fanout481 (.A(_03032_),
    .X(net481));
 sg13g2_buf_2 fanout482 (.A(_03028_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_03024_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_12672_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_11747_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_11745_),
    .X(net486));
 sg13g2_buf_2 fanout487 (.A(_11659_),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(_11444_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_11442_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_10235_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_10018_),
    .X(net491));
 sg13g2_buf_2 fanout492 (.A(_09298_),
    .X(net492));
 sg13g2_buf_2 fanout493 (.A(_09193_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_08916_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_08915_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_08777_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_08713_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_08300_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_07512_),
    .X(net499));
 sg13g2_buf_2 fanout500 (.A(_06189_),
    .X(net500));
 sg13g2_buf_2 fanout501 (.A(_06188_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_06183_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_06095_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_06094_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_06089_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_05961_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_05955_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_05941_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_05936_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_05910_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_05904_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_05890_),
    .X(net512));
 sg13g2_buf_2 fanout513 (.A(_05842_),
    .X(net513));
 sg13g2_buf_2 fanout514 (.A(_05119_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_04968_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_04961_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_04905_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_04868_),
    .X(net518));
 sg13g2_buf_2 fanout519 (.A(_04780_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_04768_),
    .X(net520));
 sg13g2_buf_4 fanout521 (.X(net521),
    .A(_04757_));
 sg13g2_buf_2 fanout522 (.A(_03678_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_03675_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_03674_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_03664_),
    .X(net525));
 sg13g2_buf_4 fanout526 (.X(net526),
    .A(_03663_));
 sg13g2_buf_2 fanout527 (.A(_03658_),
    .X(net527));
 sg13g2_buf_4 fanout528 (.X(net528),
    .A(_03654_));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_03646_));
 sg13g2_buf_2 fanout530 (.A(_03642_),
    .X(net530));
 sg13g2_buf_4 fanout531 (.X(net531),
    .A(_03628_));
 sg13g2_buf_2 fanout532 (.A(_03625_),
    .X(net532));
 sg13g2_buf_4 fanout533 (.X(net533),
    .A(_03620_));
 sg13g2_buf_1 fanout534 (.A(_03618_),
    .X(net534));
 sg13g2_buf_1 fanout535 (.A(_03616_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_03613_),
    .X(net536));
 sg13g2_buf_2 fanout537 (.A(_03611_),
    .X(net537));
 sg13g2_buf_4 fanout538 (.X(net538),
    .A(_03610_));
 sg13g2_buf_4 fanout539 (.X(net539),
    .A(_03101_));
 sg13g2_buf_4 fanout540 (.X(net540),
    .A(_03098_));
 sg13g2_buf_4 fanout541 (.X(net541),
    .A(_03086_));
 sg13g2_buf_2 fanout542 (.A(_03073_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_03046_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_03040_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_03036_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_03031_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_03027_),
    .X(net547));
 sg13g2_buf_2 fanout548 (.A(_03023_),
    .X(net548));
 sg13g2_buf_2 fanout549 (.A(_02861_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_02756_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_12518_),
    .X(net551));
 sg13g2_buf_2 fanout552 (.A(_12409_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_12109_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_11658_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_11655_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_11453_),
    .X(net556));
 sg13g2_buf_2 fanout557 (.A(_11443_),
    .X(net557));
 sg13g2_buf_2 fanout558 (.A(_10779_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_10731_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_10383_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_10270_),
    .X(net561));
 sg13g2_buf_2 fanout562 (.A(_10257_),
    .X(net562));
 sg13g2_buf_2 fanout563 (.A(_10165_),
    .X(net563));
 sg13g2_buf_2 fanout564 (.A(_10127_),
    .X(net564));
 sg13g2_buf_2 fanout565 (.A(_10041_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_10028_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_10017_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_09291_),
    .X(net568));
 sg13g2_buf_2 fanout569 (.A(_09192_),
    .X(net569));
 sg13g2_buf_4 fanout570 (.X(net570),
    .A(_08620_));
 sg13g2_buf_2 fanout571 (.A(_08533_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_08529_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_08519_),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(_08514_),
    .X(net574));
 sg13g2_buf_2 fanout575 (.A(_08512_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_08488_),
    .X(net576));
 sg13g2_buf_2 fanout577 (.A(_08479_),
    .X(net577));
 sg13g2_buf_2 fanout578 (.A(_08461_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_08459_),
    .X(net579));
 sg13g2_buf_2 fanout580 (.A(_08088_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_07965_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_07875_),
    .X(net582));
 sg13g2_buf_4 fanout583 (.X(net583),
    .A(_07835_));
 sg13g2_buf_2 fanout584 (.A(_07811_),
    .X(net584));
 sg13g2_buf_2 fanout585 (.A(_07784_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_07746_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_07712_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_07663_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_07591_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_07578_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_07299_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_06935_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_06745_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_05952_),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(_05940_),
    .X(net595));
 sg13g2_buf_2 fanout596 (.A(_05901_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_05889_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_05313_),
    .X(net598));
 sg13g2_buf_2 fanout599 (.A(_05161_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(_05152_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_05146_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_05138_),
    .X(net602));
 sg13g2_buf_2 fanout603 (.A(_05117_),
    .X(net603));
 sg13g2_buf_2 fanout604 (.A(_04861_),
    .X(net604));
 sg13g2_buf_2 fanout605 (.A(_04760_),
    .X(net605));
 sg13g2_buf_2 fanout606 (.A(_04756_),
    .X(net606));
 sg13g2_buf_2 fanout607 (.A(_04066_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_03677_),
    .X(net608));
 sg13g2_buf_2 fanout609 (.A(_03670_),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(_03669_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_03653_),
    .X(net611));
 sg13g2_buf_4 fanout612 (.X(net612),
    .A(_03651_));
 sg13g2_buf_4 fanout613 (.X(net613),
    .A(_03641_));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(_03636_));
 sg13g2_buf_4 fanout615 (.X(net615),
    .A(_03627_));
 sg13g2_buf_4 fanout616 (.X(net616),
    .A(_03624_));
 sg13g2_buf_2 fanout617 (.A(_03617_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_03615_),
    .X(net618));
 sg13g2_buf_4 fanout619 (.X(net619),
    .A(_03248_));
 sg13g2_buf_2 fanout620 (.A(_03072_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_03045_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_12563_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_12339_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_12177_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_12147_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_10954_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_10810_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_10807_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_10639_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_10291_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_10250_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_10216_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_10205_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_10201_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_10040_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_10027_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_09773_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_09641_),
    .X(net638));
 sg13g2_buf_2 fanout639 (.A(_09414_),
    .X(net639));
 sg13g2_buf_2 fanout640 (.A(_09390_),
    .X(net640));
 sg13g2_buf_2 fanout641 (.A(_09370_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_09360_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_09354_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_09349_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_09296_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_09284_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_09269_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_09191_),
    .X(net648));
 sg13g2_buf_4 fanout649 (.X(net649),
    .A(_08814_));
 sg13g2_buf_2 fanout650 (.A(_08736_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_08567_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_08532_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_08528_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_08518_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_08513_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_08487_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_08478_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_08460_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_08458_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_06966_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_06164_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_06069_),
    .X(net662));
 sg13g2_buf_4 fanout663 (.X(net663),
    .A(_05813_));
 sg13g2_buf_2 fanout664 (.A(_05160_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_04986_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_04962_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_04929_),
    .X(net667));
 sg13g2_buf_2 fanout668 (.A(_04900_),
    .X(net668));
 sg13g2_buf_2 fanout669 (.A(_04852_),
    .X(net669));
 sg13g2_buf_2 fanout670 (.A(_04843_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_04092_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_03687_),
    .X(net672));
 sg13g2_buf_2 fanout673 (.A(_03686_),
    .X(net673));
 sg13g2_buf_2 fanout674 (.A(_03051_),
    .X(net674));
 sg13g2_buf_2 fanout675 (.A(_12457_),
    .X(net675));
 sg13g2_buf_2 fanout676 (.A(_12224_),
    .X(net676));
 sg13g2_buf_2 fanout677 (.A(_12086_),
    .X(net677));
 sg13g2_buf_2 fanout678 (.A(_12085_),
    .X(net678));
 sg13g2_buf_2 fanout679 (.A(_12076_),
    .X(net679));
 sg13g2_buf_2 fanout680 (.A(_12014_),
    .X(net680));
 sg13g2_buf_2 fanout681 (.A(_10765_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(_10761_),
    .X(net682));
 sg13g2_buf_2 fanout683 (.A(_10753_),
    .X(net683));
 sg13g2_buf_2 fanout684 (.A(_10744_),
    .X(net684));
 sg13g2_buf_2 fanout685 (.A(_10737_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_10733_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_10730_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_10705_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_10655_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_10218_),
    .X(net690));
 sg13g2_buf_2 fanout691 (.A(_10197_),
    .X(net691));
 sg13g2_buf_2 fanout692 (.A(_10191_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_10188_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_10039_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_10026_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_09812_),
    .X(net696));
 sg13g2_buf_4 fanout697 (.X(net697),
    .A(_09600_));
 sg13g2_buf_2 fanout698 (.A(_09523_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_09482_),
    .X(net699));
 sg13g2_buf_4 fanout700 (.X(net700),
    .A(_09430_));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(_09398_));
 sg13g2_buf_4 fanout702 (.X(net702),
    .A(_09397_));
 sg13g2_buf_2 fanout703 (.A(_09366_),
    .X(net703));
 sg13g2_buf_2 fanout704 (.A(_09362_),
    .X(net704));
 sg13g2_buf_2 fanout705 (.A(_09353_),
    .X(net705));
 sg13g2_buf_2 fanout706 (.A(_09343_),
    .X(net706));
 sg13g2_buf_2 fanout707 (.A(_09340_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_09323_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_09315_));
 sg13g2_buf_8 fanout710 (.A(_09313_),
    .X(net710));
 sg13g2_buf_4 fanout711 (.X(net711),
    .A(_09309_));
 sg13g2_buf_4 fanout712 (.X(net712),
    .A(_09307_));
 sg13g2_buf_2 fanout713 (.A(_09304_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_09260_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_09190_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_09176_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_09107_),
    .X(net717));
 sg13g2_buf_2 fanout718 (.A(_08912_),
    .X(net718));
 sg13g2_buf_2 fanout719 (.A(_08888_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_08735_),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(_08632_),
    .X(net721));
 sg13g2_buf_4 fanout722 (.X(net722),
    .A(_08630_));
 sg13g2_buf_2 fanout723 (.A(_08624_),
    .X(net723));
 sg13g2_buf_4 fanout724 (.X(net724),
    .A(_08606_));
 sg13g2_buf_8 fanout725 (.A(_08605_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_08594_),
    .X(net726));
 sg13g2_buf_4 fanout727 (.X(net727),
    .A(_08556_));
 sg13g2_buf_8 fanout728 (.A(_08555_),
    .X(net728));
 sg13g2_buf_4 fanout729 (.X(net729),
    .A(_08547_));
 sg13g2_buf_8 fanout730 (.A(_08545_),
    .X(net730));
 sg13g2_buf_4 fanout731 (.X(net731),
    .A(_08543_));
 sg13g2_buf_4 fanout732 (.X(net732),
    .A(_08542_));
 sg13g2_buf_4 fanout733 (.X(net733),
    .A(_08494_));
 sg13g2_buf_2 fanout734 (.A(_08457_),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(_08423_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_06996_),
    .X(net736));
 sg13g2_buf_2 fanout737 (.A(_06856_),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(_06171_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_06169_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_06167_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_06166_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_06076_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_06074_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_06072_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_06071_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_05847_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_04859_),
    .X(net747));
 sg13g2_buf_2 fanout748 (.A(_03142_),
    .X(net748));
 sg13g2_buf_2 fanout749 (.A(_03102_),
    .X(net749));
 sg13g2_buf_1 fanout750 (.A(_03075_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_03066_),
    .X(net751));
 sg13g2_buf_2 fanout752 (.A(_03063_),
    .X(net752));
 sg13g2_buf_2 fanout753 (.A(_03060_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_03058_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_03050_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_02802_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_02746_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_02730_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_02727_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_02692_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_12703_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_12270_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_12266_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_12262_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_12241_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_12237_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_12122_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_12097_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_12084_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_12077_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_12075_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_12065_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_10829_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_10785_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_10757_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_10756_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_10732_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_10724_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_10680_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_10676_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_10668_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_10654_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_10650_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_10647_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_10642_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_10388_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_10248_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_10245_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_10210_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_10208_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_10200_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_10196_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_10190_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(_10187_),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_10180_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_10025_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_09971_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_09890_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_09776_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_09668_));
 sg13g2_buf_8 fanout801 (.A(_09599_),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_09526_));
 sg13g2_buf_8 fanout803 (.A(_09525_),
    .X(net803));
 sg13g2_buf_8 fanout804 (.A(_09435_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_09429_),
    .X(net805));
 sg13g2_buf_8 fanout806 (.A(_09428_),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(_09396_),
    .X(net807));
 sg13g2_buf_2 fanout808 (.A(_09320_),
    .X(net808));
 sg13g2_buf_4 fanout809 (.X(net809),
    .A(_09318_));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_09314_));
 sg13g2_buf_4 fanout811 (.X(net811),
    .A(_09312_));
 sg13g2_buf_2 fanout812 (.A(_09308_),
    .X(net812));
 sg13g2_buf_8 fanout813 (.A(_09306_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_09288_),
    .X(net814));
 sg13g2_buf_4 fanout815 (.X(net815),
    .A(_09259_));
 sg13g2_buf_2 fanout816 (.A(_09189_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_09175_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_09106_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_08972_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_08866_),
    .X(net820));
 sg13g2_buf_4 fanout821 (.X(net821),
    .A(_08636_));
 sg13g2_buf_2 fanout822 (.A(_08598_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_08593_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_08570_),
    .X(net824));
 sg13g2_buf_4 fanout825 (.X(net825),
    .A(_08560_));
 sg13g2_buf_8 fanout826 (.A(_08550_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_08520_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_08515_),
    .X(net828));
 sg13g2_buf_4 fanout829 (.X(net829),
    .A(_08493_));
 sg13g2_buf_2 fanout830 (.A(_08482_),
    .X(net830));
 sg13g2_buf_4 fanout831 (.X(net831),
    .A(_08472_));
 sg13g2_buf_2 fanout832 (.A(_08468_),
    .X(net832));
 sg13g2_buf_4 fanout833 (.X(net833),
    .A(_08464_));
 sg13g2_buf_4 fanout834 (.X(net834),
    .A(_08431_));
 sg13g2_buf_8 fanout835 (.A(_08430_),
    .X(net835));
 sg13g2_buf_4 fanout836 (.X(net836),
    .A(_08427_));
 sg13g2_buf_8 fanout837 (.A(_08426_),
    .X(net837));
 sg13g2_buf_4 fanout838 (.X(net838),
    .A(_08422_));
 sg13g2_buf_2 fanout839 (.A(_06970_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_06835_),
    .X(net840));
 sg13g2_buf_2 fanout841 (.A(_06674_),
    .X(net841));
 sg13g2_buf_2 fanout842 (.A(_06474_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_06473_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_06471_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_06469_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_06460_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_06456_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_06436_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_06431_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_06430_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_06421_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_06400_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_06394_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_06388_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_06375_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_06304_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_06174_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_06173_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_06079_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_06078_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_05965_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_05914_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_05894_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_05878_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_05877_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_05855_),
    .X(net866));
 sg13g2_buf_2 fanout867 (.A(_05818_),
    .X(net867));
 sg13g2_buf_2 fanout868 (.A(_05815_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_04845_),
    .X(net869));
 sg13g2_buf_2 fanout870 (.A(_04758_),
    .X(net870));
 sg13g2_buf_2 fanout871 (.A(_04056_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_04045_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_03665_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_03648_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_03647_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_03603_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_03141_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_03105_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_03104_),
    .X(net879));
 sg13g2_buf_1 fanout880 (.A(_03084_),
    .X(net880));
 sg13g2_buf_1 fanout881 (.A(_03083_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_03082_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_03080_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_03078_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_03071_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_03069_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_03065_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_03062_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_03059_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_03057_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_02749_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_02743_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_12269_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_12265_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_12261_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_12240_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_12236_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_12161_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_12083_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_12074_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_12064_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_10696_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_10675_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_10672_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_10667_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_10661_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_10653_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_10646_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_10644_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_10628_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_10228_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_10199_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_10195_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_10189_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_10184_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_10176_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_10169_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_10167_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_10139_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_10135_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_09986_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_09970_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_09889_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_09547_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_09500_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_09455_),
    .X(net926));
 sg13g2_buf_4 fanout927 (.X(net927),
    .A(_09427_));
 sg13g2_buf_4 fanout928 (.X(net928),
    .A(_09319_));
 sg13g2_buf_2 fanout929 (.A(_09258_),
    .X(net929));
 sg13g2_buf_4 fanout930 (.X(net930),
    .A(_09188_));
 sg13g2_buf_2 fanout931 (.A(_09179_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_09174_),
    .X(net932));
 sg13g2_buf_4 fanout933 (.X(net933),
    .A(_09105_));
 sg13g2_buf_2 fanout934 (.A(_08958_),
    .X(net934));
 sg13g2_buf_2 fanout935 (.A(_08886_),
    .X(net935));
 sg13g2_buf_4 fanout936 (.X(net936),
    .A(_08788_));
 sg13g2_buf_4 fanout937 (.X(net937),
    .A(_08637_));
 sg13g2_buf_2 fanout938 (.A(_08569_),
    .X(net938));
 sg13g2_buf_4 fanout939 (.X(net939),
    .A(_08551_));
 sg13g2_buf_2 fanout940 (.A(_08481_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_08475_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_08471_),
    .X(net942));
 sg13g2_buf_4 fanout943 (.X(net943),
    .A(_08465_));
 sg13g2_buf_4 fanout944 (.X(net944),
    .A(_08463_));
 sg13g2_buf_4 fanout945 (.X(net945),
    .A(_08438_));
 sg13g2_buf_4 fanout946 (.X(net946),
    .A(_08434_));
 sg13g2_buf_2 fanout947 (.A(_08421_),
    .X(net947));
 sg13g2_buf_4 fanout948 (.X(net948),
    .A(_08366_));
 sg13g2_buf_4 fanout949 (.X(net949),
    .A(_08360_));
 sg13g2_buf_2 fanout950 (.A(_08338_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_08244_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_07350_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_07295_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_07287_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_07272_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_07252_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_07249_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_06971_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_06776_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_06673_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_06499_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_06498_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_06497_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_06495_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_06459_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_06458_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_06439_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_06435_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_06434_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_06426_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_05954_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_05953_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_05946_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_05930_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_05929_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_05903_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_05902_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_05833_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_05820_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_05807_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_05781_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_04844_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_04765_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_04750_),
    .X(net984));
 sg13g2_buf_2 fanout985 (.A(_04713_),
    .X(net985));
 sg13g2_buf_2 fanout986 (.A(_04639_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_04611_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_04577_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_04280_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_04222_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_03747_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_03602_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_03571_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_03140_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_03081_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_03079_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_03077_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_03070_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_03068_),
    .X(net999));
 sg13g2_buf_4 fanout1000 (.X(net1000),
    .A(_03056_));
 sg13g2_buf_2 fanout1001 (.A(_03011_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_02950_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_02921_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_02674_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_12715_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_12698_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_12695_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_12668_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_12652_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_12632_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_12549_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_12509_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_12499_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_12450_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_12447_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_12434_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_12422_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_12335_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_12310_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_12304_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_12296_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_12259_),
    .X(net1022));
 sg13g2_buf_4 fanout1023 (.X(net1023),
    .A(_12251_));
 sg13g2_buf_2 fanout1024 (.A(_12246_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_12195_),
    .X(net1025));
 sg13g2_buf_4 fanout1026 (.X(net1026),
    .A(_12185_));
 sg13g2_buf_4 fanout1027 (.X(net1027),
    .A(_12168_));
 sg13g2_buf_2 fanout1028 (.A(_12150_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_12148_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_12140_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_12102_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_12068_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_12054_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_11661_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_11336_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_11334_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_11297_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_10728_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_10671_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_10666_),
    .X(net1040));
 sg13g2_buf_2 fanout1041 (.A(_10660_),
    .X(net1041));
 sg13g2_buf_2 fanout1042 (.A(_10640_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_10633_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_10557_),
    .X(net1044));
 sg13g2_buf_2 fanout1045 (.A(_10316_),
    .X(net1045));
 sg13g2_buf_2 fanout1046 (.A(_10198_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_10194_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_10183_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_10182_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_10141_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_10138_),
    .X(net1051));
 sg13g2_buf_2 fanout1052 (.A(_10132_),
    .X(net1052));
 sg13g2_buf_2 fanout1053 (.A(_10069_),
    .X(net1053));
 sg13g2_buf_2 fanout1054 (.A(_10063_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_10042_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_10016_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_10000_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_09993_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_09985_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_09979_),
    .X(net1060));
 sg13g2_buf_2 fanout1061 (.A(_09894_),
    .X(net1061));
 sg13g2_buf_2 fanout1062 (.A(_09845_),
    .X(net1062));
 sg13g2_buf_2 fanout1063 (.A(_09819_),
    .X(net1063));
 sg13g2_buf_2 fanout1064 (.A(_09453_),
    .X(net1064));
 sg13g2_buf_2 fanout1065 (.A(_09350_),
    .X(net1065));
 sg13g2_buf_2 fanout1066 (.A(_09243_),
    .X(net1066));
 sg13g2_buf_2 fanout1067 (.A(_09194_),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(_09187_),
    .X(net1068));
 sg13g2_buf_2 fanout1069 (.A(_09178_),
    .X(net1069));
 sg13g2_buf_2 fanout1070 (.A(_09173_),
    .X(net1070));
 sg13g2_buf_2 fanout1071 (.A(_09104_),
    .X(net1071));
 sg13g2_buf_2 fanout1072 (.A(_09093_),
    .X(net1072));
 sg13g2_buf_2 fanout1073 (.A(_09055_),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(_08863_),
    .X(net1074));
 sg13g2_buf_2 fanout1075 (.A(_08541_),
    .X(net1075));
 sg13g2_buf_2 fanout1076 (.A(_08525_),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(_08470_),
    .X(net1077));
 sg13g2_buf_2 fanout1078 (.A(_08462_),
    .X(net1078));
 sg13g2_buf_2 fanout1079 (.A(_08449_),
    .X(net1079));
 sg13g2_buf_2 fanout1080 (.A(_08424_),
    .X(net1080));
 sg13g2_buf_2 fanout1081 (.A(_08378_),
    .X(net1081));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(_08332_));
 sg13g2_buf_4 fanout1083 (.X(net1083),
    .A(_08315_));
 sg13g2_buf_4 fanout1084 (.X(net1084),
    .A(_08313_));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(_08311_));
 sg13g2_buf_2 fanout1086 (.A(_08278_),
    .X(net1086));
 sg13g2_buf_2 fanout1087 (.A(_08260_),
    .X(net1087));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(_08257_));
 sg13g2_buf_2 fanout1089 (.A(_08254_),
    .X(net1089));
 sg13g2_buf_4 fanout1090 (.X(net1090),
    .A(_08251_));
 sg13g2_buf_2 fanout1091 (.A(_08243_),
    .X(net1091));
 sg13g2_buf_2 fanout1092 (.A(_08053_),
    .X(net1092));
 sg13g2_buf_2 fanout1093 (.A(_08050_),
    .X(net1093));
 sg13g2_buf_2 fanout1094 (.A(_08036_),
    .X(net1094));
 sg13g2_buf_2 fanout1095 (.A(_07987_),
    .X(net1095));
 sg13g2_buf_2 fanout1096 (.A(_07349_),
    .X(net1096));
 sg13g2_buf_2 fanout1097 (.A(_07270_),
    .X(net1097));
 sg13g2_buf_2 fanout1098 (.A(_07266_),
    .X(net1098));
 sg13g2_buf_2 fanout1099 (.A(_07250_),
    .X(net1099));
 sg13g2_buf_2 fanout1100 (.A(_05797_),
    .X(net1100));
 sg13g2_buf_2 fanout1101 (.A(_02777_),
    .X(net1101));
 sg13g2_buf_2 fanout1102 (.A(_02772_),
    .X(net1102));
 sg13g2_buf_2 fanout1103 (.A(_12730_),
    .X(net1103));
 sg13g2_buf_2 fanout1104 (.A(_12691_),
    .X(net1104));
 sg13g2_buf_2 fanout1105 (.A(_12303_),
    .X(net1105));
 sg13g2_buf_2 fanout1106 (.A(_12250_),
    .X(net1106));
 sg13g2_buf_2 fanout1107 (.A(_12221_),
    .X(net1107));
 sg13g2_buf_2 fanout1108 (.A(_12214_),
    .X(net1108));
 sg13g2_buf_2 fanout1109 (.A(_12207_),
    .X(net1109));
 sg13g2_buf_2 fanout1110 (.A(_12184_),
    .X(net1110));
 sg13g2_buf_2 fanout1111 (.A(_12167_),
    .X(net1111));
 sg13g2_buf_2 fanout1112 (.A(_12151_),
    .X(net1112));
 sg13g2_buf_2 fanout1113 (.A(_12146_),
    .X(net1113));
 sg13g2_buf_2 fanout1114 (.A(_12125_),
    .X(net1114));
 sg13g2_buf_2 fanout1115 (.A(_12120_),
    .X(net1115));
 sg13g2_buf_2 fanout1116 (.A(_12104_),
    .X(net1116));
 sg13g2_buf_2 fanout1117 (.A(_12100_),
    .X(net1117));
 sg13g2_buf_2 fanout1118 (.A(_12094_),
    .X(net1118));
 sg13g2_buf_2 fanout1119 (.A(_12053_),
    .X(net1119));
 sg13g2_buf_2 fanout1120 (.A(_11874_),
    .X(net1120));
 sg13g2_buf_2 fanout1121 (.A(_11831_),
    .X(net1121));
 sg13g2_buf_2 fanout1122 (.A(_11720_),
    .X(net1122));
 sg13g2_buf_2 fanout1123 (.A(_11375_),
    .X(net1123));
 sg13g2_buf_2 fanout1124 (.A(_10798_),
    .X(net1124));
 sg13g2_buf_2 fanout1125 (.A(_10743_),
    .X(net1125));
 sg13g2_buf_2 fanout1126 (.A(_10662_),
    .X(net1126));
 sg13g2_buf_2 fanout1127 (.A(_10626_),
    .X(net1127));
 sg13g2_buf_2 fanout1128 (.A(_10613_),
    .X(net1128));
 sg13g2_buf_2 fanout1129 (.A(_10612_),
    .X(net1129));
 sg13g2_buf_2 fanout1130 (.A(_10455_),
    .X(net1130));
 sg13g2_buf_2 fanout1131 (.A(_10450_),
    .X(net1131));
 sg13g2_buf_2 fanout1132 (.A(_10376_),
    .X(net1132));
 sg13g2_buf_2 fanout1133 (.A(_10375_),
    .X(net1133));
 sg13g2_buf_2 fanout1134 (.A(_10338_),
    .X(net1134));
 sg13g2_buf_2 fanout1135 (.A(_10322_),
    .X(net1135));
 sg13g2_buf_2 fanout1136 (.A(_10312_),
    .X(net1136));
 sg13g2_buf_2 fanout1137 (.A(_10233_),
    .X(net1137));
 sg13g2_buf_2 fanout1138 (.A(_10158_),
    .X(net1138));
 sg13g2_buf_2 fanout1139 (.A(_10156_),
    .X(net1139));
 sg13g2_buf_2 fanout1140 (.A(_10154_),
    .X(net1140));
 sg13g2_buf_2 fanout1141 (.A(_10147_),
    .X(net1141));
 sg13g2_buf_2 fanout1142 (.A(_10144_),
    .X(net1142));
 sg13g2_buf_2 fanout1143 (.A(_10143_),
    .X(net1143));
 sg13g2_buf_2 fanout1144 (.A(_09992_),
    .X(net1144));
 sg13g2_buf_2 fanout1145 (.A(_09818_),
    .X(net1145));
 sg13g2_buf_2 fanout1146 (.A(_09815_),
    .X(net1146));
 sg13g2_buf_2 fanout1147 (.A(_09807_),
    .X(net1147));
 sg13g2_buf_2 fanout1148 (.A(_09785_),
    .X(net1148));
 sg13g2_buf_2 fanout1149 (.A(_09774_),
    .X(net1149));
 sg13g2_buf_2 fanout1150 (.A(_09247_),
    .X(net1150));
 sg13g2_buf_2 fanout1151 (.A(_09203_),
    .X(net1151));
 sg13g2_buf_2 fanout1152 (.A(_09200_),
    .X(net1152));
 sg13g2_buf_2 fanout1153 (.A(_09172_),
    .X(net1153));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(_09166_));
 sg13g2_buf_2 fanout1155 (.A(_09100_),
    .X(net1155));
 sg13g2_buf_2 fanout1156 (.A(_09082_),
    .X(net1156));
 sg13g2_buf_2 fanout1157 (.A(_09054_),
    .X(net1157));
 sg13g2_buf_2 fanout1158 (.A(_08452_),
    .X(net1158));
 sg13g2_buf_2 fanout1159 (.A(_08451_),
    .X(net1159));
 sg13g2_buf_2 fanout1160 (.A(_08450_),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(_08377_),
    .X(net1161));
 sg13g2_buf_2 fanout1162 (.A(_08376_),
    .X(net1162));
 sg13g2_buf_2 fanout1163 (.A(_08301_),
    .X(net1163));
 sg13g2_buf_2 fanout1164 (.A(_08273_),
    .X(net1164));
 sg13g2_buf_2 fanout1165 (.A(_08271_),
    .X(net1165));
 sg13g2_buf_2 fanout1166 (.A(_08270_),
    .X(net1166));
 sg13g2_tiehi _27592__1167 (.L_HI(net1167));
 sg13g2_tiehi _27593__1168 (.L_HI(net1168));
 sg13g2_tiehi _27594__1169 (.L_HI(net1169));
 sg13g2_tiehi _27595__1170 (.L_HI(net1170));
 sg13g2_tiehi _27596__1171 (.L_HI(net1171));
 sg13g2_tiehi \cpu.dcache.r_data[0][0]$_DFFE_PP__1172  (.L_HI(net1172));
 sg13g2_tiehi \cpu.dcache.r_data[0][10]$_DFFE_PP__1173  (.L_HI(net1173));
 sg13g2_tiehi \cpu.dcache.r_data[0][11]$_DFFE_PP__1174  (.L_HI(net1174));
 sg13g2_tiehi \cpu.dcache.r_data[0][12]$_DFFE_PP__1175  (.L_HI(net1175));
 sg13g2_tiehi \cpu.dcache.r_data[0][13]$_DFFE_PP__1176  (.L_HI(net1176));
 sg13g2_tiehi \cpu.dcache.r_data[0][14]$_DFFE_PP__1177  (.L_HI(net1177));
 sg13g2_tiehi \cpu.dcache.r_data[0][15]$_DFFE_PP__1178  (.L_HI(net1178));
 sg13g2_tiehi \cpu.dcache.r_data[0][16]$_DFFE_PP__1179  (.L_HI(net1179));
 sg13g2_tiehi \cpu.dcache.r_data[0][17]$_DFFE_PP__1180  (.L_HI(net1180));
 sg13g2_tiehi \cpu.dcache.r_data[0][18]$_DFFE_PP__1181  (.L_HI(net1181));
 sg13g2_tiehi \cpu.dcache.r_data[0][19]$_DFFE_PP__1182  (.L_HI(net1182));
 sg13g2_tiehi \cpu.dcache.r_data[0][1]$_DFFE_PP__1183  (.L_HI(net1183));
 sg13g2_tiehi \cpu.dcache.r_data[0][20]$_DFFE_PP__1184  (.L_HI(net1184));
 sg13g2_tiehi \cpu.dcache.r_data[0][21]$_DFFE_PP__1185  (.L_HI(net1185));
 sg13g2_tiehi \cpu.dcache.r_data[0][22]$_DFFE_PP__1186  (.L_HI(net1186));
 sg13g2_tiehi \cpu.dcache.r_data[0][23]$_DFFE_PP__1187  (.L_HI(net1187));
 sg13g2_tiehi \cpu.dcache.r_data[0][24]$_DFFE_PP__1188  (.L_HI(net1188));
 sg13g2_tiehi \cpu.dcache.r_data[0][25]$_DFFE_PP__1189  (.L_HI(net1189));
 sg13g2_tiehi \cpu.dcache.r_data[0][26]$_DFFE_PP__1190  (.L_HI(net1190));
 sg13g2_tiehi \cpu.dcache.r_data[0][27]$_DFFE_PP__1191  (.L_HI(net1191));
 sg13g2_tiehi \cpu.dcache.r_data[0][28]$_DFFE_PP__1192  (.L_HI(net1192));
 sg13g2_tiehi \cpu.dcache.r_data[0][29]$_DFFE_PP__1193  (.L_HI(net1193));
 sg13g2_tiehi \cpu.dcache.r_data[0][2]$_DFFE_PP__1194  (.L_HI(net1194));
 sg13g2_tiehi \cpu.dcache.r_data[0][30]$_DFFE_PP__1195  (.L_HI(net1195));
 sg13g2_tiehi \cpu.dcache.r_data[0][31]$_DFFE_PP__1196  (.L_HI(net1196));
 sg13g2_tiehi \cpu.dcache.r_data[0][3]$_DFFE_PP__1197  (.L_HI(net1197));
 sg13g2_tiehi \cpu.dcache.r_data[0][4]$_DFFE_PP__1198  (.L_HI(net1198));
 sg13g2_tiehi \cpu.dcache.r_data[0][5]$_DFFE_PP__1199  (.L_HI(net1199));
 sg13g2_tiehi \cpu.dcache.r_data[0][6]$_DFFE_PP__1200  (.L_HI(net1200));
 sg13g2_tiehi \cpu.dcache.r_data[0][7]$_DFFE_PP__1201  (.L_HI(net1201));
 sg13g2_tiehi \cpu.dcache.r_data[0][8]$_DFFE_PP__1202  (.L_HI(net1202));
 sg13g2_tiehi \cpu.dcache.r_data[0][9]$_DFFE_PP__1203  (.L_HI(net1203));
 sg13g2_tiehi \cpu.dcache.r_data[1][0]$_DFFE_PP__1204  (.L_HI(net1204));
 sg13g2_tiehi \cpu.dcache.r_data[1][10]$_DFFE_PP__1205  (.L_HI(net1205));
 sg13g2_tiehi \cpu.dcache.r_data[1][11]$_DFFE_PP__1206  (.L_HI(net1206));
 sg13g2_tiehi \cpu.dcache.r_data[1][12]$_DFFE_PP__1207  (.L_HI(net1207));
 sg13g2_tiehi \cpu.dcache.r_data[1][13]$_DFFE_PP__1208  (.L_HI(net1208));
 sg13g2_tiehi \cpu.dcache.r_data[1][14]$_DFFE_PP__1209  (.L_HI(net1209));
 sg13g2_tiehi \cpu.dcache.r_data[1][15]$_DFFE_PP__1210  (.L_HI(net1210));
 sg13g2_tiehi \cpu.dcache.r_data[1][16]$_DFFE_PP__1211  (.L_HI(net1211));
 sg13g2_tiehi \cpu.dcache.r_data[1][17]$_DFFE_PP__1212  (.L_HI(net1212));
 sg13g2_tiehi \cpu.dcache.r_data[1][18]$_DFFE_PP__1213  (.L_HI(net1213));
 sg13g2_tiehi \cpu.dcache.r_data[1][19]$_DFFE_PP__1214  (.L_HI(net1214));
 sg13g2_tiehi \cpu.dcache.r_data[1][1]$_DFFE_PP__1215  (.L_HI(net1215));
 sg13g2_tiehi \cpu.dcache.r_data[1][20]$_DFFE_PP__1216  (.L_HI(net1216));
 sg13g2_tiehi \cpu.dcache.r_data[1][21]$_DFFE_PP__1217  (.L_HI(net1217));
 sg13g2_tiehi \cpu.dcache.r_data[1][22]$_DFFE_PP__1218  (.L_HI(net1218));
 sg13g2_tiehi \cpu.dcache.r_data[1][23]$_DFFE_PP__1219  (.L_HI(net1219));
 sg13g2_tiehi \cpu.dcache.r_data[1][24]$_DFFE_PP__1220  (.L_HI(net1220));
 sg13g2_tiehi \cpu.dcache.r_data[1][25]$_DFFE_PP__1221  (.L_HI(net1221));
 sg13g2_tiehi \cpu.dcache.r_data[1][26]$_DFFE_PP__1222  (.L_HI(net1222));
 sg13g2_tiehi \cpu.dcache.r_data[1][27]$_DFFE_PP__1223  (.L_HI(net1223));
 sg13g2_tiehi \cpu.dcache.r_data[1][28]$_DFFE_PP__1224  (.L_HI(net1224));
 sg13g2_tiehi \cpu.dcache.r_data[1][29]$_DFFE_PP__1225  (.L_HI(net1225));
 sg13g2_tiehi \cpu.dcache.r_data[1][2]$_DFFE_PP__1226  (.L_HI(net1226));
 sg13g2_tiehi \cpu.dcache.r_data[1][30]$_DFFE_PP__1227  (.L_HI(net1227));
 sg13g2_tiehi \cpu.dcache.r_data[1][31]$_DFFE_PP__1228  (.L_HI(net1228));
 sg13g2_tiehi \cpu.dcache.r_data[1][3]$_DFFE_PP__1229  (.L_HI(net1229));
 sg13g2_tiehi \cpu.dcache.r_data[1][4]$_DFFE_PP__1230  (.L_HI(net1230));
 sg13g2_tiehi \cpu.dcache.r_data[1][5]$_DFFE_PP__1231  (.L_HI(net1231));
 sg13g2_tiehi \cpu.dcache.r_data[1][6]$_DFFE_PP__1232  (.L_HI(net1232));
 sg13g2_tiehi \cpu.dcache.r_data[1][7]$_DFFE_PP__1233  (.L_HI(net1233));
 sg13g2_tiehi \cpu.dcache.r_data[1][8]$_DFFE_PP__1234  (.L_HI(net1234));
 sg13g2_tiehi \cpu.dcache.r_data[1][9]$_DFFE_PP__1235  (.L_HI(net1235));
 sg13g2_tiehi \cpu.dcache.r_data[2][0]$_DFFE_PP__1236  (.L_HI(net1236));
 sg13g2_tiehi \cpu.dcache.r_data[2][10]$_DFFE_PP__1237  (.L_HI(net1237));
 sg13g2_tiehi \cpu.dcache.r_data[2][11]$_DFFE_PP__1238  (.L_HI(net1238));
 sg13g2_tiehi \cpu.dcache.r_data[2][12]$_DFFE_PP__1239  (.L_HI(net1239));
 sg13g2_tiehi \cpu.dcache.r_data[2][13]$_DFFE_PP__1240  (.L_HI(net1240));
 sg13g2_tiehi \cpu.dcache.r_data[2][14]$_DFFE_PP__1241  (.L_HI(net1241));
 sg13g2_tiehi \cpu.dcache.r_data[2][15]$_DFFE_PP__1242  (.L_HI(net1242));
 sg13g2_tiehi \cpu.dcache.r_data[2][16]$_DFFE_PP__1243  (.L_HI(net1243));
 sg13g2_tiehi \cpu.dcache.r_data[2][17]$_DFFE_PP__1244  (.L_HI(net1244));
 sg13g2_tiehi \cpu.dcache.r_data[2][18]$_DFFE_PP__1245  (.L_HI(net1245));
 sg13g2_tiehi \cpu.dcache.r_data[2][19]$_DFFE_PP__1246  (.L_HI(net1246));
 sg13g2_tiehi \cpu.dcache.r_data[2][1]$_DFFE_PP__1247  (.L_HI(net1247));
 sg13g2_tiehi \cpu.dcache.r_data[2][20]$_DFFE_PP__1248  (.L_HI(net1248));
 sg13g2_tiehi \cpu.dcache.r_data[2][21]$_DFFE_PP__1249  (.L_HI(net1249));
 sg13g2_tiehi \cpu.dcache.r_data[2][22]$_DFFE_PP__1250  (.L_HI(net1250));
 sg13g2_tiehi \cpu.dcache.r_data[2][23]$_DFFE_PP__1251  (.L_HI(net1251));
 sg13g2_tiehi \cpu.dcache.r_data[2][24]$_DFFE_PP__1252  (.L_HI(net1252));
 sg13g2_tiehi \cpu.dcache.r_data[2][25]$_DFFE_PP__1253  (.L_HI(net1253));
 sg13g2_tiehi \cpu.dcache.r_data[2][26]$_DFFE_PP__1254  (.L_HI(net1254));
 sg13g2_tiehi \cpu.dcache.r_data[2][27]$_DFFE_PP__1255  (.L_HI(net1255));
 sg13g2_tiehi \cpu.dcache.r_data[2][28]$_DFFE_PP__1256  (.L_HI(net1256));
 sg13g2_tiehi \cpu.dcache.r_data[2][29]$_DFFE_PP__1257  (.L_HI(net1257));
 sg13g2_tiehi \cpu.dcache.r_data[2][2]$_DFFE_PP__1258  (.L_HI(net1258));
 sg13g2_tiehi \cpu.dcache.r_data[2][30]$_DFFE_PP__1259  (.L_HI(net1259));
 sg13g2_tiehi \cpu.dcache.r_data[2][31]$_DFFE_PP__1260  (.L_HI(net1260));
 sg13g2_tiehi \cpu.dcache.r_data[2][3]$_DFFE_PP__1261  (.L_HI(net1261));
 sg13g2_tiehi \cpu.dcache.r_data[2][4]$_DFFE_PP__1262  (.L_HI(net1262));
 sg13g2_tiehi \cpu.dcache.r_data[2][5]$_DFFE_PP__1263  (.L_HI(net1263));
 sg13g2_tiehi \cpu.dcache.r_data[2][6]$_DFFE_PP__1264  (.L_HI(net1264));
 sg13g2_tiehi \cpu.dcache.r_data[2][7]$_DFFE_PP__1265  (.L_HI(net1265));
 sg13g2_tiehi \cpu.dcache.r_data[2][8]$_DFFE_PP__1266  (.L_HI(net1266));
 sg13g2_tiehi \cpu.dcache.r_data[2][9]$_DFFE_PP__1267  (.L_HI(net1267));
 sg13g2_tiehi \cpu.dcache.r_data[3][0]$_DFFE_PP__1268  (.L_HI(net1268));
 sg13g2_tiehi \cpu.dcache.r_data[3][10]$_DFFE_PP__1269  (.L_HI(net1269));
 sg13g2_tiehi \cpu.dcache.r_data[3][11]$_DFFE_PP__1270  (.L_HI(net1270));
 sg13g2_tiehi \cpu.dcache.r_data[3][12]$_DFFE_PP__1271  (.L_HI(net1271));
 sg13g2_tiehi \cpu.dcache.r_data[3][13]$_DFFE_PP__1272  (.L_HI(net1272));
 sg13g2_tiehi \cpu.dcache.r_data[3][14]$_DFFE_PP__1273  (.L_HI(net1273));
 sg13g2_tiehi \cpu.dcache.r_data[3][15]$_DFFE_PP__1274  (.L_HI(net1274));
 sg13g2_tiehi \cpu.dcache.r_data[3][16]$_DFFE_PP__1275  (.L_HI(net1275));
 sg13g2_tiehi \cpu.dcache.r_data[3][17]$_DFFE_PP__1276  (.L_HI(net1276));
 sg13g2_tiehi \cpu.dcache.r_data[3][18]$_DFFE_PP__1277  (.L_HI(net1277));
 sg13g2_tiehi \cpu.dcache.r_data[3][19]$_DFFE_PP__1278  (.L_HI(net1278));
 sg13g2_tiehi \cpu.dcache.r_data[3][1]$_DFFE_PP__1279  (.L_HI(net1279));
 sg13g2_tiehi \cpu.dcache.r_data[3][20]$_DFFE_PP__1280  (.L_HI(net1280));
 sg13g2_tiehi \cpu.dcache.r_data[3][21]$_DFFE_PP__1281  (.L_HI(net1281));
 sg13g2_tiehi \cpu.dcache.r_data[3][22]$_DFFE_PP__1282  (.L_HI(net1282));
 sg13g2_tiehi \cpu.dcache.r_data[3][23]$_DFFE_PP__1283  (.L_HI(net1283));
 sg13g2_tiehi \cpu.dcache.r_data[3][24]$_DFFE_PP__1284  (.L_HI(net1284));
 sg13g2_tiehi \cpu.dcache.r_data[3][25]$_DFFE_PP__1285  (.L_HI(net1285));
 sg13g2_tiehi \cpu.dcache.r_data[3][26]$_DFFE_PP__1286  (.L_HI(net1286));
 sg13g2_tiehi \cpu.dcache.r_data[3][27]$_DFFE_PP__1287  (.L_HI(net1287));
 sg13g2_tiehi \cpu.dcache.r_data[3][28]$_DFFE_PP__1288  (.L_HI(net1288));
 sg13g2_tiehi \cpu.dcache.r_data[3][29]$_DFFE_PP__1289  (.L_HI(net1289));
 sg13g2_tiehi \cpu.dcache.r_data[3][2]$_DFFE_PP__1290  (.L_HI(net1290));
 sg13g2_tiehi \cpu.dcache.r_data[3][30]$_DFFE_PP__1291  (.L_HI(net1291));
 sg13g2_tiehi \cpu.dcache.r_data[3][31]$_DFFE_PP__1292  (.L_HI(net1292));
 sg13g2_tiehi \cpu.dcache.r_data[3][3]$_DFFE_PP__1293  (.L_HI(net1293));
 sg13g2_tiehi \cpu.dcache.r_data[3][4]$_DFFE_PP__1294  (.L_HI(net1294));
 sg13g2_tiehi \cpu.dcache.r_data[3][5]$_DFFE_PP__1295  (.L_HI(net1295));
 sg13g2_tiehi \cpu.dcache.r_data[3][6]$_DFFE_PP__1296  (.L_HI(net1296));
 sg13g2_tiehi \cpu.dcache.r_data[3][7]$_DFFE_PP__1297  (.L_HI(net1297));
 sg13g2_tiehi \cpu.dcache.r_data[3][8]$_DFFE_PP__1298  (.L_HI(net1298));
 sg13g2_tiehi \cpu.dcache.r_data[3][9]$_DFFE_PP__1299  (.L_HI(net1299));
 sg13g2_tiehi \cpu.dcache.r_data[4][0]$_DFFE_PP__1300  (.L_HI(net1300));
 sg13g2_tiehi \cpu.dcache.r_data[4][10]$_DFFE_PP__1301  (.L_HI(net1301));
 sg13g2_tiehi \cpu.dcache.r_data[4][11]$_DFFE_PP__1302  (.L_HI(net1302));
 sg13g2_tiehi \cpu.dcache.r_data[4][12]$_DFFE_PP__1303  (.L_HI(net1303));
 sg13g2_tiehi \cpu.dcache.r_data[4][13]$_DFFE_PP__1304  (.L_HI(net1304));
 sg13g2_tiehi \cpu.dcache.r_data[4][14]$_DFFE_PP__1305  (.L_HI(net1305));
 sg13g2_tiehi \cpu.dcache.r_data[4][15]$_DFFE_PP__1306  (.L_HI(net1306));
 sg13g2_tiehi \cpu.dcache.r_data[4][16]$_DFFE_PP__1307  (.L_HI(net1307));
 sg13g2_tiehi \cpu.dcache.r_data[4][17]$_DFFE_PP__1308  (.L_HI(net1308));
 sg13g2_tiehi \cpu.dcache.r_data[4][18]$_DFFE_PP__1309  (.L_HI(net1309));
 sg13g2_tiehi \cpu.dcache.r_data[4][19]$_DFFE_PP__1310  (.L_HI(net1310));
 sg13g2_tiehi \cpu.dcache.r_data[4][1]$_DFFE_PP__1311  (.L_HI(net1311));
 sg13g2_tiehi \cpu.dcache.r_data[4][20]$_DFFE_PP__1312  (.L_HI(net1312));
 sg13g2_tiehi \cpu.dcache.r_data[4][21]$_DFFE_PP__1313  (.L_HI(net1313));
 sg13g2_tiehi \cpu.dcache.r_data[4][22]$_DFFE_PP__1314  (.L_HI(net1314));
 sg13g2_tiehi \cpu.dcache.r_data[4][23]$_DFFE_PP__1315  (.L_HI(net1315));
 sg13g2_tiehi \cpu.dcache.r_data[4][24]$_DFFE_PP__1316  (.L_HI(net1316));
 sg13g2_tiehi \cpu.dcache.r_data[4][25]$_DFFE_PP__1317  (.L_HI(net1317));
 sg13g2_tiehi \cpu.dcache.r_data[4][26]$_DFFE_PP__1318  (.L_HI(net1318));
 sg13g2_tiehi \cpu.dcache.r_data[4][27]$_DFFE_PP__1319  (.L_HI(net1319));
 sg13g2_tiehi \cpu.dcache.r_data[4][28]$_DFFE_PP__1320  (.L_HI(net1320));
 sg13g2_tiehi \cpu.dcache.r_data[4][29]$_DFFE_PP__1321  (.L_HI(net1321));
 sg13g2_tiehi \cpu.dcache.r_data[4][2]$_DFFE_PP__1322  (.L_HI(net1322));
 sg13g2_tiehi \cpu.dcache.r_data[4][30]$_DFFE_PP__1323  (.L_HI(net1323));
 sg13g2_tiehi \cpu.dcache.r_data[4][31]$_DFFE_PP__1324  (.L_HI(net1324));
 sg13g2_tiehi \cpu.dcache.r_data[4][3]$_DFFE_PP__1325  (.L_HI(net1325));
 sg13g2_tiehi \cpu.dcache.r_data[4][4]$_DFFE_PP__1326  (.L_HI(net1326));
 sg13g2_tiehi \cpu.dcache.r_data[4][5]$_DFFE_PP__1327  (.L_HI(net1327));
 sg13g2_tiehi \cpu.dcache.r_data[4][6]$_DFFE_PP__1328  (.L_HI(net1328));
 sg13g2_tiehi \cpu.dcache.r_data[4][7]$_DFFE_PP__1329  (.L_HI(net1329));
 sg13g2_tiehi \cpu.dcache.r_data[4][8]$_DFFE_PP__1330  (.L_HI(net1330));
 sg13g2_tiehi \cpu.dcache.r_data[4][9]$_DFFE_PP__1331  (.L_HI(net1331));
 sg13g2_tiehi \cpu.dcache.r_data[5][0]$_DFFE_PP__1332  (.L_HI(net1332));
 sg13g2_tiehi \cpu.dcache.r_data[5][10]$_DFFE_PP__1333  (.L_HI(net1333));
 sg13g2_tiehi \cpu.dcache.r_data[5][11]$_DFFE_PP__1334  (.L_HI(net1334));
 sg13g2_tiehi \cpu.dcache.r_data[5][12]$_DFFE_PP__1335  (.L_HI(net1335));
 sg13g2_tiehi \cpu.dcache.r_data[5][13]$_DFFE_PP__1336  (.L_HI(net1336));
 sg13g2_tiehi \cpu.dcache.r_data[5][14]$_DFFE_PP__1337  (.L_HI(net1337));
 sg13g2_tiehi \cpu.dcache.r_data[5][15]$_DFFE_PP__1338  (.L_HI(net1338));
 sg13g2_tiehi \cpu.dcache.r_data[5][16]$_DFFE_PP__1339  (.L_HI(net1339));
 sg13g2_tiehi \cpu.dcache.r_data[5][17]$_DFFE_PP__1340  (.L_HI(net1340));
 sg13g2_tiehi \cpu.dcache.r_data[5][18]$_DFFE_PP__1341  (.L_HI(net1341));
 sg13g2_tiehi \cpu.dcache.r_data[5][19]$_DFFE_PP__1342  (.L_HI(net1342));
 sg13g2_tiehi \cpu.dcache.r_data[5][1]$_DFFE_PP__1343  (.L_HI(net1343));
 sg13g2_tiehi \cpu.dcache.r_data[5][20]$_DFFE_PP__1344  (.L_HI(net1344));
 sg13g2_tiehi \cpu.dcache.r_data[5][21]$_DFFE_PP__1345  (.L_HI(net1345));
 sg13g2_tiehi \cpu.dcache.r_data[5][22]$_DFFE_PP__1346  (.L_HI(net1346));
 sg13g2_tiehi \cpu.dcache.r_data[5][23]$_DFFE_PP__1347  (.L_HI(net1347));
 sg13g2_tiehi \cpu.dcache.r_data[5][24]$_DFFE_PP__1348  (.L_HI(net1348));
 sg13g2_tiehi \cpu.dcache.r_data[5][25]$_DFFE_PP__1349  (.L_HI(net1349));
 sg13g2_tiehi \cpu.dcache.r_data[5][26]$_DFFE_PP__1350  (.L_HI(net1350));
 sg13g2_tiehi \cpu.dcache.r_data[5][27]$_DFFE_PP__1351  (.L_HI(net1351));
 sg13g2_tiehi \cpu.dcache.r_data[5][28]$_DFFE_PP__1352  (.L_HI(net1352));
 sg13g2_tiehi \cpu.dcache.r_data[5][29]$_DFFE_PP__1353  (.L_HI(net1353));
 sg13g2_tiehi \cpu.dcache.r_data[5][2]$_DFFE_PP__1354  (.L_HI(net1354));
 sg13g2_tiehi \cpu.dcache.r_data[5][30]$_DFFE_PP__1355  (.L_HI(net1355));
 sg13g2_tiehi \cpu.dcache.r_data[5][31]$_DFFE_PP__1356  (.L_HI(net1356));
 sg13g2_tiehi \cpu.dcache.r_data[5][3]$_DFFE_PP__1357  (.L_HI(net1357));
 sg13g2_tiehi \cpu.dcache.r_data[5][4]$_DFFE_PP__1358  (.L_HI(net1358));
 sg13g2_tiehi \cpu.dcache.r_data[5][5]$_DFFE_PP__1359  (.L_HI(net1359));
 sg13g2_tiehi \cpu.dcache.r_data[5][6]$_DFFE_PP__1360  (.L_HI(net1360));
 sg13g2_tiehi \cpu.dcache.r_data[5][7]$_DFFE_PP__1361  (.L_HI(net1361));
 sg13g2_tiehi \cpu.dcache.r_data[5][8]$_DFFE_PP__1362  (.L_HI(net1362));
 sg13g2_tiehi \cpu.dcache.r_data[5][9]$_DFFE_PP__1363  (.L_HI(net1363));
 sg13g2_tiehi \cpu.dcache.r_data[6][0]$_DFFE_PP__1364  (.L_HI(net1364));
 sg13g2_tiehi \cpu.dcache.r_data[6][10]$_DFFE_PP__1365  (.L_HI(net1365));
 sg13g2_tiehi \cpu.dcache.r_data[6][11]$_DFFE_PP__1366  (.L_HI(net1366));
 sg13g2_tiehi \cpu.dcache.r_data[6][12]$_DFFE_PP__1367  (.L_HI(net1367));
 sg13g2_tiehi \cpu.dcache.r_data[6][13]$_DFFE_PP__1368  (.L_HI(net1368));
 sg13g2_tiehi \cpu.dcache.r_data[6][14]$_DFFE_PP__1369  (.L_HI(net1369));
 sg13g2_tiehi \cpu.dcache.r_data[6][15]$_DFFE_PP__1370  (.L_HI(net1370));
 sg13g2_tiehi \cpu.dcache.r_data[6][16]$_DFFE_PP__1371  (.L_HI(net1371));
 sg13g2_tiehi \cpu.dcache.r_data[6][17]$_DFFE_PP__1372  (.L_HI(net1372));
 sg13g2_tiehi \cpu.dcache.r_data[6][18]$_DFFE_PP__1373  (.L_HI(net1373));
 sg13g2_tiehi \cpu.dcache.r_data[6][19]$_DFFE_PP__1374  (.L_HI(net1374));
 sg13g2_tiehi \cpu.dcache.r_data[6][1]$_DFFE_PP__1375  (.L_HI(net1375));
 sg13g2_tiehi \cpu.dcache.r_data[6][20]$_DFFE_PP__1376  (.L_HI(net1376));
 sg13g2_tiehi \cpu.dcache.r_data[6][21]$_DFFE_PP__1377  (.L_HI(net1377));
 sg13g2_tiehi \cpu.dcache.r_data[6][22]$_DFFE_PP__1378  (.L_HI(net1378));
 sg13g2_tiehi \cpu.dcache.r_data[6][23]$_DFFE_PP__1379  (.L_HI(net1379));
 sg13g2_tiehi \cpu.dcache.r_data[6][24]$_DFFE_PP__1380  (.L_HI(net1380));
 sg13g2_tiehi \cpu.dcache.r_data[6][25]$_DFFE_PP__1381  (.L_HI(net1381));
 sg13g2_tiehi \cpu.dcache.r_data[6][26]$_DFFE_PP__1382  (.L_HI(net1382));
 sg13g2_tiehi \cpu.dcache.r_data[6][27]$_DFFE_PP__1383  (.L_HI(net1383));
 sg13g2_tiehi \cpu.dcache.r_data[6][28]$_DFFE_PP__1384  (.L_HI(net1384));
 sg13g2_tiehi \cpu.dcache.r_data[6][29]$_DFFE_PP__1385  (.L_HI(net1385));
 sg13g2_tiehi \cpu.dcache.r_data[6][2]$_DFFE_PP__1386  (.L_HI(net1386));
 sg13g2_tiehi \cpu.dcache.r_data[6][30]$_DFFE_PP__1387  (.L_HI(net1387));
 sg13g2_tiehi \cpu.dcache.r_data[6][31]$_DFFE_PP__1388  (.L_HI(net1388));
 sg13g2_tiehi \cpu.dcache.r_data[6][3]$_DFFE_PP__1389  (.L_HI(net1389));
 sg13g2_tiehi \cpu.dcache.r_data[6][4]$_DFFE_PP__1390  (.L_HI(net1390));
 sg13g2_tiehi \cpu.dcache.r_data[6][5]$_DFFE_PP__1391  (.L_HI(net1391));
 sg13g2_tiehi \cpu.dcache.r_data[6][6]$_DFFE_PP__1392  (.L_HI(net1392));
 sg13g2_tiehi \cpu.dcache.r_data[6][7]$_DFFE_PP__1393  (.L_HI(net1393));
 sg13g2_tiehi \cpu.dcache.r_data[6][8]$_DFFE_PP__1394  (.L_HI(net1394));
 sg13g2_tiehi \cpu.dcache.r_data[6][9]$_DFFE_PP__1395  (.L_HI(net1395));
 sg13g2_tiehi \cpu.dcache.r_data[7][0]$_DFFE_PP__1396  (.L_HI(net1396));
 sg13g2_tiehi \cpu.dcache.r_data[7][10]$_DFFE_PP__1397  (.L_HI(net1397));
 sg13g2_tiehi \cpu.dcache.r_data[7][11]$_DFFE_PP__1398  (.L_HI(net1398));
 sg13g2_tiehi \cpu.dcache.r_data[7][12]$_DFFE_PP__1399  (.L_HI(net1399));
 sg13g2_tiehi \cpu.dcache.r_data[7][13]$_DFFE_PP__1400  (.L_HI(net1400));
 sg13g2_tiehi \cpu.dcache.r_data[7][14]$_DFFE_PP__1401  (.L_HI(net1401));
 sg13g2_tiehi \cpu.dcache.r_data[7][15]$_DFFE_PP__1402  (.L_HI(net1402));
 sg13g2_tiehi \cpu.dcache.r_data[7][16]$_DFFE_PP__1403  (.L_HI(net1403));
 sg13g2_tiehi \cpu.dcache.r_data[7][17]$_DFFE_PP__1404  (.L_HI(net1404));
 sg13g2_tiehi \cpu.dcache.r_data[7][18]$_DFFE_PP__1405  (.L_HI(net1405));
 sg13g2_tiehi \cpu.dcache.r_data[7][19]$_DFFE_PP__1406  (.L_HI(net1406));
 sg13g2_tiehi \cpu.dcache.r_data[7][1]$_DFFE_PP__1407  (.L_HI(net1407));
 sg13g2_tiehi \cpu.dcache.r_data[7][20]$_DFFE_PP__1408  (.L_HI(net1408));
 sg13g2_tiehi \cpu.dcache.r_data[7][21]$_DFFE_PP__1409  (.L_HI(net1409));
 sg13g2_tiehi \cpu.dcache.r_data[7][22]$_DFFE_PP__1410  (.L_HI(net1410));
 sg13g2_tiehi \cpu.dcache.r_data[7][23]$_DFFE_PP__1411  (.L_HI(net1411));
 sg13g2_tiehi \cpu.dcache.r_data[7][24]$_DFFE_PP__1412  (.L_HI(net1412));
 sg13g2_tiehi \cpu.dcache.r_data[7][25]$_DFFE_PP__1413  (.L_HI(net1413));
 sg13g2_tiehi \cpu.dcache.r_data[7][26]$_DFFE_PP__1414  (.L_HI(net1414));
 sg13g2_tiehi \cpu.dcache.r_data[7][27]$_DFFE_PP__1415  (.L_HI(net1415));
 sg13g2_tiehi \cpu.dcache.r_data[7][28]$_DFFE_PP__1416  (.L_HI(net1416));
 sg13g2_tiehi \cpu.dcache.r_data[7][29]$_DFFE_PP__1417  (.L_HI(net1417));
 sg13g2_tiehi \cpu.dcache.r_data[7][2]$_DFFE_PP__1418  (.L_HI(net1418));
 sg13g2_tiehi \cpu.dcache.r_data[7][30]$_DFFE_PP__1419  (.L_HI(net1419));
 sg13g2_tiehi \cpu.dcache.r_data[7][31]$_DFFE_PP__1420  (.L_HI(net1420));
 sg13g2_tiehi \cpu.dcache.r_data[7][3]$_DFFE_PP__1421  (.L_HI(net1421));
 sg13g2_tiehi \cpu.dcache.r_data[7][4]$_DFFE_PP__1422  (.L_HI(net1422));
 sg13g2_tiehi \cpu.dcache.r_data[7][5]$_DFFE_PP__1423  (.L_HI(net1423));
 sg13g2_tiehi \cpu.dcache.r_data[7][6]$_DFFE_PP__1424  (.L_HI(net1424));
 sg13g2_tiehi \cpu.dcache.r_data[7][7]$_DFFE_PP__1425  (.L_HI(net1425));
 sg13g2_tiehi \cpu.dcache.r_data[7][8]$_DFFE_PP__1426  (.L_HI(net1426));
 sg13g2_tiehi \cpu.dcache.r_data[7][9]$_DFFE_PP__1427  (.L_HI(net1427));
 sg13g2_tiehi \cpu.dcache.r_dirty[0]$_SDFFCE_PP1P__1428  (.L_HI(net1428));
 sg13g2_tiehi \cpu.dcache.r_dirty[1]$_SDFFCE_PP1P__1429  (.L_HI(net1429));
 sg13g2_tiehi \cpu.dcache.r_dirty[2]$_SDFFCE_PP1P__1430  (.L_HI(net1430));
 sg13g2_tiehi \cpu.dcache.r_dirty[3]$_SDFFCE_PP1P__1431  (.L_HI(net1431));
 sg13g2_tiehi \cpu.dcache.r_dirty[4]$_SDFFCE_PP1P__1432  (.L_HI(net1432));
 sg13g2_tiehi \cpu.dcache.r_dirty[5]$_SDFFCE_PP1P__1433  (.L_HI(net1433));
 sg13g2_tiehi \cpu.dcache.r_dirty[6]$_SDFFCE_PP1P__1434  (.L_HI(net1434));
 sg13g2_tiehi \cpu.dcache.r_dirty[7]$_SDFFCE_PP1P__1435  (.L_HI(net1435));
 sg13g2_tiehi \cpu.dcache.r_offset[0]$_SDFF_PN0__1436  (.L_HI(net1436));
 sg13g2_tiehi \cpu.dcache.r_offset[1]$_SDFF_PN0__1437  (.L_HI(net1437));
 sg13g2_tiehi \cpu.dcache.r_offset[2]$_SDFF_PN0__1438  (.L_HI(net1438));
 sg13g2_tiehi \cpu.dcache.r_tag[0][0]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \cpu.dcache.r_tag[0][10]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \cpu.dcache.r_tag[0][11]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \cpu.dcache.r_tag[0][12]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \cpu.dcache.r_tag[0][13]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \cpu.dcache.r_tag[0][14]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \cpu.dcache.r_tag[0][15]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \cpu.dcache.r_tag[0][16]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \cpu.dcache.r_tag[0][17]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \cpu.dcache.r_tag[0][18]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \cpu.dcache.r_tag[0][1]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \cpu.dcache.r_tag[0][2]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \cpu.dcache.r_tag[0][3]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \cpu.dcache.r_tag[0][4]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \cpu.dcache.r_tag[0][5]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \cpu.dcache.r_tag[0][6]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \cpu.dcache.r_tag[0][7]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \cpu.dcache.r_tag[0][8]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \cpu.dcache.r_tag[0][9]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \cpu.dcache.r_tag[1][0]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \cpu.dcache.r_tag[1][10]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \cpu.dcache.r_tag[1][11]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \cpu.dcache.r_tag[1][12]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \cpu.dcache.r_tag[1][13]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \cpu.dcache.r_tag[1][14]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \cpu.dcache.r_tag[1][15]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \cpu.dcache.r_tag[1][16]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \cpu.dcache.r_tag[1][17]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \cpu.dcache.r_tag[1][18]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \cpu.dcache.r_tag[1][1]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \cpu.dcache.r_tag[1][2]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \cpu.dcache.r_tag[1][3]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \cpu.dcache.r_tag[1][4]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \cpu.dcache.r_tag[1][5]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \cpu.dcache.r_tag[1][6]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \cpu.dcache.r_tag[1][7]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \cpu.dcache.r_tag[1][8]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \cpu.dcache.r_tag[1][9]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \cpu.dcache.r_tag[2][0]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \cpu.dcache.r_tag[2][10]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \cpu.dcache.r_tag[2][11]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \cpu.dcache.r_tag[2][12]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \cpu.dcache.r_tag[2][13]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \cpu.dcache.r_tag[2][14]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \cpu.dcache.r_tag[2][15]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \cpu.dcache.r_tag[2][16]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \cpu.dcache.r_tag[2][17]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \cpu.dcache.r_tag[2][18]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \cpu.dcache.r_tag[2][1]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \cpu.dcache.r_tag[2][2]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \cpu.dcache.r_tag[2][3]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \cpu.dcache.r_tag[2][4]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \cpu.dcache.r_tag[2][5]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \cpu.dcache.r_tag[2][6]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \cpu.dcache.r_tag[2][7]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \cpu.dcache.r_tag[2][8]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \cpu.dcache.r_tag[2][9]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \cpu.dcache.r_tag[3][0]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \cpu.dcache.r_tag[3][10]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \cpu.dcache.r_tag[3][11]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \cpu.dcache.r_tag[3][12]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \cpu.dcache.r_tag[3][13]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \cpu.dcache.r_tag[3][14]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \cpu.dcache.r_tag[3][15]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \cpu.dcache.r_tag[3][16]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \cpu.dcache.r_tag[3][17]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \cpu.dcache.r_tag[3][18]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \cpu.dcache.r_tag[3][1]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \cpu.dcache.r_tag[3][2]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \cpu.dcache.r_tag[3][3]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \cpu.dcache.r_tag[3][4]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \cpu.dcache.r_tag[3][5]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \cpu.dcache.r_tag[3][6]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \cpu.dcache.r_tag[3][7]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \cpu.dcache.r_tag[3][8]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \cpu.dcache.r_tag[3][9]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \cpu.dcache.r_tag[4][0]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \cpu.dcache.r_tag[4][10]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \cpu.dcache.r_tag[4][11]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \cpu.dcache.r_tag[4][12]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \cpu.dcache.r_tag[4][13]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \cpu.dcache.r_tag[4][14]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \cpu.dcache.r_tag[4][15]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \cpu.dcache.r_tag[4][16]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \cpu.dcache.r_tag[4][17]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \cpu.dcache.r_tag[4][18]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \cpu.dcache.r_tag[4][1]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \cpu.dcache.r_tag[4][2]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \cpu.dcache.r_tag[4][3]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \cpu.dcache.r_tag[4][4]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \cpu.dcache.r_tag[4][5]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \cpu.dcache.r_tag[4][6]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \cpu.dcache.r_tag[4][7]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \cpu.dcache.r_tag[4][8]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \cpu.dcache.r_tag[4][9]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \cpu.dcache.r_tag[5][0]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \cpu.dcache.r_tag[5][10]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \cpu.dcache.r_tag[5][11]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \cpu.dcache.r_tag[5][12]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \cpu.dcache.r_tag[5][13]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \cpu.dcache.r_tag[5][14]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \cpu.dcache.r_tag[5][15]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \cpu.dcache.r_tag[5][16]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \cpu.dcache.r_tag[5][17]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \cpu.dcache.r_tag[5][18]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \cpu.dcache.r_tag[5][1]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \cpu.dcache.r_tag[5][2]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \cpu.dcache.r_tag[5][3]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \cpu.dcache.r_tag[5][4]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \cpu.dcache.r_tag[5][5]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \cpu.dcache.r_tag[5][6]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \cpu.dcache.r_tag[5][7]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \cpu.dcache.r_tag[5][8]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \cpu.dcache.r_tag[5][9]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \cpu.dcache.r_tag[6][0]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \cpu.dcache.r_tag[6][10]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \cpu.dcache.r_tag[6][11]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \cpu.dcache.r_tag[6][12]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \cpu.dcache.r_tag[6][13]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \cpu.dcache.r_tag[6][14]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \cpu.dcache.r_tag[6][15]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \cpu.dcache.r_tag[6][16]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \cpu.dcache.r_tag[6][17]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \cpu.dcache.r_tag[6][18]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \cpu.dcache.r_tag[6][1]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \cpu.dcache.r_tag[6][2]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \cpu.dcache.r_tag[6][3]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \cpu.dcache.r_tag[6][4]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \cpu.dcache.r_tag[6][5]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \cpu.dcache.r_tag[6][6]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \cpu.dcache.r_tag[6][7]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \cpu.dcache.r_tag[6][8]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \cpu.dcache.r_tag[6][9]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \cpu.dcache.r_tag[7][0]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \cpu.dcache.r_tag[7][10]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \cpu.dcache.r_tag[7][11]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \cpu.dcache.r_tag[7][12]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \cpu.dcache.r_tag[7][13]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \cpu.dcache.r_tag[7][14]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \cpu.dcache.r_tag[7][15]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \cpu.dcache.r_tag[7][16]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \cpu.dcache.r_tag[7][17]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \cpu.dcache.r_tag[7][18]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \cpu.dcache.r_tag[7][1]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \cpu.dcache.r_tag[7][2]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \cpu.dcache.r_tag[7][3]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \cpu.dcache.r_tag[7][4]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \cpu.dcache.r_tag[7][5]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \cpu.dcache.r_tag[7][6]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \cpu.dcache.r_tag[7][7]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \cpu.dcache.r_tag[7][8]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \cpu.dcache.r_tag[7][9]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \cpu.dcache.r_valid[0]$_SDFFE_PP0P__1591  (.L_HI(net1591));
 sg13g2_tiehi \cpu.dcache.r_valid[1]$_SDFFE_PP0P__1592  (.L_HI(net1592));
 sg13g2_tiehi \cpu.dcache.r_valid[2]$_SDFFE_PP0P__1593  (.L_HI(net1593));
 sg13g2_tiehi \cpu.dcache.r_valid[3]$_SDFFE_PP0P__1594  (.L_HI(net1594));
 sg13g2_tiehi \cpu.dcache.r_valid[4]$_SDFFE_PP0P__1595  (.L_HI(net1595));
 sg13g2_tiehi \cpu.dcache.r_valid[5]$_SDFFE_PP0P__1596  (.L_HI(net1596));
 sg13g2_tiehi \cpu.dcache.r_valid[6]$_SDFFE_PP0P__1597  (.L_HI(net1597));
 sg13g2_tiehi \cpu.dcache.r_valid[7]$_SDFFE_PP0P__1598  (.L_HI(net1598));
 sg13g2_tiehi \cpu.dec.r_br$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \cpu.dec.r_cond[0]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \cpu.dec.r_cond[1]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \cpu.dec.r_cond[2]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \cpu.dec.r_div$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \cpu.dec.r_flush_all$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \cpu.dec.r_flush_write$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \cpu.dec.r_imm[0]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \cpu.dec.r_imm[10]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \cpu.dec.r_imm[11]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \cpu.dec.r_imm[12]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \cpu.dec.r_imm[13]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \cpu.dec.r_imm[14]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \cpu.dec.r_imm[15]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \cpu.dec.r_imm[1]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \cpu.dec.r_imm[2]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \cpu.dec.r_imm[3]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \cpu.dec.r_imm[4]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \cpu.dec.r_imm[5]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \cpu.dec.r_imm[6]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \cpu.dec.r_imm[7]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \cpu.dec.r_imm[8]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \cpu.dec.r_imm[9]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \cpu.dec.r_inv_mmu$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \cpu.dec.r_io$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \cpu.dec.r_jmp$_SDFFCE_PP0P__1624  (.L_HI(net1624));
 sg13g2_tiehi \cpu.dec.r_load$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \cpu.dec.r_mult$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \cpu.dec.r_needs_rs2$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \cpu.dec.r_op[10]$_DFF_P__1628  (.L_HI(net1628));
 sg13g2_tiehi \cpu.dec.r_op[1]$_DFF_P__1629  (.L_HI(net1629));
 sg13g2_tiehi \cpu.dec.r_op[2]$_DFF_P__1630  (.L_HI(net1630));
 sg13g2_tiehi \cpu.dec.r_op[3]$_DFF_P__1631  (.L_HI(net1631));
 sg13g2_tiehi \cpu.dec.r_op[4]$_DFF_P__1632  (.L_HI(net1632));
 sg13g2_tiehi \cpu.dec.r_op[5]$_DFF_P__1633  (.L_HI(net1633));
 sg13g2_tiehi \cpu.dec.r_op[6]$_DFF_P__1634  (.L_HI(net1634));
 sg13g2_tiehi \cpu.dec.r_op[7]$_DFF_P__1635  (.L_HI(net1635));
 sg13g2_tiehi \cpu.dec.r_op[8]$_DFF_P__1636  (.L_HI(net1636));
 sg13g2_tiehi \cpu.dec.r_op[9]$_DFF_P__1637  (.L_HI(net1637));
 sg13g2_tiehi \cpu.dec.r_rd[0]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \cpu.dec.r_rd[1]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \cpu.dec.r_rd[2]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \cpu.dec.r_rd[3]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \cpu.dec.r_ready$_DFF_P__1642  (.L_HI(net1642));
 sg13g2_tiehi \cpu.dec.r_rs1[0]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \cpu.dec.r_rs1[1]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \cpu.dec.r_rs1[2]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \cpu.dec.r_rs1[3]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \cpu.dec.r_rs2[0]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \cpu.dec.r_rs2[1]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \cpu.dec.r_rs2[2]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \cpu.dec.r_rs2[3]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \cpu.dec.r_rs2_pc$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \cpu.dec.r_set_cc$_SDFFCE_PP0P__1652  (.L_HI(net1652));
 sg13g2_tiehi \cpu.dec.r_store$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \cpu.dec.r_swapsp$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \cpu.dec.r_sys_call$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \cpu.dec.r_trap$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_d_proxy$_SDFFE_PP0P__1657  (.L_HI(net1657));
 sg13g2_tiehi \cpu.ex.genblk3.r_mmu_enable$_SDFFE_PN0P__1658  (.L_HI(net1658));
 sg13g2_tiehi \cpu.ex.genblk3.r_prev_supmode$_SDFFE_PN1P__1659  (.L_HI(net1659));
 sg13g2_tiehi \cpu.ex.genblk3.r_supmode$_DFF_P__1660  (.L_HI(net1660));
 sg13g2_tiehi \cpu.ex.genblk3.r_user_io$_SDFFE_PN0P__1661  (.L_HI(net1661));
 sg13g2_tiehi \cpu.ex.r_10[0]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \cpu.ex.r_10[10]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \cpu.ex.r_10[11]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \cpu.ex.r_10[12]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \cpu.ex.r_10[13]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \cpu.ex.r_10[14]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \cpu.ex.r_10[15]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \cpu.ex.r_10[1]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \cpu.ex.r_10[2]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \cpu.ex.r_10[3]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \cpu.ex.r_10[4]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \cpu.ex.r_10[5]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \cpu.ex.r_10[6]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \cpu.ex.r_10[7]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \cpu.ex.r_10[8]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \cpu.ex.r_10[9]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \cpu.ex.r_11[0]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \cpu.ex.r_11[10]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \cpu.ex.r_11[11]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \cpu.ex.r_11[12]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \cpu.ex.r_11[13]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \cpu.ex.r_11[14]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \cpu.ex.r_11[15]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \cpu.ex.r_11[1]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \cpu.ex.r_11[2]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \cpu.ex.r_11[3]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \cpu.ex.r_11[4]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \cpu.ex.r_11[5]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \cpu.ex.r_11[6]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \cpu.ex.r_11[7]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \cpu.ex.r_11[8]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \cpu.ex.r_11[9]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \cpu.ex.r_12[0]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \cpu.ex.r_12[10]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \cpu.ex.r_12[11]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \cpu.ex.r_12[12]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \cpu.ex.r_12[13]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \cpu.ex.r_12[14]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \cpu.ex.r_12[15]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \cpu.ex.r_12[1]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \cpu.ex.r_12[2]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \cpu.ex.r_12[3]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \cpu.ex.r_12[4]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \cpu.ex.r_12[5]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \cpu.ex.r_12[6]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \cpu.ex.r_12[7]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \cpu.ex.r_12[8]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \cpu.ex.r_12[9]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \cpu.ex.r_13[0]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \cpu.ex.r_13[10]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \cpu.ex.r_13[11]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \cpu.ex.r_13[12]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \cpu.ex.r_13[13]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \cpu.ex.r_13[14]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \cpu.ex.r_13[15]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \cpu.ex.r_13[1]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \cpu.ex.r_13[2]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \cpu.ex.r_13[3]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \cpu.ex.r_13[4]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \cpu.ex.r_13[5]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \cpu.ex.r_13[6]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \cpu.ex.r_13[7]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \cpu.ex.r_13[8]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \cpu.ex.r_13[9]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \cpu.ex.r_14[0]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \cpu.ex.r_14[10]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \cpu.ex.r_14[11]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \cpu.ex.r_14[12]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \cpu.ex.r_14[13]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \cpu.ex.r_14[14]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \cpu.ex.r_14[15]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \cpu.ex.r_14[1]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \cpu.ex.r_14[2]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \cpu.ex.r_14[3]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \cpu.ex.r_14[4]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \cpu.ex.r_14[5]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \cpu.ex.r_14[6]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \cpu.ex.r_14[7]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \cpu.ex.r_14[8]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \cpu.ex.r_14[9]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \cpu.ex.r_15[0]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \cpu.ex.r_15[10]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \cpu.ex.r_15[11]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \cpu.ex.r_15[12]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \cpu.ex.r_15[13]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \cpu.ex.r_15[14]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \cpu.ex.r_15[15]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \cpu.ex.r_15[1]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \cpu.ex.r_15[2]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \cpu.ex.r_15[3]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \cpu.ex.r_15[4]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \cpu.ex.r_15[5]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \cpu.ex.r_15[6]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \cpu.ex.r_15[7]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \cpu.ex.r_15[8]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \cpu.ex.r_15[9]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \cpu.ex.r_8[0]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \cpu.ex.r_8[10]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \cpu.ex.r_8[11]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \cpu.ex.r_8[12]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \cpu.ex.r_8[13]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \cpu.ex.r_8[14]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \cpu.ex.r_8[15]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \cpu.ex.r_8[1]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \cpu.ex.r_8[2]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \cpu.ex.r_8[3]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \cpu.ex.r_8[4]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \cpu.ex.r_8[5]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \cpu.ex.r_8[6]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \cpu.ex.r_8[7]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \cpu.ex.r_8[8]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \cpu.ex.r_8[9]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \cpu.ex.r_9[0]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \cpu.ex.r_9[10]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \cpu.ex.r_9[11]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \cpu.ex.r_9[12]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \cpu.ex.r_9[13]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \cpu.ex.r_9[14]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \cpu.ex.r_9[15]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \cpu.ex.r_9[1]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \cpu.ex.r_9[2]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \cpu.ex.r_9[3]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \cpu.ex.r_9[4]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \cpu.ex.r_9[5]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \cpu.ex.r_9[6]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \cpu.ex.r_9[7]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \cpu.ex.r_9[8]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \cpu.ex.r_9[9]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \cpu.ex.r_branch_stall$_DFF_P__1790  (.L_HI(net1790));
 sg13g2_tiehi \cpu.ex.r_d_flush_all$_SDFF_PP0__1791  (.L_HI(net1791));
 sg13g2_tiehi \cpu.ex.r_div_running$_DFF_P__1792  (.L_HI(net1792));
 sg13g2_tiehi \cpu.ex.r_epc[0]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \cpu.ex.r_epc[10]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \cpu.ex.r_epc[11]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \cpu.ex.r_epc[12]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \cpu.ex.r_epc[13]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \cpu.ex.r_epc[14]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \cpu.ex.r_epc[1]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \cpu.ex.r_epc[2]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \cpu.ex.r_epc[3]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \cpu.ex.r_epc[4]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \cpu.ex.r_epc[5]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \cpu.ex.r_epc[6]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \cpu.ex.r_epc[7]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \cpu.ex.r_epc[8]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \cpu.ex.r_epc[9]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \cpu.ex.r_fetch$_SDFF_PN1__1808  (.L_HI(net1808));
 sg13g2_tiehi \cpu.ex.r_flush_write$_SDFFE_PN0P__1809  (.L_HI(net1809));
 sg13g2_tiehi \cpu.ex.r_i_flush_all$_SDFF_PP0__1810  (.L_HI(net1810));
 sg13g2_tiehi \cpu.ex.r_ie$_SDFFE_PP0P__1811  (.L_HI(net1811));
 sg13g2_tiehi \cpu.ex.r_io_access$_SDFFE_PN0P__1812  (.L_HI(net1812));
 sg13g2_tiehi \cpu.ex.r_lr[0]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \cpu.ex.r_lr[10]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \cpu.ex.r_lr[11]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \cpu.ex.r_lr[12]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \cpu.ex.r_lr[13]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \cpu.ex.r_lr[14]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \cpu.ex.r_lr[1]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \cpu.ex.r_lr[2]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \cpu.ex.r_lr[3]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \cpu.ex.r_lr[4]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \cpu.ex.r_lr[5]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \cpu.ex.r_lr[6]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \cpu.ex.r_lr[7]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \cpu.ex.r_lr[8]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \cpu.ex.r_lr[9]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \cpu.ex.r_mult[0]$_DFF_P__1828  (.L_HI(net1828));
 sg13g2_tiehi \cpu.ex.r_mult[10]$_DFF_P__1829  (.L_HI(net1829));
 sg13g2_tiehi \cpu.ex.r_mult[11]$_DFF_P__1830  (.L_HI(net1830));
 sg13g2_tiehi \cpu.ex.r_mult[12]$_DFF_P__1831  (.L_HI(net1831));
 sg13g2_tiehi \cpu.ex.r_mult[13]$_DFF_P__1832  (.L_HI(net1832));
 sg13g2_tiehi \cpu.ex.r_mult[14]$_DFF_P__1833  (.L_HI(net1833));
 sg13g2_tiehi \cpu.ex.r_mult[15]$_DFF_P__1834  (.L_HI(net1834));
 sg13g2_tiehi \cpu.ex.r_mult[16]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \cpu.ex.r_mult[17]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \cpu.ex.r_mult[18]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \cpu.ex.r_mult[19]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \cpu.ex.r_mult[1]$_DFF_P__1839  (.L_HI(net1839));
 sg13g2_tiehi \cpu.ex.r_mult[20]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \cpu.ex.r_mult[21]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \cpu.ex.r_mult[22]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \cpu.ex.r_mult[23]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \cpu.ex.r_mult[24]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \cpu.ex.r_mult[25]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \cpu.ex.r_mult[26]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \cpu.ex.r_mult[27]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \cpu.ex.r_mult[28]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \cpu.ex.r_mult[29]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \cpu.ex.r_mult[2]$_DFF_P__1850  (.L_HI(net1850));
 sg13g2_tiehi \cpu.ex.r_mult[30]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \cpu.ex.r_mult[31]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \cpu.ex.r_mult[3]$_DFF_P__1853  (.L_HI(net1853));
 sg13g2_tiehi \cpu.ex.r_mult[4]$_DFF_P__1854  (.L_HI(net1854));
 sg13g2_tiehi \cpu.ex.r_mult[5]$_DFF_P__1855  (.L_HI(net1855));
 sg13g2_tiehi \cpu.ex.r_mult[6]$_DFF_P__1856  (.L_HI(net1856));
 sg13g2_tiehi \cpu.ex.r_mult[7]$_DFF_P__1857  (.L_HI(net1857));
 sg13g2_tiehi \cpu.ex.r_mult[8]$_DFF_P__1858  (.L_HI(net1858));
 sg13g2_tiehi \cpu.ex.r_mult[9]$_DFF_P__1859  (.L_HI(net1859));
 sg13g2_tiehi \cpu.ex.r_mult_off[0]$_DFF_P__1860  (.L_HI(net1860));
 sg13g2_tiehi \cpu.ex.r_mult_off[1]$_DFF_P__1861  (.L_HI(net1861));
 sg13g2_tiehi \cpu.ex.r_mult_off[2]$_DFF_P__1862  (.L_HI(net1862));
 sg13g2_tiehi \cpu.ex.r_mult_off[3]$_DFF_P__1863  (.L_HI(net1863));
 sg13g2_tiehi \cpu.ex.r_mult_running$_DFF_P__1864  (.L_HI(net1864));
 sg13g2_tiehi \cpu.ex.r_pc[0]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \cpu.ex.r_pc[10]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \cpu.ex.r_pc[11]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \cpu.ex.r_pc[12]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \cpu.ex.r_pc[13]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \cpu.ex.r_pc[14]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \cpu.ex.r_pc[1]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \cpu.ex.r_pc[2]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \cpu.ex.r_pc[3]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \cpu.ex.r_pc[4]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \cpu.ex.r_pc[5]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \cpu.ex.r_pc[6]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \cpu.ex.r_pc[7]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \cpu.ex.r_pc[8]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \cpu.ex.r_pc[9]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \cpu.ex.r_prev_ie$_SDFFE_PN0P__1880  (.L_HI(net1880));
 sg13g2_tiehi \cpu.ex.r_read_stall$_SDFFE_PN0P__1881  (.L_HI(net1881));
 sg13g2_tiehi \cpu.ex.r_sp[0]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \cpu.ex.r_sp[10]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \cpu.ex.r_sp[11]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \cpu.ex.r_sp[12]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \cpu.ex.r_sp[13]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \cpu.ex.r_sp[14]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \cpu.ex.r_sp[1]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \cpu.ex.r_sp[2]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \cpu.ex.r_sp[3]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \cpu.ex.r_sp[4]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \cpu.ex.r_sp[5]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \cpu.ex.r_sp[6]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \cpu.ex.r_sp[7]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \cpu.ex.r_sp[8]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \cpu.ex.r_sp[9]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \cpu.ex.r_stmp[0]$_SDFFCE_PN0P__1897  (.L_HI(net1897));
 sg13g2_tiehi \cpu.ex.r_stmp[10]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \cpu.ex.r_stmp[11]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \cpu.ex.r_stmp[12]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \cpu.ex.r_stmp[13]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \cpu.ex.r_stmp[14]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \cpu.ex.r_stmp[15]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \cpu.ex.r_stmp[1]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \cpu.ex.r_stmp[2]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \cpu.ex.r_stmp[3]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \cpu.ex.r_stmp[4]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \cpu.ex.r_stmp[5]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \cpu.ex.r_stmp[6]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \cpu.ex.r_stmp[7]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \cpu.ex.r_stmp[8]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \cpu.ex.r_stmp[9]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \cpu.ex.r_wb[0]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \cpu.ex.r_wb[10]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \cpu.ex.r_wb[11]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \cpu.ex.r_wb[12]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \cpu.ex.r_wb[13]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \cpu.ex.r_wb[14]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \cpu.ex.r_wb[15]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \cpu.ex.r_wb[1]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \cpu.ex.r_wb[2]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \cpu.ex.r_wb[3]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \cpu.ex.r_wb[4]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \cpu.ex.r_wb[5]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \cpu.ex.r_wb[6]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \cpu.ex.r_wb[7]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \cpu.ex.r_wb[8]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \cpu.ex.r_wb[9]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \cpu.ex.r_wb_addr[0]$_SDFFCE_PN0P__1929  (.L_HI(net1929));
 sg13g2_tiehi \cpu.ex.r_wb_addr[1]$_SDFFCE_PN0P__1930  (.L_HI(net1930));
 sg13g2_tiehi \cpu.ex.r_wb_addr[2]$_SDFFCE_PP0P__1931  (.L_HI(net1931));
 sg13g2_tiehi \cpu.ex.r_wb_addr[3]$_SDFFCE_PP0P__1932  (.L_HI(net1932));
 sg13g2_tiehi \cpu.ex.r_wb_swapsp$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \cpu.ex.r_wb_valid$_DFF_P__1934  (.L_HI(net1934));
 sg13g2_tiehi \cpu.ex.r_wdata[0]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \cpu.ex.r_wdata[10]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \cpu.ex.r_wdata[11]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \cpu.ex.r_wdata[12]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \cpu.ex.r_wdata[13]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \cpu.ex.r_wdata[14]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \cpu.ex.r_wdata[15]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \cpu.ex.r_wdata[1]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \cpu.ex.r_wdata[2]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \cpu.ex.r_wdata[3]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \cpu.ex.r_wdata[4]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \cpu.ex.r_wdata[5]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \cpu.ex.r_wdata[6]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \cpu.ex.r_wdata[7]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \cpu.ex.r_wdata[8]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \cpu.ex.r_wdata[9]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \cpu.ex.r_wmask[0]$_SDFFE_PP0P__1951  (.L_HI(net1951));
 sg13g2_tiehi \cpu.ex.r_wmask[1]$_SDFFE_PP0P__1952  (.L_HI(net1952));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[0]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[1]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[2]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_address[3]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_ins$_SDFFE_PN0P__1957  (.L_HI(net1957));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_sup$_SDFFE_PN0P__1958  (.L_HI(net1958));
 sg13g2_tiehi \cpu.genblk1.mmu.r_fault_type$_SDFFE_PN0P__1959  (.L_HI(net1959));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[0]$_SDFFE_PN0P__1960  (.L_HI(net1960));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[10]$_SDFFE_PN0P__1961  (.L_HI(net1961));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[11]$_SDFFE_PN0P__1962  (.L_HI(net1962));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[12]$_SDFFE_PN0P__1963  (.L_HI(net1963));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[13]$_SDFFE_PN0P__1964  (.L_HI(net1964));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[14]$_SDFFE_PN0P__1965  (.L_HI(net1965));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[15]$_SDFFE_PN0P__1966  (.L_HI(net1966));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[16]$_SDFFE_PN0P__1967  (.L_HI(net1967));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[17]$_SDFFE_PN0P__1968  (.L_HI(net1968));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[18]$_SDFFE_PN0P__1969  (.L_HI(net1969));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[19]$_SDFFE_PN0P__1970  (.L_HI(net1970));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[1]$_SDFFE_PN0P__1971  (.L_HI(net1971));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[20]$_SDFFE_PN0P__1972  (.L_HI(net1972));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[21]$_SDFFE_PN0P__1973  (.L_HI(net1973));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[22]$_SDFFE_PN0P__1974  (.L_HI(net1974));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[23]$_SDFFE_PN0P__1975  (.L_HI(net1975));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[24]$_SDFFE_PN0P__1976  (.L_HI(net1976));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[25]$_SDFFE_PN0P__1977  (.L_HI(net1977));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[26]$_SDFFE_PN0P__1978  (.L_HI(net1978));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[27]$_SDFFE_PN0P__1979  (.L_HI(net1979));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[28]$_SDFFE_PN0P__1980  (.L_HI(net1980));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[29]$_SDFFE_PN0P__1981  (.L_HI(net1981));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[2]$_SDFFE_PN0P__1982  (.L_HI(net1982));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[30]$_SDFFE_PN0P__1983  (.L_HI(net1983));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[31]$_SDFFE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[3]$_SDFFE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[4]$_SDFFE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[5]$_SDFFE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[6]$_SDFFE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[7]$_SDFFE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[8]$_SDFFE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_d[9]$_SDFFE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[0]$_SDFFE_PN0P__1992  (.L_HI(net1992));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[10]$_SDFFE_PN0P__1993  (.L_HI(net1993));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[11]$_SDFFE_PN0P__1994  (.L_HI(net1994));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[12]$_SDFFE_PN0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[13]$_SDFFE_PN0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[14]$_SDFFE_PN0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[15]$_SDFFE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[16]$_SDFFE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[17]$_SDFFE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[18]$_SDFFE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[19]$_SDFFE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[1]$_SDFFE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[20]$_SDFFE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[21]$_SDFFE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[22]$_SDFFE_PN0P__2006  (.L_HI(net2006));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[23]$_SDFFE_PN0P__2007  (.L_HI(net2007));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[24]$_SDFFE_PN0P__2008  (.L_HI(net2008));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[25]$_SDFFE_PN0P__2009  (.L_HI(net2009));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[26]$_SDFFE_PN0P__2010  (.L_HI(net2010));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[27]$_SDFFE_PN0P__2011  (.L_HI(net2011));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[28]$_SDFFE_PN0P__2012  (.L_HI(net2012));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[29]$_SDFFE_PN0P__2013  (.L_HI(net2013));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[2]$_SDFFE_PN0P__2014  (.L_HI(net2014));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[30]$_SDFFE_PN0P__2015  (.L_HI(net2015));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[31]$_SDFFE_PN0P__2016  (.L_HI(net2016));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[3]$_SDFFE_PN0P__2017  (.L_HI(net2017));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[4]$_SDFFE_PN0P__2018  (.L_HI(net2018));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[5]$_SDFFE_PN0P__2019  (.L_HI(net2019));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[6]$_SDFFE_PN0P__2020  (.L_HI(net2020));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[7]$_SDFFE_PN0P__2021  (.L_HI(net2021));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[8]$_SDFFE_PN0P__2022  (.L_HI(net2022));
 sg13g2_tiehi \cpu.genblk1.mmu.r_valid_i[9]$_SDFFE_PN0P__2023  (.L_HI(net2023));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][0]$_DFFE_PP__2024  (.L_HI(net2024));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][10]$_DFFE_PP__2025  (.L_HI(net2025));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][11]$_DFFE_PP__2026  (.L_HI(net2026));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][1]$_DFFE_PP__2027  (.L_HI(net2027));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][2]$_DFFE_PP__2028  (.L_HI(net2028));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][3]$_DFFE_PP__2029  (.L_HI(net2029));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][4]$_DFFE_PP__2030  (.L_HI(net2030));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][5]$_DFFE_PP__2031  (.L_HI(net2031));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][6]$_DFFE_PP__2032  (.L_HI(net2032));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][7]$_DFFE_PP__2033  (.L_HI(net2033));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][8]$_DFFE_PP__2034  (.L_HI(net2034));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[0][9]$_DFFE_PP__2035  (.L_HI(net2035));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][0]$_DFFE_PP__2036  (.L_HI(net2036));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][10]$_DFFE_PP__2037  (.L_HI(net2037));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][11]$_DFFE_PP__2038  (.L_HI(net2038));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][1]$_DFFE_PP__2039  (.L_HI(net2039));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][2]$_DFFE_PP__2040  (.L_HI(net2040));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][3]$_DFFE_PP__2041  (.L_HI(net2041));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][4]$_DFFE_PP__2042  (.L_HI(net2042));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][5]$_DFFE_PP__2043  (.L_HI(net2043));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][6]$_DFFE_PP__2044  (.L_HI(net2044));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][7]$_DFFE_PP__2045  (.L_HI(net2045));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][8]$_DFFE_PP__2046  (.L_HI(net2046));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[10][9]$_DFFE_PP__2047  (.L_HI(net2047));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][0]$_DFFE_PP__2048  (.L_HI(net2048));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][10]$_DFFE_PP__2049  (.L_HI(net2049));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][11]$_DFFE_PP__2050  (.L_HI(net2050));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][1]$_DFFE_PP__2051  (.L_HI(net2051));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][2]$_DFFE_PP__2052  (.L_HI(net2052));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][3]$_DFFE_PP__2053  (.L_HI(net2053));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][4]$_DFFE_PP__2054  (.L_HI(net2054));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][5]$_DFFE_PP__2055  (.L_HI(net2055));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][6]$_DFFE_PP__2056  (.L_HI(net2056));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][7]$_DFFE_PP__2057  (.L_HI(net2057));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][8]$_DFFE_PP__2058  (.L_HI(net2058));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[11][9]$_DFFE_PP__2059  (.L_HI(net2059));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][0]$_DFFE_PP__2060  (.L_HI(net2060));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][10]$_DFFE_PP__2061  (.L_HI(net2061));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][11]$_DFFE_PP__2062  (.L_HI(net2062));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][1]$_DFFE_PP__2063  (.L_HI(net2063));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][2]$_DFFE_PP__2064  (.L_HI(net2064));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][3]$_DFFE_PP__2065  (.L_HI(net2065));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][4]$_DFFE_PP__2066  (.L_HI(net2066));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][5]$_DFFE_PP__2067  (.L_HI(net2067));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][6]$_DFFE_PP__2068  (.L_HI(net2068));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][7]$_DFFE_PP__2069  (.L_HI(net2069));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][8]$_DFFE_PP__2070  (.L_HI(net2070));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[12][9]$_DFFE_PP__2071  (.L_HI(net2071));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][0]$_DFFE_PP__2072  (.L_HI(net2072));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][10]$_DFFE_PP__2073  (.L_HI(net2073));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][11]$_DFFE_PP__2074  (.L_HI(net2074));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][1]$_DFFE_PP__2075  (.L_HI(net2075));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][2]$_DFFE_PP__2076  (.L_HI(net2076));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][3]$_DFFE_PP__2077  (.L_HI(net2077));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][4]$_DFFE_PP__2078  (.L_HI(net2078));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][5]$_DFFE_PP__2079  (.L_HI(net2079));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][6]$_DFFE_PP__2080  (.L_HI(net2080));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][7]$_DFFE_PP__2081  (.L_HI(net2081));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][8]$_DFFE_PP__2082  (.L_HI(net2082));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[13][9]$_DFFE_PP__2083  (.L_HI(net2083));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][0]$_DFFE_PP__2084  (.L_HI(net2084));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][10]$_DFFE_PP__2085  (.L_HI(net2085));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][11]$_DFFE_PP__2086  (.L_HI(net2086));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][1]$_DFFE_PP__2087  (.L_HI(net2087));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][2]$_DFFE_PP__2088  (.L_HI(net2088));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][3]$_DFFE_PP__2089  (.L_HI(net2089));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][4]$_DFFE_PP__2090  (.L_HI(net2090));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][5]$_DFFE_PP__2091  (.L_HI(net2091));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][6]$_DFFE_PP__2092  (.L_HI(net2092));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][7]$_DFFE_PP__2093  (.L_HI(net2093));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][8]$_DFFE_PP__2094  (.L_HI(net2094));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[14][9]$_DFFE_PP__2095  (.L_HI(net2095));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][0]$_DFFE_PP__2096  (.L_HI(net2096));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][10]$_DFFE_PP__2097  (.L_HI(net2097));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][11]$_DFFE_PP__2098  (.L_HI(net2098));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][1]$_DFFE_PP__2099  (.L_HI(net2099));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][2]$_DFFE_PP__2100  (.L_HI(net2100));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][3]$_DFFE_PP__2101  (.L_HI(net2101));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][4]$_DFFE_PP__2102  (.L_HI(net2102));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][5]$_DFFE_PP__2103  (.L_HI(net2103));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][6]$_DFFE_PP__2104  (.L_HI(net2104));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][7]$_DFFE_PP__2105  (.L_HI(net2105));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][8]$_DFFE_PP__2106  (.L_HI(net2106));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[15][9]$_DFFE_PP__2107  (.L_HI(net2107));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][0]$_DFFE_PP__2108  (.L_HI(net2108));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][10]$_DFFE_PP__2109  (.L_HI(net2109));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][11]$_DFFE_PP__2110  (.L_HI(net2110));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][1]$_DFFE_PP__2111  (.L_HI(net2111));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][2]$_DFFE_PP__2112  (.L_HI(net2112));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][3]$_DFFE_PP__2113  (.L_HI(net2113));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][4]$_DFFE_PP__2114  (.L_HI(net2114));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][5]$_DFFE_PP__2115  (.L_HI(net2115));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][6]$_DFFE_PP__2116  (.L_HI(net2116));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][7]$_DFFE_PP__2117  (.L_HI(net2117));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][8]$_DFFE_PP__2118  (.L_HI(net2118));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[16][9]$_DFFE_PP__2119  (.L_HI(net2119));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][0]$_DFFE_PP__2120  (.L_HI(net2120));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][10]$_DFFE_PP__2121  (.L_HI(net2121));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][11]$_DFFE_PP__2122  (.L_HI(net2122));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][1]$_DFFE_PP__2123  (.L_HI(net2123));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][2]$_DFFE_PP__2124  (.L_HI(net2124));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][3]$_DFFE_PP__2125  (.L_HI(net2125));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][4]$_DFFE_PP__2126  (.L_HI(net2126));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][5]$_DFFE_PP__2127  (.L_HI(net2127));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][6]$_DFFE_PP__2128  (.L_HI(net2128));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][7]$_DFFE_PP__2129  (.L_HI(net2129));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][8]$_DFFE_PP__2130  (.L_HI(net2130));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[17][9]$_DFFE_PP__2131  (.L_HI(net2131));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][0]$_DFFE_PP__2132  (.L_HI(net2132));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][10]$_DFFE_PP__2133  (.L_HI(net2133));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][11]$_DFFE_PP__2134  (.L_HI(net2134));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][1]$_DFFE_PP__2135  (.L_HI(net2135));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][2]$_DFFE_PP__2136  (.L_HI(net2136));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][3]$_DFFE_PP__2137  (.L_HI(net2137));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][4]$_DFFE_PP__2138  (.L_HI(net2138));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][5]$_DFFE_PP__2139  (.L_HI(net2139));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][6]$_DFFE_PP__2140  (.L_HI(net2140));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][7]$_DFFE_PP__2141  (.L_HI(net2141));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][8]$_DFFE_PP__2142  (.L_HI(net2142));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[18][9]$_DFFE_PP__2143  (.L_HI(net2143));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][0]$_DFFE_PP__2144  (.L_HI(net2144));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][10]$_DFFE_PP__2145  (.L_HI(net2145));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][11]$_DFFE_PP__2146  (.L_HI(net2146));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][1]$_DFFE_PP__2147  (.L_HI(net2147));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][2]$_DFFE_PP__2148  (.L_HI(net2148));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][3]$_DFFE_PP__2149  (.L_HI(net2149));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][4]$_DFFE_PP__2150  (.L_HI(net2150));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][5]$_DFFE_PP__2151  (.L_HI(net2151));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][6]$_DFFE_PP__2152  (.L_HI(net2152));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][7]$_DFFE_PP__2153  (.L_HI(net2153));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][8]$_DFFE_PP__2154  (.L_HI(net2154));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[19][9]$_DFFE_PP__2155  (.L_HI(net2155));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][0]$_DFFE_PP__2156  (.L_HI(net2156));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][10]$_DFFE_PP__2157  (.L_HI(net2157));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][11]$_DFFE_PP__2158  (.L_HI(net2158));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][1]$_DFFE_PP__2159  (.L_HI(net2159));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][2]$_DFFE_PP__2160  (.L_HI(net2160));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][3]$_DFFE_PP__2161  (.L_HI(net2161));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][4]$_DFFE_PP__2162  (.L_HI(net2162));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][5]$_DFFE_PP__2163  (.L_HI(net2163));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][6]$_DFFE_PP__2164  (.L_HI(net2164));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][7]$_DFFE_PP__2165  (.L_HI(net2165));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][8]$_DFFE_PP__2166  (.L_HI(net2166));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[1][9]$_DFFE_PP__2167  (.L_HI(net2167));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][0]$_DFFE_PP__2168  (.L_HI(net2168));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][10]$_DFFE_PP__2169  (.L_HI(net2169));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][11]$_DFFE_PP__2170  (.L_HI(net2170));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][1]$_DFFE_PP__2171  (.L_HI(net2171));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][2]$_DFFE_PP__2172  (.L_HI(net2172));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][3]$_DFFE_PP__2173  (.L_HI(net2173));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][4]$_DFFE_PP__2174  (.L_HI(net2174));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][5]$_DFFE_PP__2175  (.L_HI(net2175));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][6]$_DFFE_PP__2176  (.L_HI(net2176));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][7]$_DFFE_PP__2177  (.L_HI(net2177));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][8]$_DFFE_PP__2178  (.L_HI(net2178));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[20][9]$_DFFE_PP__2179  (.L_HI(net2179));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][0]$_DFFE_PP__2180  (.L_HI(net2180));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][10]$_DFFE_PP__2181  (.L_HI(net2181));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][11]$_DFFE_PP__2182  (.L_HI(net2182));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][1]$_DFFE_PP__2183  (.L_HI(net2183));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][2]$_DFFE_PP__2184  (.L_HI(net2184));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][3]$_DFFE_PP__2185  (.L_HI(net2185));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][4]$_DFFE_PP__2186  (.L_HI(net2186));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][5]$_DFFE_PP__2187  (.L_HI(net2187));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][6]$_DFFE_PP__2188  (.L_HI(net2188));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][7]$_DFFE_PP__2189  (.L_HI(net2189));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][8]$_DFFE_PP__2190  (.L_HI(net2190));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[21][9]$_DFFE_PP__2191  (.L_HI(net2191));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][0]$_DFFE_PP__2192  (.L_HI(net2192));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][10]$_DFFE_PP__2193  (.L_HI(net2193));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][11]$_DFFE_PP__2194  (.L_HI(net2194));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][1]$_DFFE_PP__2195  (.L_HI(net2195));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][2]$_DFFE_PP__2196  (.L_HI(net2196));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][3]$_DFFE_PP__2197  (.L_HI(net2197));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][4]$_DFFE_PP__2198  (.L_HI(net2198));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][5]$_DFFE_PP__2199  (.L_HI(net2199));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][6]$_DFFE_PP__2200  (.L_HI(net2200));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][7]$_DFFE_PP__2201  (.L_HI(net2201));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][8]$_DFFE_PP__2202  (.L_HI(net2202));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[22][9]$_DFFE_PP__2203  (.L_HI(net2203));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][0]$_DFFE_PP__2204  (.L_HI(net2204));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][10]$_DFFE_PP__2205  (.L_HI(net2205));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][11]$_DFFE_PP__2206  (.L_HI(net2206));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][1]$_DFFE_PP__2207  (.L_HI(net2207));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][2]$_DFFE_PP__2208  (.L_HI(net2208));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][3]$_DFFE_PP__2209  (.L_HI(net2209));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][4]$_DFFE_PP__2210  (.L_HI(net2210));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][5]$_DFFE_PP__2211  (.L_HI(net2211));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][6]$_DFFE_PP__2212  (.L_HI(net2212));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][7]$_DFFE_PP__2213  (.L_HI(net2213));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][8]$_DFFE_PP__2214  (.L_HI(net2214));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[23][9]$_DFFE_PP__2215  (.L_HI(net2215));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][0]$_DFFE_PP__2216  (.L_HI(net2216));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][10]$_DFFE_PP__2217  (.L_HI(net2217));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][11]$_DFFE_PP__2218  (.L_HI(net2218));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][1]$_DFFE_PP__2219  (.L_HI(net2219));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][2]$_DFFE_PP__2220  (.L_HI(net2220));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][3]$_DFFE_PP__2221  (.L_HI(net2221));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][4]$_DFFE_PP__2222  (.L_HI(net2222));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][5]$_DFFE_PP__2223  (.L_HI(net2223));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][6]$_DFFE_PP__2224  (.L_HI(net2224));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][7]$_DFFE_PP__2225  (.L_HI(net2225));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][8]$_DFFE_PP__2226  (.L_HI(net2226));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[24][9]$_DFFE_PP__2227  (.L_HI(net2227));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][0]$_DFFE_PP__2228  (.L_HI(net2228));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][10]$_DFFE_PP__2229  (.L_HI(net2229));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][11]$_DFFE_PP__2230  (.L_HI(net2230));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][1]$_DFFE_PP__2231  (.L_HI(net2231));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][2]$_DFFE_PP__2232  (.L_HI(net2232));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][3]$_DFFE_PP__2233  (.L_HI(net2233));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][4]$_DFFE_PP__2234  (.L_HI(net2234));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][5]$_DFFE_PP__2235  (.L_HI(net2235));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][6]$_DFFE_PP__2236  (.L_HI(net2236));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][7]$_DFFE_PP__2237  (.L_HI(net2237));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][8]$_DFFE_PP__2238  (.L_HI(net2238));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[25][9]$_DFFE_PP__2239  (.L_HI(net2239));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][0]$_DFFE_PP__2240  (.L_HI(net2240));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][10]$_DFFE_PP__2241  (.L_HI(net2241));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][11]$_DFFE_PP__2242  (.L_HI(net2242));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][1]$_DFFE_PP__2243  (.L_HI(net2243));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][2]$_DFFE_PP__2244  (.L_HI(net2244));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][3]$_DFFE_PP__2245  (.L_HI(net2245));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][4]$_DFFE_PP__2246  (.L_HI(net2246));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][5]$_DFFE_PP__2247  (.L_HI(net2247));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][6]$_DFFE_PP__2248  (.L_HI(net2248));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][7]$_DFFE_PP__2249  (.L_HI(net2249));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][8]$_DFFE_PP__2250  (.L_HI(net2250));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[26][9]$_DFFE_PP__2251  (.L_HI(net2251));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][0]$_DFFE_PP__2252  (.L_HI(net2252));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][10]$_DFFE_PP__2253  (.L_HI(net2253));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][11]$_DFFE_PP__2254  (.L_HI(net2254));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][1]$_DFFE_PP__2255  (.L_HI(net2255));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][2]$_DFFE_PP__2256  (.L_HI(net2256));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][3]$_DFFE_PP__2257  (.L_HI(net2257));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][4]$_DFFE_PP__2258  (.L_HI(net2258));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][5]$_DFFE_PP__2259  (.L_HI(net2259));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][6]$_DFFE_PP__2260  (.L_HI(net2260));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][7]$_DFFE_PP__2261  (.L_HI(net2261));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][8]$_DFFE_PP__2262  (.L_HI(net2262));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[27][9]$_DFFE_PP__2263  (.L_HI(net2263));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][0]$_DFFE_PP__2264  (.L_HI(net2264));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][10]$_DFFE_PP__2265  (.L_HI(net2265));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][11]$_DFFE_PP__2266  (.L_HI(net2266));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][1]$_DFFE_PP__2267  (.L_HI(net2267));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][2]$_DFFE_PP__2268  (.L_HI(net2268));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][3]$_DFFE_PP__2269  (.L_HI(net2269));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][4]$_DFFE_PP__2270  (.L_HI(net2270));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][5]$_DFFE_PP__2271  (.L_HI(net2271));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][6]$_DFFE_PP__2272  (.L_HI(net2272));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][7]$_DFFE_PP__2273  (.L_HI(net2273));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][8]$_DFFE_PP__2274  (.L_HI(net2274));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[28][9]$_DFFE_PP__2275  (.L_HI(net2275));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][0]$_DFFE_PP__2276  (.L_HI(net2276));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][10]$_DFFE_PP__2277  (.L_HI(net2277));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][11]$_DFFE_PP__2278  (.L_HI(net2278));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][1]$_DFFE_PP__2279  (.L_HI(net2279));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][2]$_DFFE_PP__2280  (.L_HI(net2280));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][3]$_DFFE_PP__2281  (.L_HI(net2281));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][4]$_DFFE_PP__2282  (.L_HI(net2282));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][5]$_DFFE_PP__2283  (.L_HI(net2283));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][6]$_DFFE_PP__2284  (.L_HI(net2284));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][7]$_DFFE_PP__2285  (.L_HI(net2285));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][8]$_DFFE_PP__2286  (.L_HI(net2286));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[29][9]$_DFFE_PP__2287  (.L_HI(net2287));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][0]$_DFFE_PP__2288  (.L_HI(net2288));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][10]$_DFFE_PP__2289  (.L_HI(net2289));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][11]$_DFFE_PP__2290  (.L_HI(net2290));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][1]$_DFFE_PP__2291  (.L_HI(net2291));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][2]$_DFFE_PP__2292  (.L_HI(net2292));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][3]$_DFFE_PP__2293  (.L_HI(net2293));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][4]$_DFFE_PP__2294  (.L_HI(net2294));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][5]$_DFFE_PP__2295  (.L_HI(net2295));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][6]$_DFFE_PP__2296  (.L_HI(net2296));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][7]$_DFFE_PP__2297  (.L_HI(net2297));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][8]$_DFFE_PP__2298  (.L_HI(net2298));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[2][9]$_DFFE_PP__2299  (.L_HI(net2299));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][0]$_DFFE_PP__2300  (.L_HI(net2300));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][10]$_DFFE_PP__2301  (.L_HI(net2301));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][11]$_DFFE_PP__2302  (.L_HI(net2302));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][1]$_DFFE_PP__2303  (.L_HI(net2303));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][2]$_DFFE_PP__2304  (.L_HI(net2304));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][3]$_DFFE_PP__2305  (.L_HI(net2305));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][4]$_DFFE_PP__2306  (.L_HI(net2306));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][5]$_DFFE_PP__2307  (.L_HI(net2307));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][6]$_DFFE_PP__2308  (.L_HI(net2308));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][7]$_DFFE_PP__2309  (.L_HI(net2309));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][8]$_DFFE_PP__2310  (.L_HI(net2310));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[30][9]$_DFFE_PP__2311  (.L_HI(net2311));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][0]$_DFFE_PP__2312  (.L_HI(net2312));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][10]$_DFFE_PP__2313  (.L_HI(net2313));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][11]$_DFFE_PP__2314  (.L_HI(net2314));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][1]$_DFFE_PP__2315  (.L_HI(net2315));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][2]$_DFFE_PP__2316  (.L_HI(net2316));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][3]$_DFFE_PP__2317  (.L_HI(net2317));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][4]$_DFFE_PP__2318  (.L_HI(net2318));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][5]$_DFFE_PP__2319  (.L_HI(net2319));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][6]$_DFFE_PP__2320  (.L_HI(net2320));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][7]$_DFFE_PP__2321  (.L_HI(net2321));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][8]$_DFFE_PP__2322  (.L_HI(net2322));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[31][9]$_DFFE_PP__2323  (.L_HI(net2323));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][0]$_DFFE_PP__2324  (.L_HI(net2324));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][10]$_DFFE_PP__2325  (.L_HI(net2325));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][11]$_DFFE_PP__2326  (.L_HI(net2326));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][1]$_DFFE_PP__2327  (.L_HI(net2327));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][2]$_DFFE_PP__2328  (.L_HI(net2328));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][3]$_DFFE_PP__2329  (.L_HI(net2329));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][4]$_DFFE_PP__2330  (.L_HI(net2330));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][5]$_DFFE_PP__2331  (.L_HI(net2331));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][6]$_DFFE_PP__2332  (.L_HI(net2332));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][7]$_DFFE_PP__2333  (.L_HI(net2333));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][8]$_DFFE_PP__2334  (.L_HI(net2334));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[3][9]$_DFFE_PP__2335  (.L_HI(net2335));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][0]$_DFFE_PP__2336  (.L_HI(net2336));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][10]$_DFFE_PP__2337  (.L_HI(net2337));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][11]$_DFFE_PP__2338  (.L_HI(net2338));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][1]$_DFFE_PP__2339  (.L_HI(net2339));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][2]$_DFFE_PP__2340  (.L_HI(net2340));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][3]$_DFFE_PP__2341  (.L_HI(net2341));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][4]$_DFFE_PP__2342  (.L_HI(net2342));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][5]$_DFFE_PP__2343  (.L_HI(net2343));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][6]$_DFFE_PP__2344  (.L_HI(net2344));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][7]$_DFFE_PP__2345  (.L_HI(net2345));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][8]$_DFFE_PP__2346  (.L_HI(net2346));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[4][9]$_DFFE_PP__2347  (.L_HI(net2347));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][0]$_DFFE_PP__2348  (.L_HI(net2348));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][10]$_DFFE_PP__2349  (.L_HI(net2349));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][11]$_DFFE_PP__2350  (.L_HI(net2350));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][1]$_DFFE_PP__2351  (.L_HI(net2351));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][2]$_DFFE_PP__2352  (.L_HI(net2352));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][3]$_DFFE_PP__2353  (.L_HI(net2353));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][4]$_DFFE_PP__2354  (.L_HI(net2354));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][5]$_DFFE_PP__2355  (.L_HI(net2355));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][6]$_DFFE_PP__2356  (.L_HI(net2356));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][7]$_DFFE_PP__2357  (.L_HI(net2357));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][8]$_DFFE_PP__2358  (.L_HI(net2358));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[5][9]$_DFFE_PP__2359  (.L_HI(net2359));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][0]$_DFFE_PP__2360  (.L_HI(net2360));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][10]$_DFFE_PP__2361  (.L_HI(net2361));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][11]$_DFFE_PP__2362  (.L_HI(net2362));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][1]$_DFFE_PP__2363  (.L_HI(net2363));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][2]$_DFFE_PP__2364  (.L_HI(net2364));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][3]$_DFFE_PP__2365  (.L_HI(net2365));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][4]$_DFFE_PP__2366  (.L_HI(net2366));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][5]$_DFFE_PP__2367  (.L_HI(net2367));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][6]$_DFFE_PP__2368  (.L_HI(net2368));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][7]$_DFFE_PP__2369  (.L_HI(net2369));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][8]$_DFFE_PP__2370  (.L_HI(net2370));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[6][9]$_DFFE_PP__2371  (.L_HI(net2371));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][0]$_DFFE_PP__2372  (.L_HI(net2372));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][10]$_DFFE_PP__2373  (.L_HI(net2373));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][11]$_DFFE_PP__2374  (.L_HI(net2374));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][1]$_DFFE_PP__2375  (.L_HI(net2375));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][2]$_DFFE_PP__2376  (.L_HI(net2376));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][3]$_DFFE_PP__2377  (.L_HI(net2377));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][4]$_DFFE_PP__2378  (.L_HI(net2378));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][5]$_DFFE_PP__2379  (.L_HI(net2379));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][6]$_DFFE_PP__2380  (.L_HI(net2380));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][7]$_DFFE_PP__2381  (.L_HI(net2381));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][8]$_DFFE_PP__2382  (.L_HI(net2382));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[7][9]$_DFFE_PP__2383  (.L_HI(net2383));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][0]$_DFFE_PP__2384  (.L_HI(net2384));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][10]$_DFFE_PP__2385  (.L_HI(net2385));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][11]$_DFFE_PP__2386  (.L_HI(net2386));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][1]$_DFFE_PP__2387  (.L_HI(net2387));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][2]$_DFFE_PP__2388  (.L_HI(net2388));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][3]$_DFFE_PP__2389  (.L_HI(net2389));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][4]$_DFFE_PP__2390  (.L_HI(net2390));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][5]$_DFFE_PP__2391  (.L_HI(net2391));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][6]$_DFFE_PP__2392  (.L_HI(net2392));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][7]$_DFFE_PP__2393  (.L_HI(net2393));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][8]$_DFFE_PP__2394  (.L_HI(net2394));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[8][9]$_DFFE_PP__2395  (.L_HI(net2395));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][0]$_DFFE_PP__2396  (.L_HI(net2396));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][10]$_DFFE_PP__2397  (.L_HI(net2397));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][11]$_DFFE_PP__2398  (.L_HI(net2398));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][1]$_DFFE_PP__2399  (.L_HI(net2399));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][2]$_DFFE_PP__2400  (.L_HI(net2400));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][3]$_DFFE_PP__2401  (.L_HI(net2401));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][4]$_DFFE_PP__2402  (.L_HI(net2402));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][5]$_DFFE_PP__2403  (.L_HI(net2403));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][6]$_DFFE_PP__2404  (.L_HI(net2404));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][7]$_DFFE_PP__2405  (.L_HI(net2405));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][8]$_DFFE_PP__2406  (.L_HI(net2406));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_d[9][9]$_DFFE_PP__2407  (.L_HI(net2407));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][0]$_DFFE_PP__2408  (.L_HI(net2408));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][10]$_DFFE_PP__2409  (.L_HI(net2409));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][11]$_DFFE_PP__2410  (.L_HI(net2410));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][1]$_DFFE_PP__2411  (.L_HI(net2411));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][2]$_DFFE_PP__2412  (.L_HI(net2412));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][3]$_DFFE_PP__2413  (.L_HI(net2413));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][4]$_DFFE_PP__2414  (.L_HI(net2414));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][5]$_DFFE_PP__2415  (.L_HI(net2415));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][6]$_DFFE_PP__2416  (.L_HI(net2416));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][7]$_DFFE_PP__2417  (.L_HI(net2417));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][8]$_DFFE_PP__2418  (.L_HI(net2418));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[0][9]$_DFFE_PP__2419  (.L_HI(net2419));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][0]$_DFFE_PP__2420  (.L_HI(net2420));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][10]$_DFFE_PP__2421  (.L_HI(net2421));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][11]$_DFFE_PP__2422  (.L_HI(net2422));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][1]$_DFFE_PP__2423  (.L_HI(net2423));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][2]$_DFFE_PP__2424  (.L_HI(net2424));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][3]$_DFFE_PP__2425  (.L_HI(net2425));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][4]$_DFFE_PP__2426  (.L_HI(net2426));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][5]$_DFFE_PP__2427  (.L_HI(net2427));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][6]$_DFFE_PP__2428  (.L_HI(net2428));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][7]$_DFFE_PP__2429  (.L_HI(net2429));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][8]$_DFFE_PP__2430  (.L_HI(net2430));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[10][9]$_DFFE_PP__2431  (.L_HI(net2431));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][0]$_DFFE_PP__2432  (.L_HI(net2432));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][10]$_DFFE_PP__2433  (.L_HI(net2433));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][11]$_DFFE_PP__2434  (.L_HI(net2434));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][1]$_DFFE_PP__2435  (.L_HI(net2435));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][2]$_DFFE_PP__2436  (.L_HI(net2436));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][3]$_DFFE_PP__2437  (.L_HI(net2437));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][4]$_DFFE_PP__2438  (.L_HI(net2438));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][5]$_DFFE_PP__2439  (.L_HI(net2439));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][6]$_DFFE_PP__2440  (.L_HI(net2440));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][7]$_DFFE_PP__2441  (.L_HI(net2441));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][8]$_DFFE_PP__2442  (.L_HI(net2442));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[11][9]$_DFFE_PP__2443  (.L_HI(net2443));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][0]$_DFFE_PP__2444  (.L_HI(net2444));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][10]$_DFFE_PP__2445  (.L_HI(net2445));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][11]$_DFFE_PP__2446  (.L_HI(net2446));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][1]$_DFFE_PP__2447  (.L_HI(net2447));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][2]$_DFFE_PP__2448  (.L_HI(net2448));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][3]$_DFFE_PP__2449  (.L_HI(net2449));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][4]$_DFFE_PP__2450  (.L_HI(net2450));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][5]$_DFFE_PP__2451  (.L_HI(net2451));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][6]$_DFFE_PP__2452  (.L_HI(net2452));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][7]$_DFFE_PP__2453  (.L_HI(net2453));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][8]$_DFFE_PP__2454  (.L_HI(net2454));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[12][9]$_DFFE_PP__2455  (.L_HI(net2455));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][0]$_DFFE_PP__2456  (.L_HI(net2456));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][10]$_DFFE_PP__2457  (.L_HI(net2457));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][11]$_DFFE_PP__2458  (.L_HI(net2458));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][1]$_DFFE_PP__2459  (.L_HI(net2459));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][2]$_DFFE_PP__2460  (.L_HI(net2460));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][3]$_DFFE_PP__2461  (.L_HI(net2461));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][4]$_DFFE_PP__2462  (.L_HI(net2462));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][5]$_DFFE_PP__2463  (.L_HI(net2463));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][6]$_DFFE_PP__2464  (.L_HI(net2464));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][7]$_DFFE_PP__2465  (.L_HI(net2465));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][8]$_DFFE_PP__2466  (.L_HI(net2466));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[13][9]$_DFFE_PP__2467  (.L_HI(net2467));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][0]$_DFFE_PP__2468  (.L_HI(net2468));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][10]$_DFFE_PP__2469  (.L_HI(net2469));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][11]$_DFFE_PP__2470  (.L_HI(net2470));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][1]$_DFFE_PP__2471  (.L_HI(net2471));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][2]$_DFFE_PP__2472  (.L_HI(net2472));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][3]$_DFFE_PP__2473  (.L_HI(net2473));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][4]$_DFFE_PP__2474  (.L_HI(net2474));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][5]$_DFFE_PP__2475  (.L_HI(net2475));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][6]$_DFFE_PP__2476  (.L_HI(net2476));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][7]$_DFFE_PP__2477  (.L_HI(net2477));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][8]$_DFFE_PP__2478  (.L_HI(net2478));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[14][9]$_DFFE_PP__2479  (.L_HI(net2479));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][0]$_DFFE_PP__2480  (.L_HI(net2480));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][10]$_DFFE_PP__2481  (.L_HI(net2481));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][11]$_DFFE_PP__2482  (.L_HI(net2482));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][1]$_DFFE_PP__2483  (.L_HI(net2483));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][2]$_DFFE_PP__2484  (.L_HI(net2484));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][3]$_DFFE_PP__2485  (.L_HI(net2485));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][4]$_DFFE_PP__2486  (.L_HI(net2486));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][5]$_DFFE_PP__2487  (.L_HI(net2487));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][6]$_DFFE_PP__2488  (.L_HI(net2488));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][7]$_DFFE_PP__2489  (.L_HI(net2489));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][8]$_DFFE_PP__2490  (.L_HI(net2490));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[15][9]$_DFFE_PP__2491  (.L_HI(net2491));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][0]$_DFFE_PP__2492  (.L_HI(net2492));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][10]$_DFFE_PP__2493  (.L_HI(net2493));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][11]$_DFFE_PP__2494  (.L_HI(net2494));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][1]$_DFFE_PP__2495  (.L_HI(net2495));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][2]$_DFFE_PP__2496  (.L_HI(net2496));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][3]$_DFFE_PP__2497  (.L_HI(net2497));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][4]$_DFFE_PP__2498  (.L_HI(net2498));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][5]$_DFFE_PP__2499  (.L_HI(net2499));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][6]$_DFFE_PP__2500  (.L_HI(net2500));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][7]$_DFFE_PP__2501  (.L_HI(net2501));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][8]$_DFFE_PP__2502  (.L_HI(net2502));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[16][9]$_DFFE_PP__2503  (.L_HI(net2503));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][0]$_DFFE_PP__2504  (.L_HI(net2504));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][10]$_DFFE_PP__2505  (.L_HI(net2505));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][11]$_DFFE_PP__2506  (.L_HI(net2506));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][1]$_DFFE_PP__2507  (.L_HI(net2507));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][2]$_DFFE_PP__2508  (.L_HI(net2508));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][3]$_DFFE_PP__2509  (.L_HI(net2509));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][4]$_DFFE_PP__2510  (.L_HI(net2510));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][5]$_DFFE_PP__2511  (.L_HI(net2511));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][6]$_DFFE_PP__2512  (.L_HI(net2512));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][7]$_DFFE_PP__2513  (.L_HI(net2513));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][8]$_DFFE_PP__2514  (.L_HI(net2514));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[17][9]$_DFFE_PP__2515  (.L_HI(net2515));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][0]$_DFFE_PP__2516  (.L_HI(net2516));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][10]$_DFFE_PP__2517  (.L_HI(net2517));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][11]$_DFFE_PP__2518  (.L_HI(net2518));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][1]$_DFFE_PP__2519  (.L_HI(net2519));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][2]$_DFFE_PP__2520  (.L_HI(net2520));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][3]$_DFFE_PP__2521  (.L_HI(net2521));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][4]$_DFFE_PP__2522  (.L_HI(net2522));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][5]$_DFFE_PP__2523  (.L_HI(net2523));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][6]$_DFFE_PP__2524  (.L_HI(net2524));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][7]$_DFFE_PP__2525  (.L_HI(net2525));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][8]$_DFFE_PP__2526  (.L_HI(net2526));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[18][9]$_DFFE_PP__2527  (.L_HI(net2527));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][0]$_DFFE_PP__2528  (.L_HI(net2528));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][10]$_DFFE_PP__2529  (.L_HI(net2529));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][11]$_DFFE_PP__2530  (.L_HI(net2530));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][1]$_DFFE_PP__2531  (.L_HI(net2531));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][2]$_DFFE_PP__2532  (.L_HI(net2532));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][3]$_DFFE_PP__2533  (.L_HI(net2533));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][4]$_DFFE_PP__2534  (.L_HI(net2534));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][5]$_DFFE_PP__2535  (.L_HI(net2535));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][6]$_DFFE_PP__2536  (.L_HI(net2536));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][7]$_DFFE_PP__2537  (.L_HI(net2537));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][8]$_DFFE_PP__2538  (.L_HI(net2538));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[19][9]$_DFFE_PP__2539  (.L_HI(net2539));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][0]$_DFFE_PP__2540  (.L_HI(net2540));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][10]$_DFFE_PP__2541  (.L_HI(net2541));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][11]$_DFFE_PP__2542  (.L_HI(net2542));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][1]$_DFFE_PP__2543  (.L_HI(net2543));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][2]$_DFFE_PP__2544  (.L_HI(net2544));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][3]$_DFFE_PP__2545  (.L_HI(net2545));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][4]$_DFFE_PP__2546  (.L_HI(net2546));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][5]$_DFFE_PP__2547  (.L_HI(net2547));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][6]$_DFFE_PP__2548  (.L_HI(net2548));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][7]$_DFFE_PP__2549  (.L_HI(net2549));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][8]$_DFFE_PP__2550  (.L_HI(net2550));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[1][9]$_DFFE_PP__2551  (.L_HI(net2551));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][0]$_DFFE_PP__2552  (.L_HI(net2552));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][10]$_DFFE_PP__2553  (.L_HI(net2553));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][11]$_DFFE_PP__2554  (.L_HI(net2554));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][1]$_DFFE_PP__2555  (.L_HI(net2555));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][2]$_DFFE_PP__2556  (.L_HI(net2556));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][3]$_DFFE_PP__2557  (.L_HI(net2557));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][4]$_DFFE_PP__2558  (.L_HI(net2558));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][5]$_DFFE_PP__2559  (.L_HI(net2559));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][6]$_DFFE_PP__2560  (.L_HI(net2560));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][7]$_DFFE_PP__2561  (.L_HI(net2561));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][8]$_DFFE_PP__2562  (.L_HI(net2562));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[20][9]$_DFFE_PP__2563  (.L_HI(net2563));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][0]$_DFFE_PP__2564  (.L_HI(net2564));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][10]$_DFFE_PP__2565  (.L_HI(net2565));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][11]$_DFFE_PP__2566  (.L_HI(net2566));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][1]$_DFFE_PP__2567  (.L_HI(net2567));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][2]$_DFFE_PP__2568  (.L_HI(net2568));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][3]$_DFFE_PP__2569  (.L_HI(net2569));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][4]$_DFFE_PP__2570  (.L_HI(net2570));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][5]$_DFFE_PP__2571  (.L_HI(net2571));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][6]$_DFFE_PP__2572  (.L_HI(net2572));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][7]$_DFFE_PP__2573  (.L_HI(net2573));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][8]$_DFFE_PP__2574  (.L_HI(net2574));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[21][9]$_DFFE_PP__2575  (.L_HI(net2575));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][0]$_DFFE_PP__2576  (.L_HI(net2576));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][10]$_DFFE_PP__2577  (.L_HI(net2577));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][11]$_DFFE_PP__2578  (.L_HI(net2578));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][1]$_DFFE_PP__2579  (.L_HI(net2579));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][2]$_DFFE_PP__2580  (.L_HI(net2580));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][3]$_DFFE_PP__2581  (.L_HI(net2581));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][4]$_DFFE_PP__2582  (.L_HI(net2582));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][5]$_DFFE_PP__2583  (.L_HI(net2583));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][6]$_DFFE_PP__2584  (.L_HI(net2584));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][7]$_DFFE_PP__2585  (.L_HI(net2585));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][8]$_DFFE_PP__2586  (.L_HI(net2586));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[22][9]$_DFFE_PP__2587  (.L_HI(net2587));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][0]$_DFFE_PP__2588  (.L_HI(net2588));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][10]$_DFFE_PP__2589  (.L_HI(net2589));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][11]$_DFFE_PP__2590  (.L_HI(net2590));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][1]$_DFFE_PP__2591  (.L_HI(net2591));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][2]$_DFFE_PP__2592  (.L_HI(net2592));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][3]$_DFFE_PP__2593  (.L_HI(net2593));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][4]$_DFFE_PP__2594  (.L_HI(net2594));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][5]$_DFFE_PP__2595  (.L_HI(net2595));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][6]$_DFFE_PP__2596  (.L_HI(net2596));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][7]$_DFFE_PP__2597  (.L_HI(net2597));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][8]$_DFFE_PP__2598  (.L_HI(net2598));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[23][9]$_DFFE_PP__2599  (.L_HI(net2599));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][0]$_DFFE_PP__2600  (.L_HI(net2600));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][10]$_DFFE_PP__2601  (.L_HI(net2601));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][11]$_DFFE_PP__2602  (.L_HI(net2602));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][1]$_DFFE_PP__2603  (.L_HI(net2603));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][2]$_DFFE_PP__2604  (.L_HI(net2604));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][3]$_DFFE_PP__2605  (.L_HI(net2605));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][4]$_DFFE_PP__2606  (.L_HI(net2606));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][5]$_DFFE_PP__2607  (.L_HI(net2607));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][6]$_DFFE_PP__2608  (.L_HI(net2608));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][7]$_DFFE_PP__2609  (.L_HI(net2609));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][8]$_DFFE_PP__2610  (.L_HI(net2610));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[24][9]$_DFFE_PP__2611  (.L_HI(net2611));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][0]$_DFFE_PP__2612  (.L_HI(net2612));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][10]$_DFFE_PP__2613  (.L_HI(net2613));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][11]$_DFFE_PP__2614  (.L_HI(net2614));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][1]$_DFFE_PP__2615  (.L_HI(net2615));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][2]$_DFFE_PP__2616  (.L_HI(net2616));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][3]$_DFFE_PP__2617  (.L_HI(net2617));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][4]$_DFFE_PP__2618  (.L_HI(net2618));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][5]$_DFFE_PP__2619  (.L_HI(net2619));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][6]$_DFFE_PP__2620  (.L_HI(net2620));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][7]$_DFFE_PP__2621  (.L_HI(net2621));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][8]$_DFFE_PP__2622  (.L_HI(net2622));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[25][9]$_DFFE_PP__2623  (.L_HI(net2623));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][0]$_DFFE_PP__2624  (.L_HI(net2624));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][10]$_DFFE_PP__2625  (.L_HI(net2625));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][11]$_DFFE_PP__2626  (.L_HI(net2626));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][1]$_DFFE_PP__2627  (.L_HI(net2627));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][2]$_DFFE_PP__2628  (.L_HI(net2628));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][3]$_DFFE_PP__2629  (.L_HI(net2629));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][4]$_DFFE_PP__2630  (.L_HI(net2630));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][5]$_DFFE_PP__2631  (.L_HI(net2631));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][6]$_DFFE_PP__2632  (.L_HI(net2632));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][7]$_DFFE_PP__2633  (.L_HI(net2633));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][8]$_DFFE_PP__2634  (.L_HI(net2634));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[26][9]$_DFFE_PP__2635  (.L_HI(net2635));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][0]$_DFFE_PP__2636  (.L_HI(net2636));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][10]$_DFFE_PP__2637  (.L_HI(net2637));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][11]$_DFFE_PP__2638  (.L_HI(net2638));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][1]$_DFFE_PP__2639  (.L_HI(net2639));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][2]$_DFFE_PP__2640  (.L_HI(net2640));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][3]$_DFFE_PP__2641  (.L_HI(net2641));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][4]$_DFFE_PP__2642  (.L_HI(net2642));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][5]$_DFFE_PP__2643  (.L_HI(net2643));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][6]$_DFFE_PP__2644  (.L_HI(net2644));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][7]$_DFFE_PP__2645  (.L_HI(net2645));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][8]$_DFFE_PP__2646  (.L_HI(net2646));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[27][9]$_DFFE_PP__2647  (.L_HI(net2647));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][0]$_DFFE_PP__2648  (.L_HI(net2648));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][10]$_DFFE_PP__2649  (.L_HI(net2649));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][11]$_DFFE_PP__2650  (.L_HI(net2650));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][1]$_DFFE_PP__2651  (.L_HI(net2651));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][2]$_DFFE_PP__2652  (.L_HI(net2652));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][3]$_DFFE_PP__2653  (.L_HI(net2653));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][4]$_DFFE_PP__2654  (.L_HI(net2654));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][5]$_DFFE_PP__2655  (.L_HI(net2655));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][6]$_DFFE_PP__2656  (.L_HI(net2656));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][7]$_DFFE_PP__2657  (.L_HI(net2657));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][8]$_DFFE_PP__2658  (.L_HI(net2658));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[28][9]$_DFFE_PP__2659  (.L_HI(net2659));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][0]$_DFFE_PP__2660  (.L_HI(net2660));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][10]$_DFFE_PP__2661  (.L_HI(net2661));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][11]$_DFFE_PP__2662  (.L_HI(net2662));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][1]$_DFFE_PP__2663  (.L_HI(net2663));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][2]$_DFFE_PP__2664  (.L_HI(net2664));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][3]$_DFFE_PP__2665  (.L_HI(net2665));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][4]$_DFFE_PP__2666  (.L_HI(net2666));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][5]$_DFFE_PP__2667  (.L_HI(net2667));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][6]$_DFFE_PP__2668  (.L_HI(net2668));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][7]$_DFFE_PP__2669  (.L_HI(net2669));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][8]$_DFFE_PP__2670  (.L_HI(net2670));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[29][9]$_DFFE_PP__2671  (.L_HI(net2671));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][0]$_DFFE_PP__2672  (.L_HI(net2672));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][10]$_DFFE_PP__2673  (.L_HI(net2673));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][11]$_DFFE_PP__2674  (.L_HI(net2674));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][1]$_DFFE_PP__2675  (.L_HI(net2675));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][2]$_DFFE_PP__2676  (.L_HI(net2676));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][3]$_DFFE_PP__2677  (.L_HI(net2677));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][4]$_DFFE_PP__2678  (.L_HI(net2678));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][5]$_DFFE_PP__2679  (.L_HI(net2679));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][6]$_DFFE_PP__2680  (.L_HI(net2680));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][7]$_DFFE_PP__2681  (.L_HI(net2681));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][8]$_DFFE_PP__2682  (.L_HI(net2682));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[2][9]$_DFFE_PP__2683  (.L_HI(net2683));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][0]$_DFFE_PP__2684  (.L_HI(net2684));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][10]$_DFFE_PP__2685  (.L_HI(net2685));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][11]$_DFFE_PP__2686  (.L_HI(net2686));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][1]$_DFFE_PP__2687  (.L_HI(net2687));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][2]$_DFFE_PP__2688  (.L_HI(net2688));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][3]$_DFFE_PP__2689  (.L_HI(net2689));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][4]$_DFFE_PP__2690  (.L_HI(net2690));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][5]$_DFFE_PP__2691  (.L_HI(net2691));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][6]$_DFFE_PP__2692  (.L_HI(net2692));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][7]$_DFFE_PP__2693  (.L_HI(net2693));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][8]$_DFFE_PP__2694  (.L_HI(net2694));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[30][9]$_DFFE_PP__2695  (.L_HI(net2695));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][0]$_DFFE_PP__2696  (.L_HI(net2696));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][10]$_DFFE_PP__2697  (.L_HI(net2697));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][11]$_DFFE_PP__2698  (.L_HI(net2698));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][1]$_DFFE_PP__2699  (.L_HI(net2699));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][2]$_DFFE_PP__2700  (.L_HI(net2700));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][3]$_DFFE_PP__2701  (.L_HI(net2701));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][4]$_DFFE_PP__2702  (.L_HI(net2702));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][5]$_DFFE_PP__2703  (.L_HI(net2703));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][6]$_DFFE_PP__2704  (.L_HI(net2704));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][7]$_DFFE_PP__2705  (.L_HI(net2705));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][8]$_DFFE_PP__2706  (.L_HI(net2706));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[31][9]$_DFFE_PP__2707  (.L_HI(net2707));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][0]$_DFFE_PP__2708  (.L_HI(net2708));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][10]$_DFFE_PP__2709  (.L_HI(net2709));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][11]$_DFFE_PP__2710  (.L_HI(net2710));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][1]$_DFFE_PP__2711  (.L_HI(net2711));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][2]$_DFFE_PP__2712  (.L_HI(net2712));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][3]$_DFFE_PP__2713  (.L_HI(net2713));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][4]$_DFFE_PP__2714  (.L_HI(net2714));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][5]$_DFFE_PP__2715  (.L_HI(net2715));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][6]$_DFFE_PP__2716  (.L_HI(net2716));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][7]$_DFFE_PP__2717  (.L_HI(net2717));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][8]$_DFFE_PP__2718  (.L_HI(net2718));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[3][9]$_DFFE_PP__2719  (.L_HI(net2719));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][0]$_DFFE_PP__2720  (.L_HI(net2720));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][10]$_DFFE_PP__2721  (.L_HI(net2721));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][11]$_DFFE_PP__2722  (.L_HI(net2722));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][1]$_DFFE_PP__2723  (.L_HI(net2723));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][2]$_DFFE_PP__2724  (.L_HI(net2724));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][3]$_DFFE_PP__2725  (.L_HI(net2725));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][4]$_DFFE_PP__2726  (.L_HI(net2726));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][5]$_DFFE_PP__2727  (.L_HI(net2727));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][6]$_DFFE_PP__2728  (.L_HI(net2728));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][7]$_DFFE_PP__2729  (.L_HI(net2729));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][8]$_DFFE_PP__2730  (.L_HI(net2730));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[4][9]$_DFFE_PP__2731  (.L_HI(net2731));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][0]$_DFFE_PP__2732  (.L_HI(net2732));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][10]$_DFFE_PP__2733  (.L_HI(net2733));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][11]$_DFFE_PP__2734  (.L_HI(net2734));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][1]$_DFFE_PP__2735  (.L_HI(net2735));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][2]$_DFFE_PP__2736  (.L_HI(net2736));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][3]$_DFFE_PP__2737  (.L_HI(net2737));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][4]$_DFFE_PP__2738  (.L_HI(net2738));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][5]$_DFFE_PP__2739  (.L_HI(net2739));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][6]$_DFFE_PP__2740  (.L_HI(net2740));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][7]$_DFFE_PP__2741  (.L_HI(net2741));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][8]$_DFFE_PP__2742  (.L_HI(net2742));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[5][9]$_DFFE_PP__2743  (.L_HI(net2743));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][0]$_DFFE_PP__2744  (.L_HI(net2744));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][10]$_DFFE_PP__2745  (.L_HI(net2745));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][11]$_DFFE_PP__2746  (.L_HI(net2746));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][1]$_DFFE_PP__2747  (.L_HI(net2747));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][2]$_DFFE_PP__2748  (.L_HI(net2748));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][3]$_DFFE_PP__2749  (.L_HI(net2749));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][4]$_DFFE_PP__2750  (.L_HI(net2750));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][5]$_DFFE_PP__2751  (.L_HI(net2751));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][6]$_DFFE_PP__2752  (.L_HI(net2752));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][7]$_DFFE_PP__2753  (.L_HI(net2753));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][8]$_DFFE_PP__2754  (.L_HI(net2754));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[6][9]$_DFFE_PP__2755  (.L_HI(net2755));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][0]$_DFFE_PP__2756  (.L_HI(net2756));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][10]$_DFFE_PP__2757  (.L_HI(net2757));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][11]$_DFFE_PP__2758  (.L_HI(net2758));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][1]$_DFFE_PP__2759  (.L_HI(net2759));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][2]$_DFFE_PP__2760  (.L_HI(net2760));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][3]$_DFFE_PP__2761  (.L_HI(net2761));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][4]$_DFFE_PP__2762  (.L_HI(net2762));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][5]$_DFFE_PP__2763  (.L_HI(net2763));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][6]$_DFFE_PP__2764  (.L_HI(net2764));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][7]$_DFFE_PP__2765  (.L_HI(net2765));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][8]$_DFFE_PP__2766  (.L_HI(net2766));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[7][9]$_DFFE_PP__2767  (.L_HI(net2767));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][0]$_DFFE_PP__2768  (.L_HI(net2768));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][10]$_DFFE_PP__2769  (.L_HI(net2769));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][11]$_DFFE_PP__2770  (.L_HI(net2770));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][1]$_DFFE_PP__2771  (.L_HI(net2771));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][2]$_DFFE_PP__2772  (.L_HI(net2772));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][3]$_DFFE_PP__2773  (.L_HI(net2773));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][4]$_DFFE_PP__2774  (.L_HI(net2774));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][5]$_DFFE_PP__2775  (.L_HI(net2775));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][6]$_DFFE_PP__2776  (.L_HI(net2776));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][7]$_DFFE_PP__2777  (.L_HI(net2777));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][8]$_DFFE_PP__2778  (.L_HI(net2778));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[8][9]$_DFFE_PP__2779  (.L_HI(net2779));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][0]$_DFFE_PP__2780  (.L_HI(net2780));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][10]$_DFFE_PP__2781  (.L_HI(net2781));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][11]$_DFFE_PP__2782  (.L_HI(net2782));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][1]$_DFFE_PP__2783  (.L_HI(net2783));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][2]$_DFFE_PP__2784  (.L_HI(net2784));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][3]$_DFFE_PP__2785  (.L_HI(net2785));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][4]$_DFFE_PP__2786  (.L_HI(net2786));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][5]$_DFFE_PP__2787  (.L_HI(net2787));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][6]$_DFFE_PP__2788  (.L_HI(net2788));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][7]$_DFFE_PP__2789  (.L_HI(net2789));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][8]$_DFFE_PP__2790  (.L_HI(net2790));
 sg13g2_tiehi \cpu.genblk1.mmu.r_vtop_i[9][9]$_DFFE_PP__2791  (.L_HI(net2791));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[0]$_DFFE_PP__2792  (.L_HI(net2792));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[10]$_DFFE_PP__2793  (.L_HI(net2793));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[11]$_DFFE_PP__2794  (.L_HI(net2794));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[12]$_DFFE_PP__2795  (.L_HI(net2795));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[13]$_DFFE_PP__2796  (.L_HI(net2796));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[14]$_DFFE_PP__2797  (.L_HI(net2797));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[15]$_DFFE_PP__2798  (.L_HI(net2798));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[16]$_DFFE_PP__2799  (.L_HI(net2799));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[17]$_DFFE_PP__2800  (.L_HI(net2800));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[18]$_DFFE_PP__2801  (.L_HI(net2801));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[19]$_DFFE_PP__2802  (.L_HI(net2802));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[1]$_DFFE_PP__2803  (.L_HI(net2803));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[20]$_DFFE_PP__2804  (.L_HI(net2804));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[21]$_DFFE_PP__2805  (.L_HI(net2805));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[22]$_DFFE_PP__2806  (.L_HI(net2806));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[23]$_DFFE_PP__2807  (.L_HI(net2807));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[24]$_DFFE_PP__2808  (.L_HI(net2808));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[25]$_DFFE_PP__2809  (.L_HI(net2809));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[26]$_DFFE_PP__2810  (.L_HI(net2810));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[27]$_DFFE_PP__2811  (.L_HI(net2811));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[28]$_DFFE_PP__2812  (.L_HI(net2812));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[29]$_DFFE_PP__2813  (.L_HI(net2813));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[2]$_DFFE_PP__2814  (.L_HI(net2814));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[30]$_DFFE_PP__2815  (.L_HI(net2815));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[31]$_DFFE_PP__2816  (.L_HI(net2816));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[3]$_DFFE_PP__2817  (.L_HI(net2817));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[4]$_DFFE_PP__2818  (.L_HI(net2818));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[5]$_DFFE_PP__2819  (.L_HI(net2819));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[6]$_DFFE_PP__2820  (.L_HI(net2820));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[7]$_DFFE_PP__2821  (.L_HI(net2821));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[8]$_DFFE_PP__2822  (.L_HI(net2822));
 sg13g2_tiehi \cpu.genblk1.mmu.r_writeable_d[9]$_DFFE_PP__2823  (.L_HI(net2823));
 sg13g2_tiehi \cpu.gpio.r_enable_in[0]$_SDFFE_PN0P__2824  (.L_HI(net2824));
 sg13g2_tiehi \cpu.gpio.r_enable_in[1]$_SDFFE_PN0P__2825  (.L_HI(net2825));
 sg13g2_tiehi \cpu.gpio.r_enable_in[2]$_SDFFE_PN0P__2826  (.L_HI(net2826));
 sg13g2_tiehi \cpu.gpio.r_enable_in[3]$_SDFFE_PN0P__2827  (.L_HI(net2827));
 sg13g2_tiehi \cpu.gpio.r_enable_in[4]$_SDFFE_PN0P__2828  (.L_HI(net2828));
 sg13g2_tiehi \cpu.gpio.r_enable_in[5]$_SDFFE_PN0P__2829  (.L_HI(net2829));
 sg13g2_tiehi \cpu.gpio.r_enable_in[6]$_SDFFE_PN0P__2830  (.L_HI(net2830));
 sg13g2_tiehi \cpu.gpio.r_enable_in[7]$_SDFFE_PN0P__2831  (.L_HI(net2831));
 sg13g2_tiehi \cpu.gpio.r_enable_io[0]$_SDFFE_PN0P__2832  (.L_HI(net2832));
 sg13g2_tiehi \cpu.gpio.r_enable_io[1]$_SDFFE_PN0P__2833  (.L_HI(net2833));
 sg13g2_tiehi \cpu.gpio.r_enable_io[2]$_SDFFE_PN0P__2834  (.L_HI(net2834));
 sg13g2_tiehi \cpu.gpio.r_enable_io[3]$_SDFFE_PN0P__2835  (.L_HI(net2835));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[0]$_SDFFE_PN0P__2836  (.L_HI(net2836));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[1]$_SDFFE_PN0P__2837  (.L_HI(net2837));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[2]$_SDFFE_PN0P__2838  (.L_HI(net2838));
 sg13g2_tiehi \cpu.gpio.r_gpio_en[3]$_SDFFE_PN0P__2839  (.L_HI(net2839));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[0]$_DFFE_PP__2840  (.L_HI(net2840));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[1]$_DFFE_PP__2841  (.L_HI(net2841));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[2]$_DFFE_PP__2842  (.L_HI(net2842));
 sg13g2_tiehi \cpu.gpio.r_gpio_io[3]$_DFFE_PP__2843  (.L_HI(net2843));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[0]$_DFFE_PP__2844  (.L_HI(net2844));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[1]$_DFFE_PP__2845  (.L_HI(net2845));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[2]$_DFFE_PP__2846  (.L_HI(net2846));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[3]$_DFFE_PP__2847  (.L_HI(net2847));
 sg13g2_tiehi \cpu.gpio.r_gpio_o[4]$_DFFE_PP__2848  (.L_HI(net2848));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][0]$_DFFE_PP__2849  (.L_HI(net2849));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][1]$_DFFE_PP__2850  (.L_HI(net2850));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][2]$_DFFE_PP__2851  (.L_HI(net2851));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[0][3]$_DFFE_PP__2852  (.L_HI(net2852));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][0]$_DFFE_PP__2853  (.L_HI(net2853));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][1]$_DFFE_PP__2854  (.L_HI(net2854));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][2]$_DFFE_PP__2855  (.L_HI(net2855));
 sg13g2_tiehi \cpu.gpio.r_spi_miso_src[1][3]$_DFFE_PP__2856  (.L_HI(net2856));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][0]$_DFFE_PP__2857  (.L_HI(net2857));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][1]$_DFFE_PP__2858  (.L_HI(net2858));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][2]$_DFFE_PP__2859  (.L_HI(net2859));
 sg13g2_tiehi \cpu.gpio.r_src_io[4][3]$_DFFE_PP__2860  (.L_HI(net2860));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][0]$_DFFE_PP__2861  (.L_HI(net2861));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][1]$_DFFE_PP__2862  (.L_HI(net2862));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][2]$_DFFE_PP__2863  (.L_HI(net2863));
 sg13g2_tiehi \cpu.gpio.r_src_io[5][3]$_DFFE_PP__2864  (.L_HI(net2864));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][0]$_DFFE_PP__2865  (.L_HI(net2865));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][1]$_DFFE_PP__2866  (.L_HI(net2866));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][2]$_DFFE_PP__2867  (.L_HI(net2867));
 sg13g2_tiehi \cpu.gpio.r_src_io[6][3]$_DFFE_PP__2868  (.L_HI(net2868));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][0]$_DFFE_PP__2869  (.L_HI(net2869));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][1]$_DFFE_PP__2870  (.L_HI(net2870));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][2]$_DFFE_PP__2871  (.L_HI(net2871));
 sg13g2_tiehi \cpu.gpio.r_src_io[7][3]$_DFFE_PP__2872  (.L_HI(net2872));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][0]$_DFFE_PP__2873  (.L_HI(net2873));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][1]$_DFFE_PP__2874  (.L_HI(net2874));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][2]$_DFFE_PP__2875  (.L_HI(net2875));
 sg13g2_tiehi \cpu.gpio.r_src_o[3][3]$_DFFE_PP__2876  (.L_HI(net2876));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][0]$_DFFE_PP__2877  (.L_HI(net2877));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][1]$_DFFE_PP__2878  (.L_HI(net2878));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][2]$_DFFE_PP__2879  (.L_HI(net2879));
 sg13g2_tiehi \cpu.gpio.r_src_o[4][3]$_DFFE_PP__2880  (.L_HI(net2880));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][0]$_DFFE_PP__2881  (.L_HI(net2881));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][1]$_DFFE_PP__2882  (.L_HI(net2882));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][2]$_DFFE_PP__2883  (.L_HI(net2883));
 sg13g2_tiehi \cpu.gpio.r_src_o[5][3]$_DFFE_PP__2884  (.L_HI(net2884));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][0]$_SDFFE_PN1P__2885  (.L_HI(net2885));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][1]$_SDFFE_PN0P__2886  (.L_HI(net2886));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][2]$_SDFFE_PN0P__2887  (.L_HI(net2887));
 sg13g2_tiehi \cpu.gpio.r_src_o[6][3]$_SDFFE_PN0P__2888  (.L_HI(net2888));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][0]$_DFFE_PP__2889  (.L_HI(net2889));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][1]$_DFFE_PP__2890  (.L_HI(net2890));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][2]$_DFFE_PP__2891  (.L_HI(net2891));
 sg13g2_tiehi \cpu.gpio.r_src_o[7][3]$_DFFE_PP__2892  (.L_HI(net2892));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[0]$_SDFFE_PN0P__2893  (.L_HI(net2893));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[1]$_SDFFE_PN0P__2894  (.L_HI(net2894));
 sg13g2_tiehi \cpu.gpio.r_uart_rx_src[2]$_SDFFE_PN0P__2895  (.L_HI(net2895));
 sg13g2_tiehi \cpu.icache.r_data[0][0]$_DFFE_PP__2896  (.L_HI(net2896));
 sg13g2_tiehi \cpu.icache.r_data[0][10]$_DFFE_PP__2897  (.L_HI(net2897));
 sg13g2_tiehi \cpu.icache.r_data[0][11]$_DFFE_PP__2898  (.L_HI(net2898));
 sg13g2_tiehi \cpu.icache.r_data[0][12]$_DFFE_PP__2899  (.L_HI(net2899));
 sg13g2_tiehi \cpu.icache.r_data[0][13]$_DFFE_PP__2900  (.L_HI(net2900));
 sg13g2_tiehi \cpu.icache.r_data[0][14]$_DFFE_PP__2901  (.L_HI(net2901));
 sg13g2_tiehi \cpu.icache.r_data[0][15]$_DFFE_PP__2902  (.L_HI(net2902));
 sg13g2_tiehi \cpu.icache.r_data[0][16]$_DFFE_PP__2903  (.L_HI(net2903));
 sg13g2_tiehi \cpu.icache.r_data[0][17]$_DFFE_PP__2904  (.L_HI(net2904));
 sg13g2_tiehi \cpu.icache.r_data[0][18]$_DFFE_PP__2905  (.L_HI(net2905));
 sg13g2_tiehi \cpu.icache.r_data[0][19]$_DFFE_PP__2906  (.L_HI(net2906));
 sg13g2_tiehi \cpu.icache.r_data[0][1]$_DFFE_PP__2907  (.L_HI(net2907));
 sg13g2_tiehi \cpu.icache.r_data[0][20]$_DFFE_PP__2908  (.L_HI(net2908));
 sg13g2_tiehi \cpu.icache.r_data[0][21]$_DFFE_PP__2909  (.L_HI(net2909));
 sg13g2_tiehi \cpu.icache.r_data[0][22]$_DFFE_PP__2910  (.L_HI(net2910));
 sg13g2_tiehi \cpu.icache.r_data[0][23]$_DFFE_PP__2911  (.L_HI(net2911));
 sg13g2_tiehi \cpu.icache.r_data[0][24]$_DFFE_PP__2912  (.L_HI(net2912));
 sg13g2_tiehi \cpu.icache.r_data[0][25]$_DFFE_PP__2913  (.L_HI(net2913));
 sg13g2_tiehi \cpu.icache.r_data[0][26]$_DFFE_PP__2914  (.L_HI(net2914));
 sg13g2_tiehi \cpu.icache.r_data[0][27]$_DFFE_PP__2915  (.L_HI(net2915));
 sg13g2_tiehi \cpu.icache.r_data[0][28]$_DFFE_PP__2916  (.L_HI(net2916));
 sg13g2_tiehi \cpu.icache.r_data[0][29]$_DFFE_PP__2917  (.L_HI(net2917));
 sg13g2_tiehi \cpu.icache.r_data[0][2]$_DFFE_PP__2918  (.L_HI(net2918));
 sg13g2_tiehi \cpu.icache.r_data[0][30]$_DFFE_PP__2919  (.L_HI(net2919));
 sg13g2_tiehi \cpu.icache.r_data[0][31]$_DFFE_PP__2920  (.L_HI(net2920));
 sg13g2_tiehi \cpu.icache.r_data[0][3]$_DFFE_PP__2921  (.L_HI(net2921));
 sg13g2_tiehi \cpu.icache.r_data[0][4]$_DFFE_PP__2922  (.L_HI(net2922));
 sg13g2_tiehi \cpu.icache.r_data[0][5]$_DFFE_PP__2923  (.L_HI(net2923));
 sg13g2_tiehi \cpu.icache.r_data[0][6]$_DFFE_PP__2924  (.L_HI(net2924));
 sg13g2_tiehi \cpu.icache.r_data[0][7]$_DFFE_PP__2925  (.L_HI(net2925));
 sg13g2_tiehi \cpu.icache.r_data[0][8]$_DFFE_PP__2926  (.L_HI(net2926));
 sg13g2_tiehi \cpu.icache.r_data[0][9]$_DFFE_PP__2927  (.L_HI(net2927));
 sg13g2_tiehi \cpu.icache.r_data[1][0]$_DFFE_PP__2928  (.L_HI(net2928));
 sg13g2_tiehi \cpu.icache.r_data[1][10]$_DFFE_PP__2929  (.L_HI(net2929));
 sg13g2_tiehi \cpu.icache.r_data[1][11]$_DFFE_PP__2930  (.L_HI(net2930));
 sg13g2_tiehi \cpu.icache.r_data[1][12]$_DFFE_PP__2931  (.L_HI(net2931));
 sg13g2_tiehi \cpu.icache.r_data[1][13]$_DFFE_PP__2932  (.L_HI(net2932));
 sg13g2_tiehi \cpu.icache.r_data[1][14]$_DFFE_PP__2933  (.L_HI(net2933));
 sg13g2_tiehi \cpu.icache.r_data[1][15]$_DFFE_PP__2934  (.L_HI(net2934));
 sg13g2_tiehi \cpu.icache.r_data[1][16]$_DFFE_PP__2935  (.L_HI(net2935));
 sg13g2_tiehi \cpu.icache.r_data[1][17]$_DFFE_PP__2936  (.L_HI(net2936));
 sg13g2_tiehi \cpu.icache.r_data[1][18]$_DFFE_PP__2937  (.L_HI(net2937));
 sg13g2_tiehi \cpu.icache.r_data[1][19]$_DFFE_PP__2938  (.L_HI(net2938));
 sg13g2_tiehi \cpu.icache.r_data[1][1]$_DFFE_PP__2939  (.L_HI(net2939));
 sg13g2_tiehi \cpu.icache.r_data[1][20]$_DFFE_PP__2940  (.L_HI(net2940));
 sg13g2_tiehi \cpu.icache.r_data[1][21]$_DFFE_PP__2941  (.L_HI(net2941));
 sg13g2_tiehi \cpu.icache.r_data[1][22]$_DFFE_PP__2942  (.L_HI(net2942));
 sg13g2_tiehi \cpu.icache.r_data[1][23]$_DFFE_PP__2943  (.L_HI(net2943));
 sg13g2_tiehi \cpu.icache.r_data[1][24]$_DFFE_PP__2944  (.L_HI(net2944));
 sg13g2_tiehi \cpu.icache.r_data[1][25]$_DFFE_PP__2945  (.L_HI(net2945));
 sg13g2_tiehi \cpu.icache.r_data[1][26]$_DFFE_PP__2946  (.L_HI(net2946));
 sg13g2_tiehi \cpu.icache.r_data[1][27]$_DFFE_PP__2947  (.L_HI(net2947));
 sg13g2_tiehi \cpu.icache.r_data[1][28]$_DFFE_PP__2948  (.L_HI(net2948));
 sg13g2_tiehi \cpu.icache.r_data[1][29]$_DFFE_PP__2949  (.L_HI(net2949));
 sg13g2_tiehi \cpu.icache.r_data[1][2]$_DFFE_PP__2950  (.L_HI(net2950));
 sg13g2_tiehi \cpu.icache.r_data[1][30]$_DFFE_PP__2951  (.L_HI(net2951));
 sg13g2_tiehi \cpu.icache.r_data[1][31]$_DFFE_PP__2952  (.L_HI(net2952));
 sg13g2_tiehi \cpu.icache.r_data[1][3]$_DFFE_PP__2953  (.L_HI(net2953));
 sg13g2_tiehi \cpu.icache.r_data[1][4]$_DFFE_PP__2954  (.L_HI(net2954));
 sg13g2_tiehi \cpu.icache.r_data[1][5]$_DFFE_PP__2955  (.L_HI(net2955));
 sg13g2_tiehi \cpu.icache.r_data[1][6]$_DFFE_PP__2956  (.L_HI(net2956));
 sg13g2_tiehi \cpu.icache.r_data[1][7]$_DFFE_PP__2957  (.L_HI(net2957));
 sg13g2_tiehi \cpu.icache.r_data[1][8]$_DFFE_PP__2958  (.L_HI(net2958));
 sg13g2_tiehi \cpu.icache.r_data[1][9]$_DFFE_PP__2959  (.L_HI(net2959));
 sg13g2_tiehi \cpu.icache.r_data[2][0]$_DFFE_PP__2960  (.L_HI(net2960));
 sg13g2_tiehi \cpu.icache.r_data[2][10]$_DFFE_PP__2961  (.L_HI(net2961));
 sg13g2_tiehi \cpu.icache.r_data[2][11]$_DFFE_PP__2962  (.L_HI(net2962));
 sg13g2_tiehi \cpu.icache.r_data[2][12]$_DFFE_PP__2963  (.L_HI(net2963));
 sg13g2_tiehi \cpu.icache.r_data[2][13]$_DFFE_PP__2964  (.L_HI(net2964));
 sg13g2_tiehi \cpu.icache.r_data[2][14]$_DFFE_PP__2965  (.L_HI(net2965));
 sg13g2_tiehi \cpu.icache.r_data[2][15]$_DFFE_PP__2966  (.L_HI(net2966));
 sg13g2_tiehi \cpu.icache.r_data[2][16]$_DFFE_PP__2967  (.L_HI(net2967));
 sg13g2_tiehi \cpu.icache.r_data[2][17]$_DFFE_PP__2968  (.L_HI(net2968));
 sg13g2_tiehi \cpu.icache.r_data[2][18]$_DFFE_PP__2969  (.L_HI(net2969));
 sg13g2_tiehi \cpu.icache.r_data[2][19]$_DFFE_PP__2970  (.L_HI(net2970));
 sg13g2_tiehi \cpu.icache.r_data[2][1]$_DFFE_PP__2971  (.L_HI(net2971));
 sg13g2_tiehi \cpu.icache.r_data[2][20]$_DFFE_PP__2972  (.L_HI(net2972));
 sg13g2_tiehi \cpu.icache.r_data[2][21]$_DFFE_PP__2973  (.L_HI(net2973));
 sg13g2_tiehi \cpu.icache.r_data[2][22]$_DFFE_PP__2974  (.L_HI(net2974));
 sg13g2_tiehi \cpu.icache.r_data[2][23]$_DFFE_PP__2975  (.L_HI(net2975));
 sg13g2_tiehi \cpu.icache.r_data[2][24]$_DFFE_PP__2976  (.L_HI(net2976));
 sg13g2_tiehi \cpu.icache.r_data[2][25]$_DFFE_PP__2977  (.L_HI(net2977));
 sg13g2_tiehi \cpu.icache.r_data[2][26]$_DFFE_PP__2978  (.L_HI(net2978));
 sg13g2_tiehi \cpu.icache.r_data[2][27]$_DFFE_PP__2979  (.L_HI(net2979));
 sg13g2_tiehi \cpu.icache.r_data[2][28]$_DFFE_PP__2980  (.L_HI(net2980));
 sg13g2_tiehi \cpu.icache.r_data[2][29]$_DFFE_PP__2981  (.L_HI(net2981));
 sg13g2_tiehi \cpu.icache.r_data[2][2]$_DFFE_PP__2982  (.L_HI(net2982));
 sg13g2_tiehi \cpu.icache.r_data[2][30]$_DFFE_PP__2983  (.L_HI(net2983));
 sg13g2_tiehi \cpu.icache.r_data[2][31]$_DFFE_PP__2984  (.L_HI(net2984));
 sg13g2_tiehi \cpu.icache.r_data[2][3]$_DFFE_PP__2985  (.L_HI(net2985));
 sg13g2_tiehi \cpu.icache.r_data[2][4]$_DFFE_PP__2986  (.L_HI(net2986));
 sg13g2_tiehi \cpu.icache.r_data[2][5]$_DFFE_PP__2987  (.L_HI(net2987));
 sg13g2_tiehi \cpu.icache.r_data[2][6]$_DFFE_PP__2988  (.L_HI(net2988));
 sg13g2_tiehi \cpu.icache.r_data[2][7]$_DFFE_PP__2989  (.L_HI(net2989));
 sg13g2_tiehi \cpu.icache.r_data[2][8]$_DFFE_PP__2990  (.L_HI(net2990));
 sg13g2_tiehi \cpu.icache.r_data[2][9]$_DFFE_PP__2991  (.L_HI(net2991));
 sg13g2_tiehi \cpu.icache.r_data[3][0]$_DFFE_PP__2992  (.L_HI(net2992));
 sg13g2_tiehi \cpu.icache.r_data[3][10]$_DFFE_PP__2993  (.L_HI(net2993));
 sg13g2_tiehi \cpu.icache.r_data[3][11]$_DFFE_PP__2994  (.L_HI(net2994));
 sg13g2_tiehi \cpu.icache.r_data[3][12]$_DFFE_PP__2995  (.L_HI(net2995));
 sg13g2_tiehi \cpu.icache.r_data[3][13]$_DFFE_PP__2996  (.L_HI(net2996));
 sg13g2_tiehi \cpu.icache.r_data[3][14]$_DFFE_PP__2997  (.L_HI(net2997));
 sg13g2_tiehi \cpu.icache.r_data[3][15]$_DFFE_PP__2998  (.L_HI(net2998));
 sg13g2_tiehi \cpu.icache.r_data[3][16]$_DFFE_PP__2999  (.L_HI(net2999));
 sg13g2_tiehi \cpu.icache.r_data[3][17]$_DFFE_PP__3000  (.L_HI(net3000));
 sg13g2_tiehi \cpu.icache.r_data[3][18]$_DFFE_PP__3001  (.L_HI(net3001));
 sg13g2_tiehi \cpu.icache.r_data[3][19]$_DFFE_PP__3002  (.L_HI(net3002));
 sg13g2_tiehi \cpu.icache.r_data[3][1]$_DFFE_PP__3003  (.L_HI(net3003));
 sg13g2_tiehi \cpu.icache.r_data[3][20]$_DFFE_PP__3004  (.L_HI(net3004));
 sg13g2_tiehi \cpu.icache.r_data[3][21]$_DFFE_PP__3005  (.L_HI(net3005));
 sg13g2_tiehi \cpu.icache.r_data[3][22]$_DFFE_PP__3006  (.L_HI(net3006));
 sg13g2_tiehi \cpu.icache.r_data[3][23]$_DFFE_PP__3007  (.L_HI(net3007));
 sg13g2_tiehi \cpu.icache.r_data[3][24]$_DFFE_PP__3008  (.L_HI(net3008));
 sg13g2_tiehi \cpu.icache.r_data[3][25]$_DFFE_PP__3009  (.L_HI(net3009));
 sg13g2_tiehi \cpu.icache.r_data[3][26]$_DFFE_PP__3010  (.L_HI(net3010));
 sg13g2_tiehi \cpu.icache.r_data[3][27]$_DFFE_PP__3011  (.L_HI(net3011));
 sg13g2_tiehi \cpu.icache.r_data[3][28]$_DFFE_PP__3012  (.L_HI(net3012));
 sg13g2_tiehi \cpu.icache.r_data[3][29]$_DFFE_PP__3013  (.L_HI(net3013));
 sg13g2_tiehi \cpu.icache.r_data[3][2]$_DFFE_PP__3014  (.L_HI(net3014));
 sg13g2_tiehi \cpu.icache.r_data[3][30]$_DFFE_PP__3015  (.L_HI(net3015));
 sg13g2_tiehi \cpu.icache.r_data[3][31]$_DFFE_PP__3016  (.L_HI(net3016));
 sg13g2_tiehi \cpu.icache.r_data[3][3]$_DFFE_PP__3017  (.L_HI(net3017));
 sg13g2_tiehi \cpu.icache.r_data[3][4]$_DFFE_PP__3018  (.L_HI(net3018));
 sg13g2_tiehi \cpu.icache.r_data[3][5]$_DFFE_PP__3019  (.L_HI(net3019));
 sg13g2_tiehi \cpu.icache.r_data[3][6]$_DFFE_PP__3020  (.L_HI(net3020));
 sg13g2_tiehi \cpu.icache.r_data[3][7]$_DFFE_PP__3021  (.L_HI(net3021));
 sg13g2_tiehi \cpu.icache.r_data[3][8]$_DFFE_PP__3022  (.L_HI(net3022));
 sg13g2_tiehi \cpu.icache.r_data[3][9]$_DFFE_PP__3023  (.L_HI(net3023));
 sg13g2_tiehi \cpu.icache.r_data[4][0]$_DFFE_PP__3024  (.L_HI(net3024));
 sg13g2_tiehi \cpu.icache.r_data[4][10]$_DFFE_PP__3025  (.L_HI(net3025));
 sg13g2_tiehi \cpu.icache.r_data[4][11]$_DFFE_PP__3026  (.L_HI(net3026));
 sg13g2_tiehi \cpu.icache.r_data[4][12]$_DFFE_PP__3027  (.L_HI(net3027));
 sg13g2_tiehi \cpu.icache.r_data[4][13]$_DFFE_PP__3028  (.L_HI(net3028));
 sg13g2_tiehi \cpu.icache.r_data[4][14]$_DFFE_PP__3029  (.L_HI(net3029));
 sg13g2_tiehi \cpu.icache.r_data[4][15]$_DFFE_PP__3030  (.L_HI(net3030));
 sg13g2_tiehi \cpu.icache.r_data[4][16]$_DFFE_PP__3031  (.L_HI(net3031));
 sg13g2_tiehi \cpu.icache.r_data[4][17]$_DFFE_PP__3032  (.L_HI(net3032));
 sg13g2_tiehi \cpu.icache.r_data[4][18]$_DFFE_PP__3033  (.L_HI(net3033));
 sg13g2_tiehi \cpu.icache.r_data[4][19]$_DFFE_PP__3034  (.L_HI(net3034));
 sg13g2_tiehi \cpu.icache.r_data[4][1]$_DFFE_PP__3035  (.L_HI(net3035));
 sg13g2_tiehi \cpu.icache.r_data[4][20]$_DFFE_PP__3036  (.L_HI(net3036));
 sg13g2_tiehi \cpu.icache.r_data[4][21]$_DFFE_PP__3037  (.L_HI(net3037));
 sg13g2_tiehi \cpu.icache.r_data[4][22]$_DFFE_PP__3038  (.L_HI(net3038));
 sg13g2_tiehi \cpu.icache.r_data[4][23]$_DFFE_PP__3039  (.L_HI(net3039));
 sg13g2_tiehi \cpu.icache.r_data[4][24]$_DFFE_PP__3040  (.L_HI(net3040));
 sg13g2_tiehi \cpu.icache.r_data[4][25]$_DFFE_PP__3041  (.L_HI(net3041));
 sg13g2_tiehi \cpu.icache.r_data[4][26]$_DFFE_PP__3042  (.L_HI(net3042));
 sg13g2_tiehi \cpu.icache.r_data[4][27]$_DFFE_PP__3043  (.L_HI(net3043));
 sg13g2_tiehi \cpu.icache.r_data[4][28]$_DFFE_PP__3044  (.L_HI(net3044));
 sg13g2_tiehi \cpu.icache.r_data[4][29]$_DFFE_PP__3045  (.L_HI(net3045));
 sg13g2_tiehi \cpu.icache.r_data[4][2]$_DFFE_PP__3046  (.L_HI(net3046));
 sg13g2_tiehi \cpu.icache.r_data[4][30]$_DFFE_PP__3047  (.L_HI(net3047));
 sg13g2_tiehi \cpu.icache.r_data[4][31]$_DFFE_PP__3048  (.L_HI(net3048));
 sg13g2_tiehi \cpu.icache.r_data[4][3]$_DFFE_PP__3049  (.L_HI(net3049));
 sg13g2_tiehi \cpu.icache.r_data[4][4]$_DFFE_PP__3050  (.L_HI(net3050));
 sg13g2_tiehi \cpu.icache.r_data[4][5]$_DFFE_PP__3051  (.L_HI(net3051));
 sg13g2_tiehi \cpu.icache.r_data[4][6]$_DFFE_PP__3052  (.L_HI(net3052));
 sg13g2_tiehi \cpu.icache.r_data[4][7]$_DFFE_PP__3053  (.L_HI(net3053));
 sg13g2_tiehi \cpu.icache.r_data[4][8]$_DFFE_PP__3054  (.L_HI(net3054));
 sg13g2_tiehi \cpu.icache.r_data[4][9]$_DFFE_PP__3055  (.L_HI(net3055));
 sg13g2_tiehi \cpu.icache.r_data[5][0]$_DFFE_PP__3056  (.L_HI(net3056));
 sg13g2_tiehi \cpu.icache.r_data[5][10]$_DFFE_PP__3057  (.L_HI(net3057));
 sg13g2_tiehi \cpu.icache.r_data[5][11]$_DFFE_PP__3058  (.L_HI(net3058));
 sg13g2_tiehi \cpu.icache.r_data[5][12]$_DFFE_PP__3059  (.L_HI(net3059));
 sg13g2_tiehi \cpu.icache.r_data[5][13]$_DFFE_PP__3060  (.L_HI(net3060));
 sg13g2_tiehi \cpu.icache.r_data[5][14]$_DFFE_PP__3061  (.L_HI(net3061));
 sg13g2_tiehi \cpu.icache.r_data[5][15]$_DFFE_PP__3062  (.L_HI(net3062));
 sg13g2_tiehi \cpu.icache.r_data[5][16]$_DFFE_PP__3063  (.L_HI(net3063));
 sg13g2_tiehi \cpu.icache.r_data[5][17]$_DFFE_PP__3064  (.L_HI(net3064));
 sg13g2_tiehi \cpu.icache.r_data[5][18]$_DFFE_PP__3065  (.L_HI(net3065));
 sg13g2_tiehi \cpu.icache.r_data[5][19]$_DFFE_PP__3066  (.L_HI(net3066));
 sg13g2_tiehi \cpu.icache.r_data[5][1]$_DFFE_PP__3067  (.L_HI(net3067));
 sg13g2_tiehi \cpu.icache.r_data[5][20]$_DFFE_PP__3068  (.L_HI(net3068));
 sg13g2_tiehi \cpu.icache.r_data[5][21]$_DFFE_PP__3069  (.L_HI(net3069));
 sg13g2_tiehi \cpu.icache.r_data[5][22]$_DFFE_PP__3070  (.L_HI(net3070));
 sg13g2_tiehi \cpu.icache.r_data[5][23]$_DFFE_PP__3071  (.L_HI(net3071));
 sg13g2_tiehi \cpu.icache.r_data[5][24]$_DFFE_PP__3072  (.L_HI(net3072));
 sg13g2_tiehi \cpu.icache.r_data[5][25]$_DFFE_PP__3073  (.L_HI(net3073));
 sg13g2_tiehi \cpu.icache.r_data[5][26]$_DFFE_PP__3074  (.L_HI(net3074));
 sg13g2_tiehi \cpu.icache.r_data[5][27]$_DFFE_PP__3075  (.L_HI(net3075));
 sg13g2_tiehi \cpu.icache.r_data[5][28]$_DFFE_PP__3076  (.L_HI(net3076));
 sg13g2_tiehi \cpu.icache.r_data[5][29]$_DFFE_PP__3077  (.L_HI(net3077));
 sg13g2_tiehi \cpu.icache.r_data[5][2]$_DFFE_PP__3078  (.L_HI(net3078));
 sg13g2_tiehi \cpu.icache.r_data[5][30]$_DFFE_PP__3079  (.L_HI(net3079));
 sg13g2_tiehi \cpu.icache.r_data[5][31]$_DFFE_PP__3080  (.L_HI(net3080));
 sg13g2_tiehi \cpu.icache.r_data[5][3]$_DFFE_PP__3081  (.L_HI(net3081));
 sg13g2_tiehi \cpu.icache.r_data[5][4]$_DFFE_PP__3082  (.L_HI(net3082));
 sg13g2_tiehi \cpu.icache.r_data[5][5]$_DFFE_PP__3083  (.L_HI(net3083));
 sg13g2_tiehi \cpu.icache.r_data[5][6]$_DFFE_PP__3084  (.L_HI(net3084));
 sg13g2_tiehi \cpu.icache.r_data[5][7]$_DFFE_PP__3085  (.L_HI(net3085));
 sg13g2_tiehi \cpu.icache.r_data[5][8]$_DFFE_PP__3086  (.L_HI(net3086));
 sg13g2_tiehi \cpu.icache.r_data[5][9]$_DFFE_PP__3087  (.L_HI(net3087));
 sg13g2_tiehi \cpu.icache.r_data[6][0]$_DFFE_PP__3088  (.L_HI(net3088));
 sg13g2_tiehi \cpu.icache.r_data[6][10]$_DFFE_PP__3089  (.L_HI(net3089));
 sg13g2_tiehi \cpu.icache.r_data[6][11]$_DFFE_PP__3090  (.L_HI(net3090));
 sg13g2_tiehi \cpu.icache.r_data[6][12]$_DFFE_PP__3091  (.L_HI(net3091));
 sg13g2_tiehi \cpu.icache.r_data[6][13]$_DFFE_PP__3092  (.L_HI(net3092));
 sg13g2_tiehi \cpu.icache.r_data[6][14]$_DFFE_PP__3093  (.L_HI(net3093));
 sg13g2_tiehi \cpu.icache.r_data[6][15]$_DFFE_PP__3094  (.L_HI(net3094));
 sg13g2_tiehi \cpu.icache.r_data[6][16]$_DFFE_PP__3095  (.L_HI(net3095));
 sg13g2_tiehi \cpu.icache.r_data[6][17]$_DFFE_PP__3096  (.L_HI(net3096));
 sg13g2_tiehi \cpu.icache.r_data[6][18]$_DFFE_PP__3097  (.L_HI(net3097));
 sg13g2_tiehi \cpu.icache.r_data[6][19]$_DFFE_PP__3098  (.L_HI(net3098));
 sg13g2_tiehi \cpu.icache.r_data[6][1]$_DFFE_PP__3099  (.L_HI(net3099));
 sg13g2_tiehi \cpu.icache.r_data[6][20]$_DFFE_PP__3100  (.L_HI(net3100));
 sg13g2_tiehi \cpu.icache.r_data[6][21]$_DFFE_PP__3101  (.L_HI(net3101));
 sg13g2_tiehi \cpu.icache.r_data[6][22]$_DFFE_PP__3102  (.L_HI(net3102));
 sg13g2_tiehi \cpu.icache.r_data[6][23]$_DFFE_PP__3103  (.L_HI(net3103));
 sg13g2_tiehi \cpu.icache.r_data[6][24]$_DFFE_PP__3104  (.L_HI(net3104));
 sg13g2_tiehi \cpu.icache.r_data[6][25]$_DFFE_PP__3105  (.L_HI(net3105));
 sg13g2_tiehi \cpu.icache.r_data[6][26]$_DFFE_PP__3106  (.L_HI(net3106));
 sg13g2_tiehi \cpu.icache.r_data[6][27]$_DFFE_PP__3107  (.L_HI(net3107));
 sg13g2_tiehi \cpu.icache.r_data[6][28]$_DFFE_PP__3108  (.L_HI(net3108));
 sg13g2_tiehi \cpu.icache.r_data[6][29]$_DFFE_PP__3109  (.L_HI(net3109));
 sg13g2_tiehi \cpu.icache.r_data[6][2]$_DFFE_PP__3110  (.L_HI(net3110));
 sg13g2_tiehi \cpu.icache.r_data[6][30]$_DFFE_PP__3111  (.L_HI(net3111));
 sg13g2_tiehi \cpu.icache.r_data[6][31]$_DFFE_PP__3112  (.L_HI(net3112));
 sg13g2_tiehi \cpu.icache.r_data[6][3]$_DFFE_PP__3113  (.L_HI(net3113));
 sg13g2_tiehi \cpu.icache.r_data[6][4]$_DFFE_PP__3114  (.L_HI(net3114));
 sg13g2_tiehi \cpu.icache.r_data[6][5]$_DFFE_PP__3115  (.L_HI(net3115));
 sg13g2_tiehi \cpu.icache.r_data[6][6]$_DFFE_PP__3116  (.L_HI(net3116));
 sg13g2_tiehi \cpu.icache.r_data[6][7]$_DFFE_PP__3117  (.L_HI(net3117));
 sg13g2_tiehi \cpu.icache.r_data[6][8]$_DFFE_PP__3118  (.L_HI(net3118));
 sg13g2_tiehi \cpu.icache.r_data[6][9]$_DFFE_PP__3119  (.L_HI(net3119));
 sg13g2_tiehi \cpu.icache.r_data[7][0]$_DFFE_PP__3120  (.L_HI(net3120));
 sg13g2_tiehi \cpu.icache.r_data[7][10]$_DFFE_PP__3121  (.L_HI(net3121));
 sg13g2_tiehi \cpu.icache.r_data[7][11]$_DFFE_PP__3122  (.L_HI(net3122));
 sg13g2_tiehi \cpu.icache.r_data[7][12]$_DFFE_PP__3123  (.L_HI(net3123));
 sg13g2_tiehi \cpu.icache.r_data[7][13]$_DFFE_PP__3124  (.L_HI(net3124));
 sg13g2_tiehi \cpu.icache.r_data[7][14]$_DFFE_PP__3125  (.L_HI(net3125));
 sg13g2_tiehi \cpu.icache.r_data[7][15]$_DFFE_PP__3126  (.L_HI(net3126));
 sg13g2_tiehi \cpu.icache.r_data[7][16]$_DFFE_PP__3127  (.L_HI(net3127));
 sg13g2_tiehi \cpu.icache.r_data[7][17]$_DFFE_PP__3128  (.L_HI(net3128));
 sg13g2_tiehi \cpu.icache.r_data[7][18]$_DFFE_PP__3129  (.L_HI(net3129));
 sg13g2_tiehi \cpu.icache.r_data[7][19]$_DFFE_PP__3130  (.L_HI(net3130));
 sg13g2_tiehi \cpu.icache.r_data[7][1]$_DFFE_PP__3131  (.L_HI(net3131));
 sg13g2_tiehi \cpu.icache.r_data[7][20]$_DFFE_PP__3132  (.L_HI(net3132));
 sg13g2_tiehi \cpu.icache.r_data[7][21]$_DFFE_PP__3133  (.L_HI(net3133));
 sg13g2_tiehi \cpu.icache.r_data[7][22]$_DFFE_PP__3134  (.L_HI(net3134));
 sg13g2_tiehi \cpu.icache.r_data[7][23]$_DFFE_PP__3135  (.L_HI(net3135));
 sg13g2_tiehi \cpu.icache.r_data[7][24]$_DFFE_PP__3136  (.L_HI(net3136));
 sg13g2_tiehi \cpu.icache.r_data[7][25]$_DFFE_PP__3137  (.L_HI(net3137));
 sg13g2_tiehi \cpu.icache.r_data[7][26]$_DFFE_PP__3138  (.L_HI(net3138));
 sg13g2_tiehi \cpu.icache.r_data[7][27]$_DFFE_PP__3139  (.L_HI(net3139));
 sg13g2_tiehi \cpu.icache.r_data[7][28]$_DFFE_PP__3140  (.L_HI(net3140));
 sg13g2_tiehi \cpu.icache.r_data[7][29]$_DFFE_PP__3141  (.L_HI(net3141));
 sg13g2_tiehi \cpu.icache.r_data[7][2]$_DFFE_PP__3142  (.L_HI(net3142));
 sg13g2_tiehi \cpu.icache.r_data[7][30]$_DFFE_PP__3143  (.L_HI(net3143));
 sg13g2_tiehi \cpu.icache.r_data[7][31]$_DFFE_PP__3144  (.L_HI(net3144));
 sg13g2_tiehi \cpu.icache.r_data[7][3]$_DFFE_PP__3145  (.L_HI(net3145));
 sg13g2_tiehi \cpu.icache.r_data[7][4]$_DFFE_PP__3146  (.L_HI(net3146));
 sg13g2_tiehi \cpu.icache.r_data[7][5]$_DFFE_PP__3147  (.L_HI(net3147));
 sg13g2_tiehi \cpu.icache.r_data[7][6]$_DFFE_PP__3148  (.L_HI(net3148));
 sg13g2_tiehi \cpu.icache.r_data[7][7]$_DFFE_PP__3149  (.L_HI(net3149));
 sg13g2_tiehi \cpu.icache.r_data[7][8]$_DFFE_PP__3150  (.L_HI(net3150));
 sg13g2_tiehi \cpu.icache.r_data[7][9]$_DFFE_PP__3151  (.L_HI(net3151));
 sg13g2_tiehi \cpu.icache.r_offset[0]$_SDFF_PN0__3152  (.L_HI(net3152));
 sg13g2_tiehi \cpu.icache.r_offset[1]$_SDFF_PN0__3153  (.L_HI(net3153));
 sg13g2_tiehi \cpu.icache.r_offset[2]$_SDFF_PN0__3154  (.L_HI(net3154));
 sg13g2_tiehi \cpu.icache.r_tag[0][0]$_DFFE_PP__3155  (.L_HI(net3155));
 sg13g2_tiehi \cpu.icache.r_tag[0][10]$_DFFE_PP__3156  (.L_HI(net3156));
 sg13g2_tiehi \cpu.icache.r_tag[0][11]$_DFFE_PP__3157  (.L_HI(net3157));
 sg13g2_tiehi \cpu.icache.r_tag[0][12]$_DFFE_PP__3158  (.L_HI(net3158));
 sg13g2_tiehi \cpu.icache.r_tag[0][13]$_DFFE_PP__3159  (.L_HI(net3159));
 sg13g2_tiehi \cpu.icache.r_tag[0][14]$_DFFE_PP__3160  (.L_HI(net3160));
 sg13g2_tiehi \cpu.icache.r_tag[0][15]$_DFFE_PP__3161  (.L_HI(net3161));
 sg13g2_tiehi \cpu.icache.r_tag[0][16]$_DFFE_PP__3162  (.L_HI(net3162));
 sg13g2_tiehi \cpu.icache.r_tag[0][17]$_DFFE_PP__3163  (.L_HI(net3163));
 sg13g2_tiehi \cpu.icache.r_tag[0][18]$_DFFE_PP__3164  (.L_HI(net3164));
 sg13g2_tiehi \cpu.icache.r_tag[0][1]$_DFFE_PP__3165  (.L_HI(net3165));
 sg13g2_tiehi \cpu.icache.r_tag[0][2]$_DFFE_PP__3166  (.L_HI(net3166));
 sg13g2_tiehi \cpu.icache.r_tag[0][3]$_DFFE_PP__3167  (.L_HI(net3167));
 sg13g2_tiehi \cpu.icache.r_tag[0][4]$_DFFE_PP__3168  (.L_HI(net3168));
 sg13g2_tiehi \cpu.icache.r_tag[0][5]$_DFFE_PP__3169  (.L_HI(net3169));
 sg13g2_tiehi \cpu.icache.r_tag[0][6]$_DFFE_PP__3170  (.L_HI(net3170));
 sg13g2_tiehi \cpu.icache.r_tag[0][7]$_DFFE_PP__3171  (.L_HI(net3171));
 sg13g2_tiehi \cpu.icache.r_tag[0][8]$_DFFE_PP__3172  (.L_HI(net3172));
 sg13g2_tiehi \cpu.icache.r_tag[0][9]$_DFFE_PP__3173  (.L_HI(net3173));
 sg13g2_tiehi \cpu.icache.r_tag[1][0]$_DFFE_PP__3174  (.L_HI(net3174));
 sg13g2_tiehi \cpu.icache.r_tag[1][10]$_DFFE_PP__3175  (.L_HI(net3175));
 sg13g2_tiehi \cpu.icache.r_tag[1][11]$_DFFE_PP__3176  (.L_HI(net3176));
 sg13g2_tiehi \cpu.icache.r_tag[1][12]$_DFFE_PP__3177  (.L_HI(net3177));
 sg13g2_tiehi \cpu.icache.r_tag[1][13]$_DFFE_PP__3178  (.L_HI(net3178));
 sg13g2_tiehi \cpu.icache.r_tag[1][14]$_DFFE_PP__3179  (.L_HI(net3179));
 sg13g2_tiehi \cpu.icache.r_tag[1][15]$_DFFE_PP__3180  (.L_HI(net3180));
 sg13g2_tiehi \cpu.icache.r_tag[1][16]$_DFFE_PP__3181  (.L_HI(net3181));
 sg13g2_tiehi \cpu.icache.r_tag[1][17]$_DFFE_PP__3182  (.L_HI(net3182));
 sg13g2_tiehi \cpu.icache.r_tag[1][18]$_DFFE_PP__3183  (.L_HI(net3183));
 sg13g2_tiehi \cpu.icache.r_tag[1][1]$_DFFE_PP__3184  (.L_HI(net3184));
 sg13g2_tiehi \cpu.icache.r_tag[1][2]$_DFFE_PP__3185  (.L_HI(net3185));
 sg13g2_tiehi \cpu.icache.r_tag[1][3]$_DFFE_PP__3186  (.L_HI(net3186));
 sg13g2_tiehi \cpu.icache.r_tag[1][4]$_DFFE_PP__3187  (.L_HI(net3187));
 sg13g2_tiehi \cpu.icache.r_tag[1][5]$_DFFE_PP__3188  (.L_HI(net3188));
 sg13g2_tiehi \cpu.icache.r_tag[1][6]$_DFFE_PP__3189  (.L_HI(net3189));
 sg13g2_tiehi \cpu.icache.r_tag[1][7]$_DFFE_PP__3190  (.L_HI(net3190));
 sg13g2_tiehi \cpu.icache.r_tag[1][8]$_DFFE_PP__3191  (.L_HI(net3191));
 sg13g2_tiehi \cpu.icache.r_tag[1][9]$_DFFE_PP__3192  (.L_HI(net3192));
 sg13g2_tiehi \cpu.icache.r_tag[2][0]$_DFFE_PP__3193  (.L_HI(net3193));
 sg13g2_tiehi \cpu.icache.r_tag[2][10]$_DFFE_PP__3194  (.L_HI(net3194));
 sg13g2_tiehi \cpu.icache.r_tag[2][11]$_DFFE_PP__3195  (.L_HI(net3195));
 sg13g2_tiehi \cpu.icache.r_tag[2][12]$_DFFE_PP__3196  (.L_HI(net3196));
 sg13g2_tiehi \cpu.icache.r_tag[2][13]$_DFFE_PP__3197  (.L_HI(net3197));
 sg13g2_tiehi \cpu.icache.r_tag[2][14]$_DFFE_PP__3198  (.L_HI(net3198));
 sg13g2_tiehi \cpu.icache.r_tag[2][15]$_DFFE_PP__3199  (.L_HI(net3199));
 sg13g2_tiehi \cpu.icache.r_tag[2][16]$_DFFE_PP__3200  (.L_HI(net3200));
 sg13g2_tiehi \cpu.icache.r_tag[2][17]$_DFFE_PP__3201  (.L_HI(net3201));
 sg13g2_tiehi \cpu.icache.r_tag[2][18]$_DFFE_PP__3202  (.L_HI(net3202));
 sg13g2_tiehi \cpu.icache.r_tag[2][1]$_DFFE_PP__3203  (.L_HI(net3203));
 sg13g2_tiehi \cpu.icache.r_tag[2][2]$_DFFE_PP__3204  (.L_HI(net3204));
 sg13g2_tiehi \cpu.icache.r_tag[2][3]$_DFFE_PP__3205  (.L_HI(net3205));
 sg13g2_tiehi \cpu.icache.r_tag[2][4]$_DFFE_PP__3206  (.L_HI(net3206));
 sg13g2_tiehi \cpu.icache.r_tag[2][5]$_DFFE_PP__3207  (.L_HI(net3207));
 sg13g2_tiehi \cpu.icache.r_tag[2][6]$_DFFE_PP__3208  (.L_HI(net3208));
 sg13g2_tiehi \cpu.icache.r_tag[2][7]$_DFFE_PP__3209  (.L_HI(net3209));
 sg13g2_tiehi \cpu.icache.r_tag[2][8]$_DFFE_PP__3210  (.L_HI(net3210));
 sg13g2_tiehi \cpu.icache.r_tag[2][9]$_DFFE_PP__3211  (.L_HI(net3211));
 sg13g2_tiehi \cpu.icache.r_tag[3][0]$_DFFE_PP__3212  (.L_HI(net3212));
 sg13g2_tiehi \cpu.icache.r_tag[3][10]$_DFFE_PP__3213  (.L_HI(net3213));
 sg13g2_tiehi \cpu.icache.r_tag[3][11]$_DFFE_PP__3214  (.L_HI(net3214));
 sg13g2_tiehi \cpu.icache.r_tag[3][12]$_DFFE_PP__3215  (.L_HI(net3215));
 sg13g2_tiehi \cpu.icache.r_tag[3][13]$_DFFE_PP__3216  (.L_HI(net3216));
 sg13g2_tiehi \cpu.icache.r_tag[3][14]$_DFFE_PP__3217  (.L_HI(net3217));
 sg13g2_tiehi \cpu.icache.r_tag[3][15]$_DFFE_PP__3218  (.L_HI(net3218));
 sg13g2_tiehi \cpu.icache.r_tag[3][16]$_DFFE_PP__3219  (.L_HI(net3219));
 sg13g2_tiehi \cpu.icache.r_tag[3][17]$_DFFE_PP__3220  (.L_HI(net3220));
 sg13g2_tiehi \cpu.icache.r_tag[3][18]$_DFFE_PP__3221  (.L_HI(net3221));
 sg13g2_tiehi \cpu.icache.r_tag[3][1]$_DFFE_PP__3222  (.L_HI(net3222));
 sg13g2_tiehi \cpu.icache.r_tag[3][2]$_DFFE_PP__3223  (.L_HI(net3223));
 sg13g2_tiehi \cpu.icache.r_tag[3][3]$_DFFE_PP__3224  (.L_HI(net3224));
 sg13g2_tiehi \cpu.icache.r_tag[3][4]$_DFFE_PP__3225  (.L_HI(net3225));
 sg13g2_tiehi \cpu.icache.r_tag[3][5]$_DFFE_PP__3226  (.L_HI(net3226));
 sg13g2_tiehi \cpu.icache.r_tag[3][6]$_DFFE_PP__3227  (.L_HI(net3227));
 sg13g2_tiehi \cpu.icache.r_tag[3][7]$_DFFE_PP__3228  (.L_HI(net3228));
 sg13g2_tiehi \cpu.icache.r_tag[3][8]$_DFFE_PP__3229  (.L_HI(net3229));
 sg13g2_tiehi \cpu.icache.r_tag[3][9]$_DFFE_PP__3230  (.L_HI(net3230));
 sg13g2_tiehi \cpu.icache.r_tag[4][0]$_DFFE_PP__3231  (.L_HI(net3231));
 sg13g2_tiehi \cpu.icache.r_tag[4][10]$_DFFE_PP__3232  (.L_HI(net3232));
 sg13g2_tiehi \cpu.icache.r_tag[4][11]$_DFFE_PP__3233  (.L_HI(net3233));
 sg13g2_tiehi \cpu.icache.r_tag[4][12]$_DFFE_PP__3234  (.L_HI(net3234));
 sg13g2_tiehi \cpu.icache.r_tag[4][13]$_DFFE_PP__3235  (.L_HI(net3235));
 sg13g2_tiehi \cpu.icache.r_tag[4][14]$_DFFE_PP__3236  (.L_HI(net3236));
 sg13g2_tiehi \cpu.icache.r_tag[4][15]$_DFFE_PP__3237  (.L_HI(net3237));
 sg13g2_tiehi \cpu.icache.r_tag[4][16]$_DFFE_PP__3238  (.L_HI(net3238));
 sg13g2_tiehi \cpu.icache.r_tag[4][17]$_DFFE_PP__3239  (.L_HI(net3239));
 sg13g2_tiehi \cpu.icache.r_tag[4][18]$_DFFE_PP__3240  (.L_HI(net3240));
 sg13g2_tiehi \cpu.icache.r_tag[4][1]$_DFFE_PP__3241  (.L_HI(net3241));
 sg13g2_tiehi \cpu.icache.r_tag[4][2]$_DFFE_PP__3242  (.L_HI(net3242));
 sg13g2_tiehi \cpu.icache.r_tag[4][3]$_DFFE_PP__3243  (.L_HI(net3243));
 sg13g2_tiehi \cpu.icache.r_tag[4][4]$_DFFE_PP__3244  (.L_HI(net3244));
 sg13g2_tiehi \cpu.icache.r_tag[4][5]$_DFFE_PP__3245  (.L_HI(net3245));
 sg13g2_tiehi \cpu.icache.r_tag[4][6]$_DFFE_PP__3246  (.L_HI(net3246));
 sg13g2_tiehi \cpu.icache.r_tag[4][7]$_DFFE_PP__3247  (.L_HI(net3247));
 sg13g2_tiehi \cpu.icache.r_tag[4][8]$_DFFE_PP__3248  (.L_HI(net3248));
 sg13g2_tiehi \cpu.icache.r_tag[4][9]$_DFFE_PP__3249  (.L_HI(net3249));
 sg13g2_tiehi \cpu.icache.r_tag[5][0]$_DFFE_PP__3250  (.L_HI(net3250));
 sg13g2_tiehi \cpu.icache.r_tag[5][10]$_DFFE_PP__3251  (.L_HI(net3251));
 sg13g2_tiehi \cpu.icache.r_tag[5][11]$_DFFE_PP__3252  (.L_HI(net3252));
 sg13g2_tiehi \cpu.icache.r_tag[5][12]$_DFFE_PP__3253  (.L_HI(net3253));
 sg13g2_tiehi \cpu.icache.r_tag[5][13]$_DFFE_PP__3254  (.L_HI(net3254));
 sg13g2_tiehi \cpu.icache.r_tag[5][14]$_DFFE_PP__3255  (.L_HI(net3255));
 sg13g2_tiehi \cpu.icache.r_tag[5][15]$_DFFE_PP__3256  (.L_HI(net3256));
 sg13g2_tiehi \cpu.icache.r_tag[5][16]$_DFFE_PP__3257  (.L_HI(net3257));
 sg13g2_tiehi \cpu.icache.r_tag[5][17]$_DFFE_PP__3258  (.L_HI(net3258));
 sg13g2_tiehi \cpu.icache.r_tag[5][18]$_DFFE_PP__3259  (.L_HI(net3259));
 sg13g2_tiehi \cpu.icache.r_tag[5][1]$_DFFE_PP__3260  (.L_HI(net3260));
 sg13g2_tiehi \cpu.icache.r_tag[5][2]$_DFFE_PP__3261  (.L_HI(net3261));
 sg13g2_tiehi \cpu.icache.r_tag[5][3]$_DFFE_PP__3262  (.L_HI(net3262));
 sg13g2_tiehi \cpu.icache.r_tag[5][4]$_DFFE_PP__3263  (.L_HI(net3263));
 sg13g2_tiehi \cpu.icache.r_tag[5][5]$_DFFE_PP__3264  (.L_HI(net3264));
 sg13g2_tiehi \cpu.icache.r_tag[5][6]$_DFFE_PP__3265  (.L_HI(net3265));
 sg13g2_tiehi \cpu.icache.r_tag[5][7]$_DFFE_PP__3266  (.L_HI(net3266));
 sg13g2_tiehi \cpu.icache.r_tag[5][8]$_DFFE_PP__3267  (.L_HI(net3267));
 sg13g2_tiehi \cpu.icache.r_tag[5][9]$_DFFE_PP__3268  (.L_HI(net3268));
 sg13g2_tiehi \cpu.icache.r_tag[6][0]$_DFFE_PP__3269  (.L_HI(net3269));
 sg13g2_tiehi \cpu.icache.r_tag[6][10]$_DFFE_PP__3270  (.L_HI(net3270));
 sg13g2_tiehi \cpu.icache.r_tag[6][11]$_DFFE_PP__3271  (.L_HI(net3271));
 sg13g2_tiehi \cpu.icache.r_tag[6][12]$_DFFE_PP__3272  (.L_HI(net3272));
 sg13g2_tiehi \cpu.icache.r_tag[6][13]$_DFFE_PP__3273  (.L_HI(net3273));
 sg13g2_tiehi \cpu.icache.r_tag[6][14]$_DFFE_PP__3274  (.L_HI(net3274));
 sg13g2_tiehi \cpu.icache.r_tag[6][15]$_DFFE_PP__3275  (.L_HI(net3275));
 sg13g2_tiehi \cpu.icache.r_tag[6][16]$_DFFE_PP__3276  (.L_HI(net3276));
 sg13g2_tiehi \cpu.icache.r_tag[6][17]$_DFFE_PP__3277  (.L_HI(net3277));
 sg13g2_tiehi \cpu.icache.r_tag[6][18]$_DFFE_PP__3278  (.L_HI(net3278));
 sg13g2_tiehi \cpu.icache.r_tag[6][1]$_DFFE_PP__3279  (.L_HI(net3279));
 sg13g2_tiehi \cpu.icache.r_tag[6][2]$_DFFE_PP__3280  (.L_HI(net3280));
 sg13g2_tiehi \cpu.icache.r_tag[6][3]$_DFFE_PP__3281  (.L_HI(net3281));
 sg13g2_tiehi \cpu.icache.r_tag[6][4]$_DFFE_PP__3282  (.L_HI(net3282));
 sg13g2_tiehi \cpu.icache.r_tag[6][5]$_DFFE_PP__3283  (.L_HI(net3283));
 sg13g2_tiehi \cpu.icache.r_tag[6][6]$_DFFE_PP__3284  (.L_HI(net3284));
 sg13g2_tiehi \cpu.icache.r_tag[6][7]$_DFFE_PP__3285  (.L_HI(net3285));
 sg13g2_tiehi \cpu.icache.r_tag[6][8]$_DFFE_PP__3286  (.L_HI(net3286));
 sg13g2_tiehi \cpu.icache.r_tag[6][9]$_DFFE_PP__3287  (.L_HI(net3287));
 sg13g2_tiehi \cpu.icache.r_tag[7][0]$_DFFE_PP__3288  (.L_HI(net3288));
 sg13g2_tiehi \cpu.icache.r_tag[7][10]$_DFFE_PP__3289  (.L_HI(net3289));
 sg13g2_tiehi \cpu.icache.r_tag[7][11]$_DFFE_PP__3290  (.L_HI(net3290));
 sg13g2_tiehi \cpu.icache.r_tag[7][12]$_DFFE_PP__3291  (.L_HI(net3291));
 sg13g2_tiehi \cpu.icache.r_tag[7][13]$_DFFE_PP__3292  (.L_HI(net3292));
 sg13g2_tiehi \cpu.icache.r_tag[7][14]$_DFFE_PP__3293  (.L_HI(net3293));
 sg13g2_tiehi \cpu.icache.r_tag[7][15]$_DFFE_PP__3294  (.L_HI(net3294));
 sg13g2_tiehi \cpu.icache.r_tag[7][16]$_DFFE_PP__3295  (.L_HI(net3295));
 sg13g2_tiehi \cpu.icache.r_tag[7][17]$_DFFE_PP__3296  (.L_HI(net3296));
 sg13g2_tiehi \cpu.icache.r_tag[7][18]$_DFFE_PP__3297  (.L_HI(net3297));
 sg13g2_tiehi \cpu.icache.r_tag[7][1]$_DFFE_PP__3298  (.L_HI(net3298));
 sg13g2_tiehi \cpu.icache.r_tag[7][2]$_DFFE_PP__3299  (.L_HI(net3299));
 sg13g2_tiehi \cpu.icache.r_tag[7][3]$_DFFE_PP__3300  (.L_HI(net3300));
 sg13g2_tiehi \cpu.icache.r_tag[7][4]$_DFFE_PP__3301  (.L_HI(net3301));
 sg13g2_tiehi \cpu.icache.r_tag[7][5]$_DFFE_PP__3302  (.L_HI(net3302));
 sg13g2_tiehi \cpu.icache.r_tag[7][6]$_DFFE_PP__3303  (.L_HI(net3303));
 sg13g2_tiehi \cpu.icache.r_tag[7][7]$_DFFE_PP__3304  (.L_HI(net3304));
 sg13g2_tiehi \cpu.icache.r_tag[7][8]$_DFFE_PP__3305  (.L_HI(net3305));
 sg13g2_tiehi \cpu.icache.r_tag[7][9]$_DFFE_PP__3306  (.L_HI(net3306));
 sg13g2_tiehi \cpu.icache.r_valid[0]$_SDFFE_PP0P__3307  (.L_HI(net3307));
 sg13g2_tiehi \cpu.icache.r_valid[1]$_SDFFE_PP0P__3308  (.L_HI(net3308));
 sg13g2_tiehi \cpu.icache.r_valid[2]$_SDFFE_PP0P__3309  (.L_HI(net3309));
 sg13g2_tiehi \cpu.icache.r_valid[3]$_SDFFE_PP0P__3310  (.L_HI(net3310));
 sg13g2_tiehi \cpu.icache.r_valid[4]$_SDFFE_PP0P__3311  (.L_HI(net3311));
 sg13g2_tiehi \cpu.icache.r_valid[5]$_SDFFE_PP0P__3312  (.L_HI(net3312));
 sg13g2_tiehi \cpu.icache.r_valid[6]$_SDFFE_PP0P__3313  (.L_HI(net3313));
 sg13g2_tiehi \cpu.icache.r_valid[7]$_SDFFE_PP0P__3314  (.L_HI(net3314));
 sg13g2_tiehi \cpu.intr.r_clock$_SDFFE_PN0P__3315  (.L_HI(net3315));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[0]$_DFFE_PP__3316  (.L_HI(net3316));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[10]$_DFFE_PP__3317  (.L_HI(net3317));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[11]$_DFFE_PP__3318  (.L_HI(net3318));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[12]$_DFFE_PP__3319  (.L_HI(net3319));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[13]$_DFFE_PP__3320  (.L_HI(net3320));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[14]$_DFFE_PP__3321  (.L_HI(net3321));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[15]$_DFFE_PP__3322  (.L_HI(net3322));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[16]$_DFFE_PP__3323  (.L_HI(net3323));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[17]$_DFFE_PP__3324  (.L_HI(net3324));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[18]$_DFFE_PP__3325  (.L_HI(net3325));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[19]$_DFFE_PP__3326  (.L_HI(net3326));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[1]$_DFFE_PP__3327  (.L_HI(net3327));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[20]$_DFFE_PP__3328  (.L_HI(net3328));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[21]$_DFFE_PP__3329  (.L_HI(net3329));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[22]$_DFFE_PP__3330  (.L_HI(net3330));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[23]$_DFFE_PP__3331  (.L_HI(net3331));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[24]$_DFFE_PP__3332  (.L_HI(net3332));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[25]$_DFFE_PP__3333  (.L_HI(net3333));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[26]$_DFFE_PP__3334  (.L_HI(net3334));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[27]$_DFFE_PP__3335  (.L_HI(net3335));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[28]$_DFFE_PP__3336  (.L_HI(net3336));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[29]$_DFFE_PP__3337  (.L_HI(net3337));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[2]$_DFFE_PP__3338  (.L_HI(net3338));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[30]$_DFFE_PP__3339  (.L_HI(net3339));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[31]$_DFFE_PP__3340  (.L_HI(net3340));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[3]$_DFFE_PP__3341  (.L_HI(net3341));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[4]$_DFFE_PP__3342  (.L_HI(net3342));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[5]$_DFFE_PP__3343  (.L_HI(net3343));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[6]$_DFFE_PP__3344  (.L_HI(net3344));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[7]$_DFFE_PP__3345  (.L_HI(net3345));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[8]$_DFFE_PP__3346  (.L_HI(net3346));
 sg13g2_tiehi \cpu.intr.r_clock_cmp[9]$_DFFE_PP__3347  (.L_HI(net3347));
 sg13g2_tiehi \cpu.intr.r_clock_count[0]$_DFF_P__3348  (.L_HI(net3348));
 sg13g2_tiehi \cpu.intr.r_clock_count[10]$_DFF_P__3349  (.L_HI(net3349));
 sg13g2_tiehi \cpu.intr.r_clock_count[11]$_DFF_P__3350  (.L_HI(net3350));
 sg13g2_tiehi \cpu.intr.r_clock_count[12]$_DFF_P__3351  (.L_HI(net3351));
 sg13g2_tiehi \cpu.intr.r_clock_count[13]$_DFF_P__3352  (.L_HI(net3352));
 sg13g2_tiehi \cpu.intr.r_clock_count[14]$_DFF_P__3353  (.L_HI(net3353));
 sg13g2_tiehi \cpu.intr.r_clock_count[15]$_DFF_P__3354  (.L_HI(net3354));
 sg13g2_tiehi \cpu.intr.r_clock_count[16]$_DFFE_PN__3355  (.L_HI(net3355));
 sg13g2_tiehi \cpu.intr.r_clock_count[17]$_DFFE_PN__3356  (.L_HI(net3356));
 sg13g2_tiehi \cpu.intr.r_clock_count[18]$_DFFE_PN__3357  (.L_HI(net3357));
 sg13g2_tiehi \cpu.intr.r_clock_count[19]$_DFFE_PN__3358  (.L_HI(net3358));
 sg13g2_tiehi \cpu.intr.r_clock_count[1]$_DFF_P__3359  (.L_HI(net3359));
 sg13g2_tiehi \cpu.intr.r_clock_count[20]$_DFFE_PN__3360  (.L_HI(net3360));
 sg13g2_tiehi \cpu.intr.r_clock_count[21]$_DFFE_PN__3361  (.L_HI(net3361));
 sg13g2_tiehi \cpu.intr.r_clock_count[22]$_DFFE_PN__3362  (.L_HI(net3362));
 sg13g2_tiehi \cpu.intr.r_clock_count[23]$_DFFE_PN__3363  (.L_HI(net3363));
 sg13g2_tiehi \cpu.intr.r_clock_count[24]$_DFFE_PN__3364  (.L_HI(net3364));
 sg13g2_tiehi \cpu.intr.r_clock_count[25]$_DFFE_PN__3365  (.L_HI(net3365));
 sg13g2_tiehi \cpu.intr.r_clock_count[26]$_DFFE_PN__3366  (.L_HI(net3366));
 sg13g2_tiehi \cpu.intr.r_clock_count[27]$_DFFE_PN__3367  (.L_HI(net3367));
 sg13g2_tiehi \cpu.intr.r_clock_count[28]$_DFFE_PN__3368  (.L_HI(net3368));
 sg13g2_tiehi \cpu.intr.r_clock_count[29]$_DFFE_PN__3369  (.L_HI(net3369));
 sg13g2_tiehi \cpu.intr.r_clock_count[2]$_DFF_P__3370  (.L_HI(net3370));
 sg13g2_tiehi \cpu.intr.r_clock_count[30]$_DFFE_PN__3371  (.L_HI(net3371));
 sg13g2_tiehi \cpu.intr.r_clock_count[31]$_DFFE_PN__3372  (.L_HI(net3372));
 sg13g2_tiehi \cpu.intr.r_clock_count[3]$_DFF_P__3373  (.L_HI(net3373));
 sg13g2_tiehi \cpu.intr.r_clock_count[4]$_DFF_P__3374  (.L_HI(net3374));
 sg13g2_tiehi \cpu.intr.r_clock_count[5]$_DFF_P__3375  (.L_HI(net3375));
 sg13g2_tiehi \cpu.intr.r_clock_count[6]$_DFF_P__3376  (.L_HI(net3376));
 sg13g2_tiehi \cpu.intr.r_clock_count[7]$_DFF_P__3377  (.L_HI(net3377));
 sg13g2_tiehi \cpu.intr.r_clock_count[8]$_DFF_P__3378  (.L_HI(net3378));
 sg13g2_tiehi \cpu.intr.r_clock_count[9]$_DFF_P__3379  (.L_HI(net3379));
 sg13g2_tiehi \cpu.intr.r_enable[0]$_SDFFE_PN0P__3380  (.L_HI(net3380));
 sg13g2_tiehi \cpu.intr.r_enable[1]$_SDFFE_PN0P__3381  (.L_HI(net3381));
 sg13g2_tiehi \cpu.intr.r_enable[2]$_SDFFE_PN0P__3382  (.L_HI(net3382));
 sg13g2_tiehi \cpu.intr.r_enable[3]$_SDFFE_PN0P__3383  (.L_HI(net3383));
 sg13g2_tiehi \cpu.intr.r_enable[4]$_SDFFE_PN0P__3384  (.L_HI(net3384));
 sg13g2_tiehi \cpu.intr.r_enable[5]$_SDFFE_PN0P__3385  (.L_HI(net3385));
 sg13g2_tiehi \cpu.intr.r_timer$_SDFFE_PN0P__3386  (.L_HI(net3386));
 sg13g2_tiehi \cpu.intr.r_timer_count[0]$_DFF_P__3387  (.L_HI(net3387));
 sg13g2_tiehi \cpu.intr.r_timer_count[10]$_DFF_P__3388  (.L_HI(net3388));
 sg13g2_tiehi \cpu.intr.r_timer_count[11]$_DFF_P__3389  (.L_HI(net3389));
 sg13g2_tiehi \cpu.intr.r_timer_count[12]$_DFF_P__3390  (.L_HI(net3390));
 sg13g2_tiehi \cpu.intr.r_timer_count[13]$_DFF_P__3391  (.L_HI(net3391));
 sg13g2_tiehi \cpu.intr.r_timer_count[14]$_DFF_P__3392  (.L_HI(net3392));
 sg13g2_tiehi \cpu.intr.r_timer_count[15]$_DFF_P__3393  (.L_HI(net3393));
 sg13g2_tiehi \cpu.intr.r_timer_count[16]$_DFF_P__3394  (.L_HI(net3394));
 sg13g2_tiehi \cpu.intr.r_timer_count[17]$_DFF_P__3395  (.L_HI(net3395));
 sg13g2_tiehi \cpu.intr.r_timer_count[18]$_DFF_P__3396  (.L_HI(net3396));
 sg13g2_tiehi \cpu.intr.r_timer_count[19]$_DFF_P__3397  (.L_HI(net3397));
 sg13g2_tiehi \cpu.intr.r_timer_count[1]$_DFF_P__3398  (.L_HI(net3398));
 sg13g2_tiehi \cpu.intr.r_timer_count[20]$_DFF_P__3399  (.L_HI(net3399));
 sg13g2_tiehi \cpu.intr.r_timer_count[21]$_DFF_P__3400  (.L_HI(net3400));
 sg13g2_tiehi \cpu.intr.r_timer_count[22]$_DFF_P__3401  (.L_HI(net3401));
 sg13g2_tiehi \cpu.intr.r_timer_count[23]$_DFF_P__3402  (.L_HI(net3402));
 sg13g2_tiehi \cpu.intr.r_timer_count[2]$_DFF_P__3403  (.L_HI(net3403));
 sg13g2_tiehi \cpu.intr.r_timer_count[3]$_DFF_P__3404  (.L_HI(net3404));
 sg13g2_tiehi \cpu.intr.r_timer_count[4]$_DFF_P__3405  (.L_HI(net3405));
 sg13g2_tiehi \cpu.intr.r_timer_count[5]$_DFF_P__3406  (.L_HI(net3406));
 sg13g2_tiehi \cpu.intr.r_timer_count[6]$_DFF_P__3407  (.L_HI(net3407));
 sg13g2_tiehi \cpu.intr.r_timer_count[7]$_DFF_P__3408  (.L_HI(net3408));
 sg13g2_tiehi \cpu.intr.r_timer_count[8]$_DFF_P__3409  (.L_HI(net3409));
 sg13g2_tiehi \cpu.intr.r_timer_count[9]$_DFF_P__3410  (.L_HI(net3410));
 sg13g2_tiehi \cpu.intr.r_timer_reload[0]$_DFFE_PP__3411  (.L_HI(net3411));
 sg13g2_tiehi \cpu.intr.r_timer_reload[10]$_DFFE_PP__3412  (.L_HI(net3412));
 sg13g2_tiehi \cpu.intr.r_timer_reload[11]$_DFFE_PP__3413  (.L_HI(net3413));
 sg13g2_tiehi \cpu.intr.r_timer_reload[12]$_DFFE_PP__3414  (.L_HI(net3414));
 sg13g2_tiehi \cpu.intr.r_timer_reload[13]$_DFFE_PP__3415  (.L_HI(net3415));
 sg13g2_tiehi \cpu.intr.r_timer_reload[14]$_DFFE_PP__3416  (.L_HI(net3416));
 sg13g2_tiehi \cpu.intr.r_timer_reload[15]$_DFFE_PP__3417  (.L_HI(net3417));
 sg13g2_tiehi \cpu.intr.r_timer_reload[16]$_DFFE_PP__3418  (.L_HI(net3418));
 sg13g2_tiehi \cpu.intr.r_timer_reload[17]$_DFFE_PP__3419  (.L_HI(net3419));
 sg13g2_tiehi \cpu.intr.r_timer_reload[18]$_DFFE_PP__3420  (.L_HI(net3420));
 sg13g2_tiehi \cpu.intr.r_timer_reload[19]$_DFFE_PP__3421  (.L_HI(net3421));
 sg13g2_tiehi \cpu.intr.r_timer_reload[1]$_DFFE_PP__3422  (.L_HI(net3422));
 sg13g2_tiehi \cpu.intr.r_timer_reload[20]$_DFFE_PP__3423  (.L_HI(net3423));
 sg13g2_tiehi \cpu.intr.r_timer_reload[21]$_DFFE_PP__3424  (.L_HI(net3424));
 sg13g2_tiehi \cpu.intr.r_timer_reload[22]$_DFFE_PP__3425  (.L_HI(net3425));
 sg13g2_tiehi \cpu.intr.r_timer_reload[23]$_DFFE_PP__3426  (.L_HI(net3426));
 sg13g2_tiehi \cpu.intr.r_timer_reload[2]$_DFFE_PP__3427  (.L_HI(net3427));
 sg13g2_tiehi \cpu.intr.r_timer_reload[3]$_DFFE_PP__3428  (.L_HI(net3428));
 sg13g2_tiehi \cpu.intr.r_timer_reload[4]$_DFFE_PP__3429  (.L_HI(net3429));
 sg13g2_tiehi \cpu.intr.r_timer_reload[5]$_DFFE_PP__3430  (.L_HI(net3430));
 sg13g2_tiehi \cpu.intr.r_timer_reload[6]$_DFFE_PP__3431  (.L_HI(net3431));
 sg13g2_tiehi \cpu.intr.r_timer_reload[7]$_DFFE_PP__3432  (.L_HI(net3432));
 sg13g2_tiehi \cpu.intr.r_timer_reload[8]$_DFFE_PP__3433  (.L_HI(net3433));
 sg13g2_tiehi \cpu.intr.r_timer_reload[9]$_DFFE_PP__3434  (.L_HI(net3434));
 sg13g2_tiehi \cpu.qspi.r_count[0]$_DFFE_PP__3435  (.L_HI(net3435));
 sg13g2_tiehi \cpu.qspi.r_count[1]$_DFFE_PP__3436  (.L_HI(net3436));
 sg13g2_tiehi \cpu.qspi.r_count[2]$_DFFE_PP__3437  (.L_HI(net3437));
 sg13g2_tiehi \cpu.qspi.r_count[3]$_DFFE_PP__3438  (.L_HI(net3438));
 sg13g2_tiehi \cpu.qspi.r_count[4]$_DFFE_PP__3439  (.L_HI(net3439));
 sg13g2_tiehi \cpu.qspi.r_cs[0]$_SDFFE_PN1P__3440  (.L_HI(net3440));
 sg13g2_tiehi \cpu.qspi.r_cs[1]$_SDFFE_PN1P__3441  (.L_HI(net3441));
 sg13g2_tiehi \cpu.qspi.r_cs[2]$_SDFFE_PN1P__3442  (.L_HI(net3442));
 sg13g2_tiehi \cpu.qspi.r_ind$_SDFFE_PN0N__3443  (.L_HI(net3443));
 sg13g2_tiehi \cpu.qspi.r_mask[0]$_SDFFE_PN0P__3444  (.L_HI(net3444));
 sg13g2_tiehi \cpu.qspi.r_mask[1]$_SDFFE_PN1P__3445  (.L_HI(net3445));
 sg13g2_tiehi \cpu.qspi.r_mask[2]$_SDFFE_PN0P__3446  (.L_HI(net3446));
 sg13g2_tiehi \cpu.qspi.r_quad[0]$_SDFFE_PN1P__3447  (.L_HI(net3447));
 sg13g2_tiehi \cpu.qspi.r_quad[1]$_SDFFE_PN0P__3448  (.L_HI(net3448));
 sg13g2_tiehi \cpu.qspi.r_quad[2]$_SDFFE_PN1P__3449  (.L_HI(net3449));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][0]$_SDFFCE_PN0P__3450  (.L_HI(net3450));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][1]$_SDFFCE_PN0P__3451  (.L_HI(net3451));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][2]$_SDFFCE_PN1P__3452  (.L_HI(net3452));
 sg13g2_tiehi \cpu.qspi.r_read_delay[0][3]$_SDFFCE_PN0P__3453  (.L_HI(net3453));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][0]$_SDFFCE_PN0P__3454  (.L_HI(net3454));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][1]$_SDFFCE_PN0P__3455  (.L_HI(net3455));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][2]$_SDFFCE_PN1P__3456  (.L_HI(net3456));
 sg13g2_tiehi \cpu.qspi.r_read_delay[1][3]$_SDFFCE_PN0P__3457  (.L_HI(net3457));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][0]$_SDFFCE_PN0P__3458  (.L_HI(net3458));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][1]$_SDFFCE_PN0P__3459  (.L_HI(net3459));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][2]$_SDFFCE_PN1P__3460  (.L_HI(net3460));
 sg13g2_tiehi \cpu.qspi.r_read_delay[2][3]$_SDFFCE_PN0P__3461  (.L_HI(net3461));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[0]$_SDFFE_PN1P__3462  (.L_HI(net3462));
 sg13g2_tiehi \cpu.qspi.r_rom_mode[1]$_SDFFE_PN1P__3463  (.L_HI(net3463));
 sg13g2_tiehi \cpu.qspi.r_rstrobe_d$_DFF_P__3464  (.L_HI(net3464));
 sg13g2_tiehi \cpu.qspi.r_state[0]$_DFF_P__3465  (.L_HI(net3465));
 sg13g2_tiehi \cpu.qspi.r_state[10]$_DFF_P__3466  (.L_HI(net3466));
 sg13g2_tiehi \cpu.qspi.r_state[11]$_DFF_P__3467  (.L_HI(net3467));
 sg13g2_tiehi \cpu.qspi.r_state[12]$_DFF_P__3468  (.L_HI(net3468));
 sg13g2_tiehi \cpu.qspi.r_state[13]$_DFF_P__3469  (.L_HI(net3469));
 sg13g2_tiehi \cpu.qspi.r_state[14]$_DFF_P__3470  (.L_HI(net3470));
 sg13g2_tiehi \cpu.qspi.r_state[15]$_DFF_P__3471  (.L_HI(net3471));
 sg13g2_tiehi \cpu.qspi.r_state[16]$_DFF_P__3472  (.L_HI(net3472));
 sg13g2_tiehi \cpu.qspi.r_state[17]$_DFF_P__3473  (.L_HI(net3473));
 sg13g2_tiehi \cpu.qspi.r_state[1]$_DFF_P__3474  (.L_HI(net3474));
 sg13g2_tiehi \cpu.qspi.r_state[2]$_DFF_P__3475  (.L_HI(net3475));
 sg13g2_tiehi \cpu.qspi.r_state[3]$_DFF_P__3476  (.L_HI(net3476));
 sg13g2_tiehi \cpu.qspi.r_state[4]$_DFF_P__3477  (.L_HI(net3477));
 sg13g2_tiehi \cpu.qspi.r_state[5]$_DFF_P__3478  (.L_HI(net3478));
 sg13g2_tiehi \cpu.qspi.r_state[6]$_DFF_P__3479  (.L_HI(net3479));
 sg13g2_tiehi \cpu.qspi.r_state[7]$_DFF_P__3480  (.L_HI(net3480));
 sg13g2_tiehi \cpu.qspi.r_state[8]$_DFF_P__3481  (.L_HI(net3481));
 sg13g2_tiehi \cpu.qspi.r_state[9]$_DFF_P__3482  (.L_HI(net3482));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[0]$_SDFFE_PN0P__3483  (.L_HI(net3483));
 sg13g2_tiehi \cpu.qspi.r_uio_oe[1]$_SDFFE_PN0P__3484  (.L_HI(net3484));
 sg13g2_tiehi \cpu.qspi.r_uio_out[0]$_DFFE_PP__3485  (.L_HI(net3485));
 sg13g2_tiehi \cpu.qspi.r_uio_out[1]$_DFFE_PP__3486  (.L_HI(net3486));
 sg13g2_tiehi \cpu.qspi.r_uio_out[2]$_DFFE_PP__3487  (.L_HI(net3487));
 sg13g2_tiehi \cpu.qspi.r_uio_out[3]$_DFFE_PP__3488  (.L_HI(net3488));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_d$_DFF_P__3489  (.L_HI(net3489));
 sg13g2_tiehi \cpu.qspi.r_wstrobe_i$_DFF_P__3490  (.L_HI(net3490));
 sg13g2_tiehi \cpu.r_clk_invert$_DFFE_PN__3491  (.L_HI(net3491));
 sg13g2_tiehi \cpu.spi.r_bits[0]$_SDFFE_PN1P__3492  (.L_HI(net3492));
 sg13g2_tiehi \cpu.spi.r_bits[1]$_SDFFE_PN1P__3493  (.L_HI(net3493));
 sg13g2_tiehi \cpu.spi.r_bits[2]$_SDFFE_PN1P__3494  (.L_HI(net3494));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][0]$_DFFE_PP__3495  (.L_HI(net3495));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][1]$_DFFE_PP__3496  (.L_HI(net3496));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][2]$_DFFE_PP__3497  (.L_HI(net3497));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][3]$_DFFE_PP__3498  (.L_HI(net3498));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][4]$_DFFE_PP__3499  (.L_HI(net3499));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][5]$_DFFE_PP__3500  (.L_HI(net3500));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][6]$_DFFE_PP__3501  (.L_HI(net3501));
 sg13g2_tiehi \cpu.spi.r_clk_count[0][7]$_DFFE_PP__3502  (.L_HI(net3502));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][0]$_DFFE_PP__3503  (.L_HI(net3503));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][1]$_DFFE_PP__3504  (.L_HI(net3504));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][2]$_DFFE_PP__3505  (.L_HI(net3505));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][3]$_DFFE_PP__3506  (.L_HI(net3506));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][4]$_DFFE_PP__3507  (.L_HI(net3507));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][5]$_DFFE_PP__3508  (.L_HI(net3508));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][6]$_DFFE_PP__3509  (.L_HI(net3509));
 sg13g2_tiehi \cpu.spi.r_clk_count[1][7]$_DFFE_PP__3510  (.L_HI(net3510));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][0]$_DFFE_PP__3511  (.L_HI(net3511));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][1]$_DFFE_PP__3512  (.L_HI(net3512));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][2]$_DFFE_PP__3513  (.L_HI(net3513));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][3]$_DFFE_PP__3514  (.L_HI(net3514));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][4]$_DFFE_PP__3515  (.L_HI(net3515));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][5]$_DFFE_PP__3516  (.L_HI(net3516));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][6]$_DFFE_PP__3517  (.L_HI(net3517));
 sg13g2_tiehi \cpu.spi.r_clk_count[2][7]$_DFFE_PP__3518  (.L_HI(net3518));
 sg13g2_tiehi \cpu.spi.r_count[0]$_DFFE_PP__3519  (.L_HI(net3519));
 sg13g2_tiehi \cpu.spi.r_count[1]$_DFFE_PP__3520  (.L_HI(net3520));
 sg13g2_tiehi \cpu.spi.r_count[2]$_DFFE_PP__3521  (.L_HI(net3521));
 sg13g2_tiehi \cpu.spi.r_count[3]$_DFFE_PP__3522  (.L_HI(net3522));
 sg13g2_tiehi \cpu.spi.r_count[4]$_DFFE_PP__3523  (.L_HI(net3523));
 sg13g2_tiehi \cpu.spi.r_count[5]$_DFFE_PP__3524  (.L_HI(net3524));
 sg13g2_tiehi \cpu.spi.r_count[6]$_DFFE_PP__3525  (.L_HI(net3525));
 sg13g2_tiehi \cpu.spi.r_count[7]$_DFFE_PP__3526  (.L_HI(net3526));
 sg13g2_tiehi \cpu.spi.r_cs[0]$_SDFFE_PN1P__3527  (.L_HI(net3527));
 sg13g2_tiehi \cpu.spi.r_cs[1]$_SDFFE_PN1P__3528  (.L_HI(net3528));
 sg13g2_tiehi \cpu.spi.r_cs[2]$_SDFFE_PN1P__3529  (.L_HI(net3529));
 sg13g2_tiehi \cpu.spi.r_in[0]$_DFFE_PP__3530  (.L_HI(net3530));
 sg13g2_tiehi \cpu.spi.r_in[1]$_DFFE_PP__3531  (.L_HI(net3531));
 sg13g2_tiehi \cpu.spi.r_in[2]$_DFFE_PP__3532  (.L_HI(net3532));
 sg13g2_tiehi \cpu.spi.r_in[3]$_DFFE_PP__3533  (.L_HI(net3533));
 sg13g2_tiehi \cpu.spi.r_in[4]$_DFFE_PP__3534  (.L_HI(net3534));
 sg13g2_tiehi \cpu.spi.r_in[5]$_DFFE_PP__3535  (.L_HI(net3535));
 sg13g2_tiehi \cpu.spi.r_in[6]$_DFFE_PP__3536  (.L_HI(net3536));
 sg13g2_tiehi \cpu.spi.r_in[7]$_DFFE_PP__3537  (.L_HI(net3537));
 sg13g2_tiehi \cpu.spi.r_interrupt$_SDFFE_PN0P__3538  (.L_HI(net3538));
 sg13g2_tiehi \cpu.spi.r_mode[0][0]$_DFFE_PP__3539  (.L_HI(net3539));
 sg13g2_tiehi \cpu.spi.r_mode[0][1]$_DFFE_PP__3540  (.L_HI(net3540));
 sg13g2_tiehi \cpu.spi.r_mode[1][0]$_DFFE_PP__3541  (.L_HI(net3541));
 sg13g2_tiehi \cpu.spi.r_mode[1][1]$_DFFE_PP__3542  (.L_HI(net3542));
 sg13g2_tiehi \cpu.spi.r_mode[2][0]$_DFFE_PP__3543  (.L_HI(net3543));
 sg13g2_tiehi \cpu.spi.r_mode[2][1]$_DFFE_PP__3544  (.L_HI(net3544));
 sg13g2_tiehi \cpu.spi.r_out[0]$_DFFE_PP__3545  (.L_HI(net3545));
 sg13g2_tiehi \cpu.spi.r_out[1]$_DFFE_PP__3546  (.L_HI(net3546));
 sg13g2_tiehi \cpu.spi.r_out[2]$_DFFE_PP__3547  (.L_HI(net3547));
 sg13g2_tiehi \cpu.spi.r_out[3]$_DFFE_PP__3548  (.L_HI(net3548));
 sg13g2_tiehi \cpu.spi.r_out[4]$_DFFE_PP__3549  (.L_HI(net3549));
 sg13g2_tiehi \cpu.spi.r_out[5]$_DFFE_PP__3550  (.L_HI(net3550));
 sg13g2_tiehi \cpu.spi.r_out[6]$_DFFE_PP__3551  (.L_HI(net3551));
 sg13g2_tiehi \cpu.spi.r_out[7]$_DFFE_PP__3552  (.L_HI(net3552));
 sg13g2_tiehi \cpu.spi.r_ready$_SDFFE_PN1P__3553  (.L_HI(net3553));
 sg13g2_tiehi \cpu.spi.r_searching$_SDFFE_PN0P__3554  (.L_HI(net3554));
 sg13g2_tiehi \cpu.spi.r_sel[0]$_DFFE_PP__3555  (.L_HI(net3555));
 sg13g2_tiehi \cpu.spi.r_sel[1]$_DFFE_PP__3556  (.L_HI(net3556));
 sg13g2_tiehi \cpu.spi.r_src[0]$_DFFE_PP__3557  (.L_HI(net3557));
 sg13g2_tiehi \cpu.spi.r_src[1]$_DFFE_PP__3558  (.L_HI(net3558));
 sg13g2_tiehi \cpu.spi.r_src[2]$_DFFE_PP__3559  (.L_HI(net3559));
 sg13g2_tiehi \cpu.spi.r_state[0]$_DFF_P__3560  (.L_HI(net3560));
 sg13g2_tiehi \cpu.spi.r_state[1]$_DFF_P__3561  (.L_HI(net3561));
 sg13g2_tiehi \cpu.spi.r_state[2]$_DFF_P__3562  (.L_HI(net3562));
 sg13g2_tiehi \cpu.spi.r_state[3]$_DFF_P__3563  (.L_HI(net3563));
 sg13g2_tiehi \cpu.spi.r_state[4]$_DFF_P__3564  (.L_HI(net3564));
 sg13g2_tiehi \cpu.spi.r_state[5]$_DFF_P__3565  (.L_HI(net3565));
 sg13g2_tiehi \cpu.spi.r_state[6]$_DFF_P__3566  (.L_HI(net3566));
 sg13g2_tiehi \cpu.spi.r_timeout[0]$_DFFE_PP__3567  (.L_HI(net3567));
 sg13g2_tiehi \cpu.spi.r_timeout[1]$_DFFE_PP__3568  (.L_HI(net3568));
 sg13g2_tiehi \cpu.spi.r_timeout[2]$_DFFE_PP__3569  (.L_HI(net3569));
 sg13g2_tiehi \cpu.spi.r_timeout[3]$_DFFE_PP__3570  (.L_HI(net3570));
 sg13g2_tiehi \cpu.spi.r_timeout[4]$_DFFE_PP__3571  (.L_HI(net3571));
 sg13g2_tiehi \cpu.spi.r_timeout[5]$_DFFE_PP__3572  (.L_HI(net3572));
 sg13g2_tiehi \cpu.spi.r_timeout[6]$_DFFE_PP__3573  (.L_HI(net3573));
 sg13g2_tiehi \cpu.spi.r_timeout[7]$_DFFE_PP__3574  (.L_HI(net3574));
 sg13g2_tiehi \cpu.spi.r_timeout_count[0]$_DFFE_PP__3575  (.L_HI(net3575));
 sg13g2_tiehi \cpu.spi.r_timeout_count[1]$_DFFE_PP__3576  (.L_HI(net3576));
 sg13g2_tiehi \cpu.spi.r_timeout_count[2]$_DFFE_PP__3577  (.L_HI(net3577));
 sg13g2_tiehi \cpu.spi.r_timeout_count[3]$_DFFE_PP__3578  (.L_HI(net3578));
 sg13g2_tiehi \cpu.spi.r_timeout_count[4]$_DFFE_PP__3579  (.L_HI(net3579));
 sg13g2_tiehi \cpu.spi.r_timeout_count[5]$_DFFE_PP__3580  (.L_HI(net3580));
 sg13g2_tiehi \cpu.spi.r_timeout_count[6]$_DFFE_PP__3581  (.L_HI(net3581));
 sg13g2_tiehi \cpu.spi.r_timeout_count[7]$_DFFE_PP__3582  (.L_HI(net3582));
 sg13g2_tiehi \cpu.uart.r_div[0]$_DFF_P__3583  (.L_HI(net3583));
 sg13g2_tiehi \cpu.uart.r_div[10]$_DFF_P__3584  (.L_HI(net3584));
 sg13g2_tiehi \cpu.uart.r_div[11]$_DFF_P__3585  (.L_HI(net3585));
 sg13g2_tiehi \cpu.uart.r_div[1]$_DFF_P__3586  (.L_HI(net3586));
 sg13g2_tiehi \cpu.uart.r_div[2]$_DFF_P__3587  (.L_HI(net3587));
 sg13g2_tiehi \cpu.uart.r_div[3]$_DFF_P__3588  (.L_HI(net3588));
 sg13g2_tiehi \cpu.uart.r_div[4]$_DFF_P__3589  (.L_HI(net3589));
 sg13g2_tiehi \cpu.uart.r_div[5]$_DFF_P__3590  (.L_HI(net3590));
 sg13g2_tiehi \cpu.uart.r_div[6]$_DFF_P__3591  (.L_HI(net3591));
 sg13g2_tiehi \cpu.uart.r_div[7]$_DFF_P__3592  (.L_HI(net3592));
 sg13g2_tiehi \cpu.uart.r_div[8]$_DFF_P__3593  (.L_HI(net3593));
 sg13g2_tiehi \cpu.uart.r_div[9]$_DFF_P__3594  (.L_HI(net3594));
 sg13g2_tiehi \cpu.uart.r_div_value[0]$_SDFFE_PN1P__3595  (.L_HI(net3595));
 sg13g2_tiehi \cpu.uart.r_div_value[10]$_SDFFE_PN0P__3596  (.L_HI(net3596));
 sg13g2_tiehi \cpu.uart.r_div_value[11]$_SDFFE_PN0P__3597  (.L_HI(net3597));
 sg13g2_tiehi \cpu.uart.r_div_value[1]$_SDFFE_PN0P__3598  (.L_HI(net3598));
 sg13g2_tiehi \cpu.uart.r_div_value[2]$_SDFFE_PN0P__3599  (.L_HI(net3599));
 sg13g2_tiehi \cpu.uart.r_div_value[3]$_SDFFE_PN0P__3600  (.L_HI(net3600));
 sg13g2_tiehi \cpu.uart.r_div_value[4]$_SDFFE_PN0P__3601  (.L_HI(net3601));
 sg13g2_tiehi \cpu.uart.r_div_value[5]$_SDFFE_PN0P__3602  (.L_HI(net3602));
 sg13g2_tiehi \cpu.uart.r_div_value[6]$_SDFFE_PN0P__3603  (.L_HI(net3603));
 sg13g2_tiehi \cpu.uart.r_div_value[7]$_SDFFE_PN0P__3604  (.L_HI(net3604));
 sg13g2_tiehi \cpu.uart.r_div_value[8]$_SDFFE_PN0P__3605  (.L_HI(net3605));
 sg13g2_tiehi \cpu.uart.r_div_value[9]$_SDFFE_PN0P__3606  (.L_HI(net3606));
 sg13g2_tiehi \cpu.uart.r_ib[0]$_DFFE_PP__3607  (.L_HI(net3607));
 sg13g2_tiehi \cpu.uart.r_ib[1]$_DFFE_PP__3608  (.L_HI(net3608));
 sg13g2_tiehi \cpu.uart.r_ib[2]$_DFFE_PP__3609  (.L_HI(net3609));
 sg13g2_tiehi \cpu.uart.r_ib[3]$_DFFE_PP__3610  (.L_HI(net3610));
 sg13g2_tiehi \cpu.uart.r_ib[4]$_DFFE_PP__3611  (.L_HI(net3611));
 sg13g2_tiehi \cpu.uart.r_ib[5]$_DFFE_PP__3612  (.L_HI(net3612));
 sg13g2_tiehi \cpu.uart.r_ib[6]$_DFFE_PP__3613  (.L_HI(net3613));
 sg13g2_tiehi \cpu.uart.r_in[0]$_DFFE_PP__3614  (.L_HI(net3614));
 sg13g2_tiehi \cpu.uart.r_in[1]$_DFFE_PP__3615  (.L_HI(net3615));
 sg13g2_tiehi \cpu.uart.r_in[2]$_DFFE_PP__3616  (.L_HI(net3616));
 sg13g2_tiehi \cpu.uart.r_in[3]$_DFFE_PP__3617  (.L_HI(net3617));
 sg13g2_tiehi \cpu.uart.r_in[4]$_DFFE_PP__3618  (.L_HI(net3618));
 sg13g2_tiehi \cpu.uart.r_in[5]$_DFFE_PP__3619  (.L_HI(net3619));
 sg13g2_tiehi \cpu.uart.r_in[6]$_DFFE_PP__3620  (.L_HI(net3620));
 sg13g2_tiehi \cpu.uart.r_in[7]$_DFFE_PP__3621  (.L_HI(net3621));
 sg13g2_tiehi \cpu.uart.r_out[0]$_DFFE_PP__3622  (.L_HI(net3622));
 sg13g2_tiehi \cpu.uart.r_out[1]$_DFFE_PP__3623  (.L_HI(net3623));
 sg13g2_tiehi \cpu.uart.r_out[2]$_DFFE_PP__3624  (.L_HI(net3624));
 sg13g2_tiehi \cpu.uart.r_out[3]$_DFFE_PP__3625  (.L_HI(net3625));
 sg13g2_tiehi \cpu.uart.r_out[4]$_DFFE_PP__3626  (.L_HI(net3626));
 sg13g2_tiehi \cpu.uart.r_out[5]$_DFFE_PP__3627  (.L_HI(net3627));
 sg13g2_tiehi \cpu.uart.r_out[6]$_DFFE_PP__3628  (.L_HI(net3628));
 sg13g2_tiehi \cpu.uart.r_out[7]$_DFFE_PP__3629  (.L_HI(net3629));
 sg13g2_tiehi \cpu.uart.r_r$_DFF_P__3630  (.L_HI(net3630));
 sg13g2_tiehi \cpu.uart.r_r_int$_SDFFE_PN0P__3631  (.L_HI(net3631));
 sg13g2_tiehi \cpu.uart.r_r_invert$_SDFFE_PN0P__3632  (.L_HI(net3632));
 sg13g2_tiehi \cpu.uart.r_rcnt[0]$_DFFE_PP__3633  (.L_HI(net3633));
 sg13g2_tiehi \cpu.uart.r_rcnt[1]$_DFFE_PP__3634  (.L_HI(net3634));
 sg13g2_tiehi \cpu.uart.r_rstate[0]$_SDFFE_PN0P__3635  (.L_HI(net3635));
 sg13g2_tiehi \cpu.uart.r_rstate[1]$_SDFFE_PN0P__3636  (.L_HI(net3636));
 sg13g2_tiehi \cpu.uart.r_rstate[2]$_SDFFE_PN0P__3637  (.L_HI(net3637));
 sg13g2_tiehi \cpu.uart.r_rstate[3]$_SDFFE_PN0P__3638  (.L_HI(net3638));
 sg13g2_tiehi \cpu.uart.r_x$_DFFE_PP__3639  (.L_HI(net3639));
 sg13g2_tiehi \cpu.uart.r_x_int$_SDFFE_PN0P__3640  (.L_HI(net3640));
 sg13g2_tiehi \cpu.uart.r_x_invert$_SDFFE_PN0P__3641  (.L_HI(net3641));
 sg13g2_tiehi \cpu.uart.r_xcnt[0]$_DFFE_PP__3642  (.L_HI(net3642));
 sg13g2_tiehi \cpu.uart.r_xcnt[1]$_DFFE_PP__3643  (.L_HI(net3643));
 sg13g2_tiehi \cpu.uart.r_xstate[0]$_SDFFE_PN0P__3644  (.L_HI(net3644));
 sg13g2_tiehi \cpu.uart.r_xstate[1]$_SDFFE_PN0P__3645  (.L_HI(net3645));
 sg13g2_tiehi \cpu.uart.r_xstate[2]$_SDFFE_PN0P__3646  (.L_HI(net3646));
 sg13g2_tiehi \cpu.uart.r_xstate[3]$_SDFFE_PN0P__3647  (.L_HI(net3647));
 sg13g2_tiehi \r_reset$_DFF_P__3648  (.L_HI(net3648));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_55__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_63__leaf_clk));
 sg13g2_buf_16 clkload7 (.A(clknet_leaf_312_clk));
 sg13g2_inv_2 clkload8 (.A(clknet_leaf_253_clk));
 sg13g2_inv_4 clkload9 (.A(clknet_leaf_258_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_leaf_120_clk));
 sg13g2_inv_2 clkload11 (.A(clknet_leaf_178_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_119_clk));
 sg13g2_inv_2 clkload13 (.A(clknet_leaf_122_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00054_));
 sg13g2_antennanp ANTENNA_2 (.A(_00054_));
 sg13g2_antennanp ANTENNA_3 (.A(_00741_));
 sg13g2_antennanp ANTENNA_4 (.A(_00743_));
 sg13g2_antennanp ANTENNA_5 (.A(_00783_));
 sg13g2_antennanp ANTENNA_6 (.A(_00788_));
 sg13g2_antennanp ANTENNA_7 (.A(_00788_));
 sg13g2_antennanp ANTENNA_8 (.A(_00919_));
 sg13g2_antennanp ANTENNA_9 (.A(_01062_));
 sg13g2_antennanp ANTENNA_10 (.A(_02921_));
 sg13g2_antennanp ANTENNA_11 (.A(_02921_));
 sg13g2_antennanp ANTENNA_12 (.A(_02921_));
 sg13g2_antennanp ANTENNA_13 (.A(_02921_));
 sg13g2_antennanp ANTENNA_14 (.A(_02950_));
 sg13g2_antennanp ANTENNA_15 (.A(_02950_));
 sg13g2_antennanp ANTENNA_16 (.A(_02950_));
 sg13g2_antennanp ANTENNA_17 (.A(_02950_));
 sg13g2_antennanp ANTENNA_18 (.A(_03050_));
 sg13g2_antennanp ANTENNA_19 (.A(_03050_));
 sg13g2_antennanp ANTENNA_20 (.A(_03050_));
 sg13g2_antennanp ANTENNA_21 (.A(_03050_));
 sg13g2_antennanp ANTENNA_22 (.A(_03056_));
 sg13g2_antennanp ANTENNA_23 (.A(_03056_));
 sg13g2_antennanp ANTENNA_24 (.A(_03056_));
 sg13g2_antennanp ANTENNA_25 (.A(_03056_));
 sg13g2_antennanp ANTENNA_26 (.A(_03057_));
 sg13g2_antennanp ANTENNA_27 (.A(_03057_));
 sg13g2_antennanp ANTENNA_28 (.A(_03057_));
 sg13g2_antennanp ANTENNA_29 (.A(_03072_));
 sg13g2_antennanp ANTENNA_30 (.A(_03072_));
 sg13g2_antennanp ANTENNA_31 (.A(_03072_));
 sg13g2_antennanp ANTENNA_32 (.A(_03072_));
 sg13g2_antennanp ANTENNA_33 (.A(_03072_));
 sg13g2_antennanp ANTENNA_34 (.A(_03072_));
 sg13g2_antennanp ANTENNA_35 (.A(_03072_));
 sg13g2_antennanp ANTENNA_36 (.A(_03072_));
 sg13g2_antennanp ANTENNA_37 (.A(_03072_));
 sg13g2_antennanp ANTENNA_38 (.A(_03073_));
 sg13g2_antennanp ANTENNA_39 (.A(_03073_));
 sg13g2_antennanp ANTENNA_40 (.A(_03073_));
 sg13g2_antennanp ANTENNA_41 (.A(_03073_));
 sg13g2_antennanp ANTENNA_42 (.A(_03073_));
 sg13g2_antennanp ANTENNA_43 (.A(_03073_));
 sg13g2_antennanp ANTENNA_44 (.A(_03077_));
 sg13g2_antennanp ANTENNA_45 (.A(_03077_));
 sg13g2_antennanp ANTENNA_46 (.A(_03077_));
 sg13g2_antennanp ANTENNA_47 (.A(_03077_));
 sg13g2_antennanp ANTENNA_48 (.A(_03077_));
 sg13g2_antennanp ANTENNA_49 (.A(_03077_));
 sg13g2_antennanp ANTENNA_50 (.A(_03077_));
 sg13g2_antennanp ANTENNA_51 (.A(_03077_));
 sg13g2_antennanp ANTENNA_52 (.A(_03077_));
 sg13g2_antennanp ANTENNA_53 (.A(_03078_));
 sg13g2_antennanp ANTENNA_54 (.A(_03078_));
 sg13g2_antennanp ANTENNA_55 (.A(_03078_));
 sg13g2_antennanp ANTENNA_56 (.A(_03078_));
 sg13g2_antennanp ANTENNA_57 (.A(_03078_));
 sg13g2_antennanp ANTENNA_58 (.A(_03078_));
 sg13g2_antennanp ANTENNA_59 (.A(_03080_));
 sg13g2_antennanp ANTENNA_60 (.A(_03080_));
 sg13g2_antennanp ANTENNA_61 (.A(_03080_));
 sg13g2_antennanp ANTENNA_62 (.A(_03080_));
 sg13g2_antennanp ANTENNA_63 (.A(_03102_));
 sg13g2_antennanp ANTENNA_64 (.A(_03102_));
 sg13g2_antennanp ANTENNA_65 (.A(_03102_));
 sg13g2_antennanp ANTENNA_66 (.A(_03115_));
 sg13g2_antennanp ANTENNA_67 (.A(_03115_));
 sg13g2_antennanp ANTENNA_68 (.A(_03228_));
 sg13g2_antennanp ANTENNA_69 (.A(_03252_));
 sg13g2_antennanp ANTENNA_70 (.A(_03354_));
 sg13g2_antennanp ANTENNA_71 (.A(_03615_));
 sg13g2_antennanp ANTENNA_72 (.A(_03615_));
 sg13g2_antennanp ANTENNA_73 (.A(_03615_));
 sg13g2_antennanp ANTENNA_74 (.A(_03615_));
 sg13g2_antennanp ANTENNA_75 (.A(_03620_));
 sg13g2_antennanp ANTENNA_76 (.A(_03620_));
 sg13g2_antennanp ANTENNA_77 (.A(_03620_));
 sg13g2_antennanp ANTENNA_78 (.A(_03620_));
 sg13g2_antennanp ANTENNA_79 (.A(_03620_));
 sg13g2_antennanp ANTENNA_80 (.A(_03620_));
 sg13g2_antennanp ANTENNA_81 (.A(_03622_));
 sg13g2_antennanp ANTENNA_82 (.A(_03622_));
 sg13g2_antennanp ANTENNA_83 (.A(_03622_));
 sg13g2_antennanp ANTENNA_84 (.A(_03622_));
 sg13g2_antennanp ANTENNA_85 (.A(_03622_));
 sg13g2_antennanp ANTENNA_86 (.A(_03622_));
 sg13g2_antennanp ANTENNA_87 (.A(_03624_));
 sg13g2_antennanp ANTENNA_88 (.A(_03624_));
 sg13g2_antennanp ANTENNA_89 (.A(_03624_));
 sg13g2_antennanp ANTENNA_90 (.A(_03624_));
 sg13g2_antennanp ANTENNA_91 (.A(_03624_));
 sg13g2_antennanp ANTENNA_92 (.A(_03624_));
 sg13g2_antennanp ANTENNA_93 (.A(_03624_));
 sg13g2_antennanp ANTENNA_94 (.A(_03624_));
 sg13g2_antennanp ANTENNA_95 (.A(_03625_));
 sg13g2_antennanp ANTENNA_96 (.A(_03625_));
 sg13g2_antennanp ANTENNA_97 (.A(_03625_));
 sg13g2_antennanp ANTENNA_98 (.A(_03625_));
 sg13g2_antennanp ANTENNA_99 (.A(_04758_));
 sg13g2_antennanp ANTENNA_100 (.A(_04758_));
 sg13g2_antennanp ANTENNA_101 (.A(_04758_));
 sg13g2_antennanp ANTENNA_102 (.A(_04758_));
 sg13g2_antennanp ANTENNA_103 (.A(_05150_));
 sg13g2_antennanp ANTENNA_104 (.A(_05213_));
 sg13g2_antennanp ANTENNA_105 (.A(_05278_));
 sg13g2_antennanp ANTENNA_106 (.A(_05287_));
 sg13g2_antennanp ANTENNA_107 (.A(_05297_));
 sg13g2_antennanp ANTENNA_108 (.A(_05447_));
 sg13g2_antennanp ANTENNA_109 (.A(_05453_));
 sg13g2_antennanp ANTENNA_110 (.A(_05580_));
 sg13g2_antennanp ANTENNA_111 (.A(_05584_));
 sg13g2_antennanp ANTENNA_112 (.A(_05760_));
 sg13g2_antennanp ANTENNA_113 (.A(_05760_));
 sg13g2_antennanp ANTENNA_114 (.A(_05764_));
 sg13g2_antennanp ANTENNA_115 (.A(_05769_));
 sg13g2_antennanp ANTENNA_116 (.A(_05772_));
 sg13g2_antennanp ANTENNA_117 (.A(_05778_));
 sg13g2_antennanp ANTENNA_118 (.A(_05779_));
 sg13g2_antennanp ANTENNA_119 (.A(_05780_));
 sg13g2_antennanp ANTENNA_120 (.A(_05783_));
 sg13g2_antennanp ANTENNA_121 (.A(_05813_));
 sg13g2_antennanp ANTENNA_122 (.A(_05813_));
 sg13g2_antennanp ANTENNA_123 (.A(_05813_));
 sg13g2_antennanp ANTENNA_124 (.A(_05813_));
 sg13g2_antennanp ANTENNA_125 (.A(_05813_));
 sg13g2_antennanp ANTENNA_126 (.A(_05813_));
 sg13g2_antennanp ANTENNA_127 (.A(_06004_));
 sg13g2_antennanp ANTENNA_128 (.A(_06495_));
 sg13g2_antennanp ANTENNA_129 (.A(_06495_));
 sg13g2_antennanp ANTENNA_130 (.A(_06495_));
 sg13g2_antennanp ANTENNA_131 (.A(_06495_));
 sg13g2_antennanp ANTENNA_132 (.A(_06495_));
 sg13g2_antennanp ANTENNA_133 (.A(_06495_));
 sg13g2_antennanp ANTENNA_134 (.A(_06495_));
 sg13g2_antennanp ANTENNA_135 (.A(_06495_));
 sg13g2_antennanp ANTENNA_136 (.A(_06495_));
 sg13g2_antennanp ANTENNA_137 (.A(_06498_));
 sg13g2_antennanp ANTENNA_138 (.A(_06498_));
 sg13g2_antennanp ANTENNA_139 (.A(_06498_));
 sg13g2_antennanp ANTENNA_140 (.A(_06498_));
 sg13g2_antennanp ANTENNA_141 (.A(_06745_));
 sg13g2_antennanp ANTENNA_142 (.A(_06745_));
 sg13g2_antennanp ANTENNA_143 (.A(_06745_));
 sg13g2_antennanp ANTENNA_144 (.A(_07591_));
 sg13g2_antennanp ANTENNA_145 (.A(_07591_));
 sg13g2_antennanp ANTENNA_146 (.A(_07591_));
 sg13g2_antennanp ANTENNA_147 (.A(_07591_));
 sg13g2_antennanp ANTENNA_148 (.A(_08276_));
 sg13g2_antennanp ANTENNA_149 (.A(_08278_));
 sg13g2_antennanp ANTENNA_150 (.A(_08278_));
 sg13g2_antennanp ANTENNA_151 (.A(_08278_));
 sg13g2_antennanp ANTENNA_152 (.A(_08278_));
 sg13g2_antennanp ANTENNA_153 (.A(_08290_));
 sg13g2_antennanp ANTENNA_154 (.A(_08290_));
 sg13g2_antennanp ANTENNA_155 (.A(_08290_));
 sg13g2_antennanp ANTENNA_156 (.A(_08290_));
 sg13g2_antennanp ANTENNA_157 (.A(_08290_));
 sg13g2_antennanp ANTENNA_158 (.A(_08290_));
 sg13g2_antennanp ANTENNA_159 (.A(_08290_));
 sg13g2_antennanp ANTENNA_160 (.A(_08290_));
 sg13g2_antennanp ANTENNA_161 (.A(_08290_));
 sg13g2_antennanp ANTENNA_162 (.A(_08290_));
 sg13g2_antennanp ANTENNA_163 (.A(_08290_));
 sg13g2_antennanp ANTENNA_164 (.A(_08292_));
 sg13g2_antennanp ANTENNA_165 (.A(_08301_));
 sg13g2_antennanp ANTENNA_166 (.A(_08301_));
 sg13g2_antennanp ANTENNA_167 (.A(_08336_));
 sg13g2_antennanp ANTENNA_168 (.A(_08336_));
 sg13g2_antennanp ANTENNA_169 (.A(_08336_));
 sg13g2_antennanp ANTENNA_170 (.A(_08336_));
 sg13g2_antennanp ANTENNA_171 (.A(_08336_));
 sg13g2_antennanp ANTENNA_172 (.A(_08336_));
 sg13g2_antennanp ANTENNA_173 (.A(_08336_));
 sg13g2_antennanp ANTENNA_174 (.A(_08336_));
 sg13g2_antennanp ANTENNA_175 (.A(_08336_));
 sg13g2_antennanp ANTENNA_176 (.A(_08459_));
 sg13g2_antennanp ANTENNA_177 (.A(_08459_));
 sg13g2_antennanp ANTENNA_178 (.A(_08459_));
 sg13g2_antennanp ANTENNA_179 (.A(_08529_));
 sg13g2_antennanp ANTENNA_180 (.A(_08529_));
 sg13g2_antennanp ANTENNA_181 (.A(_08529_));
 sg13g2_antennanp ANTENNA_182 (.A(_08529_));
 sg13g2_antennanp ANTENNA_183 (.A(_08561_));
 sg13g2_antennanp ANTENNA_184 (.A(_08570_));
 sg13g2_antennanp ANTENNA_185 (.A(_08570_));
 sg13g2_antennanp ANTENNA_186 (.A(_08570_));
 sg13g2_antennanp ANTENNA_187 (.A(_08590_));
 sg13g2_antennanp ANTENNA_188 (.A(_08670_));
 sg13g2_antennanp ANTENNA_189 (.A(_08670_));
 sg13g2_antennanp ANTENNA_190 (.A(_08670_));
 sg13g2_antennanp ANTENNA_191 (.A(_08690_));
 sg13g2_antennanp ANTENNA_192 (.A(_08777_));
 sg13g2_antennanp ANTENNA_193 (.A(_08777_));
 sg13g2_antennanp ANTENNA_194 (.A(_08777_));
 sg13g2_antennanp ANTENNA_195 (.A(_08906_));
 sg13g2_antennanp ANTENNA_196 (.A(_08930_));
 sg13g2_antennanp ANTENNA_197 (.A(_08930_));
 sg13g2_antennanp ANTENNA_198 (.A(_08968_));
 sg13g2_antennanp ANTENNA_199 (.A(_08968_));
 sg13g2_antennanp ANTENNA_200 (.A(_09006_));
 sg13g2_antennanp ANTENNA_201 (.A(_09072_));
 sg13g2_antennanp ANTENNA_202 (.A(_09104_));
 sg13g2_antennanp ANTENNA_203 (.A(_09104_));
 sg13g2_antennanp ANTENNA_204 (.A(_09104_));
 sg13g2_antennanp ANTENNA_205 (.A(_09104_));
 sg13g2_antennanp ANTENNA_206 (.A(_09157_));
 sg13g2_antennanp ANTENNA_207 (.A(_09164_));
 sg13g2_antennanp ANTENNA_208 (.A(_09164_));
 sg13g2_antennanp ANTENNA_209 (.A(_09164_));
 sg13g2_antennanp ANTENNA_210 (.A(_09164_));
 sg13g2_antennanp ANTENNA_211 (.A(_09164_));
 sg13g2_antennanp ANTENNA_212 (.A(_09164_));
 sg13g2_antennanp ANTENNA_213 (.A(_09164_));
 sg13g2_antennanp ANTENNA_214 (.A(_09164_));
 sg13g2_antennanp ANTENNA_215 (.A(_09256_));
 sg13g2_antennanp ANTENNA_216 (.A(_09260_));
 sg13g2_antennanp ANTENNA_217 (.A(_09260_));
 sg13g2_antennanp ANTENNA_218 (.A(_09260_));
 sg13g2_antennanp ANTENNA_219 (.A(_09260_));
 sg13g2_antennanp ANTENNA_220 (.A(_09269_));
 sg13g2_antennanp ANTENNA_221 (.A(_09269_));
 sg13g2_antennanp ANTENNA_222 (.A(_09269_));
 sg13g2_antennanp ANTENNA_223 (.A(_09269_));
 sg13g2_antennanp ANTENNA_224 (.A(_09330_));
 sg13g2_antennanp ANTENNA_225 (.A(_09360_));
 sg13g2_antennanp ANTENNA_226 (.A(_09360_));
 sg13g2_antennanp ANTENNA_227 (.A(_09360_));
 sg13g2_antennanp ANTENNA_228 (.A(_09386_));
 sg13g2_antennanp ANTENNA_229 (.A(_09411_));
 sg13g2_antennanp ANTENNA_230 (.A(_09440_));
 sg13g2_antennanp ANTENNA_231 (.A(_09455_));
 sg13g2_antennanp ANTENNA_232 (.A(_09455_));
 sg13g2_antennanp ANTENNA_233 (.A(_09455_));
 sg13g2_antennanp ANTENNA_234 (.A(_09455_));
 sg13g2_antennanp ANTENNA_235 (.A(_09478_));
 sg13g2_antennanp ANTENNA_236 (.A(_09538_));
 sg13g2_antennanp ANTENNA_237 (.A(_09613_));
 sg13g2_antennanp ANTENNA_238 (.A(_09634_));
 sg13g2_antennanp ANTENNA_239 (.A(_09657_));
 sg13g2_antennanp ANTENNA_240 (.A(_09657_));
 sg13g2_antennanp ANTENNA_241 (.A(_09699_));
 sg13g2_antennanp ANTENNA_242 (.A(_09726_));
 sg13g2_antennanp ANTENNA_243 (.A(_09757_));
 sg13g2_antennanp ANTENNA_244 (.A(_09757_));
 sg13g2_antennanp ANTENNA_245 (.A(_09757_));
 sg13g2_antennanp ANTENNA_246 (.A(_09757_));
 sg13g2_antennanp ANTENNA_247 (.A(_09893_));
 sg13g2_antennanp ANTENNA_248 (.A(_09893_));
 sg13g2_antennanp ANTENNA_249 (.A(_09893_));
 sg13g2_antennanp ANTENNA_250 (.A(_09893_));
 sg13g2_antennanp ANTENNA_251 (.A(_09893_));
 sg13g2_antennanp ANTENNA_252 (.A(_09893_));
 sg13g2_antennanp ANTENNA_253 (.A(_10028_));
 sg13g2_antennanp ANTENNA_254 (.A(_10028_));
 sg13g2_antennanp ANTENNA_255 (.A(_10028_));
 sg13g2_antennanp ANTENNA_256 (.A(_10028_));
 sg13g2_antennanp ANTENNA_257 (.A(_10039_));
 sg13g2_antennanp ANTENNA_258 (.A(_10039_));
 sg13g2_antennanp ANTENNA_259 (.A(_10039_));
 sg13g2_antennanp ANTENNA_260 (.A(_10040_));
 sg13g2_antennanp ANTENNA_261 (.A(_10040_));
 sg13g2_antennanp ANTENNA_262 (.A(_10040_));
 sg13g2_antennanp ANTENNA_263 (.A(_10040_));
 sg13g2_antennanp ANTENNA_264 (.A(_10143_));
 sg13g2_antennanp ANTENNA_265 (.A(_10143_));
 sg13g2_antennanp ANTENNA_266 (.A(_10143_));
 sg13g2_antennanp ANTENNA_267 (.A(_10143_));
 sg13g2_antennanp ANTENNA_268 (.A(_10312_));
 sg13g2_antennanp ANTENNA_269 (.A(_10312_));
 sg13g2_antennanp ANTENNA_270 (.A(_10312_));
 sg13g2_antennanp ANTENNA_271 (.A(_10312_));
 sg13g2_antennanp ANTENNA_272 (.A(_10312_));
 sg13g2_antennanp ANTENNA_273 (.A(_10322_));
 sg13g2_antennanp ANTENNA_274 (.A(_10322_));
 sg13g2_antennanp ANTENNA_275 (.A(_10322_));
 sg13g2_antennanp ANTENNA_276 (.A(_10322_));
 sg13g2_antennanp ANTENNA_277 (.A(_10615_));
 sg13g2_antennanp ANTENNA_278 (.A(_10616_));
 sg13g2_antennanp ANTENNA_279 (.A(_10812_));
 sg13g2_antennanp ANTENNA_280 (.A(_10812_));
 sg13g2_antennanp ANTENNA_281 (.A(_10812_));
 sg13g2_antennanp ANTENNA_282 (.A(_10812_));
 sg13g2_antennanp ANTENNA_283 (.A(_10812_));
 sg13g2_antennanp ANTENNA_284 (.A(_10984_));
 sg13g2_antennanp ANTENNA_285 (.A(_10984_));
 sg13g2_antennanp ANTENNA_286 (.A(_10984_));
 sg13g2_antennanp ANTENNA_287 (.A(_10984_));
 sg13g2_antennanp ANTENNA_288 (.A(_10984_));
 sg13g2_antennanp ANTENNA_289 (.A(_10984_));
 sg13g2_antennanp ANTENNA_290 (.A(_10984_));
 sg13g2_antennanp ANTENNA_291 (.A(_11080_));
 sg13g2_antennanp ANTENNA_292 (.A(_11080_));
 sg13g2_antennanp ANTENNA_293 (.A(_11080_));
 sg13g2_antennanp ANTENNA_294 (.A(_11080_));
 sg13g2_antennanp ANTENNA_295 (.A(_11080_));
 sg13g2_antennanp ANTENNA_296 (.A(_11080_));
 sg13g2_antennanp ANTENNA_297 (.A(_11080_));
 sg13g2_antennanp ANTENNA_298 (.A(_11080_));
 sg13g2_antennanp ANTENNA_299 (.A(_11080_));
 sg13g2_antennanp ANTENNA_300 (.A(_12014_));
 sg13g2_antennanp ANTENNA_301 (.A(_12014_));
 sg13g2_antennanp ANTENNA_302 (.A(_12014_));
 sg13g2_antennanp ANTENNA_303 (.A(_12014_));
 sg13g2_antennanp ANTENNA_304 (.A(_12074_));
 sg13g2_antennanp ANTENNA_305 (.A(_12074_));
 sg13g2_antennanp ANTENNA_306 (.A(_12074_));
 sg13g2_antennanp ANTENNA_307 (.A(_12074_));
 sg13g2_antennanp ANTENNA_308 (.A(_12074_));
 sg13g2_antennanp ANTENNA_309 (.A(_12074_));
 sg13g2_antennanp ANTENNA_310 (.A(_12074_));
 sg13g2_antennanp ANTENNA_311 (.A(_12074_));
 sg13g2_antennanp ANTENNA_312 (.A(_12074_));
 sg13g2_antennanp ANTENNA_313 (.A(_12074_));
 sg13g2_antennanp ANTENNA_314 (.A(_12074_));
 sg13g2_antennanp ANTENNA_315 (.A(_12074_));
 sg13g2_antennanp ANTENNA_316 (.A(_12140_));
 sg13g2_antennanp ANTENNA_317 (.A(_12140_));
 sg13g2_antennanp ANTENNA_318 (.A(_12140_));
 sg13g2_antennanp ANTENNA_319 (.A(_12140_));
 sg13g2_antennanp ANTENNA_320 (.A(_12140_));
 sg13g2_antennanp ANTENNA_321 (.A(_12140_));
 sg13g2_antennanp ANTENNA_322 (.A(_12140_));
 sg13g2_antennanp ANTENNA_323 (.A(_12140_));
 sg13g2_antennanp ANTENNA_324 (.A(_12140_));
 sg13g2_antennanp ANTENNA_325 (.A(_12140_));
 sg13g2_antennanp ANTENNA_326 (.A(_12161_));
 sg13g2_antennanp ANTENNA_327 (.A(_12161_));
 sg13g2_antennanp ANTENNA_328 (.A(_12161_));
 sg13g2_antennanp ANTENNA_329 (.A(_12161_));
 sg13g2_antennanp ANTENNA_330 (.A(_12161_));
 sg13g2_antennanp ANTENNA_331 (.A(_12161_));
 sg13g2_antennanp ANTENNA_332 (.A(_12161_));
 sg13g2_antennanp ANTENNA_333 (.A(_12161_));
 sg13g2_antennanp ANTENNA_334 (.A(_12161_));
 sg13g2_antennanp ANTENNA_335 (.A(_12161_));
 sg13g2_antennanp ANTENNA_336 (.A(_12185_));
 sg13g2_antennanp ANTENNA_337 (.A(_12185_));
 sg13g2_antennanp ANTENNA_338 (.A(_12185_));
 sg13g2_antennanp ANTENNA_339 (.A(_12185_));
 sg13g2_antennanp ANTENNA_340 (.A(_12185_));
 sg13g2_antennanp ANTENNA_341 (.A(_12185_));
 sg13g2_antennanp ANTENNA_342 (.A(_12185_));
 sg13g2_antennanp ANTENNA_343 (.A(_12185_));
 sg13g2_antennanp ANTENNA_344 (.A(_12185_));
 sg13g2_antennanp ANTENNA_345 (.A(_12207_));
 sg13g2_antennanp ANTENNA_346 (.A(_12207_));
 sg13g2_antennanp ANTENNA_347 (.A(_12207_));
 sg13g2_antennanp ANTENNA_348 (.A(_12207_));
 sg13g2_antennanp ANTENNA_349 (.A(_12207_));
 sg13g2_antennanp ANTENNA_350 (.A(_12207_));
 sg13g2_antennanp ANTENNA_351 (.A(_12207_));
 sg13g2_antennanp ANTENNA_352 (.A(_12207_));
 sg13g2_antennanp ANTENNA_353 (.A(_12207_));
 sg13g2_antennanp ANTENNA_354 (.A(_12207_));
 sg13g2_antennanp ANTENNA_355 (.A(_12214_));
 sg13g2_antennanp ANTENNA_356 (.A(_12214_));
 sg13g2_antennanp ANTENNA_357 (.A(_12214_));
 sg13g2_antennanp ANTENNA_358 (.A(_12214_));
 sg13g2_antennanp ANTENNA_359 (.A(_12214_));
 sg13g2_antennanp ANTENNA_360 (.A(_12214_));
 sg13g2_antennanp ANTENNA_361 (.A(_12214_));
 sg13g2_antennanp ANTENNA_362 (.A(_12214_));
 sg13g2_antennanp ANTENNA_363 (.A(_12214_));
 sg13g2_antennanp ANTENNA_364 (.A(_12251_));
 sg13g2_antennanp ANTENNA_365 (.A(_12251_));
 sg13g2_antennanp ANTENNA_366 (.A(_12251_));
 sg13g2_antennanp ANTENNA_367 (.A(_12251_));
 sg13g2_antennanp ANTENNA_368 (.A(_12251_));
 sg13g2_antennanp ANTENNA_369 (.A(_12251_));
 sg13g2_antennanp ANTENNA_370 (.A(_12251_));
 sg13g2_antennanp ANTENNA_371 (.A(_12251_));
 sg13g2_antennanp ANTENNA_372 (.A(_12251_));
 sg13g2_antennanp ANTENNA_373 (.A(_12269_));
 sg13g2_antennanp ANTENNA_374 (.A(_12269_));
 sg13g2_antennanp ANTENNA_375 (.A(_12269_));
 sg13g2_antennanp ANTENNA_376 (.A(_12335_));
 sg13g2_antennanp ANTENNA_377 (.A(_12335_));
 sg13g2_antennanp ANTENNA_378 (.A(_12335_));
 sg13g2_antennanp ANTENNA_379 (.A(_12335_));
 sg13g2_antennanp ANTENNA_380 (.A(_12335_));
 sg13g2_antennanp ANTENNA_381 (.A(_12335_));
 sg13g2_antennanp ANTENNA_382 (.A(_12335_));
 sg13g2_antennanp ANTENNA_383 (.A(_12335_));
 sg13g2_antennanp ANTENNA_384 (.A(_12335_));
 sg13g2_antennanp ANTENNA_385 (.A(_12632_));
 sg13g2_antennanp ANTENNA_386 (.A(_12632_));
 sg13g2_antennanp ANTENNA_387 (.A(_12632_));
 sg13g2_antennanp ANTENNA_388 (.A(_12632_));
 sg13g2_antennanp ANTENNA_389 (.A(_12632_));
 sg13g2_antennanp ANTENNA_390 (.A(_12632_));
 sg13g2_antennanp ANTENNA_391 (.A(_12632_));
 sg13g2_antennanp ANTENNA_392 (.A(_12632_));
 sg13g2_antennanp ANTENNA_393 (.A(_12632_));
 sg13g2_antennanp ANTENNA_394 (.A(_12632_));
 sg13g2_antennanp ANTENNA_395 (.A(_12632_));
 sg13g2_antennanp ANTENNA_396 (.A(_12632_));
 sg13g2_antennanp ANTENNA_397 (.A(_12632_));
 sg13g2_antennanp ANTENNA_398 (.A(_12632_));
 sg13g2_antennanp ANTENNA_399 (.A(_12632_));
 sg13g2_antennanp ANTENNA_400 (.A(_12632_));
 sg13g2_antennanp ANTENNA_401 (.A(_12632_));
 sg13g2_antennanp ANTENNA_402 (.A(_12632_));
 sg13g2_antennanp ANTENNA_403 (.A(_12668_));
 sg13g2_antennanp ANTENNA_404 (.A(_12668_));
 sg13g2_antennanp ANTENNA_405 (.A(_12668_));
 sg13g2_antennanp ANTENNA_406 (.A(_12668_));
 sg13g2_antennanp ANTENNA_407 (.A(_12668_));
 sg13g2_antennanp ANTENNA_408 (.A(_12668_));
 sg13g2_antennanp ANTENNA_409 (.A(_12668_));
 sg13g2_antennanp ANTENNA_410 (.A(_12668_));
 sg13g2_antennanp ANTENNA_411 (.A(_12668_));
 sg13g2_antennanp ANTENNA_412 (.A(clk));
 sg13g2_antennanp ANTENNA_413 (.A(clk));
 sg13g2_antennanp ANTENNA_414 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_415 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_416 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_417 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_418 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_419 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_420 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_421 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_422 (.A(net3));
 sg13g2_antennanp ANTENNA_423 (.A(net3));
 sg13g2_antennanp ANTENNA_424 (.A(net3));
 sg13g2_antennanp ANTENNA_425 (.A(net11));
 sg13g2_antennanp ANTENNA_426 (.A(net11));
 sg13g2_antennanp ANTENNA_427 (.A(net11));
 sg13g2_antennanp ANTENNA_428 (.A(net12));
 sg13g2_antennanp ANTENNA_429 (.A(net12));
 sg13g2_antennanp ANTENNA_430 (.A(net12));
 sg13g2_antennanp ANTENNA_431 (.A(net13));
 sg13g2_antennanp ANTENNA_432 (.A(net13));
 sg13g2_antennanp ANTENNA_433 (.A(net13));
 sg13g2_antennanp ANTENNA_434 (.A(net14));
 sg13g2_antennanp ANTENNA_435 (.A(net14));
 sg13g2_antennanp ANTENNA_436 (.A(net14));
 sg13g2_antennanp ANTENNA_437 (.A(net131));
 sg13g2_antennanp ANTENNA_438 (.A(net131));
 sg13g2_antennanp ANTENNA_439 (.A(net131));
 sg13g2_antennanp ANTENNA_440 (.A(net131));
 sg13g2_antennanp ANTENNA_441 (.A(net131));
 sg13g2_antennanp ANTENNA_442 (.A(net131));
 sg13g2_antennanp ANTENNA_443 (.A(net131));
 sg13g2_antennanp ANTENNA_444 (.A(net131));
 sg13g2_antennanp ANTENNA_445 (.A(net131));
 sg13g2_antennanp ANTENNA_446 (.A(net467));
 sg13g2_antennanp ANTENNA_447 (.A(net467));
 sg13g2_antennanp ANTENNA_448 (.A(net467));
 sg13g2_antennanp ANTENNA_449 (.A(net467));
 sg13g2_antennanp ANTENNA_450 (.A(net467));
 sg13g2_antennanp ANTENNA_451 (.A(net467));
 sg13g2_antennanp ANTENNA_452 (.A(net467));
 sg13g2_antennanp ANTENNA_453 (.A(net467));
 sg13g2_antennanp ANTENNA_454 (.A(net467));
 sg13g2_antennanp ANTENNA_455 (.A(net533));
 sg13g2_antennanp ANTENNA_456 (.A(net533));
 sg13g2_antennanp ANTENNA_457 (.A(net533));
 sg13g2_antennanp ANTENNA_458 (.A(net533));
 sg13g2_antennanp ANTENNA_459 (.A(net533));
 sg13g2_antennanp ANTENNA_460 (.A(net533));
 sg13g2_antennanp ANTENNA_461 (.A(net533));
 sg13g2_antennanp ANTENNA_462 (.A(net533));
 sg13g2_antennanp ANTENNA_463 (.A(net533));
 sg13g2_antennanp ANTENNA_464 (.A(net533));
 sg13g2_antennanp ANTENNA_465 (.A(net533));
 sg13g2_antennanp ANTENNA_466 (.A(net533));
 sg13g2_antennanp ANTENNA_467 (.A(net533));
 sg13g2_antennanp ANTENNA_468 (.A(net583));
 sg13g2_antennanp ANTENNA_469 (.A(net583));
 sg13g2_antennanp ANTENNA_470 (.A(net583));
 sg13g2_antennanp ANTENNA_471 (.A(net583));
 sg13g2_antennanp ANTENNA_472 (.A(net583));
 sg13g2_antennanp ANTENNA_473 (.A(net583));
 sg13g2_antennanp ANTENNA_474 (.A(net583));
 sg13g2_antennanp ANTENNA_475 (.A(net583));
 sg13g2_antennanp ANTENNA_476 (.A(net616));
 sg13g2_antennanp ANTENNA_477 (.A(net616));
 sg13g2_antennanp ANTENNA_478 (.A(net616));
 sg13g2_antennanp ANTENNA_479 (.A(net616));
 sg13g2_antennanp ANTENNA_480 (.A(net616));
 sg13g2_antennanp ANTENNA_481 (.A(net616));
 sg13g2_antennanp ANTENNA_482 (.A(net616));
 sg13g2_antennanp ANTENNA_483 (.A(net616));
 sg13g2_antennanp ANTENNA_484 (.A(net616));
 sg13g2_antennanp ANTENNA_485 (.A(net616));
 sg13g2_antennanp ANTENNA_486 (.A(net616));
 sg13g2_antennanp ANTENNA_487 (.A(net616));
 sg13g2_antennanp ANTENNA_488 (.A(net616));
 sg13g2_antennanp ANTENNA_489 (.A(net616));
 sg13g2_antennanp ANTENNA_490 (.A(net680));
 sg13g2_antennanp ANTENNA_491 (.A(net680));
 sg13g2_antennanp ANTENNA_492 (.A(net680));
 sg13g2_antennanp ANTENNA_493 (.A(net680));
 sg13g2_antennanp ANTENNA_494 (.A(net680));
 sg13g2_antennanp ANTENNA_495 (.A(net680));
 sg13g2_antennanp ANTENNA_496 (.A(net680));
 sg13g2_antennanp ANTENNA_497 (.A(net680));
 sg13g2_antennanp ANTENNA_498 (.A(net680));
 sg13g2_antennanp ANTENNA_499 (.A(net680));
 sg13g2_antennanp ANTENNA_500 (.A(net680));
 sg13g2_antennanp ANTENNA_501 (.A(net680));
 sg13g2_antennanp ANTENNA_502 (.A(net680));
 sg13g2_antennanp ANTENNA_503 (.A(net680));
 sg13g2_antennanp ANTENNA_504 (.A(net680));
 sg13g2_antennanp ANTENNA_505 (.A(net702));
 sg13g2_antennanp ANTENNA_506 (.A(net702));
 sg13g2_antennanp ANTENNA_507 (.A(net702));
 sg13g2_antennanp ANTENNA_508 (.A(net702));
 sg13g2_antennanp ANTENNA_509 (.A(net702));
 sg13g2_antennanp ANTENNA_510 (.A(net702));
 sg13g2_antennanp ANTENNA_511 (.A(net702));
 sg13g2_antennanp ANTENNA_512 (.A(net702));
 sg13g2_antennanp ANTENNA_513 (.A(net702));
 sg13g2_antennanp ANTENNA_514 (.A(net749));
 sg13g2_antennanp ANTENNA_515 (.A(net749));
 sg13g2_antennanp ANTENNA_516 (.A(net749));
 sg13g2_antennanp ANTENNA_517 (.A(net749));
 sg13g2_antennanp ANTENNA_518 (.A(net749));
 sg13g2_antennanp ANTENNA_519 (.A(net749));
 sg13g2_antennanp ANTENNA_520 (.A(net749));
 sg13g2_antennanp ANTENNA_521 (.A(net749));
 sg13g2_antennanp ANTENNA_522 (.A(net749));
 sg13g2_antennanp ANTENNA_523 (.A(net875));
 sg13g2_antennanp ANTENNA_524 (.A(net875));
 sg13g2_antennanp ANTENNA_525 (.A(net875));
 sg13g2_antennanp ANTENNA_526 (.A(net875));
 sg13g2_antennanp ANTENNA_527 (.A(net875));
 sg13g2_antennanp ANTENNA_528 (.A(net875));
 sg13g2_antennanp ANTENNA_529 (.A(net875));
 sg13g2_antennanp ANTENNA_530 (.A(net875));
 sg13g2_antennanp ANTENNA_531 (.A(net875));
 sg13g2_antennanp ANTENNA_532 (.A(net882));
 sg13g2_antennanp ANTENNA_533 (.A(net882));
 sg13g2_antennanp ANTENNA_534 (.A(net882));
 sg13g2_antennanp ANTENNA_535 (.A(net882));
 sg13g2_antennanp ANTENNA_536 (.A(net882));
 sg13g2_antennanp ANTENNA_537 (.A(net882));
 sg13g2_antennanp ANTENNA_538 (.A(net882));
 sg13g2_antennanp ANTENNA_539 (.A(net882));
 sg13g2_antennanp ANTENNA_540 (.A(net882));
 sg13g2_antennanp ANTENNA_541 (.A(net883));
 sg13g2_antennanp ANTENNA_542 (.A(net883));
 sg13g2_antennanp ANTENNA_543 (.A(net883));
 sg13g2_antennanp ANTENNA_544 (.A(net883));
 sg13g2_antennanp ANTENNA_545 (.A(net883));
 sg13g2_antennanp ANTENNA_546 (.A(net883));
 sg13g2_antennanp ANTENNA_547 (.A(net883));
 sg13g2_antennanp ANTENNA_548 (.A(net883));
 sg13g2_antennanp ANTENNA_549 (.A(net883));
 sg13g2_antennanp ANTENNA_550 (.A(net890));
 sg13g2_antennanp ANTENNA_551 (.A(net890));
 sg13g2_antennanp ANTENNA_552 (.A(net890));
 sg13g2_antennanp ANTENNA_553 (.A(net890));
 sg13g2_antennanp ANTENNA_554 (.A(net890));
 sg13g2_antennanp ANTENNA_555 (.A(net890));
 sg13g2_antennanp ANTENNA_556 (.A(net890));
 sg13g2_antennanp ANTENNA_557 (.A(net890));
 sg13g2_antennanp ANTENNA_558 (.A(net890));
 sg13g2_antennanp ANTENNA_559 (.A(net890));
 sg13g2_antennanp ANTENNA_560 (.A(net890));
 sg13g2_antennanp ANTENNA_561 (.A(net929));
 sg13g2_antennanp ANTENNA_562 (.A(net929));
 sg13g2_antennanp ANTENNA_563 (.A(net929));
 sg13g2_antennanp ANTENNA_564 (.A(net929));
 sg13g2_antennanp ANTENNA_565 (.A(net929));
 sg13g2_antennanp ANTENNA_566 (.A(net929));
 sg13g2_antennanp ANTENNA_567 (.A(net929));
 sg13g2_antennanp ANTENNA_568 (.A(net929));
 sg13g2_antennanp ANTENNA_569 (.A(net929));
 sg13g2_antennanp ANTENNA_570 (.A(net929));
 sg13g2_antennanp ANTENNA_571 (.A(net929));
 sg13g2_antennanp ANTENNA_572 (.A(net929));
 sg13g2_antennanp ANTENNA_573 (.A(net929));
 sg13g2_antennanp ANTENNA_574 (.A(net929));
 sg13g2_antennanp ANTENNA_575 (.A(net929));
 sg13g2_antennanp ANTENNA_576 (.A(net929));
 sg13g2_antennanp ANTENNA_577 (.A(net929));
 sg13g2_antennanp ANTENNA_578 (.A(net929));
 sg13g2_antennanp ANTENNA_579 (.A(net929));
 sg13g2_antennanp ANTENNA_580 (.A(net929));
 sg13g2_antennanp ANTENNA_581 (.A(net942));
 sg13g2_antennanp ANTENNA_582 (.A(net942));
 sg13g2_antennanp ANTENNA_583 (.A(net942));
 sg13g2_antennanp ANTENNA_584 (.A(net942));
 sg13g2_antennanp ANTENNA_585 (.A(net942));
 sg13g2_antennanp ANTENNA_586 (.A(net942));
 sg13g2_antennanp ANTENNA_587 (.A(net942));
 sg13g2_antennanp ANTENNA_588 (.A(net942));
 sg13g2_antennanp ANTENNA_589 (.A(net993));
 sg13g2_antennanp ANTENNA_590 (.A(net993));
 sg13g2_antennanp ANTENNA_591 (.A(net993));
 sg13g2_antennanp ANTENNA_592 (.A(net993));
 sg13g2_antennanp ANTENNA_593 (.A(net993));
 sg13g2_antennanp ANTENNA_594 (.A(net993));
 sg13g2_antennanp ANTENNA_595 (.A(net993));
 sg13g2_antennanp ANTENNA_596 (.A(net993));
 sg13g2_antennanp ANTENNA_597 (.A(net993));
 sg13g2_antennanp ANTENNA_598 (.A(net1000));
 sg13g2_antennanp ANTENNA_599 (.A(net1000));
 sg13g2_antennanp ANTENNA_600 (.A(net1000));
 sg13g2_antennanp ANTENNA_601 (.A(net1000));
 sg13g2_antennanp ANTENNA_602 (.A(net1000));
 sg13g2_antennanp ANTENNA_603 (.A(net1000));
 sg13g2_antennanp ANTENNA_604 (.A(net1000));
 sg13g2_antennanp ANTENNA_605 (.A(net1000));
 sg13g2_antennanp ANTENNA_606 (.A(net1000));
 sg13g2_antennanp ANTENNA_607 (.A(net1000));
 sg13g2_antennanp ANTENNA_608 (.A(net1023));
 sg13g2_antennanp ANTENNA_609 (.A(net1023));
 sg13g2_antennanp ANTENNA_610 (.A(net1023));
 sg13g2_antennanp ANTENNA_611 (.A(net1023));
 sg13g2_antennanp ANTENNA_612 (.A(net1023));
 sg13g2_antennanp ANTENNA_613 (.A(net1023));
 sg13g2_antennanp ANTENNA_614 (.A(net1023));
 sg13g2_antennanp ANTENNA_615 (.A(net1023));
 sg13g2_antennanp ANTENNA_616 (.A(net1023));
 sg13g2_antennanp ANTENNA_617 (.A(net1023));
 sg13g2_antennanp ANTENNA_618 (.A(net1023));
 sg13g2_antennanp ANTENNA_619 (.A(net1023));
 sg13g2_antennanp ANTENNA_620 (.A(net1023));
 sg13g2_antennanp ANTENNA_621 (.A(net1023));
 sg13g2_antennanp ANTENNA_622 (.A(net1023));
 sg13g2_antennanp ANTENNA_623 (.A(net1023));
 sg13g2_antennanp ANTENNA_624 (.A(net1023));
 sg13g2_antennanp ANTENNA_625 (.A(net1023));
 sg13g2_antennanp ANTENNA_626 (.A(net1023));
 sg13g2_antennanp ANTENNA_627 (.A(net1023));
 sg13g2_antennanp ANTENNA_628 (.A(net1023));
 sg13g2_antennanp ANTENNA_629 (.A(net1023));
 sg13g2_antennanp ANTENNA_630 (.A(net1023));
 sg13g2_antennanp ANTENNA_631 (.A(net1023));
 sg13g2_antennanp ANTENNA_632 (.A(net1023));
 sg13g2_antennanp ANTENNA_633 (.A(net1023));
 sg13g2_antennanp ANTENNA_634 (.A(net1023));
 sg13g2_antennanp ANTENNA_635 (.A(net1023));
 sg13g2_antennanp ANTENNA_636 (.A(net1023));
 sg13g2_antennanp ANTENNA_637 (.A(net1023));
 sg13g2_antennanp ANTENNA_638 (.A(net1023));
 sg13g2_antennanp ANTENNA_639 (.A(net1023));
 sg13g2_antennanp ANTENNA_640 (.A(net1023));
 sg13g2_antennanp ANTENNA_641 (.A(net1023));
 sg13g2_antennanp ANTENNA_642 (.A(net1023));
 sg13g2_antennanp ANTENNA_643 (.A(net1023));
 sg13g2_antennanp ANTENNA_644 (.A(net1026));
 sg13g2_antennanp ANTENNA_645 (.A(net1026));
 sg13g2_antennanp ANTENNA_646 (.A(net1026));
 sg13g2_antennanp ANTENNA_647 (.A(net1026));
 sg13g2_antennanp ANTENNA_648 (.A(net1026));
 sg13g2_antennanp ANTENNA_649 (.A(net1026));
 sg13g2_antennanp ANTENNA_650 (.A(net1026));
 sg13g2_antennanp ANTENNA_651 (.A(net1026));
 sg13g2_antennanp ANTENNA_652 (.A(net1026));
 sg13g2_antennanp ANTENNA_653 (.A(net1026));
 sg13g2_antennanp ANTENNA_654 (.A(net1026));
 sg13g2_antennanp ANTENNA_655 (.A(net1026));
 sg13g2_antennanp ANTENNA_656 (.A(net1027));
 sg13g2_antennanp ANTENNA_657 (.A(net1027));
 sg13g2_antennanp ANTENNA_658 (.A(net1027));
 sg13g2_antennanp ANTENNA_659 (.A(net1027));
 sg13g2_antennanp ANTENNA_660 (.A(net1027));
 sg13g2_antennanp ANTENNA_661 (.A(net1027));
 sg13g2_antennanp ANTENNA_662 (.A(net1027));
 sg13g2_antennanp ANTENNA_663 (.A(net1027));
 sg13g2_antennanp ANTENNA_664 (.A(net1027));
 sg13g2_antennanp ANTENNA_665 (.A(net1027));
 sg13g2_antennanp ANTENNA_666 (.A(net1027));
 sg13g2_antennanp ANTENNA_667 (.A(net1027));
 sg13g2_antennanp ANTENNA_668 (.A(net1027));
 sg13g2_antennanp ANTENNA_669 (.A(net1027));
 sg13g2_antennanp ANTENNA_670 (.A(net1027));
 sg13g2_antennanp ANTENNA_671 (.A(net1027));
 sg13g2_antennanp ANTENNA_672 (.A(net1027));
 sg13g2_antennanp ANTENNA_673 (.A(net1027));
 sg13g2_antennanp ANTENNA_674 (.A(net1027));
 sg13g2_antennanp ANTENNA_675 (.A(net1027));
 sg13g2_antennanp ANTENNA_676 (.A(net1027));
 sg13g2_antennanp ANTENNA_677 (.A(net1108));
 sg13g2_antennanp ANTENNA_678 (.A(net1108));
 sg13g2_antennanp ANTENNA_679 (.A(net1108));
 sg13g2_antennanp ANTENNA_680 (.A(net1108));
 sg13g2_antennanp ANTENNA_681 (.A(net1108));
 sg13g2_antennanp ANTENNA_682 (.A(net1108));
 sg13g2_antennanp ANTENNA_683 (.A(net1108));
 sg13g2_antennanp ANTENNA_684 (.A(net1108));
 sg13g2_antennanp ANTENNA_685 (.A(net1108));
 sg13g2_antennanp ANTENNA_686 (.A(net1108));
 sg13g2_antennanp ANTENNA_687 (.A(net1108));
 sg13g2_antennanp ANTENNA_688 (.A(net1108));
 sg13g2_antennanp ANTENNA_689 (.A(net1108));
 sg13g2_antennanp ANTENNA_690 (.A(net1108));
 sg13g2_antennanp ANTENNA_691 (.A(net1108));
 sg13g2_antennanp ANTENNA_692 (.A(net1108));
 sg13g2_antennanp ANTENNA_693 (.A(net1108));
 sg13g2_antennanp ANTENNA_694 (.A(net1108));
 sg13g2_antennanp ANTENNA_695 (.A(net1108));
 sg13g2_antennanp ANTENNA_696 (.A(net1108));
 sg13g2_antennanp ANTENNA_697 (.A(net1108));
 sg13g2_antennanp ANTENNA_698 (.A(net1108));
 sg13g2_antennanp ANTENNA_699 (.A(net1108));
 sg13g2_antennanp ANTENNA_700 (.A(net1108));
 sg13g2_antennanp ANTENNA_701 (.A(net1109));
 sg13g2_antennanp ANTENNA_702 (.A(net1109));
 sg13g2_antennanp ANTENNA_703 (.A(net1109));
 sg13g2_antennanp ANTENNA_704 (.A(net1109));
 sg13g2_antennanp ANTENNA_705 (.A(net1109));
 sg13g2_antennanp ANTENNA_706 (.A(net1109));
 sg13g2_antennanp ANTENNA_707 (.A(net1109));
 sg13g2_antennanp ANTENNA_708 (.A(net1109));
 sg13g2_antennanp ANTENNA_709 (.A(net1109));
 sg13g2_antennanp ANTENNA_710 (.A(net1109));
 sg13g2_antennanp ANTENNA_711 (.A(net1109));
 sg13g2_antennanp ANTENNA_712 (.A(net1109));
 sg13g2_antennanp ANTENNA_713 (.A(net1109));
 sg13g2_antennanp ANTENNA_714 (.A(net1143));
 sg13g2_antennanp ANTENNA_715 (.A(net1143));
 sg13g2_antennanp ANTENNA_716 (.A(net1143));
 sg13g2_antennanp ANTENNA_717 (.A(net1143));
 sg13g2_antennanp ANTENNA_718 (.A(net1143));
 sg13g2_antennanp ANTENNA_719 (.A(net1143));
 sg13g2_antennanp ANTENNA_720 (.A(net1143));
 sg13g2_antennanp ANTENNA_721 (.A(net1143));
 sg13g2_antennanp ANTENNA_722 (.A(net1143));
 sg13g2_antennanp ANTENNA_723 (.A(net1154));
 sg13g2_antennanp ANTENNA_724 (.A(net1154));
 sg13g2_antennanp ANTENNA_725 (.A(net1154));
 sg13g2_antennanp ANTENNA_726 (.A(net1154));
 sg13g2_antennanp ANTENNA_727 (.A(net1154));
 sg13g2_antennanp ANTENNA_728 (.A(net1154));
 sg13g2_antennanp ANTENNA_729 (.A(net1154));
 sg13g2_antennanp ANTENNA_730 (.A(net1154));
 sg13g2_antennanp ANTENNA_731 (.A(net1154));
 sg13g2_antennanp ANTENNA_732 (.A(net1154));
 sg13g2_antennanp ANTENNA_733 (.A(net1154));
 sg13g2_antennanp ANTENNA_734 (.A(net1154));
 sg13g2_antennanp ANTENNA_735 (.A(net1154));
 sg13g2_antennanp ANTENNA_736 (.A(net1154));
 sg13g2_antennanp ANTENNA_737 (.A(net1166));
 sg13g2_antennanp ANTENNA_738 (.A(net1166));
 sg13g2_antennanp ANTENNA_739 (.A(net1166));
 sg13g2_antennanp ANTENNA_740 (.A(net1166));
 sg13g2_antennanp ANTENNA_741 (.A(net1166));
 sg13g2_antennanp ANTENNA_742 (.A(net1166));
 sg13g2_antennanp ANTENNA_743 (.A(net1166));
 sg13g2_antennanp ANTENNA_744 (.A(net1166));
 sg13g2_antennanp ANTENNA_745 (.A(net1166));
 sg13g2_antennanp ANTENNA_746 (.A(net1166));
 sg13g2_antennanp ANTENNA_747 (.A(net1166));
 sg13g2_antennanp ANTENNA_748 (.A(net1166));
 sg13g2_antennanp ANTENNA_749 (.A(_00741_));
 sg13g2_antennanp ANTENNA_750 (.A(_00743_));
 sg13g2_antennanp ANTENNA_751 (.A(_00783_));
 sg13g2_antennanp ANTENNA_752 (.A(_00788_));
 sg13g2_antennanp ANTENNA_753 (.A(_00788_));
 sg13g2_antennanp ANTENNA_754 (.A(_00919_));
 sg13g2_antennanp ANTENNA_755 (.A(_02921_));
 sg13g2_antennanp ANTENNA_756 (.A(_02921_));
 sg13g2_antennanp ANTENNA_757 (.A(_02921_));
 sg13g2_antennanp ANTENNA_758 (.A(_02921_));
 sg13g2_antennanp ANTENNA_759 (.A(_02950_));
 sg13g2_antennanp ANTENNA_760 (.A(_02950_));
 sg13g2_antennanp ANTENNA_761 (.A(_02950_));
 sg13g2_antennanp ANTENNA_762 (.A(_02950_));
 sg13g2_antennanp ANTENNA_763 (.A(_02950_));
 sg13g2_antennanp ANTENNA_764 (.A(_03050_));
 sg13g2_antennanp ANTENNA_765 (.A(_03050_));
 sg13g2_antennanp ANTENNA_766 (.A(_03050_));
 sg13g2_antennanp ANTENNA_767 (.A(_03050_));
 sg13g2_antennanp ANTENNA_768 (.A(_03056_));
 sg13g2_antennanp ANTENNA_769 (.A(_03056_));
 sg13g2_antennanp ANTENNA_770 (.A(_03056_));
 sg13g2_antennanp ANTENNA_771 (.A(_03056_));
 sg13g2_antennanp ANTENNA_772 (.A(_03072_));
 sg13g2_antennanp ANTENNA_773 (.A(_03072_));
 sg13g2_antennanp ANTENNA_774 (.A(_03072_));
 sg13g2_antennanp ANTENNA_775 (.A(_03072_));
 sg13g2_antennanp ANTENNA_776 (.A(_03073_));
 sg13g2_antennanp ANTENNA_777 (.A(_03073_));
 sg13g2_antennanp ANTENNA_778 (.A(_03073_));
 sg13g2_antennanp ANTENNA_779 (.A(_03073_));
 sg13g2_antennanp ANTENNA_780 (.A(_03077_));
 sg13g2_antennanp ANTENNA_781 (.A(_03077_));
 sg13g2_antennanp ANTENNA_782 (.A(_03077_));
 sg13g2_antennanp ANTENNA_783 (.A(_03077_));
 sg13g2_antennanp ANTENNA_784 (.A(_03077_));
 sg13g2_antennanp ANTENNA_785 (.A(_03077_));
 sg13g2_antennanp ANTENNA_786 (.A(_03077_));
 sg13g2_antennanp ANTENNA_787 (.A(_03077_));
 sg13g2_antennanp ANTENNA_788 (.A(_03077_));
 sg13g2_antennanp ANTENNA_789 (.A(_03078_));
 sg13g2_antennanp ANTENNA_790 (.A(_03078_));
 sg13g2_antennanp ANTENNA_791 (.A(_03078_));
 sg13g2_antennanp ANTENNA_792 (.A(_03078_));
 sg13g2_antennanp ANTENNA_793 (.A(_03078_));
 sg13g2_antennanp ANTENNA_794 (.A(_03078_));
 sg13g2_antennanp ANTENNA_795 (.A(_03080_));
 sg13g2_antennanp ANTENNA_796 (.A(_03080_));
 sg13g2_antennanp ANTENNA_797 (.A(_03080_));
 sg13g2_antennanp ANTENNA_798 (.A(_03080_));
 sg13g2_antennanp ANTENNA_799 (.A(_03102_));
 sg13g2_antennanp ANTENNA_800 (.A(_03102_));
 sg13g2_antennanp ANTENNA_801 (.A(_03102_));
 sg13g2_antennanp ANTENNA_802 (.A(_03115_));
 sg13g2_antennanp ANTENNA_803 (.A(_03115_));
 sg13g2_antennanp ANTENNA_804 (.A(_03228_));
 sg13g2_antennanp ANTENNA_805 (.A(_03252_));
 sg13g2_antennanp ANTENNA_806 (.A(_03354_));
 sg13g2_antennanp ANTENNA_807 (.A(_03615_));
 sg13g2_antennanp ANTENNA_808 (.A(_03615_));
 sg13g2_antennanp ANTENNA_809 (.A(_03615_));
 sg13g2_antennanp ANTENNA_810 (.A(_03615_));
 sg13g2_antennanp ANTENNA_811 (.A(_03620_));
 sg13g2_antennanp ANTENNA_812 (.A(_03620_));
 sg13g2_antennanp ANTENNA_813 (.A(_03620_));
 sg13g2_antennanp ANTENNA_814 (.A(_03620_));
 sg13g2_antennanp ANTENNA_815 (.A(_03620_));
 sg13g2_antennanp ANTENNA_816 (.A(_03620_));
 sg13g2_antennanp ANTENNA_817 (.A(_03624_));
 sg13g2_antennanp ANTENNA_818 (.A(_03624_));
 sg13g2_antennanp ANTENNA_819 (.A(_03624_));
 sg13g2_antennanp ANTENNA_820 (.A(_03624_));
 sg13g2_antennanp ANTENNA_821 (.A(_03624_));
 sg13g2_antennanp ANTENNA_822 (.A(_03624_));
 sg13g2_antennanp ANTENNA_823 (.A(_03624_));
 sg13g2_antennanp ANTENNA_824 (.A(_03624_));
 sg13g2_antennanp ANTENNA_825 (.A(_03625_));
 sg13g2_antennanp ANTENNA_826 (.A(_03625_));
 sg13g2_antennanp ANTENNA_827 (.A(_03625_));
 sg13g2_antennanp ANTENNA_828 (.A(_03625_));
 sg13g2_antennanp ANTENNA_829 (.A(_05213_));
 sg13g2_antennanp ANTENNA_830 (.A(_05278_));
 sg13g2_antennanp ANTENNA_831 (.A(_05287_));
 sg13g2_antennanp ANTENNA_832 (.A(_05297_));
 sg13g2_antennanp ANTENNA_833 (.A(_05297_));
 sg13g2_antennanp ANTENNA_834 (.A(_05447_));
 sg13g2_antennanp ANTENNA_835 (.A(_05453_));
 sg13g2_antennanp ANTENNA_836 (.A(_05453_));
 sg13g2_antennanp ANTENNA_837 (.A(_05580_));
 sg13g2_antennanp ANTENNA_838 (.A(_05584_));
 sg13g2_antennanp ANTENNA_839 (.A(_05760_));
 sg13g2_antennanp ANTENNA_840 (.A(_05760_));
 sg13g2_antennanp ANTENNA_841 (.A(_05764_));
 sg13g2_antennanp ANTENNA_842 (.A(_05769_));
 sg13g2_antennanp ANTENNA_843 (.A(_05772_));
 sg13g2_antennanp ANTENNA_844 (.A(_05778_));
 sg13g2_antennanp ANTENNA_845 (.A(_05779_));
 sg13g2_antennanp ANTENNA_846 (.A(_05780_));
 sg13g2_antennanp ANTENNA_847 (.A(_05783_));
 sg13g2_antennanp ANTENNA_848 (.A(_06004_));
 sg13g2_antennanp ANTENNA_849 (.A(_06495_));
 sg13g2_antennanp ANTENNA_850 (.A(_06495_));
 sg13g2_antennanp ANTENNA_851 (.A(_06495_));
 sg13g2_antennanp ANTENNA_852 (.A(_06495_));
 sg13g2_antennanp ANTENNA_853 (.A(_06495_));
 sg13g2_antennanp ANTENNA_854 (.A(_06495_));
 sg13g2_antennanp ANTENNA_855 (.A(_06495_));
 sg13g2_antennanp ANTENNA_856 (.A(_06495_));
 sg13g2_antennanp ANTENNA_857 (.A(_06495_));
 sg13g2_antennanp ANTENNA_858 (.A(_06498_));
 sg13g2_antennanp ANTENNA_859 (.A(_06498_));
 sg13g2_antennanp ANTENNA_860 (.A(_06498_));
 sg13g2_antennanp ANTENNA_861 (.A(_06498_));
 sg13g2_antennanp ANTENNA_862 (.A(_07528_));
 sg13g2_antennanp ANTENNA_863 (.A(_07528_));
 sg13g2_antennanp ANTENNA_864 (.A(_07528_));
 sg13g2_antennanp ANTENNA_865 (.A(_08276_));
 sg13g2_antennanp ANTENNA_866 (.A(_08290_));
 sg13g2_antennanp ANTENNA_867 (.A(_08290_));
 sg13g2_antennanp ANTENNA_868 (.A(_08290_));
 sg13g2_antennanp ANTENNA_869 (.A(_08290_));
 sg13g2_antennanp ANTENNA_870 (.A(_08290_));
 sg13g2_antennanp ANTENNA_871 (.A(_08292_));
 sg13g2_antennanp ANTENNA_872 (.A(_08301_));
 sg13g2_antennanp ANTENNA_873 (.A(_08301_));
 sg13g2_antennanp ANTENNA_874 (.A(_08301_));
 sg13g2_antennanp ANTENNA_875 (.A(_08336_));
 sg13g2_antennanp ANTENNA_876 (.A(_08336_));
 sg13g2_antennanp ANTENNA_877 (.A(_08336_));
 sg13g2_antennanp ANTENNA_878 (.A(_08336_));
 sg13g2_antennanp ANTENNA_879 (.A(_08336_));
 sg13g2_antennanp ANTENNA_880 (.A(_08336_));
 sg13g2_antennanp ANTENNA_881 (.A(_08336_));
 sg13g2_antennanp ANTENNA_882 (.A(_08336_));
 sg13g2_antennanp ANTENNA_883 (.A(_08336_));
 sg13g2_antennanp ANTENNA_884 (.A(_08459_));
 sg13g2_antennanp ANTENNA_885 (.A(_08459_));
 sg13g2_antennanp ANTENNA_886 (.A(_08459_));
 sg13g2_antennanp ANTENNA_887 (.A(_08529_));
 sg13g2_antennanp ANTENNA_888 (.A(_08529_));
 sg13g2_antennanp ANTENNA_889 (.A(_08529_));
 sg13g2_antennanp ANTENNA_890 (.A(_08529_));
 sg13g2_antennanp ANTENNA_891 (.A(_08561_));
 sg13g2_antennanp ANTENNA_892 (.A(_08570_));
 sg13g2_antennanp ANTENNA_893 (.A(_08570_));
 sg13g2_antennanp ANTENNA_894 (.A(_08570_));
 sg13g2_antennanp ANTENNA_895 (.A(_08590_));
 sg13g2_antennanp ANTENNA_896 (.A(_08690_));
 sg13g2_antennanp ANTENNA_897 (.A(_08777_));
 sg13g2_antennanp ANTENNA_898 (.A(_08777_));
 sg13g2_antennanp ANTENNA_899 (.A(_08777_));
 sg13g2_antennanp ANTENNA_900 (.A(_08906_));
 sg13g2_antennanp ANTENNA_901 (.A(_08930_));
 sg13g2_antennanp ANTENNA_902 (.A(_08930_));
 sg13g2_antennanp ANTENNA_903 (.A(_08968_));
 sg13g2_antennanp ANTENNA_904 (.A(_08968_));
 sg13g2_antennanp ANTENNA_905 (.A(_09006_));
 sg13g2_antennanp ANTENNA_906 (.A(_09072_));
 sg13g2_antennanp ANTENNA_907 (.A(_09104_));
 sg13g2_antennanp ANTENNA_908 (.A(_09104_));
 sg13g2_antennanp ANTENNA_909 (.A(_09104_));
 sg13g2_antennanp ANTENNA_910 (.A(_09104_));
 sg13g2_antennanp ANTENNA_911 (.A(_09157_));
 sg13g2_antennanp ANTENNA_912 (.A(_09164_));
 sg13g2_antennanp ANTENNA_913 (.A(_09164_));
 sg13g2_antennanp ANTENNA_914 (.A(_09164_));
 sg13g2_antennanp ANTENNA_915 (.A(_09164_));
 sg13g2_antennanp ANTENNA_916 (.A(_09164_));
 sg13g2_antennanp ANTENNA_917 (.A(_09164_));
 sg13g2_antennanp ANTENNA_918 (.A(_09164_));
 sg13g2_antennanp ANTENNA_919 (.A(_09164_));
 sg13g2_antennanp ANTENNA_920 (.A(_09164_));
 sg13g2_antennanp ANTENNA_921 (.A(_09164_));
 sg13g2_antennanp ANTENNA_922 (.A(_09164_));
 sg13g2_antennanp ANTENNA_923 (.A(_09164_));
 sg13g2_antennanp ANTENNA_924 (.A(_09164_));
 sg13g2_antennanp ANTENNA_925 (.A(_09164_));
 sg13g2_antennanp ANTENNA_926 (.A(_09164_));
 sg13g2_antennanp ANTENNA_927 (.A(_09164_));
 sg13g2_antennanp ANTENNA_928 (.A(_09164_));
 sg13g2_antennanp ANTENNA_929 (.A(_09164_));
 sg13g2_antennanp ANTENNA_930 (.A(_09164_));
 sg13g2_antennanp ANTENNA_931 (.A(_09164_));
 sg13g2_antennanp ANTENNA_932 (.A(_09164_));
 sg13g2_antennanp ANTENNA_933 (.A(_09164_));
 sg13g2_antennanp ANTENNA_934 (.A(_09164_));
 sg13g2_antennanp ANTENNA_935 (.A(_09164_));
 sg13g2_antennanp ANTENNA_936 (.A(_09164_));
 sg13g2_antennanp ANTENNA_937 (.A(_09164_));
 sg13g2_antennanp ANTENNA_938 (.A(_09164_));
 sg13g2_antennanp ANTENNA_939 (.A(_09164_));
 sg13g2_antennanp ANTENNA_940 (.A(_09164_));
 sg13g2_antennanp ANTENNA_941 (.A(_09164_));
 sg13g2_antennanp ANTENNA_942 (.A(_09260_));
 sg13g2_antennanp ANTENNA_943 (.A(_09260_));
 sg13g2_antennanp ANTENNA_944 (.A(_09260_));
 sg13g2_antennanp ANTENNA_945 (.A(_09260_));
 sg13g2_antennanp ANTENNA_946 (.A(_09269_));
 sg13g2_antennanp ANTENNA_947 (.A(_09269_));
 sg13g2_antennanp ANTENNA_948 (.A(_09269_));
 sg13g2_antennanp ANTENNA_949 (.A(_09269_));
 sg13g2_antennanp ANTENNA_950 (.A(_09330_));
 sg13g2_antennanp ANTENNA_951 (.A(_09330_));
 sg13g2_antennanp ANTENNA_952 (.A(_09330_));
 sg13g2_antennanp ANTENNA_953 (.A(_09360_));
 sg13g2_antennanp ANTENNA_954 (.A(_09360_));
 sg13g2_antennanp ANTENNA_955 (.A(_09360_));
 sg13g2_antennanp ANTENNA_956 (.A(_09386_));
 sg13g2_antennanp ANTENNA_957 (.A(_09386_));
 sg13g2_antennanp ANTENNA_958 (.A(_09411_));
 sg13g2_antennanp ANTENNA_959 (.A(_09440_));
 sg13g2_antennanp ANTENNA_960 (.A(_09455_));
 sg13g2_antennanp ANTENNA_961 (.A(_09455_));
 sg13g2_antennanp ANTENNA_962 (.A(_09455_));
 sg13g2_antennanp ANTENNA_963 (.A(_09455_));
 sg13g2_antennanp ANTENNA_964 (.A(_09478_));
 sg13g2_antennanp ANTENNA_965 (.A(_09538_));
 sg13g2_antennanp ANTENNA_966 (.A(_09613_));
 sg13g2_antennanp ANTENNA_967 (.A(_09634_));
 sg13g2_antennanp ANTENNA_968 (.A(_09657_));
 sg13g2_antennanp ANTENNA_969 (.A(_09657_));
 sg13g2_antennanp ANTENNA_970 (.A(_09699_));
 sg13g2_antennanp ANTENNA_971 (.A(_09726_));
 sg13g2_antennanp ANTENNA_972 (.A(_09726_));
 sg13g2_antennanp ANTENNA_973 (.A(_09757_));
 sg13g2_antennanp ANTENNA_974 (.A(_09757_));
 sg13g2_antennanp ANTENNA_975 (.A(_09757_));
 sg13g2_antennanp ANTENNA_976 (.A(_09893_));
 sg13g2_antennanp ANTENNA_977 (.A(_09893_));
 sg13g2_antennanp ANTENNA_978 (.A(_09893_));
 sg13g2_antennanp ANTENNA_979 (.A(_09893_));
 sg13g2_antennanp ANTENNA_980 (.A(_09893_));
 sg13g2_antennanp ANTENNA_981 (.A(_09893_));
 sg13g2_antennanp ANTENNA_982 (.A(_10322_));
 sg13g2_antennanp ANTENNA_983 (.A(_10322_));
 sg13g2_antennanp ANTENNA_984 (.A(_10322_));
 sg13g2_antennanp ANTENNA_985 (.A(_10322_));
 sg13g2_antennanp ANTENNA_986 (.A(_10616_));
 sg13g2_antennanp ANTENNA_987 (.A(_10984_));
 sg13g2_antennanp ANTENNA_988 (.A(_10984_));
 sg13g2_antennanp ANTENNA_989 (.A(_10984_));
 sg13g2_antennanp ANTENNA_990 (.A(_10984_));
 sg13g2_antennanp ANTENNA_991 (.A(_10984_));
 sg13g2_antennanp ANTENNA_992 (.A(_10984_));
 sg13g2_antennanp ANTENNA_993 (.A(_10984_));
 sg13g2_antennanp ANTENNA_994 (.A(_11080_));
 sg13g2_antennanp ANTENNA_995 (.A(_11080_));
 sg13g2_antennanp ANTENNA_996 (.A(_11080_));
 sg13g2_antennanp ANTENNA_997 (.A(_11080_));
 sg13g2_antennanp ANTENNA_998 (.A(_11080_));
 sg13g2_antennanp ANTENNA_999 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1000 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1001 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1002 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1003 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1004 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1005 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1006 (.A(_12014_));
 sg13g2_antennanp ANTENNA_1007 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1008 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1009 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1010 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1011 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1012 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1013 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1014 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1015 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1016 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1017 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1018 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1019 (.A(_12161_));
 sg13g2_antennanp ANTENNA_1020 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1021 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1022 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1023 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1024 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1025 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1026 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1027 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1028 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1029 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1030 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1031 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1032 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1033 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1034 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1035 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1036 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1037 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1038 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1039 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1040 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1041 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1042 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1043 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1044 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1045 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1046 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1047 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1048 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1049 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1050 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1051 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1052 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1053 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1054 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1055 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1056 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1057 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1058 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1059 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1060 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1061 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1062 (.A(_12269_));
 sg13g2_antennanp ANTENNA_1063 (.A(_12269_));
 sg13g2_antennanp ANTENNA_1064 (.A(_12269_));
 sg13g2_antennanp ANTENNA_1065 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1066 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1067 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1068 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1069 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1070 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1071 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1072 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1073 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1074 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1075 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1076 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1077 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1078 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1079 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1080 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1081 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1082 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1083 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1084 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1085 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1086 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1087 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1088 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1089 (.A(clk));
 sg13g2_antennanp ANTENNA_1090 (.A(clk));
 sg13g2_antennanp ANTENNA_1091 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1092 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1093 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1094 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_1095 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1096 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_1097 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1098 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1099 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1100 (.A(net3));
 sg13g2_antennanp ANTENNA_1101 (.A(net3));
 sg13g2_antennanp ANTENNA_1102 (.A(net3));
 sg13g2_antennanp ANTENNA_1103 (.A(net11));
 sg13g2_antennanp ANTENNA_1104 (.A(net11));
 sg13g2_antennanp ANTENNA_1105 (.A(net11));
 sg13g2_antennanp ANTENNA_1106 (.A(net12));
 sg13g2_antennanp ANTENNA_1107 (.A(net12));
 sg13g2_antennanp ANTENNA_1108 (.A(net12));
 sg13g2_antennanp ANTENNA_1109 (.A(net13));
 sg13g2_antennanp ANTENNA_1110 (.A(net13));
 sg13g2_antennanp ANTENNA_1111 (.A(net13));
 sg13g2_antennanp ANTENNA_1112 (.A(net14));
 sg13g2_antennanp ANTENNA_1113 (.A(net14));
 sg13g2_antennanp ANTENNA_1114 (.A(net14));
 sg13g2_antennanp ANTENNA_1115 (.A(net467));
 sg13g2_antennanp ANTENNA_1116 (.A(net467));
 sg13g2_antennanp ANTENNA_1117 (.A(net467));
 sg13g2_antennanp ANTENNA_1118 (.A(net467));
 sg13g2_antennanp ANTENNA_1119 (.A(net467));
 sg13g2_antennanp ANTENNA_1120 (.A(net467));
 sg13g2_antennanp ANTENNA_1121 (.A(net467));
 sg13g2_antennanp ANTENNA_1122 (.A(net467));
 sg13g2_antennanp ANTENNA_1123 (.A(net467));
 sg13g2_antennanp ANTENNA_1124 (.A(net533));
 sg13g2_antennanp ANTENNA_1125 (.A(net533));
 sg13g2_antennanp ANTENNA_1126 (.A(net533));
 sg13g2_antennanp ANTENNA_1127 (.A(net533));
 sg13g2_antennanp ANTENNA_1128 (.A(net533));
 sg13g2_antennanp ANTENNA_1129 (.A(net533));
 sg13g2_antennanp ANTENNA_1130 (.A(net533));
 sg13g2_antennanp ANTENNA_1131 (.A(net533));
 sg13g2_antennanp ANTENNA_1132 (.A(net533));
 sg13g2_antennanp ANTENNA_1133 (.A(net533));
 sg13g2_antennanp ANTENNA_1134 (.A(net533));
 sg13g2_antennanp ANTENNA_1135 (.A(net533));
 sg13g2_antennanp ANTENNA_1136 (.A(net533));
 sg13g2_antennanp ANTENNA_1137 (.A(net533));
 sg13g2_antennanp ANTENNA_1138 (.A(net533));
 sg13g2_antennanp ANTENNA_1139 (.A(net533));
 sg13g2_antennanp ANTENNA_1140 (.A(net616));
 sg13g2_antennanp ANTENNA_1141 (.A(net616));
 sg13g2_antennanp ANTENNA_1142 (.A(net616));
 sg13g2_antennanp ANTENNA_1143 (.A(net616));
 sg13g2_antennanp ANTENNA_1144 (.A(net616));
 sg13g2_antennanp ANTENNA_1145 (.A(net616));
 sg13g2_antennanp ANTENNA_1146 (.A(net616));
 sg13g2_antennanp ANTENNA_1147 (.A(net616));
 sg13g2_antennanp ANTENNA_1148 (.A(net616));
 sg13g2_antennanp ANTENNA_1149 (.A(net616));
 sg13g2_antennanp ANTENNA_1150 (.A(net616));
 sg13g2_antennanp ANTENNA_1151 (.A(net616));
 sg13g2_antennanp ANTENNA_1152 (.A(net616));
 sg13g2_antennanp ANTENNA_1153 (.A(net616));
 sg13g2_antennanp ANTENNA_1154 (.A(net680));
 sg13g2_antennanp ANTENNA_1155 (.A(net680));
 sg13g2_antennanp ANTENNA_1156 (.A(net680));
 sg13g2_antennanp ANTENNA_1157 (.A(net680));
 sg13g2_antennanp ANTENNA_1158 (.A(net680));
 sg13g2_antennanp ANTENNA_1159 (.A(net680));
 sg13g2_antennanp ANTENNA_1160 (.A(net680));
 sg13g2_antennanp ANTENNA_1161 (.A(net680));
 sg13g2_antennanp ANTENNA_1162 (.A(net702));
 sg13g2_antennanp ANTENNA_1163 (.A(net702));
 sg13g2_antennanp ANTENNA_1164 (.A(net702));
 sg13g2_antennanp ANTENNA_1165 (.A(net702));
 sg13g2_antennanp ANTENNA_1166 (.A(net702));
 sg13g2_antennanp ANTENNA_1167 (.A(net702));
 sg13g2_antennanp ANTENNA_1168 (.A(net702));
 sg13g2_antennanp ANTENNA_1169 (.A(net702));
 sg13g2_antennanp ANTENNA_1170 (.A(net702));
 sg13g2_antennanp ANTENNA_1171 (.A(net749));
 sg13g2_antennanp ANTENNA_1172 (.A(net749));
 sg13g2_antennanp ANTENNA_1173 (.A(net749));
 sg13g2_antennanp ANTENNA_1174 (.A(net749));
 sg13g2_antennanp ANTENNA_1175 (.A(net749));
 sg13g2_antennanp ANTENNA_1176 (.A(net749));
 sg13g2_antennanp ANTENNA_1177 (.A(net749));
 sg13g2_antennanp ANTENNA_1178 (.A(net749));
 sg13g2_antennanp ANTENNA_1179 (.A(net749));
 sg13g2_antennanp ANTENNA_1180 (.A(net882));
 sg13g2_antennanp ANTENNA_1181 (.A(net882));
 sg13g2_antennanp ANTENNA_1182 (.A(net882));
 sg13g2_antennanp ANTENNA_1183 (.A(net882));
 sg13g2_antennanp ANTENNA_1184 (.A(net882));
 sg13g2_antennanp ANTENNA_1185 (.A(net882));
 sg13g2_antennanp ANTENNA_1186 (.A(net882));
 sg13g2_antennanp ANTENNA_1187 (.A(net882));
 sg13g2_antennanp ANTENNA_1188 (.A(net882));
 sg13g2_antennanp ANTENNA_1189 (.A(net884));
 sg13g2_antennanp ANTENNA_1190 (.A(net884));
 sg13g2_antennanp ANTENNA_1191 (.A(net884));
 sg13g2_antennanp ANTENNA_1192 (.A(net884));
 sg13g2_antennanp ANTENNA_1193 (.A(net884));
 sg13g2_antennanp ANTENNA_1194 (.A(net884));
 sg13g2_antennanp ANTENNA_1195 (.A(net884));
 sg13g2_antennanp ANTENNA_1196 (.A(net884));
 sg13g2_antennanp ANTENNA_1197 (.A(net884));
 sg13g2_antennanp ANTENNA_1198 (.A(net929));
 sg13g2_antennanp ANTENNA_1199 (.A(net929));
 sg13g2_antennanp ANTENNA_1200 (.A(net929));
 sg13g2_antennanp ANTENNA_1201 (.A(net929));
 sg13g2_antennanp ANTENNA_1202 (.A(net929));
 sg13g2_antennanp ANTENNA_1203 (.A(net929));
 sg13g2_antennanp ANTENNA_1204 (.A(net929));
 sg13g2_antennanp ANTENNA_1205 (.A(net929));
 sg13g2_antennanp ANTENNA_1206 (.A(net929));
 sg13g2_antennanp ANTENNA_1207 (.A(net929));
 sg13g2_antennanp ANTENNA_1208 (.A(net929));
 sg13g2_antennanp ANTENNA_1209 (.A(net929));
 sg13g2_antennanp ANTENNA_1210 (.A(net929));
 sg13g2_antennanp ANTENNA_1211 (.A(net929));
 sg13g2_antennanp ANTENNA_1212 (.A(net929));
 sg13g2_antennanp ANTENNA_1213 (.A(net929));
 sg13g2_antennanp ANTENNA_1214 (.A(net929));
 sg13g2_antennanp ANTENNA_1215 (.A(net929));
 sg13g2_antennanp ANTENNA_1216 (.A(net929));
 sg13g2_antennanp ANTENNA_1217 (.A(net929));
 sg13g2_antennanp ANTENNA_1218 (.A(net942));
 sg13g2_antennanp ANTENNA_1219 (.A(net942));
 sg13g2_antennanp ANTENNA_1220 (.A(net942));
 sg13g2_antennanp ANTENNA_1221 (.A(net942));
 sg13g2_antennanp ANTENNA_1222 (.A(net942));
 sg13g2_antennanp ANTENNA_1223 (.A(net942));
 sg13g2_antennanp ANTENNA_1224 (.A(net942));
 sg13g2_antennanp ANTENNA_1225 (.A(net942));
 sg13g2_antennanp ANTENNA_1226 (.A(net1000));
 sg13g2_antennanp ANTENNA_1227 (.A(net1000));
 sg13g2_antennanp ANTENNA_1228 (.A(net1000));
 sg13g2_antennanp ANTENNA_1229 (.A(net1000));
 sg13g2_antennanp ANTENNA_1230 (.A(net1000));
 sg13g2_antennanp ANTENNA_1231 (.A(net1000));
 sg13g2_antennanp ANTENNA_1232 (.A(net1000));
 sg13g2_antennanp ANTENNA_1233 (.A(net1000));
 sg13g2_antennanp ANTENNA_1234 (.A(net1000));
 sg13g2_antennanp ANTENNA_1235 (.A(net1000));
 sg13g2_antennanp ANTENNA_1236 (.A(net1000));
 sg13g2_antennanp ANTENNA_1237 (.A(net1000));
 sg13g2_antennanp ANTENNA_1238 (.A(net1000));
 sg13g2_antennanp ANTENNA_1239 (.A(net1000));
 sg13g2_antennanp ANTENNA_1240 (.A(net1000));
 sg13g2_antennanp ANTENNA_1241 (.A(net1000));
 sg13g2_antennanp ANTENNA_1242 (.A(net1000));
 sg13g2_antennanp ANTENNA_1243 (.A(net1000));
 sg13g2_antennanp ANTENNA_1244 (.A(net1000));
 sg13g2_antennanp ANTENNA_1245 (.A(net1000));
 sg13g2_antennanp ANTENNA_1246 (.A(net1027));
 sg13g2_antennanp ANTENNA_1247 (.A(net1027));
 sg13g2_antennanp ANTENNA_1248 (.A(net1027));
 sg13g2_antennanp ANTENNA_1249 (.A(net1027));
 sg13g2_antennanp ANTENNA_1250 (.A(net1027));
 sg13g2_antennanp ANTENNA_1251 (.A(net1027));
 sg13g2_antennanp ANTENNA_1252 (.A(net1027));
 sg13g2_antennanp ANTENNA_1253 (.A(net1027));
 sg13g2_antennanp ANTENNA_1254 (.A(net1071));
 sg13g2_antennanp ANTENNA_1255 (.A(net1071));
 sg13g2_antennanp ANTENNA_1256 (.A(net1071));
 sg13g2_antennanp ANTENNA_1257 (.A(net1071));
 sg13g2_antennanp ANTENNA_1258 (.A(net1071));
 sg13g2_antennanp ANTENNA_1259 (.A(net1071));
 sg13g2_antennanp ANTENNA_1260 (.A(net1071));
 sg13g2_antennanp ANTENNA_1261 (.A(net1071));
 sg13g2_antennanp ANTENNA_1262 (.A(net1071));
 sg13g2_antennanp ANTENNA_1263 (.A(net1071));
 sg13g2_antennanp ANTENNA_1264 (.A(net1071));
 sg13g2_antennanp ANTENNA_1265 (.A(net1071));
 sg13g2_antennanp ANTENNA_1266 (.A(net1071));
 sg13g2_antennanp ANTENNA_1267 (.A(net1071));
 sg13g2_antennanp ANTENNA_1268 (.A(net1135));
 sg13g2_antennanp ANTENNA_1269 (.A(net1135));
 sg13g2_antennanp ANTENNA_1270 (.A(net1135));
 sg13g2_antennanp ANTENNA_1271 (.A(net1135));
 sg13g2_antennanp ANTENNA_1272 (.A(net1135));
 sg13g2_antennanp ANTENNA_1273 (.A(net1135));
 sg13g2_antennanp ANTENNA_1274 (.A(net1135));
 sg13g2_antennanp ANTENNA_1275 (.A(net1135));
 sg13g2_antennanp ANTENNA_1276 (.A(net1143));
 sg13g2_antennanp ANTENNA_1277 (.A(net1143));
 sg13g2_antennanp ANTENNA_1278 (.A(net1143));
 sg13g2_antennanp ANTENNA_1279 (.A(net1143));
 sg13g2_antennanp ANTENNA_1280 (.A(net1143));
 sg13g2_antennanp ANTENNA_1281 (.A(net1143));
 sg13g2_antennanp ANTENNA_1282 (.A(net1143));
 sg13g2_antennanp ANTENNA_1283 (.A(net1143));
 sg13g2_antennanp ANTENNA_1284 (.A(net1143));
 sg13g2_antennanp ANTENNA_1285 (.A(net1166));
 sg13g2_antennanp ANTENNA_1286 (.A(net1166));
 sg13g2_antennanp ANTENNA_1287 (.A(net1166));
 sg13g2_antennanp ANTENNA_1288 (.A(net1166));
 sg13g2_antennanp ANTENNA_1289 (.A(net1166));
 sg13g2_antennanp ANTENNA_1290 (.A(net1166));
 sg13g2_antennanp ANTENNA_1291 (.A(net1166));
 sg13g2_antennanp ANTENNA_1292 (.A(net1166));
 sg13g2_antennanp ANTENNA_1293 (.A(net1166));
 sg13g2_antennanp ANTENNA_1294 (.A(_00741_));
 sg13g2_antennanp ANTENNA_1295 (.A(_00743_));
 sg13g2_antennanp ANTENNA_1296 (.A(_00783_));
 sg13g2_antennanp ANTENNA_1297 (.A(_00919_));
 sg13g2_antennanp ANTENNA_1298 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1299 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1300 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1301 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1302 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1303 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1304 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1305 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1306 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1307 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1308 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1309 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1310 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1311 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1312 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1313 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1314 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1315 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1316 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1317 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1318 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1319 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1320 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1321 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1322 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1323 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1324 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1325 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1326 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1327 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1328 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1329 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1330 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1331 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1332 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1333 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1334 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1335 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1336 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1337 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1338 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1339 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1340 (.A(_03078_));
 sg13g2_antennanp ANTENNA_1341 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1342 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1343 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1344 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1345 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1346 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1347 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1348 (.A(_03115_));
 sg13g2_antennanp ANTENNA_1349 (.A(_03228_));
 sg13g2_antennanp ANTENNA_1350 (.A(_03252_));
 sg13g2_antennanp ANTENNA_1351 (.A(_03354_));
 sg13g2_antennanp ANTENNA_1352 (.A(_03615_));
 sg13g2_antennanp ANTENNA_1353 (.A(_03615_));
 sg13g2_antennanp ANTENNA_1354 (.A(_03615_));
 sg13g2_antennanp ANTENNA_1355 (.A(_03615_));
 sg13g2_antennanp ANTENNA_1356 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1357 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1358 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1359 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1360 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1361 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1362 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1363 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1364 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1365 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1366 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1367 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1368 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1369 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1370 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1371 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1372 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1373 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1374 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1375 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1376 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1377 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1378 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1379 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1380 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1381 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1382 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1383 (.A(_05213_));
 sg13g2_antennanp ANTENNA_1384 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1385 (.A(_05287_));
 sg13g2_antennanp ANTENNA_1386 (.A(_05297_));
 sg13g2_antennanp ANTENNA_1387 (.A(_05447_));
 sg13g2_antennanp ANTENNA_1388 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1389 (.A(_05580_));
 sg13g2_antennanp ANTENNA_1390 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1391 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1392 (.A(_05764_));
 sg13g2_antennanp ANTENNA_1393 (.A(_05764_));
 sg13g2_antennanp ANTENNA_1394 (.A(_05769_));
 sg13g2_antennanp ANTENNA_1395 (.A(_05772_));
 sg13g2_antennanp ANTENNA_1396 (.A(_05778_));
 sg13g2_antennanp ANTENNA_1397 (.A(_05779_));
 sg13g2_antennanp ANTENNA_1398 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1399 (.A(_05783_));
 sg13g2_antennanp ANTENNA_1400 (.A(_06004_));
 sg13g2_antennanp ANTENNA_1401 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1402 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1403 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1404 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1405 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1406 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1407 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1408 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1409 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1410 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1411 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1412 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1413 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1414 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1415 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1416 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1417 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1418 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1419 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1420 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1421 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1422 (.A(_08276_));
 sg13g2_antennanp ANTENNA_1423 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1424 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1425 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1426 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1427 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1428 (.A(_08292_));
 sg13g2_antennanp ANTENNA_1429 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1430 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1431 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1432 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1433 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1434 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1435 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1436 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1437 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1438 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1439 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1440 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1441 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1442 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1443 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1444 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1445 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1446 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1447 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1448 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1449 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1450 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1451 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1452 (.A(_08561_));
 sg13g2_antennanp ANTENNA_1453 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1454 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1455 (.A(_08570_));
 sg13g2_antennanp ANTENNA_1456 (.A(_08590_));
 sg13g2_antennanp ANTENNA_1457 (.A(_08690_));
 sg13g2_antennanp ANTENNA_1458 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1459 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1460 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1461 (.A(_08906_));
 sg13g2_antennanp ANTENNA_1462 (.A(_08906_));
 sg13g2_antennanp ANTENNA_1463 (.A(_08930_));
 sg13g2_antennanp ANTENNA_1464 (.A(_08930_));
 sg13g2_antennanp ANTENNA_1465 (.A(_08968_));
 sg13g2_antennanp ANTENNA_1466 (.A(_08968_));
 sg13g2_antennanp ANTENNA_1467 (.A(_09006_));
 sg13g2_antennanp ANTENNA_1468 (.A(_09072_));
 sg13g2_antennanp ANTENNA_1469 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1470 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1471 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1472 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1473 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1474 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1475 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1476 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1477 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1478 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1479 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1480 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1481 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1482 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1483 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1484 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1485 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1486 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1487 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1488 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1489 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1490 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1491 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1492 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1493 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1494 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1495 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1496 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1497 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1498 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1499 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1500 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1501 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1502 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1503 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1504 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1505 (.A(_09330_));
 sg13g2_antennanp ANTENNA_1506 (.A(_09330_));
 sg13g2_antennanp ANTENNA_1507 (.A(_09330_));
 sg13g2_antennanp ANTENNA_1508 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1509 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1510 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1511 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1512 (.A(_09411_));
 sg13g2_antennanp ANTENNA_1513 (.A(_09440_));
 sg13g2_antennanp ANTENNA_1514 (.A(_09455_));
 sg13g2_antennanp ANTENNA_1515 (.A(_09455_));
 sg13g2_antennanp ANTENNA_1516 (.A(_09455_));
 sg13g2_antennanp ANTENNA_1517 (.A(_09455_));
 sg13g2_antennanp ANTENNA_1518 (.A(_09478_));
 sg13g2_antennanp ANTENNA_1519 (.A(_09538_));
 sg13g2_antennanp ANTENNA_1520 (.A(_09613_));
 sg13g2_antennanp ANTENNA_1521 (.A(_09613_));
 sg13g2_antennanp ANTENNA_1522 (.A(_09634_));
 sg13g2_antennanp ANTENNA_1523 (.A(_09657_));
 sg13g2_antennanp ANTENNA_1524 (.A(_09657_));
 sg13g2_antennanp ANTENNA_1525 (.A(_09699_));
 sg13g2_antennanp ANTENNA_1526 (.A(_09726_));
 sg13g2_antennanp ANTENNA_1527 (.A(_09726_));
 sg13g2_antennanp ANTENNA_1528 (.A(_09757_));
 sg13g2_antennanp ANTENNA_1529 (.A(_09757_));
 sg13g2_antennanp ANTENNA_1530 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1531 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1532 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1533 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1534 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1535 (.A(_09893_));
 sg13g2_antennanp ANTENNA_1536 (.A(_10143_));
 sg13g2_antennanp ANTENNA_1537 (.A(_10143_));
 sg13g2_antennanp ANTENNA_1538 (.A(_10143_));
 sg13g2_antennanp ANTENNA_1539 (.A(_10143_));
 sg13g2_antennanp ANTENNA_1540 (.A(_10616_));
 sg13g2_antennanp ANTENNA_1541 (.A(_10616_));
 sg13g2_antennanp ANTENNA_1542 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1543 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1544 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1545 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1546 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1547 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1548 (.A(_10984_));
 sg13g2_antennanp ANTENNA_1549 (.A(_11080_));
 sg13g2_antennanp ANTENNA_1550 (.A(_11080_));
 sg13g2_antennanp ANTENNA_1551 (.A(_11080_));
 sg13g2_antennanp ANTENNA_1552 (.A(_11080_));
 sg13g2_antennanp ANTENNA_1553 (.A(_11080_));
 sg13g2_antennanp ANTENNA_1554 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1555 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1556 (.A(_12140_));
 sg13g2_antennanp ANTENNA_1557 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1558 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1559 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1560 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1561 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1562 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1563 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1564 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1565 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1566 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1567 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1568 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1569 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1570 (.A(_12168_));
 sg13g2_antennanp ANTENNA_1571 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1572 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1573 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1574 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1575 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1576 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1577 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1578 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1579 (.A(_12185_));
 sg13g2_antennanp ANTENNA_1580 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1581 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1582 (.A(_12207_));
 sg13g2_antennanp ANTENNA_1583 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1584 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1585 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1586 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1587 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1588 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1589 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1590 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1591 (.A(_12214_));
 sg13g2_antennanp ANTENNA_1592 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1593 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1594 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1595 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1596 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1597 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1598 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1599 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1600 (.A(_12251_));
 sg13g2_antennanp ANTENNA_1601 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1602 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1603 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1604 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1605 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1606 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1607 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1608 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1609 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1610 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1611 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1612 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1613 (.A(_12335_));
 sg13g2_antennanp ANTENNA_1614 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1615 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1616 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1617 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1618 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1619 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1620 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1621 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1622 (.A(_12632_));
 sg13g2_antennanp ANTENNA_1623 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1624 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1625 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1626 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1627 (.A(_12668_));
 sg13g2_antennanp ANTENNA_1628 (.A(clk));
 sg13g2_antennanp ANTENNA_1629 (.A(clk));
 sg13g2_antennanp ANTENNA_1630 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1631 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1632 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_1633 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_1634 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_1635 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_1636 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_1637 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1638 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_1639 (.A(net467));
 sg13g2_antennanp ANTENNA_1640 (.A(net467));
 sg13g2_antennanp ANTENNA_1641 (.A(net467));
 sg13g2_antennanp ANTENNA_1642 (.A(net467));
 sg13g2_antennanp ANTENNA_1643 (.A(net467));
 sg13g2_antennanp ANTENNA_1644 (.A(net467));
 sg13g2_antennanp ANTENNA_1645 (.A(net467));
 sg13g2_antennanp ANTENNA_1646 (.A(net467));
 sg13g2_antennanp ANTENNA_1647 (.A(net467));
 sg13g2_antennanp ANTENNA_1648 (.A(net533));
 sg13g2_antennanp ANTENNA_1649 (.A(net533));
 sg13g2_antennanp ANTENNA_1650 (.A(net533));
 sg13g2_antennanp ANTENNA_1651 (.A(net533));
 sg13g2_antennanp ANTENNA_1652 (.A(net533));
 sg13g2_antennanp ANTENNA_1653 (.A(net533));
 sg13g2_antennanp ANTENNA_1654 (.A(net533));
 sg13g2_antennanp ANTENNA_1655 (.A(net533));
 sg13g2_antennanp ANTENNA_1656 (.A(net616));
 sg13g2_antennanp ANTENNA_1657 (.A(net616));
 sg13g2_antennanp ANTENNA_1658 (.A(net616));
 sg13g2_antennanp ANTENNA_1659 (.A(net616));
 sg13g2_antennanp ANTENNA_1660 (.A(net616));
 sg13g2_antennanp ANTENNA_1661 (.A(net616));
 sg13g2_antennanp ANTENNA_1662 (.A(net616));
 sg13g2_antennanp ANTENNA_1663 (.A(net616));
 sg13g2_antennanp ANTENNA_1664 (.A(net680));
 sg13g2_antennanp ANTENNA_1665 (.A(net680));
 sg13g2_antennanp ANTENNA_1666 (.A(net680));
 sg13g2_antennanp ANTENNA_1667 (.A(net680));
 sg13g2_antennanp ANTENNA_1668 (.A(net680));
 sg13g2_antennanp ANTENNA_1669 (.A(net680));
 sg13g2_antennanp ANTENNA_1670 (.A(net680));
 sg13g2_antennanp ANTENNA_1671 (.A(net680));
 sg13g2_antennanp ANTENNA_1672 (.A(net702));
 sg13g2_antennanp ANTENNA_1673 (.A(net702));
 sg13g2_antennanp ANTENNA_1674 (.A(net702));
 sg13g2_antennanp ANTENNA_1675 (.A(net702));
 sg13g2_antennanp ANTENNA_1676 (.A(net702));
 sg13g2_antennanp ANTENNA_1677 (.A(net702));
 sg13g2_antennanp ANTENNA_1678 (.A(net702));
 sg13g2_antennanp ANTENNA_1679 (.A(net702));
 sg13g2_antennanp ANTENNA_1680 (.A(net702));
 sg13g2_antennanp ANTENNA_1681 (.A(net749));
 sg13g2_antennanp ANTENNA_1682 (.A(net749));
 sg13g2_antennanp ANTENNA_1683 (.A(net749));
 sg13g2_antennanp ANTENNA_1684 (.A(net749));
 sg13g2_antennanp ANTENNA_1685 (.A(net749));
 sg13g2_antennanp ANTENNA_1686 (.A(net749));
 sg13g2_antennanp ANTENNA_1687 (.A(net749));
 sg13g2_antennanp ANTENNA_1688 (.A(net749));
 sg13g2_antennanp ANTENNA_1689 (.A(net749));
 sg13g2_antennanp ANTENNA_1690 (.A(net882));
 sg13g2_antennanp ANTENNA_1691 (.A(net882));
 sg13g2_antennanp ANTENNA_1692 (.A(net882));
 sg13g2_antennanp ANTENNA_1693 (.A(net882));
 sg13g2_antennanp ANTENNA_1694 (.A(net882));
 sg13g2_antennanp ANTENNA_1695 (.A(net882));
 sg13g2_antennanp ANTENNA_1696 (.A(net882));
 sg13g2_antennanp ANTENNA_1697 (.A(net882));
 sg13g2_antennanp ANTENNA_1698 (.A(net882));
 sg13g2_antennanp ANTENNA_1699 (.A(net884));
 sg13g2_antennanp ANTENNA_1700 (.A(net884));
 sg13g2_antennanp ANTENNA_1701 (.A(net884));
 sg13g2_antennanp ANTENNA_1702 (.A(net884));
 sg13g2_antennanp ANTENNA_1703 (.A(net884));
 sg13g2_antennanp ANTENNA_1704 (.A(net884));
 sg13g2_antennanp ANTENNA_1705 (.A(net884));
 sg13g2_antennanp ANTENNA_1706 (.A(net884));
 sg13g2_antennanp ANTENNA_1707 (.A(net884));
 sg13g2_antennanp ANTENNA_1708 (.A(net929));
 sg13g2_antennanp ANTENNA_1709 (.A(net929));
 sg13g2_antennanp ANTENNA_1710 (.A(net929));
 sg13g2_antennanp ANTENNA_1711 (.A(net929));
 sg13g2_antennanp ANTENNA_1712 (.A(net929));
 sg13g2_antennanp ANTENNA_1713 (.A(net929));
 sg13g2_antennanp ANTENNA_1714 (.A(net929));
 sg13g2_antennanp ANTENNA_1715 (.A(net929));
 sg13g2_antennanp ANTENNA_1716 (.A(net929));
 sg13g2_antennanp ANTENNA_1717 (.A(net929));
 sg13g2_antennanp ANTENNA_1718 (.A(net929));
 sg13g2_antennanp ANTENNA_1719 (.A(net929));
 sg13g2_antennanp ANTENNA_1720 (.A(net929));
 sg13g2_antennanp ANTENNA_1721 (.A(net929));
 sg13g2_antennanp ANTENNA_1722 (.A(net929));
 sg13g2_antennanp ANTENNA_1723 (.A(net929));
 sg13g2_antennanp ANTENNA_1724 (.A(net929));
 sg13g2_antennanp ANTENNA_1725 (.A(net929));
 sg13g2_antennanp ANTENNA_1726 (.A(net929));
 sg13g2_antennanp ANTENNA_1727 (.A(net929));
 sg13g2_antennanp ANTENNA_1728 (.A(net942));
 sg13g2_antennanp ANTENNA_1729 (.A(net942));
 sg13g2_antennanp ANTENNA_1730 (.A(net942));
 sg13g2_antennanp ANTENNA_1731 (.A(net942));
 sg13g2_antennanp ANTENNA_1732 (.A(net942));
 sg13g2_antennanp ANTENNA_1733 (.A(net942));
 sg13g2_antennanp ANTENNA_1734 (.A(net942));
 sg13g2_antennanp ANTENNA_1735 (.A(net942));
 sg13g2_antennanp ANTENNA_1736 (.A(net1000));
 sg13g2_antennanp ANTENNA_1737 (.A(net1000));
 sg13g2_antennanp ANTENNA_1738 (.A(net1000));
 sg13g2_antennanp ANTENNA_1739 (.A(net1000));
 sg13g2_antennanp ANTENNA_1740 (.A(net1000));
 sg13g2_antennanp ANTENNA_1741 (.A(net1000));
 sg13g2_antennanp ANTENNA_1742 (.A(net1000));
 sg13g2_antennanp ANTENNA_1743 (.A(net1000));
 sg13g2_antennanp ANTENNA_1744 (.A(net1000));
 sg13g2_antennanp ANTENNA_1745 (.A(net1000));
 sg13g2_antennanp ANTENNA_1746 (.A(net1000));
 sg13g2_antennanp ANTENNA_1747 (.A(net1000));
 sg13g2_antennanp ANTENNA_1748 (.A(net1000));
 sg13g2_antennanp ANTENNA_1749 (.A(net1000));
 sg13g2_antennanp ANTENNA_1750 (.A(net1000));
 sg13g2_antennanp ANTENNA_1751 (.A(net1000));
 sg13g2_antennanp ANTENNA_1752 (.A(net1000));
 sg13g2_antennanp ANTENNA_1753 (.A(net1000));
 sg13g2_antennanp ANTENNA_1754 (.A(net1000));
 sg13g2_antennanp ANTENNA_1755 (.A(net1000));
 sg13g2_antennanp ANTENNA_1756 (.A(net1000));
 sg13g2_antennanp ANTENNA_1757 (.A(net1023));
 sg13g2_antennanp ANTENNA_1758 (.A(net1023));
 sg13g2_antennanp ANTENNA_1759 (.A(net1023));
 sg13g2_antennanp ANTENNA_1760 (.A(net1023));
 sg13g2_antennanp ANTENNA_1761 (.A(net1023));
 sg13g2_antennanp ANTENNA_1762 (.A(net1023));
 sg13g2_antennanp ANTENNA_1763 (.A(net1023));
 sg13g2_antennanp ANTENNA_1764 (.A(net1023));
 sg13g2_antennanp ANTENNA_1765 (.A(net1023));
 sg13g2_antennanp ANTENNA_1766 (.A(net1026));
 sg13g2_antennanp ANTENNA_1767 (.A(net1026));
 sg13g2_antennanp ANTENNA_1768 (.A(net1026));
 sg13g2_antennanp ANTENNA_1769 (.A(net1026));
 sg13g2_antennanp ANTENNA_1770 (.A(net1026));
 sg13g2_antennanp ANTENNA_1771 (.A(net1026));
 sg13g2_antennanp ANTENNA_1772 (.A(net1026));
 sg13g2_antennanp ANTENNA_1773 (.A(net1026));
 sg13g2_antennanp ANTENNA_1774 (.A(net1027));
 sg13g2_antennanp ANTENNA_1775 (.A(net1027));
 sg13g2_antennanp ANTENNA_1776 (.A(net1027));
 sg13g2_antennanp ANTENNA_1777 (.A(net1027));
 sg13g2_antennanp ANTENNA_1778 (.A(net1027));
 sg13g2_antennanp ANTENNA_1779 (.A(net1027));
 sg13g2_antennanp ANTENNA_1780 (.A(net1027));
 sg13g2_antennanp ANTENNA_1781 (.A(net1027));
 sg13g2_antennanp ANTENNA_1782 (.A(net1109));
 sg13g2_antennanp ANTENNA_1783 (.A(net1109));
 sg13g2_antennanp ANTENNA_1784 (.A(net1109));
 sg13g2_antennanp ANTENNA_1785 (.A(net1109));
 sg13g2_antennanp ANTENNA_1786 (.A(net1109));
 sg13g2_antennanp ANTENNA_1787 (.A(net1109));
 sg13g2_antennanp ANTENNA_1788 (.A(net1109));
 sg13g2_antennanp ANTENNA_1789 (.A(net1109));
 sg13g2_antennanp ANTENNA_1790 (.A(net1143));
 sg13g2_antennanp ANTENNA_1791 (.A(net1143));
 sg13g2_antennanp ANTENNA_1792 (.A(net1143));
 sg13g2_antennanp ANTENNA_1793 (.A(net1143));
 sg13g2_antennanp ANTENNA_1794 (.A(net1143));
 sg13g2_antennanp ANTENNA_1795 (.A(net1143));
 sg13g2_antennanp ANTENNA_1796 (.A(net1143));
 sg13g2_antennanp ANTENNA_1797 (.A(net1143));
 sg13g2_antennanp ANTENNA_1798 (.A(net1143));
 sg13g2_antennanp ANTENNA_1799 (.A(net1166));
 sg13g2_antennanp ANTENNA_1800 (.A(net1166));
 sg13g2_antennanp ANTENNA_1801 (.A(net1166));
 sg13g2_antennanp ANTENNA_1802 (.A(net1166));
 sg13g2_antennanp ANTENNA_1803 (.A(net1166));
 sg13g2_antennanp ANTENNA_1804 (.A(net1166));
 sg13g2_antennanp ANTENNA_1805 (.A(net1166));
 sg13g2_antennanp ANTENNA_1806 (.A(net1166));
 sg13g2_antennanp ANTENNA_1807 (.A(net1166));
 sg13g2_antennanp ANTENNA_1808 (.A(_00741_));
 sg13g2_antennanp ANTENNA_1809 (.A(_00743_));
 sg13g2_antennanp ANTENNA_1810 (.A(_00783_));
 sg13g2_antennanp ANTENNA_1811 (.A(_00919_));
 sg13g2_antennanp ANTENNA_1812 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1813 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1814 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1815 (.A(_02921_));
 sg13g2_antennanp ANTENNA_1816 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1817 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1818 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1819 (.A(_02950_));
 sg13g2_antennanp ANTENNA_1820 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1821 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1822 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1823 (.A(_03050_));
 sg13g2_antennanp ANTENNA_1824 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1825 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1826 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1827 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1828 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1829 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1830 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1831 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1832 (.A(_03056_));
 sg13g2_antennanp ANTENNA_1833 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1834 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1835 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1836 (.A(_03072_));
 sg13g2_antennanp ANTENNA_1837 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1838 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1839 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1840 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1841 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1842 (.A(_03073_));
 sg13g2_antennanp ANTENNA_1843 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1844 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1845 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1846 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1847 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1848 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1849 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1850 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1851 (.A(_03077_));
 sg13g2_antennanp ANTENNA_1852 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1853 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1854 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1855 (.A(_03080_));
 sg13g2_antennanp ANTENNA_1856 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1857 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1858 (.A(_03102_));
 sg13g2_antennanp ANTENNA_1859 (.A(_03115_));
 sg13g2_antennanp ANTENNA_1860 (.A(_03228_));
 sg13g2_antennanp ANTENNA_1861 (.A(_03252_));
 sg13g2_antennanp ANTENNA_1862 (.A(_03354_));
 sg13g2_antennanp ANTENNA_1863 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1864 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1865 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1866 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1867 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1868 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1869 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1870 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1871 (.A(_03620_));
 sg13g2_antennanp ANTENNA_1872 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1873 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1874 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1875 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1876 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1877 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1878 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1879 (.A(_03624_));
 sg13g2_antennanp ANTENNA_1880 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1881 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1882 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1883 (.A(_03625_));
 sg13g2_antennanp ANTENNA_1884 (.A(_05150_));
 sg13g2_antennanp ANTENNA_1885 (.A(_05213_));
 sg13g2_antennanp ANTENNA_1886 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1887 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1888 (.A(_05287_));
 sg13g2_antennanp ANTENNA_1889 (.A(_05297_));
 sg13g2_antennanp ANTENNA_1890 (.A(_05447_));
 sg13g2_antennanp ANTENNA_1891 (.A(_05453_));
 sg13g2_antennanp ANTENNA_1892 (.A(_05580_));
 sg13g2_antennanp ANTENNA_1893 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1894 (.A(_05760_));
 sg13g2_antennanp ANTENNA_1895 (.A(_05764_));
 sg13g2_antennanp ANTENNA_1896 (.A(_05764_));
 sg13g2_antennanp ANTENNA_1897 (.A(_05769_));
 sg13g2_antennanp ANTENNA_1898 (.A(_05772_));
 sg13g2_antennanp ANTENNA_1899 (.A(_05778_));
 sg13g2_antennanp ANTENNA_1900 (.A(_05779_));
 sg13g2_antennanp ANTENNA_1901 (.A(_05780_));
 sg13g2_antennanp ANTENNA_1902 (.A(_05783_));
 sg13g2_antennanp ANTENNA_1903 (.A(_06004_));
 sg13g2_antennanp ANTENNA_1904 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1905 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1906 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1907 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1908 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1909 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1910 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1911 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1912 (.A(_06495_));
 sg13g2_antennanp ANTENNA_1913 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1914 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1915 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1916 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1917 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1918 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1919 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1920 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1921 (.A(_06498_));
 sg13g2_antennanp ANTENNA_1922 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1923 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1924 (.A(_06745_));
 sg13g2_antennanp ANTENNA_1925 (.A(_08276_));
 sg13g2_antennanp ANTENNA_1926 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1927 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1928 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1929 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1930 (.A(_08290_));
 sg13g2_antennanp ANTENNA_1931 (.A(_08292_));
 sg13g2_antennanp ANTENNA_1932 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1933 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1934 (.A(_08301_));
 sg13g2_antennanp ANTENNA_1935 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1936 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1937 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1938 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1939 (.A(_08336_));
 sg13g2_antennanp ANTENNA_1940 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1941 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1942 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1943 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1944 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1945 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1946 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1947 (.A(_08355_));
 sg13g2_antennanp ANTENNA_1948 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1949 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1950 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1951 (.A(_08459_));
 sg13g2_antennanp ANTENNA_1952 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1953 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1954 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1955 (.A(_08529_));
 sg13g2_antennanp ANTENNA_1956 (.A(_08561_));
 sg13g2_antennanp ANTENNA_1957 (.A(_08590_));
 sg13g2_antennanp ANTENNA_1958 (.A(_08670_));
 sg13g2_antennanp ANTENNA_1959 (.A(_08670_));
 sg13g2_antennanp ANTENNA_1960 (.A(_08670_));
 sg13g2_antennanp ANTENNA_1961 (.A(_08690_));
 sg13g2_antennanp ANTENNA_1962 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1963 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1964 (.A(_08777_));
 sg13g2_antennanp ANTENNA_1965 (.A(_08906_));
 sg13g2_antennanp ANTENNA_1966 (.A(_08906_));
 sg13g2_antennanp ANTENNA_1967 (.A(_08930_));
 sg13g2_antennanp ANTENNA_1968 (.A(_08930_));
 sg13g2_antennanp ANTENNA_1969 (.A(_08968_));
 sg13g2_antennanp ANTENNA_1970 (.A(_08968_));
 sg13g2_antennanp ANTENNA_1971 (.A(_09006_));
 sg13g2_antennanp ANTENNA_1972 (.A(_09072_));
 sg13g2_antennanp ANTENNA_1973 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1974 (.A(_09104_));
 sg13g2_antennanp ANTENNA_1975 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1976 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1977 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1978 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1979 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1980 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1981 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1982 (.A(_09164_));
 sg13g2_antennanp ANTENNA_1983 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1984 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1985 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1986 (.A(_09269_));
 sg13g2_antennanp ANTENNA_1987 (.A(_09330_));
 sg13g2_antennanp ANTENNA_1988 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1989 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1990 (.A(_09360_));
 sg13g2_antennanp ANTENNA_1991 (.A(_09386_));
 sg13g2_antennanp ANTENNA_1992 (.A(_09411_));
 sg13g2_antennanp ANTENNA_1993 (.A(_09411_));
 sg13g2_antennanp ANTENNA_1994 (.A(_09411_));
 sg13g2_antennanp ANTENNA_1995 (.A(_09440_));
 sg13g2_antennanp ANTENNA_1996 (.A(_09478_));
 sg13g2_antennanp ANTENNA_1997 (.A(_09538_));
 sg13g2_antennanp ANTENNA_1998 (.A(_09613_));
 sg13g2_antennanp ANTENNA_1999 (.A(_09613_));
 sg13g2_antennanp ANTENNA_2000 (.A(_09634_));
 sg13g2_antennanp ANTENNA_2001 (.A(_09657_));
 sg13g2_antennanp ANTENNA_2002 (.A(_09657_));
 sg13g2_antennanp ANTENNA_2003 (.A(_09699_));
 sg13g2_antennanp ANTENNA_2004 (.A(_09726_));
 sg13g2_antennanp ANTENNA_2005 (.A(_09726_));
 sg13g2_antennanp ANTENNA_2006 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2007 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2008 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2009 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2010 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2011 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2012 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2013 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2014 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2015 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2016 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2017 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2018 (.A(_10616_));
 sg13g2_antennanp ANTENNA_2019 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2020 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2021 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2022 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2023 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2024 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2025 (.A(_10984_));
 sg13g2_antennanp ANTENNA_2026 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2027 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2028 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2029 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2030 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2031 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2032 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2033 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2034 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2035 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2036 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2037 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2038 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2039 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2040 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2041 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2042 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2043 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2044 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2045 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2046 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2047 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2048 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2049 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2050 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2051 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2052 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2053 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2054 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2055 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2056 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2057 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2058 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2059 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2060 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2061 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2062 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2063 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2064 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2065 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2066 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2067 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2068 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2069 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2070 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2071 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2072 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2073 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2074 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2075 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2076 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2077 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2078 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2079 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2080 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2081 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2082 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2083 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2084 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2085 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2086 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2087 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2088 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2089 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2090 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2091 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2092 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2093 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2094 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2095 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2096 (.A(clk));
 sg13g2_antennanp ANTENNA_2097 (.A(clk));
 sg13g2_antennanp ANTENNA_2098 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2099 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2100 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2101 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2102 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_2103 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2104 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_2105 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2106 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2107 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2108 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2109 (.A(net11));
 sg13g2_antennanp ANTENNA_2110 (.A(net11));
 sg13g2_antennanp ANTENNA_2111 (.A(net11));
 sg13g2_antennanp ANTENNA_2112 (.A(net68));
 sg13g2_antennanp ANTENNA_2113 (.A(net68));
 sg13g2_antennanp ANTENNA_2114 (.A(net68));
 sg13g2_antennanp ANTENNA_2115 (.A(net68));
 sg13g2_antennanp ANTENNA_2116 (.A(net68));
 sg13g2_antennanp ANTENNA_2117 (.A(net68));
 sg13g2_antennanp ANTENNA_2118 (.A(net68));
 sg13g2_antennanp ANTENNA_2119 (.A(net68));
 sg13g2_antennanp ANTENNA_2120 (.A(net533));
 sg13g2_antennanp ANTENNA_2121 (.A(net533));
 sg13g2_antennanp ANTENNA_2122 (.A(net533));
 sg13g2_antennanp ANTENNA_2123 (.A(net533));
 sg13g2_antennanp ANTENNA_2124 (.A(net533));
 sg13g2_antennanp ANTENNA_2125 (.A(net533));
 sg13g2_antennanp ANTENNA_2126 (.A(net533));
 sg13g2_antennanp ANTENNA_2127 (.A(net533));
 sg13g2_antennanp ANTENNA_2128 (.A(net616));
 sg13g2_antennanp ANTENNA_2129 (.A(net616));
 sg13g2_antennanp ANTENNA_2130 (.A(net616));
 sg13g2_antennanp ANTENNA_2131 (.A(net616));
 sg13g2_antennanp ANTENNA_2132 (.A(net616));
 sg13g2_antennanp ANTENNA_2133 (.A(net616));
 sg13g2_antennanp ANTENNA_2134 (.A(net616));
 sg13g2_antennanp ANTENNA_2135 (.A(net616));
 sg13g2_antennanp ANTENNA_2136 (.A(net680));
 sg13g2_antennanp ANTENNA_2137 (.A(net680));
 sg13g2_antennanp ANTENNA_2138 (.A(net680));
 sg13g2_antennanp ANTENNA_2139 (.A(net680));
 sg13g2_antennanp ANTENNA_2140 (.A(net680));
 sg13g2_antennanp ANTENNA_2141 (.A(net680));
 sg13g2_antennanp ANTENNA_2142 (.A(net680));
 sg13g2_antennanp ANTENNA_2143 (.A(net680));
 sg13g2_antennanp ANTENNA_2144 (.A(net680));
 sg13g2_antennanp ANTENNA_2145 (.A(net680));
 sg13g2_antennanp ANTENNA_2146 (.A(net680));
 sg13g2_antennanp ANTENNA_2147 (.A(net680));
 sg13g2_antennanp ANTENNA_2148 (.A(net680));
 sg13g2_antennanp ANTENNA_2149 (.A(net680));
 sg13g2_antennanp ANTENNA_2150 (.A(net680));
 sg13g2_antennanp ANTENNA_2151 (.A(net702));
 sg13g2_antennanp ANTENNA_2152 (.A(net702));
 sg13g2_antennanp ANTENNA_2153 (.A(net702));
 sg13g2_antennanp ANTENNA_2154 (.A(net702));
 sg13g2_antennanp ANTENNA_2155 (.A(net702));
 sg13g2_antennanp ANTENNA_2156 (.A(net702));
 sg13g2_antennanp ANTENNA_2157 (.A(net702));
 sg13g2_antennanp ANTENNA_2158 (.A(net702));
 sg13g2_antennanp ANTENNA_2159 (.A(net702));
 sg13g2_antennanp ANTENNA_2160 (.A(net749));
 sg13g2_antennanp ANTENNA_2161 (.A(net749));
 sg13g2_antennanp ANTENNA_2162 (.A(net749));
 sg13g2_antennanp ANTENNA_2163 (.A(net749));
 sg13g2_antennanp ANTENNA_2164 (.A(net749));
 sg13g2_antennanp ANTENNA_2165 (.A(net749));
 sg13g2_antennanp ANTENNA_2166 (.A(net749));
 sg13g2_antennanp ANTENNA_2167 (.A(net749));
 sg13g2_antennanp ANTENNA_2168 (.A(net749));
 sg13g2_antennanp ANTENNA_2169 (.A(net882));
 sg13g2_antennanp ANTENNA_2170 (.A(net882));
 sg13g2_antennanp ANTENNA_2171 (.A(net882));
 sg13g2_antennanp ANTENNA_2172 (.A(net882));
 sg13g2_antennanp ANTENNA_2173 (.A(net882));
 sg13g2_antennanp ANTENNA_2174 (.A(net882));
 sg13g2_antennanp ANTENNA_2175 (.A(net882));
 sg13g2_antennanp ANTENNA_2176 (.A(net882));
 sg13g2_antennanp ANTENNA_2177 (.A(net882));
 sg13g2_antennanp ANTENNA_2178 (.A(net884));
 sg13g2_antennanp ANTENNA_2179 (.A(net884));
 sg13g2_antennanp ANTENNA_2180 (.A(net884));
 sg13g2_antennanp ANTENNA_2181 (.A(net884));
 sg13g2_antennanp ANTENNA_2182 (.A(net884));
 sg13g2_antennanp ANTENNA_2183 (.A(net884));
 sg13g2_antennanp ANTENNA_2184 (.A(net884));
 sg13g2_antennanp ANTENNA_2185 (.A(net884));
 sg13g2_antennanp ANTENNA_2186 (.A(net884));
 sg13g2_antennanp ANTENNA_2187 (.A(net929));
 sg13g2_antennanp ANTENNA_2188 (.A(net929));
 sg13g2_antennanp ANTENNA_2189 (.A(net929));
 sg13g2_antennanp ANTENNA_2190 (.A(net929));
 sg13g2_antennanp ANTENNA_2191 (.A(net929));
 sg13g2_antennanp ANTENNA_2192 (.A(net929));
 sg13g2_antennanp ANTENNA_2193 (.A(net929));
 sg13g2_antennanp ANTENNA_2194 (.A(net929));
 sg13g2_antennanp ANTENNA_2195 (.A(net929));
 sg13g2_antennanp ANTENNA_2196 (.A(net929));
 sg13g2_antennanp ANTENNA_2197 (.A(net929));
 sg13g2_antennanp ANTENNA_2198 (.A(net929));
 sg13g2_antennanp ANTENNA_2199 (.A(net929));
 sg13g2_antennanp ANTENNA_2200 (.A(net929));
 sg13g2_antennanp ANTENNA_2201 (.A(net929));
 sg13g2_antennanp ANTENNA_2202 (.A(net929));
 sg13g2_antennanp ANTENNA_2203 (.A(net929));
 sg13g2_antennanp ANTENNA_2204 (.A(net929));
 sg13g2_antennanp ANTENNA_2205 (.A(net929));
 sg13g2_antennanp ANTENNA_2206 (.A(net929));
 sg13g2_antennanp ANTENNA_2207 (.A(net942));
 sg13g2_antennanp ANTENNA_2208 (.A(net942));
 sg13g2_antennanp ANTENNA_2209 (.A(net942));
 sg13g2_antennanp ANTENNA_2210 (.A(net942));
 sg13g2_antennanp ANTENNA_2211 (.A(net942));
 sg13g2_antennanp ANTENNA_2212 (.A(net942));
 sg13g2_antennanp ANTENNA_2213 (.A(net942));
 sg13g2_antennanp ANTENNA_2214 (.A(net942));
 sg13g2_antennanp ANTENNA_2215 (.A(net1000));
 sg13g2_antennanp ANTENNA_2216 (.A(net1000));
 sg13g2_antennanp ANTENNA_2217 (.A(net1000));
 sg13g2_antennanp ANTENNA_2218 (.A(net1000));
 sg13g2_antennanp ANTENNA_2219 (.A(net1000));
 sg13g2_antennanp ANTENNA_2220 (.A(net1000));
 sg13g2_antennanp ANTENNA_2221 (.A(net1000));
 sg13g2_antennanp ANTENNA_2222 (.A(net1000));
 sg13g2_antennanp ANTENNA_2223 (.A(net1000));
 sg13g2_antennanp ANTENNA_2224 (.A(net1000));
 sg13g2_antennanp ANTENNA_2225 (.A(net1000));
 sg13g2_antennanp ANTENNA_2226 (.A(net1000));
 sg13g2_antennanp ANTENNA_2227 (.A(net1000));
 sg13g2_antennanp ANTENNA_2228 (.A(net1023));
 sg13g2_antennanp ANTENNA_2229 (.A(net1023));
 sg13g2_antennanp ANTENNA_2230 (.A(net1023));
 sg13g2_antennanp ANTENNA_2231 (.A(net1023));
 sg13g2_antennanp ANTENNA_2232 (.A(net1023));
 sg13g2_antennanp ANTENNA_2233 (.A(net1023));
 sg13g2_antennanp ANTENNA_2234 (.A(net1023));
 sg13g2_antennanp ANTENNA_2235 (.A(net1023));
 sg13g2_antennanp ANTENNA_2236 (.A(net1023));
 sg13g2_antennanp ANTENNA_2237 (.A(net1023));
 sg13g2_antennanp ANTENNA_2238 (.A(net1023));
 sg13g2_antennanp ANTENNA_2239 (.A(net1023));
 sg13g2_antennanp ANTENNA_2240 (.A(net1023));
 sg13g2_antennanp ANTENNA_2241 (.A(net1026));
 sg13g2_antennanp ANTENNA_2242 (.A(net1026));
 sg13g2_antennanp ANTENNA_2243 (.A(net1026));
 sg13g2_antennanp ANTENNA_2244 (.A(net1026));
 sg13g2_antennanp ANTENNA_2245 (.A(net1026));
 sg13g2_antennanp ANTENNA_2246 (.A(net1026));
 sg13g2_antennanp ANTENNA_2247 (.A(net1026));
 sg13g2_antennanp ANTENNA_2248 (.A(net1026));
 sg13g2_antennanp ANTENNA_2249 (.A(net1027));
 sg13g2_antennanp ANTENNA_2250 (.A(net1027));
 sg13g2_antennanp ANTENNA_2251 (.A(net1027));
 sg13g2_antennanp ANTENNA_2252 (.A(net1027));
 sg13g2_antennanp ANTENNA_2253 (.A(net1027));
 sg13g2_antennanp ANTENNA_2254 (.A(net1027));
 sg13g2_antennanp ANTENNA_2255 (.A(net1027));
 sg13g2_antennanp ANTENNA_2256 (.A(net1027));
 sg13g2_antennanp ANTENNA_2257 (.A(net1166));
 sg13g2_antennanp ANTENNA_2258 (.A(net1166));
 sg13g2_antennanp ANTENNA_2259 (.A(net1166));
 sg13g2_antennanp ANTENNA_2260 (.A(net1166));
 sg13g2_antennanp ANTENNA_2261 (.A(net1166));
 sg13g2_antennanp ANTENNA_2262 (.A(net1166));
 sg13g2_antennanp ANTENNA_2263 (.A(net1166));
 sg13g2_antennanp ANTENNA_2264 (.A(net1166));
 sg13g2_antennanp ANTENNA_2265 (.A(net1166));
 sg13g2_antennanp ANTENNA_2266 (.A(_00741_));
 sg13g2_antennanp ANTENNA_2267 (.A(_00743_));
 sg13g2_antennanp ANTENNA_2268 (.A(_00783_));
 sg13g2_antennanp ANTENNA_2269 (.A(_00919_));
 sg13g2_antennanp ANTENNA_2270 (.A(_02921_));
 sg13g2_antennanp ANTENNA_2271 (.A(_02921_));
 sg13g2_antennanp ANTENNA_2272 (.A(_02921_));
 sg13g2_antennanp ANTENNA_2273 (.A(_02921_));
 sg13g2_antennanp ANTENNA_2274 (.A(_02950_));
 sg13g2_antennanp ANTENNA_2275 (.A(_02950_));
 sg13g2_antennanp ANTENNA_2276 (.A(_02950_));
 sg13g2_antennanp ANTENNA_2277 (.A(_02950_));
 sg13g2_antennanp ANTENNA_2278 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2279 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2280 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2281 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2282 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2283 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2284 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2285 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2286 (.A(_03056_));
 sg13g2_antennanp ANTENNA_2287 (.A(_03072_));
 sg13g2_antennanp ANTENNA_2288 (.A(_03072_));
 sg13g2_antennanp ANTENNA_2289 (.A(_03072_));
 sg13g2_antennanp ANTENNA_2290 (.A(_03072_));
 sg13g2_antennanp ANTENNA_2291 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2292 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2293 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2294 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2295 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2296 (.A(_03073_));
 sg13g2_antennanp ANTENNA_2297 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2298 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2299 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2300 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2301 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2302 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2303 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2304 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2305 (.A(_03077_));
 sg13g2_antennanp ANTENNA_2306 (.A(_03080_));
 sg13g2_antennanp ANTENNA_2307 (.A(_03080_));
 sg13g2_antennanp ANTENNA_2308 (.A(_03080_));
 sg13g2_antennanp ANTENNA_2309 (.A(_03080_));
 sg13g2_antennanp ANTENNA_2310 (.A(_03228_));
 sg13g2_antennanp ANTENNA_2311 (.A(_03252_));
 sg13g2_antennanp ANTENNA_2312 (.A(_03354_));
 sg13g2_antennanp ANTENNA_2313 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2314 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2315 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2316 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2317 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2318 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2319 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2320 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2321 (.A(_03620_));
 sg13g2_antennanp ANTENNA_2322 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2323 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2324 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2325 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2326 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2327 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2328 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2329 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2330 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2331 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2332 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2333 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2334 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2335 (.A(_03624_));
 sg13g2_antennanp ANTENNA_2336 (.A(_05150_));
 sg13g2_antennanp ANTENNA_2337 (.A(_05150_));
 sg13g2_antennanp ANTENNA_2338 (.A(_05213_));
 sg13g2_antennanp ANTENNA_2339 (.A(_05278_));
 sg13g2_antennanp ANTENNA_2340 (.A(_05287_));
 sg13g2_antennanp ANTENNA_2341 (.A(_05297_));
 sg13g2_antennanp ANTENNA_2342 (.A(_05447_));
 sg13g2_antennanp ANTENNA_2343 (.A(_05453_));
 sg13g2_antennanp ANTENNA_2344 (.A(_05580_));
 sg13g2_antennanp ANTENNA_2345 (.A(_05760_));
 sg13g2_antennanp ANTENNA_2346 (.A(_05760_));
 sg13g2_antennanp ANTENNA_2347 (.A(_05764_));
 sg13g2_antennanp ANTENNA_2348 (.A(_05769_));
 sg13g2_antennanp ANTENNA_2349 (.A(_05772_));
 sg13g2_antennanp ANTENNA_2350 (.A(_05778_));
 sg13g2_antennanp ANTENNA_2351 (.A(_05779_));
 sg13g2_antennanp ANTENNA_2352 (.A(_05780_));
 sg13g2_antennanp ANTENNA_2353 (.A(_05783_));
 sg13g2_antennanp ANTENNA_2354 (.A(_06004_));
 sg13g2_antennanp ANTENNA_2355 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2356 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2357 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2358 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2359 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2360 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2361 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2362 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2363 (.A(_06495_));
 sg13g2_antennanp ANTENNA_2364 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2365 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2366 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2367 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2368 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2369 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2370 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2371 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2372 (.A(_06498_));
 sg13g2_antennanp ANTENNA_2373 (.A(_06745_));
 sg13g2_antennanp ANTENNA_2374 (.A(_06745_));
 sg13g2_antennanp ANTENNA_2375 (.A(_06745_));
 sg13g2_antennanp ANTENNA_2376 (.A(_08276_));
 sg13g2_antennanp ANTENNA_2377 (.A(_08292_));
 sg13g2_antennanp ANTENNA_2378 (.A(_08301_));
 sg13g2_antennanp ANTENNA_2379 (.A(_08301_));
 sg13g2_antennanp ANTENNA_2380 (.A(_08301_));
 sg13g2_antennanp ANTENNA_2381 (.A(_08336_));
 sg13g2_antennanp ANTENNA_2382 (.A(_08336_));
 sg13g2_antennanp ANTENNA_2383 (.A(_08336_));
 sg13g2_antennanp ANTENNA_2384 (.A(_08336_));
 sg13g2_antennanp ANTENNA_2385 (.A(_08336_));
 sg13g2_antennanp ANTENNA_2386 (.A(_08511_));
 sg13g2_antennanp ANTENNA_2387 (.A(_08511_));
 sg13g2_antennanp ANTENNA_2388 (.A(_08511_));
 sg13g2_antennanp ANTENNA_2389 (.A(_08529_));
 sg13g2_antennanp ANTENNA_2390 (.A(_08529_));
 sg13g2_antennanp ANTENNA_2391 (.A(_08529_));
 sg13g2_antennanp ANTENNA_2392 (.A(_08529_));
 sg13g2_antennanp ANTENNA_2393 (.A(_08561_));
 sg13g2_antennanp ANTENNA_2394 (.A(_08590_));
 sg13g2_antennanp ANTENNA_2395 (.A(_08690_));
 sg13g2_antennanp ANTENNA_2396 (.A(_08777_));
 sg13g2_antennanp ANTENNA_2397 (.A(_08777_));
 sg13g2_antennanp ANTENNA_2398 (.A(_08777_));
 sg13g2_antennanp ANTENNA_2399 (.A(_08906_));
 sg13g2_antennanp ANTENNA_2400 (.A(_08906_));
 sg13g2_antennanp ANTENNA_2401 (.A(_08930_));
 sg13g2_antennanp ANTENNA_2402 (.A(_08968_));
 sg13g2_antennanp ANTENNA_2403 (.A(_08968_));
 sg13g2_antennanp ANTENNA_2404 (.A(_09006_));
 sg13g2_antennanp ANTENNA_2405 (.A(_09072_));
 sg13g2_antennanp ANTENNA_2406 (.A(_09072_));
 sg13g2_antennanp ANTENNA_2407 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2408 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2409 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2410 (.A(_09104_));
 sg13g2_antennanp ANTENNA_2411 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2412 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2413 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2414 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2415 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2416 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2417 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2418 (.A(_09164_));
 sg13g2_antennanp ANTENNA_2419 (.A(_09269_));
 sg13g2_antennanp ANTENNA_2420 (.A(_09269_));
 sg13g2_antennanp ANTENNA_2421 (.A(_09269_));
 sg13g2_antennanp ANTENNA_2422 (.A(_09269_));
 sg13g2_antennanp ANTENNA_2423 (.A(_09330_));
 sg13g2_antennanp ANTENNA_2424 (.A(_09330_));
 sg13g2_antennanp ANTENNA_2425 (.A(_09330_));
 sg13g2_antennanp ANTENNA_2426 (.A(_09360_));
 sg13g2_antennanp ANTENNA_2427 (.A(_09360_));
 sg13g2_antennanp ANTENNA_2428 (.A(_09360_));
 sg13g2_antennanp ANTENNA_2429 (.A(_09386_));
 sg13g2_antennanp ANTENNA_2430 (.A(_09411_));
 sg13g2_antennanp ANTENNA_2431 (.A(_09440_));
 sg13g2_antennanp ANTENNA_2432 (.A(_09440_));
 sg13g2_antennanp ANTENNA_2433 (.A(_09455_));
 sg13g2_antennanp ANTENNA_2434 (.A(_09455_));
 sg13g2_antennanp ANTENNA_2435 (.A(_09455_));
 sg13g2_antennanp ANTENNA_2436 (.A(_09455_));
 sg13g2_antennanp ANTENNA_2437 (.A(_09478_));
 sg13g2_antennanp ANTENNA_2438 (.A(_09538_));
 sg13g2_antennanp ANTENNA_2439 (.A(_09538_));
 sg13g2_antennanp ANTENNA_2440 (.A(_09613_));
 sg13g2_antennanp ANTENNA_2441 (.A(_09613_));
 sg13g2_antennanp ANTENNA_2442 (.A(_09613_));
 sg13g2_antennanp ANTENNA_2443 (.A(_09634_));
 sg13g2_antennanp ANTENNA_2444 (.A(_09657_));
 sg13g2_antennanp ANTENNA_2445 (.A(_09657_));
 sg13g2_antennanp ANTENNA_2446 (.A(_09699_));
 sg13g2_antennanp ANTENNA_2447 (.A(_09699_));
 sg13g2_antennanp ANTENNA_2448 (.A(_09726_));
 sg13g2_antennanp ANTENNA_2449 (.A(_09726_));
 sg13g2_antennanp ANTENNA_2450 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2451 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2452 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2453 (.A(_09757_));
 sg13g2_antennanp ANTENNA_2454 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2455 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2456 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2457 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2458 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2459 (.A(_09893_));
 sg13g2_antennanp ANTENNA_2460 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2461 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2462 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2463 (.A(_10040_));
 sg13g2_antennanp ANTENNA_2464 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2465 (.A(_10143_));
 sg13g2_antennanp ANTENNA_2466 (.A(_10322_));
 sg13g2_antennanp ANTENNA_2467 (.A(_10322_));
 sg13g2_antennanp ANTENNA_2468 (.A(_10616_));
 sg13g2_antennanp ANTENNA_2469 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2470 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2471 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2472 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2473 (.A(_11080_));
 sg13g2_antennanp ANTENNA_2474 (.A(_12014_));
 sg13g2_antennanp ANTENNA_2475 (.A(_12014_));
 sg13g2_antennanp ANTENNA_2476 (.A(_12014_));
 sg13g2_antennanp ANTENNA_2477 (.A(_12074_));
 sg13g2_antennanp ANTENNA_2478 (.A(_12074_));
 sg13g2_antennanp ANTENNA_2479 (.A(_12074_));
 sg13g2_antennanp ANTENNA_2480 (.A(_12074_));
 sg13g2_antennanp ANTENNA_2481 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2482 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2483 (.A(_12140_));
 sg13g2_antennanp ANTENNA_2484 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2485 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2486 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2487 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2488 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2489 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2490 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2491 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2492 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2493 (.A(_12161_));
 sg13g2_antennanp ANTENNA_2494 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2495 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2496 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2497 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2498 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2499 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2500 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2501 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2502 (.A(_12168_));
 sg13g2_antennanp ANTENNA_2503 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2504 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2505 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2506 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2507 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2508 (.A(_12185_));
 sg13g2_antennanp ANTENNA_2509 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2510 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2511 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2512 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2513 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2514 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2515 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2516 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2517 (.A(_12207_));
 sg13g2_antennanp ANTENNA_2518 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2519 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2520 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2521 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2522 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2523 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2524 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2525 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2526 (.A(_12214_));
 sg13g2_antennanp ANTENNA_2527 (.A(_12251_));
 sg13g2_antennanp ANTENNA_2528 (.A(_12251_));
 sg13g2_antennanp ANTENNA_2529 (.A(_12251_));
 sg13g2_antennanp ANTENNA_2530 (.A(_12251_));
 sg13g2_antennanp ANTENNA_2531 (.A(_12251_));
 sg13g2_antennanp ANTENNA_2532 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2533 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2534 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2535 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2536 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2537 (.A(_12335_));
 sg13g2_antennanp ANTENNA_2538 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2539 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2540 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2541 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2542 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2543 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2544 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2545 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2546 (.A(_12632_));
 sg13g2_antennanp ANTENNA_2547 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2548 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2549 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2550 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2551 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2552 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2553 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2554 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2555 (.A(_12668_));
 sg13g2_antennanp ANTENNA_2556 (.A(clk));
 sg13g2_antennanp ANTENNA_2557 (.A(clk));
 sg13g2_antennanp ANTENNA_2558 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2559 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2560 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2561 (.A(\cpu.ex.c_mult[0] ));
 sg13g2_antennanp ANTENNA_2562 (.A(\cpu.ex.pc[1] ));
 sg13g2_antennanp ANTENNA_2563 (.A(\cpu.ex.pc[2] ));
 sg13g2_antennanp ANTENNA_2564 (.A(\cpu.ex.pc[3] ));
 sg13g2_antennanp ANTENNA_2565 (.A(\cpu.qspi.c_wstrobe_i ));
 sg13g2_antennanp ANTENNA_2566 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2567 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2568 (.A(uio_in[3]));
 sg13g2_antennanp ANTENNA_2569 (.A(net11));
 sg13g2_antennanp ANTENNA_2570 (.A(net11));
 sg13g2_antennanp ANTENNA_2571 (.A(net467));
 sg13g2_antennanp ANTENNA_2572 (.A(net467));
 sg13g2_antennanp ANTENNA_2573 (.A(net467));
 sg13g2_antennanp ANTENNA_2574 (.A(net467));
 sg13g2_antennanp ANTENNA_2575 (.A(net467));
 sg13g2_antennanp ANTENNA_2576 (.A(net467));
 sg13g2_antennanp ANTENNA_2577 (.A(net467));
 sg13g2_antennanp ANTENNA_2578 (.A(net467));
 sg13g2_antennanp ANTENNA_2579 (.A(net467));
 sg13g2_antennanp ANTENNA_2580 (.A(net533));
 sg13g2_antennanp ANTENNA_2581 (.A(net533));
 sg13g2_antennanp ANTENNA_2582 (.A(net533));
 sg13g2_antennanp ANTENNA_2583 (.A(net533));
 sg13g2_antennanp ANTENNA_2584 (.A(net533));
 sg13g2_antennanp ANTENNA_2585 (.A(net533));
 sg13g2_antennanp ANTENNA_2586 (.A(net533));
 sg13g2_antennanp ANTENNA_2587 (.A(net533));
 sg13g2_antennanp ANTENNA_2588 (.A(net616));
 sg13g2_antennanp ANTENNA_2589 (.A(net616));
 sg13g2_antennanp ANTENNA_2590 (.A(net616));
 sg13g2_antennanp ANTENNA_2591 (.A(net616));
 sg13g2_antennanp ANTENNA_2592 (.A(net616));
 sg13g2_antennanp ANTENNA_2593 (.A(net616));
 sg13g2_antennanp ANTENNA_2594 (.A(net616));
 sg13g2_antennanp ANTENNA_2595 (.A(net616));
 sg13g2_antennanp ANTENNA_2596 (.A(net680));
 sg13g2_antennanp ANTENNA_2597 (.A(net680));
 sg13g2_antennanp ANTENNA_2598 (.A(net680));
 sg13g2_antennanp ANTENNA_2599 (.A(net680));
 sg13g2_antennanp ANTENNA_2600 (.A(net680));
 sg13g2_antennanp ANTENNA_2601 (.A(net680));
 sg13g2_antennanp ANTENNA_2602 (.A(net680));
 sg13g2_antennanp ANTENNA_2603 (.A(net680));
 sg13g2_antennanp ANTENNA_2604 (.A(net680));
 sg13g2_antennanp ANTENNA_2605 (.A(net680));
 sg13g2_antennanp ANTENNA_2606 (.A(net680));
 sg13g2_antennanp ANTENNA_2607 (.A(net680));
 sg13g2_antennanp ANTENNA_2608 (.A(net680));
 sg13g2_antennanp ANTENNA_2609 (.A(net680));
 sg13g2_antennanp ANTENNA_2610 (.A(net680));
 sg13g2_antennanp ANTENNA_2611 (.A(net702));
 sg13g2_antennanp ANTENNA_2612 (.A(net702));
 sg13g2_antennanp ANTENNA_2613 (.A(net702));
 sg13g2_antennanp ANTENNA_2614 (.A(net702));
 sg13g2_antennanp ANTENNA_2615 (.A(net702));
 sg13g2_antennanp ANTENNA_2616 (.A(net702));
 sg13g2_antennanp ANTENNA_2617 (.A(net702));
 sg13g2_antennanp ANTENNA_2618 (.A(net702));
 sg13g2_antennanp ANTENNA_2619 (.A(net702));
 sg13g2_antennanp ANTENNA_2620 (.A(net749));
 sg13g2_antennanp ANTENNA_2621 (.A(net749));
 sg13g2_antennanp ANTENNA_2622 (.A(net749));
 sg13g2_antennanp ANTENNA_2623 (.A(net749));
 sg13g2_antennanp ANTENNA_2624 (.A(net749));
 sg13g2_antennanp ANTENNA_2625 (.A(net749));
 sg13g2_antennanp ANTENNA_2626 (.A(net749));
 sg13g2_antennanp ANTENNA_2627 (.A(net749));
 sg13g2_antennanp ANTENNA_2628 (.A(net749));
 sg13g2_antennanp ANTENNA_2629 (.A(net882));
 sg13g2_antennanp ANTENNA_2630 (.A(net882));
 sg13g2_antennanp ANTENNA_2631 (.A(net882));
 sg13g2_antennanp ANTENNA_2632 (.A(net882));
 sg13g2_antennanp ANTENNA_2633 (.A(net882));
 sg13g2_antennanp ANTENNA_2634 (.A(net882));
 sg13g2_antennanp ANTENNA_2635 (.A(net882));
 sg13g2_antennanp ANTENNA_2636 (.A(net882));
 sg13g2_antennanp ANTENNA_2637 (.A(net882));
 sg13g2_antennanp ANTENNA_2638 (.A(net884));
 sg13g2_antennanp ANTENNA_2639 (.A(net884));
 sg13g2_antennanp ANTENNA_2640 (.A(net884));
 sg13g2_antennanp ANTENNA_2641 (.A(net884));
 sg13g2_antennanp ANTENNA_2642 (.A(net884));
 sg13g2_antennanp ANTENNA_2643 (.A(net884));
 sg13g2_antennanp ANTENNA_2644 (.A(net884));
 sg13g2_antennanp ANTENNA_2645 (.A(net884));
 sg13g2_antennanp ANTENNA_2646 (.A(net884));
 sg13g2_antennanp ANTENNA_2647 (.A(net929));
 sg13g2_antennanp ANTENNA_2648 (.A(net929));
 sg13g2_antennanp ANTENNA_2649 (.A(net929));
 sg13g2_antennanp ANTENNA_2650 (.A(net929));
 sg13g2_antennanp ANTENNA_2651 (.A(net929));
 sg13g2_antennanp ANTENNA_2652 (.A(net929));
 sg13g2_antennanp ANTENNA_2653 (.A(net929));
 sg13g2_antennanp ANTENNA_2654 (.A(net929));
 sg13g2_antennanp ANTENNA_2655 (.A(net929));
 sg13g2_antennanp ANTENNA_2656 (.A(net929));
 sg13g2_antennanp ANTENNA_2657 (.A(net929));
 sg13g2_antennanp ANTENNA_2658 (.A(net929));
 sg13g2_antennanp ANTENNA_2659 (.A(net929));
 sg13g2_antennanp ANTENNA_2660 (.A(net929));
 sg13g2_antennanp ANTENNA_2661 (.A(net929));
 sg13g2_antennanp ANTENNA_2662 (.A(net929));
 sg13g2_antennanp ANTENNA_2663 (.A(net929));
 sg13g2_antennanp ANTENNA_2664 (.A(net929));
 sg13g2_antennanp ANTENNA_2665 (.A(net929));
 sg13g2_antennanp ANTENNA_2666 (.A(net929));
 sg13g2_antennanp ANTENNA_2667 (.A(net1023));
 sg13g2_antennanp ANTENNA_2668 (.A(net1023));
 sg13g2_antennanp ANTENNA_2669 (.A(net1023));
 sg13g2_antennanp ANTENNA_2670 (.A(net1023));
 sg13g2_antennanp ANTENNA_2671 (.A(net1023));
 sg13g2_antennanp ANTENNA_2672 (.A(net1023));
 sg13g2_antennanp ANTENNA_2673 (.A(net1023));
 sg13g2_antennanp ANTENNA_2674 (.A(net1023));
 sg13g2_antennanp ANTENNA_2675 (.A(net1023));
 sg13g2_antennanp ANTENNA_2676 (.A(net1026));
 sg13g2_antennanp ANTENNA_2677 (.A(net1026));
 sg13g2_antennanp ANTENNA_2678 (.A(net1026));
 sg13g2_antennanp ANTENNA_2679 (.A(net1026));
 sg13g2_antennanp ANTENNA_2680 (.A(net1026));
 sg13g2_antennanp ANTENNA_2681 (.A(net1026));
 sg13g2_antennanp ANTENNA_2682 (.A(net1026));
 sg13g2_antennanp ANTENNA_2683 (.A(net1026));
 sg13g2_antennanp ANTENNA_2684 (.A(net1166));
 sg13g2_antennanp ANTENNA_2685 (.A(net1166));
 sg13g2_antennanp ANTENNA_2686 (.A(net1166));
 sg13g2_antennanp ANTENNA_2687 (.A(net1166));
 sg13g2_antennanp ANTENNA_2688 (.A(net1166));
 sg13g2_antennanp ANTENNA_2689 (.A(net1166));
 sg13g2_antennanp ANTENNA_2690 (.A(net1166));
 sg13g2_antennanp ANTENNA_2691 (.A(net1166));
 sg13g2_antennanp ANTENNA_2692 (.A(net1166));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_4 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_58 ();
 sg13g2_decap_4 FILLER_0_65 ();
 sg13g2_fill_1 FILLER_0_69 ();
 sg13g2_fill_1 FILLER_0_74 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_1 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_110 ();
 sg13g2_decap_8 FILLER_0_120 ();
 sg13g2_decap_8 FILLER_0_127 ();
 sg13g2_decap_8 FILLER_0_134 ();
 sg13g2_decap_8 FILLER_0_145 ();
 sg13g2_decap_8 FILLER_0_152 ();
 sg13g2_decap_8 FILLER_0_159 ();
 sg13g2_decap_8 FILLER_0_166 ();
 sg13g2_decap_8 FILLER_0_173 ();
 sg13g2_fill_1 FILLER_0_180 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_fill_1 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_4 FILLER_0_270 ();
 sg13g2_fill_2 FILLER_0_274 ();
 sg13g2_decap_8 FILLER_0_302 ();
 sg13g2_decap_8 FILLER_0_309 ();
 sg13g2_decap_8 FILLER_0_316 ();
 sg13g2_decap_8 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_330 ();
 sg13g2_decap_8 FILLER_0_337 ();
 sg13g2_decap_8 FILLER_0_344 ();
 sg13g2_decap_4 FILLER_0_351 ();
 sg13g2_fill_2 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_366 ();
 sg13g2_fill_2 FILLER_0_373 ();
 sg13g2_fill_1 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_380 ();
 sg13g2_decap_8 FILLER_0_387 ();
 sg13g2_decap_8 FILLER_0_394 ();
 sg13g2_fill_1 FILLER_0_401 ();
 sg13g2_decap_8 FILLER_0_407 ();
 sg13g2_decap_4 FILLER_0_414 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_fill_2 FILLER_0_504 ();
 sg13g2_fill_1 FILLER_0_506 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_522 ();
 sg13g2_decap_4 FILLER_0_529 ();
 sg13g2_fill_2 FILLER_0_533 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_fill_2 FILLER_0_560 ();
 sg13g2_fill_2 FILLER_0_592 ();
 sg13g2_fill_1 FILLER_0_594 ();
 sg13g2_fill_1 FILLER_0_599 ();
 sg13g2_decap_8 FILLER_0_604 ();
 sg13g2_decap_8 FILLER_0_611 ();
 sg13g2_decap_4 FILLER_0_618 ();
 sg13g2_fill_2 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_628 ();
 sg13g2_decap_8 FILLER_0_635 ();
 sg13g2_decap_8 FILLER_0_642 ();
 sg13g2_decap_8 FILLER_0_649 ();
 sg13g2_decap_8 FILLER_0_656 ();
 sg13g2_fill_2 FILLER_0_663 ();
 sg13g2_fill_1 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_670 ();
 sg13g2_decap_8 FILLER_0_677 ();
 sg13g2_decap_8 FILLER_0_684 ();
 sg13g2_decap_8 FILLER_0_691 ();
 sg13g2_decap_4 FILLER_0_698 ();
 sg13g2_fill_1 FILLER_0_702 ();
 sg13g2_decap_8 FILLER_0_729 ();
 sg13g2_decap_4 FILLER_0_736 ();
 sg13g2_fill_1 FILLER_0_740 ();
 sg13g2_decap_8 FILLER_0_767 ();
 sg13g2_decap_8 FILLER_0_774 ();
 sg13g2_decap_8 FILLER_0_781 ();
 sg13g2_decap_8 FILLER_0_788 ();
 sg13g2_decap_8 FILLER_0_795 ();
 sg13g2_fill_2 FILLER_0_802 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_4 FILLER_0_836 ();
 sg13g2_fill_2 FILLER_0_840 ();
 sg13g2_fill_1 FILLER_0_852 ();
 sg13g2_fill_2 FILLER_0_879 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_4 FILLER_0_892 ();
 sg13g2_decap_8 FILLER_0_900 ();
 sg13g2_decap_8 FILLER_0_907 ();
 sg13g2_decap_8 FILLER_0_914 ();
 sg13g2_decap_8 FILLER_0_921 ();
 sg13g2_decap_4 FILLER_0_928 ();
 sg13g2_decap_8 FILLER_0_958 ();
 sg13g2_decap_8 FILLER_0_965 ();
 sg13g2_decap_8 FILLER_0_972 ();
 sg13g2_fill_2 FILLER_0_979 ();
 sg13g2_decap_8 FILLER_0_985 ();
 sg13g2_decap_8 FILLER_0_992 ();
 sg13g2_decap_4 FILLER_0_999 ();
 sg13g2_fill_1 FILLER_0_1070 ();
 sg13g2_decap_8 FILLER_0_1079 ();
 sg13g2_decap_8 FILLER_0_1086 ();
 sg13g2_decap_4 FILLER_0_1093 ();
 sg13g2_decap_8 FILLER_0_1123 ();
 sg13g2_decap_8 FILLER_0_1130 ();
 sg13g2_decap_8 FILLER_0_1137 ();
 sg13g2_decap_8 FILLER_0_1144 ();
 sg13g2_decap_8 FILLER_0_1151 ();
 sg13g2_decap_4 FILLER_0_1158 ();
 sg13g2_fill_2 FILLER_0_1162 ();
 sg13g2_decap_8 FILLER_0_1190 ();
 sg13g2_decap_8 FILLER_0_1197 ();
 sg13g2_decap_8 FILLER_0_1204 ();
 sg13g2_fill_1 FILLER_0_1211 ();
 sg13g2_decap_4 FILLER_0_1238 ();
 sg13g2_decap_8 FILLER_0_1268 ();
 sg13g2_decap_4 FILLER_0_1275 ();
 sg13g2_fill_2 FILLER_0_1279 ();
 sg13g2_decap_4 FILLER_0_1307 ();
 sg13g2_fill_2 FILLER_0_1311 ();
 sg13g2_decap_8 FILLER_0_1323 ();
 sg13g2_decap_8 FILLER_0_1330 ();
 sg13g2_decap_8 FILLER_0_1337 ();
 sg13g2_decap_8 FILLER_0_1344 ();
 sg13g2_decap_8 FILLER_0_1351 ();
 sg13g2_fill_1 FILLER_0_1358 ();
 sg13g2_decap_4 FILLER_0_1369 ();
 sg13g2_fill_1 FILLER_0_1373 ();
 sg13g2_decap_8 FILLER_0_1400 ();
 sg13g2_decap_8 FILLER_0_1407 ();
 sg13g2_fill_2 FILLER_0_1414 ();
 sg13g2_decap_8 FILLER_0_1420 ();
 sg13g2_decap_8 FILLER_0_1427 ();
 sg13g2_decap_8 FILLER_0_1434 ();
 sg13g2_fill_1 FILLER_0_1441 ();
 sg13g2_decap_4 FILLER_0_1446 ();
 sg13g2_fill_2 FILLER_0_1450 ();
 sg13g2_decap_8 FILLER_0_1462 ();
 sg13g2_decap_4 FILLER_0_1469 ();
 sg13g2_fill_1 FILLER_0_1473 ();
 sg13g2_decap_8 FILLER_0_1512 ();
 sg13g2_fill_2 FILLER_0_1519 ();
 sg13g2_fill_1 FILLER_0_1521 ();
 sg13g2_fill_1 FILLER_0_1526 ();
 sg13g2_decap_8 FILLER_0_1553 ();
 sg13g2_decap_4 FILLER_0_1560 ();
 sg13g2_fill_1 FILLER_0_1564 ();
 sg13g2_decap_8 FILLER_0_1569 ();
 sg13g2_decap_8 FILLER_0_1576 ();
 sg13g2_decap_8 FILLER_0_1583 ();
 sg13g2_fill_1 FILLER_0_1594 ();
 sg13g2_decap_8 FILLER_0_1625 ();
 sg13g2_decap_8 FILLER_0_1632 ();
 sg13g2_fill_1 FILLER_0_1639 ();
 sg13g2_decap_8 FILLER_0_1670 ();
 sg13g2_decap_4 FILLER_0_1677 ();
 sg13g2_fill_1 FILLER_0_1681 ();
 sg13g2_decap_8 FILLER_0_1692 ();
 sg13g2_decap_8 FILLER_0_1725 ();
 sg13g2_decap_8 FILLER_0_1732 ();
 sg13g2_fill_1 FILLER_0_1739 ();
 sg13g2_decap_8 FILLER_0_1770 ();
 sg13g2_decap_8 FILLER_0_1777 ();
 sg13g2_decap_8 FILLER_0_1784 ();
 sg13g2_fill_2 FILLER_0_1791 ();
 sg13g2_fill_1 FILLER_0_1793 ();
 sg13g2_decap_8 FILLER_0_1798 ();
 sg13g2_decap_8 FILLER_0_1805 ();
 sg13g2_decap_8 FILLER_0_1812 ();
 sg13g2_decap_8 FILLER_0_1819 ();
 sg13g2_decap_4 FILLER_0_1826 ();
 sg13g2_decap_8 FILLER_0_1838 ();
 sg13g2_decap_8 FILLER_0_1845 ();
 sg13g2_fill_1 FILLER_0_1852 ();
 sg13g2_decap_4 FILLER_0_1857 ();
 sg13g2_decap_8 FILLER_0_1873 ();
 sg13g2_decap_8 FILLER_0_1880 ();
 sg13g2_decap_8 FILLER_0_1887 ();
 sg13g2_decap_8 FILLER_0_1894 ();
 sg13g2_decap_8 FILLER_0_1901 ();
 sg13g2_decap_8 FILLER_0_1908 ();
 sg13g2_decap_8 FILLER_0_1915 ();
 sg13g2_decap_8 FILLER_0_1922 ();
 sg13g2_decap_8 FILLER_0_1929 ();
 sg13g2_decap_4 FILLER_0_1936 ();
 sg13g2_decap_8 FILLER_0_1950 ();
 sg13g2_decap_8 FILLER_0_1957 ();
 sg13g2_decap_8 FILLER_0_1964 ();
 sg13g2_decap_8 FILLER_0_1971 ();
 sg13g2_decap_8 FILLER_0_1978 ();
 sg13g2_decap_8 FILLER_0_2011 ();
 sg13g2_fill_1 FILLER_0_2018 ();
 sg13g2_decap_8 FILLER_0_2027 ();
 sg13g2_decap_8 FILLER_0_2034 ();
 sg13g2_fill_1 FILLER_0_2041 ();
 sg13g2_decap_8 FILLER_0_2068 ();
 sg13g2_decap_8 FILLER_0_2075 ();
 sg13g2_fill_2 FILLER_0_2082 ();
 sg13g2_fill_1 FILLER_0_2084 ();
 sg13g2_decap_8 FILLER_0_2089 ();
 sg13g2_decap_8 FILLER_0_2096 ();
 sg13g2_fill_2 FILLER_0_2103 ();
 sg13g2_decap_4 FILLER_0_2115 ();
 sg13g2_fill_2 FILLER_0_2119 ();
 sg13g2_decap_8 FILLER_0_2125 ();
 sg13g2_decap_8 FILLER_0_2132 ();
 sg13g2_decap_8 FILLER_0_2139 ();
 sg13g2_decap_4 FILLER_0_2150 ();
 sg13g2_decap_8 FILLER_0_2158 ();
 sg13g2_fill_1 FILLER_0_2165 ();
 sg13g2_decap_4 FILLER_0_2174 ();
 sg13g2_fill_2 FILLER_0_2178 ();
 sg13g2_fill_2 FILLER_0_2184 ();
 sg13g2_fill_1 FILLER_0_2186 ();
 sg13g2_decap_8 FILLER_0_2197 ();
 sg13g2_decap_8 FILLER_0_2204 ();
 sg13g2_decap_8 FILLER_0_2211 ();
 sg13g2_decap_8 FILLER_0_2218 ();
 sg13g2_fill_2 FILLER_0_2225 ();
 sg13g2_fill_2 FILLER_0_2237 ();
 sg13g2_fill_1 FILLER_0_2239 ();
 sg13g2_decap_8 FILLER_0_2267 ();
 sg13g2_decap_8 FILLER_0_2274 ();
 sg13g2_decap_8 FILLER_0_2281 ();
 sg13g2_fill_1 FILLER_0_2288 ();
 sg13g2_decap_4 FILLER_0_2309 ();
 sg13g2_decap_8 FILLER_0_2327 ();
 sg13g2_decap_8 FILLER_0_2334 ();
 sg13g2_decap_8 FILLER_0_2341 ();
 sg13g2_decap_8 FILLER_0_2348 ();
 sg13g2_decap_8 FILLER_0_2355 ();
 sg13g2_decap_4 FILLER_0_2362 ();
 sg13g2_fill_1 FILLER_0_2366 ();
 sg13g2_decap_4 FILLER_0_2375 ();
 sg13g2_fill_2 FILLER_0_2379 ();
 sg13g2_decap_8 FILLER_0_2395 ();
 sg13g2_fill_2 FILLER_0_2402 ();
 sg13g2_decap_8 FILLER_0_2408 ();
 sg13g2_decap_8 FILLER_0_2415 ();
 sg13g2_decap_8 FILLER_0_2432 ();
 sg13g2_decap_8 FILLER_0_2439 ();
 sg13g2_decap_8 FILLER_0_2446 ();
 sg13g2_decap_8 FILLER_0_2453 ();
 sg13g2_decap_8 FILLER_0_2460 ();
 sg13g2_decap_8 FILLER_0_2467 ();
 sg13g2_decap_8 FILLER_0_2474 ();
 sg13g2_decap_8 FILLER_0_2481 ();
 sg13g2_decap_8 FILLER_0_2488 ();
 sg13g2_decap_8 FILLER_0_2495 ();
 sg13g2_decap_8 FILLER_0_2506 ();
 sg13g2_decap_8 FILLER_0_2513 ();
 sg13g2_decap_8 FILLER_0_2520 ();
 sg13g2_decap_8 FILLER_0_2527 ();
 sg13g2_decap_8 FILLER_0_2534 ();
 sg13g2_decap_8 FILLER_0_2541 ();
 sg13g2_decap_8 FILLER_0_2548 ();
 sg13g2_decap_8 FILLER_0_2555 ();
 sg13g2_decap_8 FILLER_0_2562 ();
 sg13g2_decap_8 FILLER_0_2569 ();
 sg13g2_decap_8 FILLER_0_2576 ();
 sg13g2_decap_8 FILLER_0_2583 ();
 sg13g2_decap_8 FILLER_0_2590 ();
 sg13g2_decap_8 FILLER_0_2597 ();
 sg13g2_decap_8 FILLER_0_2604 ();
 sg13g2_decap_8 FILLER_0_2611 ();
 sg13g2_decap_8 FILLER_0_2618 ();
 sg13g2_decap_8 FILLER_0_2625 ();
 sg13g2_decap_8 FILLER_0_2632 ();
 sg13g2_decap_8 FILLER_0_2639 ();
 sg13g2_decap_8 FILLER_0_2646 ();
 sg13g2_decap_8 FILLER_0_2653 ();
 sg13g2_decap_8 FILLER_0_2660 ();
 sg13g2_fill_2 FILLER_0_2667 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_4 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_32 ();
 sg13g2_fill_2 FILLER_1_63 ();
 sg13g2_decap_4 FILLER_1_91 ();
 sg13g2_fill_1 FILLER_1_95 ();
 sg13g2_fill_2 FILLER_1_129 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_fill_2 FILLER_1_168 ();
 sg13g2_fill_1 FILLER_1_170 ();
 sg13g2_fill_1 FILLER_1_181 ();
 sg13g2_decap_8 FILLER_1_212 ();
 sg13g2_decap_4 FILLER_1_219 ();
 sg13g2_fill_2 FILLER_1_223 ();
 sg13g2_decap_4 FILLER_1_269 ();
 sg13g2_fill_1 FILLER_1_273 ();
 sg13g2_fill_1 FILLER_1_282 ();
 sg13g2_decap_4 FILLER_1_313 ();
 sg13g2_fill_2 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_4 FILLER_1_388 ();
 sg13g2_fill_2 FILLER_1_392 ();
 sg13g2_decap_4 FILLER_1_463 ();
 sg13g2_fill_1 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_554 ();
 sg13g2_decap_8 FILLER_1_561 ();
 sg13g2_fill_1 FILLER_1_568 ();
 sg13g2_fill_2 FILLER_1_630 ();
 sg13g2_fill_2 FILLER_1_636 ();
 sg13g2_fill_1 FILLER_1_638 ();
 sg13g2_fill_1 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_671 ();
 sg13g2_decap_8 FILLER_1_678 ();
 sg13g2_decap_4 FILLER_1_685 ();
 sg13g2_fill_2 FILLER_1_689 ();
 sg13g2_decap_8 FILLER_1_696 ();
 sg13g2_decap_8 FILLER_1_712 ();
 sg13g2_fill_2 FILLER_1_719 ();
 sg13g2_fill_1 FILLER_1_721 ();
 sg13g2_decap_4 FILLER_1_731 ();
 sg13g2_fill_1 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_759 ();
 sg13g2_decap_4 FILLER_1_766 ();
 sg13g2_fill_1 FILLER_1_770 ();
 sg13g2_decap_4 FILLER_1_775 ();
 sg13g2_fill_2 FILLER_1_779 ();
 sg13g2_fill_2 FILLER_1_817 ();
 sg13g2_fill_2 FILLER_1_829 ();
 sg13g2_fill_1 FILLER_1_831 ();
 sg13g2_fill_1 FILLER_1_855 ();
 sg13g2_decap_4 FILLER_1_866 ();
 sg13g2_fill_2 FILLER_1_870 ();
 sg13g2_fill_1 FILLER_1_907 ();
 sg13g2_fill_1 FILLER_1_912 ();
 sg13g2_fill_1 FILLER_1_918 ();
 sg13g2_fill_2 FILLER_1_923 ();
 sg13g2_fill_2 FILLER_1_961 ();
 sg13g2_fill_2 FILLER_1_989 ();
 sg13g2_fill_1 FILLER_1_991 ();
 sg13g2_fill_2 FILLER_1_1018 ();
 sg13g2_fill_1 FILLER_1_1020 ();
 sg13g2_fill_2 FILLER_1_1025 ();
 sg13g2_fill_1 FILLER_1_1027 ();
 sg13g2_fill_2 FILLER_1_1038 ();
 sg13g2_fill_1 FILLER_1_1053 ();
 sg13g2_decap_8 FILLER_1_1098 ();
 sg13g2_decap_8 FILLER_1_1105 ();
 sg13g2_decap_8 FILLER_1_1112 ();
 sg13g2_fill_1 FILLER_1_1119 ();
 sg13g2_fill_2 FILLER_1_1124 ();
 sg13g2_fill_2 FILLER_1_1161 ();
 sg13g2_fill_1 FILLER_1_1163 ();
 sg13g2_decap_8 FILLER_1_1200 ();
 sg13g2_fill_1 FILLER_1_1207 ();
 sg13g2_fill_2 FILLER_1_1234 ();
 sg13g2_fill_1 FILLER_1_1244 ();
 sg13g2_decap_8 FILLER_1_1276 ();
 sg13g2_fill_1 FILLER_1_1293 ();
 sg13g2_decap_4 FILLER_1_1346 ();
 sg13g2_fill_1 FILLER_1_1350 ();
 sg13g2_decap_4 FILLER_1_1355 ();
 sg13g2_fill_2 FILLER_1_1395 ();
 sg13g2_fill_2 FILLER_1_1433 ();
 sg13g2_fill_1 FILLER_1_1435 ();
 sg13g2_decap_4 FILLER_1_1462 ();
 sg13g2_fill_2 FILLER_1_1466 ();
 sg13g2_decap_4 FILLER_1_1498 ();
 sg13g2_fill_2 FILLER_1_1512 ();
 sg13g2_fill_1 FILLER_1_1540 ();
 sg13g2_decap_8 FILLER_1_1545 ();
 sg13g2_decap_4 FILLER_1_1552 ();
 sg13g2_fill_2 FILLER_1_1582 ();
 sg13g2_fill_1 FILLER_1_1584 ();
 sg13g2_decap_4 FILLER_1_1641 ();
 sg13g2_decap_8 FILLER_1_1674 ();
 sg13g2_fill_1 FILLER_1_1681 ();
 sg13g2_decap_8 FILLER_1_1711 ();
 sg13g2_decap_8 FILLER_1_1718 ();
 sg13g2_decap_8 FILLER_1_1725 ();
 sg13g2_decap_8 FILLER_1_1762 ();
 sg13g2_fill_2 FILLER_1_1803 ();
 sg13g2_decap_8 FILLER_1_1815 ();
 sg13g2_fill_2 FILLER_1_1822 ();
 sg13g2_fill_1 FILLER_1_1824 ();
 sg13g2_fill_1 FILLER_1_1856 ();
 sg13g2_decap_8 FILLER_1_1909 ();
 sg13g2_fill_2 FILLER_1_1916 ();
 sg13g2_fill_1 FILLER_1_1918 ();
 sg13g2_fill_2 FILLER_1_1971 ();
 sg13g2_fill_1 FILLER_1_2003 ();
 sg13g2_fill_2 FILLER_1_2040 ();
 sg13g2_decap_8 FILLER_1_2062 ();
 sg13g2_decap_4 FILLER_1_2069 ();
 sg13g2_fill_2 FILLER_1_2139 ();
 sg13g2_fill_1 FILLER_1_2145 ();
 sg13g2_decap_4 FILLER_1_2232 ();
 sg13g2_fill_2 FILLER_1_2266 ();
 sg13g2_decap_4 FILLER_1_2276 ();
 sg13g2_decap_4 FILLER_1_2310 ();
 sg13g2_fill_1 FILLER_1_2314 ();
 sg13g2_decap_4 FILLER_1_2345 ();
 sg13g2_fill_1 FILLER_1_2349 ();
 sg13g2_fill_1 FILLER_1_2381 ();
 sg13g2_fill_2 FILLER_1_2392 ();
 sg13g2_fill_1 FILLER_1_2394 ();
 sg13g2_decap_4 FILLER_1_2421 ();
 sg13g2_fill_2 FILLER_1_2451 ();
 sg13g2_fill_2 FILLER_1_2483 ();
 sg13g2_decap_8 FILLER_1_2525 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_4 FILLER_1_2665 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_fill_2 FILLER_2_35 ();
 sg13g2_fill_1 FILLER_2_37 ();
 sg13g2_fill_1 FILLER_2_48 ();
 sg13g2_fill_2 FILLER_2_69 ();
 sg13g2_fill_1 FILLER_2_90 ();
 sg13g2_decap_4 FILLER_2_156 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_decap_4 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_186 ();
 sg13g2_fill_1 FILLER_2_257 ();
 sg13g2_decap_8 FILLER_2_262 ();
 sg13g2_decap_4 FILLER_2_269 ();
 sg13g2_fill_1 FILLER_2_368 ();
 sg13g2_fill_1 FILLER_2_395 ();
 sg13g2_fill_2 FILLER_2_440 ();
 sg13g2_fill_2 FILLER_2_468 ();
 sg13g2_fill_2 FILLER_2_475 ();
 sg13g2_fill_1 FILLER_2_477 ();
 sg13g2_fill_1 FILLER_2_504 ();
 sg13g2_fill_2 FILLER_2_520 ();
 sg13g2_fill_1 FILLER_2_532 ();
 sg13g2_decap_8 FILLER_2_559 ();
 sg13g2_fill_1 FILLER_2_566 ();
 sg13g2_fill_1 FILLER_2_595 ();
 sg13g2_fill_2 FILLER_2_656 ();
 sg13g2_fill_1 FILLER_2_684 ();
 sg13g2_fill_1 FILLER_2_711 ();
 sg13g2_fill_2 FILLER_2_759 ();
 sg13g2_fill_2 FILLER_2_787 ();
 sg13g2_fill_2 FILLER_2_927 ();
 sg13g2_decap_4 FILLER_2_985 ();
 sg13g2_fill_1 FILLER_2_989 ();
 sg13g2_fill_2 FILLER_2_999 ();
 sg13g2_fill_1 FILLER_2_1001 ();
 sg13g2_decap_4 FILLER_2_1006 ();
 sg13g2_fill_1 FILLER_2_1010 ();
 sg13g2_decap_4 FILLER_2_1015 ();
 sg13g2_fill_1 FILLER_2_1019 ();
 sg13g2_fill_1 FILLER_2_1046 ();
 sg13g2_fill_2 FILLER_2_1105 ();
 sg13g2_fill_2 FILLER_2_1159 ();
 sg13g2_fill_1 FILLER_2_1161 ();
 sg13g2_fill_2 FILLER_2_1202 ();
 sg13g2_fill_1 FILLER_2_1204 ();
 sg13g2_decap_4 FILLER_2_1251 ();
 sg13g2_fill_2 FILLER_2_1255 ();
 sg13g2_decap_4 FILLER_2_1297 ();
 sg13g2_fill_2 FILLER_2_1305 ();
 sg13g2_fill_1 FILLER_2_1307 ();
 sg13g2_fill_2 FILLER_2_1380 ();
 sg13g2_fill_1 FILLER_2_1412 ();
 sg13g2_fill_1 FILLER_2_1439 ();
 sg13g2_decap_4 FILLER_2_1499 ();
 sg13g2_fill_2 FILLER_2_1503 ();
 sg13g2_fill_2 FILLER_2_1519 ();
 sg13g2_fill_1 FILLER_2_1521 ();
 sg13g2_fill_1 FILLER_2_1558 ();
 sg13g2_decap_8 FILLER_2_1585 ();
 sg13g2_decap_4 FILLER_2_1592 ();
 sg13g2_fill_1 FILLER_2_1615 ();
 sg13g2_fill_1 FILLER_2_1645 ();
 sg13g2_fill_2 FILLER_2_1650 ();
 sg13g2_fill_1 FILLER_2_1652 ();
 sg13g2_decap_8 FILLER_2_1660 ();
 sg13g2_decap_4 FILLER_2_1667 ();
 sg13g2_fill_1 FILLER_2_1681 ();
 sg13g2_fill_2 FILLER_2_1690 ();
 sg13g2_decap_4 FILLER_2_1718 ();
 sg13g2_fill_1 FILLER_2_1726 ();
 sg13g2_decap_8 FILLER_2_1769 ();
 sg13g2_fill_2 FILLER_2_1794 ();
 sg13g2_fill_1 FILLER_2_1796 ();
 sg13g2_fill_1 FILLER_2_1895 ();
 sg13g2_decap_8 FILLER_2_1900 ();
 sg13g2_decap_4 FILLER_2_1907 ();
 sg13g2_fill_2 FILLER_2_2002 ();
 sg13g2_decap_8 FILLER_2_2057 ();
 sg13g2_decap_4 FILLER_2_2068 ();
 sg13g2_fill_1 FILLER_2_2072 ();
 sg13g2_fill_2 FILLER_2_2099 ();
 sg13g2_fill_1 FILLER_2_2127 ();
 sg13g2_fill_2 FILLER_2_2158 ();
 sg13g2_fill_1 FILLER_2_2185 ();
 sg13g2_fill_2 FILLER_2_2248 ();
 sg13g2_decap_4 FILLER_2_2276 ();
 sg13g2_fill_2 FILLER_2_2280 ();
 sg13g2_fill_2 FILLER_2_2286 ();
 sg13g2_fill_1 FILLER_2_2288 ();
 sg13g2_fill_2 FILLER_2_2390 ();
 sg13g2_fill_2 FILLER_2_2418 ();
 sg13g2_fill_2 FILLER_2_2498 ();
 sg13g2_fill_1 FILLER_2_2500 ();
 sg13g2_fill_2 FILLER_2_2531 ();
 sg13g2_decap_8 FILLER_2_2546 ();
 sg13g2_decap_8 FILLER_2_2553 ();
 sg13g2_decap_8 FILLER_2_2560 ();
 sg13g2_decap_8 FILLER_2_2567 ();
 sg13g2_decap_8 FILLER_2_2574 ();
 sg13g2_decap_8 FILLER_2_2581 ();
 sg13g2_decap_8 FILLER_2_2588 ();
 sg13g2_decap_8 FILLER_2_2595 ();
 sg13g2_decap_8 FILLER_2_2602 ();
 sg13g2_decap_8 FILLER_2_2609 ();
 sg13g2_decap_8 FILLER_2_2616 ();
 sg13g2_decap_8 FILLER_2_2623 ();
 sg13g2_decap_8 FILLER_2_2630 ();
 sg13g2_decap_8 FILLER_2_2637 ();
 sg13g2_decap_8 FILLER_2_2644 ();
 sg13g2_decap_8 FILLER_2_2651 ();
 sg13g2_decap_8 FILLER_2_2658 ();
 sg13g2_decap_4 FILLER_2_2665 ();
 sg13g2_fill_1 FILLER_2_2669 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_fill_1 FILLER_3_30 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_4 FILLER_3_42 ();
 sg13g2_fill_1 FILLER_3_46 ();
 sg13g2_fill_1 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_4 FILLER_3_151 ();
 sg13g2_fill_2 FILLER_3_155 ();
 sg13g2_decap_4 FILLER_3_193 ();
 sg13g2_fill_2 FILLER_3_197 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_fill_2 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_216 ();
 sg13g2_decap_4 FILLER_3_271 ();
 sg13g2_fill_2 FILLER_3_275 ();
 sg13g2_fill_2 FILLER_3_304 ();
 sg13g2_fill_1 FILLER_3_332 ();
 sg13g2_fill_1 FILLER_3_343 ();
 sg13g2_fill_2 FILLER_3_363 ();
 sg13g2_decap_4 FILLER_3_384 ();
 sg13g2_fill_2 FILLER_3_388 ();
 sg13g2_decap_4 FILLER_3_435 ();
 sg13g2_fill_1 FILLER_3_439 ();
 sg13g2_fill_1 FILLER_3_445 ();
 sg13g2_fill_2 FILLER_3_460 ();
 sg13g2_fill_1 FILLER_3_462 ();
 sg13g2_fill_2 FILLER_3_493 ();
 sg13g2_fill_2 FILLER_3_544 ();
 sg13g2_decap_4 FILLER_3_550 ();
 sg13g2_fill_1 FILLER_3_580 ();
 sg13g2_fill_1 FILLER_3_613 ();
 sg13g2_fill_2 FILLER_3_629 ();
 sg13g2_fill_2 FILLER_3_720 ();
 sg13g2_decap_8 FILLER_3_766 ();
 sg13g2_decap_8 FILLER_3_773 ();
 sg13g2_decap_4 FILLER_3_780 ();
 sg13g2_fill_2 FILLER_3_784 ();
 sg13g2_fill_2 FILLER_3_822 ();
 sg13g2_fill_1 FILLER_3_897 ();
 sg13g2_fill_2 FILLER_3_945 ();
 sg13g2_fill_1 FILLER_3_964 ();
 sg13g2_decap_8 FILLER_3_974 ();
 sg13g2_decap_4 FILLER_3_1012 ();
 sg13g2_fill_1 FILLER_3_1016 ();
 sg13g2_fill_2 FILLER_3_1043 ();
 sg13g2_fill_1 FILLER_3_1045 ();
 sg13g2_decap_4 FILLER_3_1076 ();
 sg13g2_fill_2 FILLER_3_1089 ();
 sg13g2_fill_1 FILLER_3_1091 ();
 sg13g2_fill_2 FILLER_3_1122 ();
 sg13g2_decap_4 FILLER_3_1198 ();
 sg13g2_fill_2 FILLER_3_1212 ();
 sg13g2_fill_1 FILLER_3_1218 ();
 sg13g2_fill_1 FILLER_3_1255 ();
 sg13g2_decap_4 FILLER_3_1287 ();
 sg13g2_fill_1 FILLER_3_1291 ();
 sg13g2_decap_8 FILLER_3_1313 ();
 sg13g2_decap_8 FILLER_3_1320 ();
 sg13g2_decap_4 FILLER_3_1335 ();
 sg13g2_decap_8 FILLER_3_1349 ();
 sg13g2_fill_1 FILLER_3_1356 ();
 sg13g2_fill_1 FILLER_3_1393 ();
 sg13g2_fill_1 FILLER_3_1420 ();
 sg13g2_fill_1 FILLER_3_1425 ();
 sg13g2_decap_8 FILLER_3_1514 ();
 sg13g2_fill_1 FILLER_3_1521 ();
 sg13g2_fill_1 FILLER_3_1587 ();
 sg13g2_fill_1 FILLER_3_1615 ();
 sg13g2_decap_8 FILLER_3_1676 ();
 sg13g2_decap_8 FILLER_3_1683 ();
 sg13g2_decap_8 FILLER_3_1690 ();
 sg13g2_fill_1 FILLER_3_1697 ();
 sg13g2_fill_2 FILLER_3_1702 ();
 sg13g2_fill_1 FILLER_3_1704 ();
 sg13g2_fill_2 FILLER_3_1718 ();
 sg13g2_decap_4 FILLER_3_1733 ();
 sg13g2_decap_8 FILLER_3_1773 ();
 sg13g2_fill_2 FILLER_3_1791 ();
 sg13g2_fill_1 FILLER_3_1793 ();
 sg13g2_fill_1 FILLER_3_1820 ();
 sg13g2_decap_8 FILLER_3_1884 ();
 sg13g2_fill_2 FILLER_3_1891 ();
 sg13g2_fill_1 FILLER_3_1893 ();
 sg13g2_decap_8 FILLER_3_1907 ();
 sg13g2_fill_2 FILLER_3_1914 ();
 sg13g2_fill_2 FILLER_3_1934 ();
 sg13g2_fill_1 FILLER_3_1936 ();
 sg13g2_fill_1 FILLER_3_1958 ();
 sg13g2_decap_8 FILLER_3_1999 ();
 sg13g2_fill_2 FILLER_3_2006 ();
 sg13g2_fill_1 FILLER_3_2008 ();
 sg13g2_fill_1 FILLER_3_2019 ();
 sg13g2_fill_2 FILLER_3_2041 ();
 sg13g2_fill_2 FILLER_3_2099 ();
 sg13g2_fill_1 FILLER_3_2178 ();
 sg13g2_fill_1 FILLER_3_2238 ();
 sg13g2_fill_1 FILLER_3_2265 ();
 sg13g2_fill_2 FILLER_3_2309 ();
 sg13g2_decap_8 FILLER_3_2321 ();
 sg13g2_decap_8 FILLER_3_2328 ();
 sg13g2_decap_8 FILLER_3_2335 ();
 sg13g2_fill_2 FILLER_3_2342 ();
 sg13g2_fill_1 FILLER_3_2344 ();
 sg13g2_decap_4 FILLER_3_2440 ();
 sg13g2_fill_1 FILLER_3_2467 ();
 sg13g2_fill_2 FILLER_3_2498 ();
 sg13g2_decap_8 FILLER_3_2544 ();
 sg13g2_fill_1 FILLER_3_2551 ();
 sg13g2_decap_8 FILLER_3_2556 ();
 sg13g2_decap_8 FILLER_3_2563 ();
 sg13g2_decap_8 FILLER_3_2570 ();
 sg13g2_decap_8 FILLER_3_2577 ();
 sg13g2_decap_8 FILLER_3_2584 ();
 sg13g2_decap_8 FILLER_3_2591 ();
 sg13g2_decap_8 FILLER_3_2598 ();
 sg13g2_decap_8 FILLER_3_2605 ();
 sg13g2_decap_8 FILLER_3_2612 ();
 sg13g2_decap_8 FILLER_3_2619 ();
 sg13g2_decap_8 FILLER_3_2626 ();
 sg13g2_decap_8 FILLER_3_2633 ();
 sg13g2_decap_8 FILLER_3_2640 ();
 sg13g2_decap_8 FILLER_3_2647 ();
 sg13g2_decap_8 FILLER_3_2654 ();
 sg13g2_decap_8 FILLER_3_2661 ();
 sg13g2_fill_2 FILLER_3_2668 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_fill_2 FILLER_4_21 ();
 sg13g2_fill_1 FILLER_4_23 ();
 sg13g2_decap_4 FILLER_4_50 ();
 sg13g2_fill_2 FILLER_4_101 ();
 sg13g2_fill_1 FILLER_4_119 ();
 sg13g2_fill_2 FILLER_4_124 ();
 sg13g2_fill_1 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_157 ();
 sg13g2_decap_8 FILLER_4_164 ();
 sg13g2_decap_8 FILLER_4_171 ();
 sg13g2_decap_4 FILLER_4_178 ();
 sg13g2_decap_4 FILLER_4_192 ();
 sg13g2_fill_1 FILLER_4_196 ();
 sg13g2_decap_4 FILLER_4_209 ();
 sg13g2_fill_1 FILLER_4_213 ();
 sg13g2_fill_2 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_4 FILLER_4_232 ();
 sg13g2_decap_8 FILLER_4_250 ();
 sg13g2_decap_8 FILLER_4_257 ();
 sg13g2_fill_2 FILLER_4_264 ();
 sg13g2_fill_1 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_302 ();
 sg13g2_decap_4 FILLER_4_309 ();
 sg13g2_fill_1 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_323 ();
 sg13g2_fill_2 FILLER_4_341 ();
 sg13g2_fill_1 FILLER_4_343 ();
 sg13g2_fill_1 FILLER_4_349 ();
 sg13g2_fill_1 FILLER_4_364 ();
 sg13g2_fill_2 FILLER_4_402 ();
 sg13g2_fill_1 FILLER_4_404 ();
 sg13g2_fill_2 FILLER_4_409 ();
 sg13g2_fill_2 FILLER_4_421 ();
 sg13g2_fill_1 FILLER_4_428 ();
 sg13g2_decap_4 FILLER_4_433 ();
 sg13g2_decap_4 FILLER_4_447 ();
 sg13g2_decap_8 FILLER_4_456 ();
 sg13g2_decap_4 FILLER_4_463 ();
 sg13g2_fill_1 FILLER_4_504 ();
 sg13g2_fill_2 FILLER_4_537 ();
 sg13g2_fill_1 FILLER_4_539 ();
 sg13g2_decap_4 FILLER_4_544 ();
 sg13g2_fill_2 FILLER_4_558 ();
 sg13g2_fill_1 FILLER_4_560 ();
 sg13g2_fill_2 FILLER_4_565 ();
 sg13g2_fill_1 FILLER_4_567 ();
 sg13g2_fill_2 FILLER_4_598 ();
 sg13g2_fill_2 FILLER_4_631 ();
 sg13g2_fill_1 FILLER_4_633 ();
 sg13g2_fill_2 FILLER_4_643 ();
 sg13g2_fill_1 FILLER_4_645 ();
 sg13g2_decap_4 FILLER_4_672 ();
 sg13g2_fill_2 FILLER_4_676 ();
 sg13g2_decap_4 FILLER_4_682 ();
 sg13g2_fill_1 FILLER_4_691 ();
 sg13g2_fill_1 FILLER_4_697 ();
 sg13g2_fill_1 FILLER_4_726 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_fill_1 FILLER_4_784 ();
 sg13g2_fill_1 FILLER_4_836 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_fill_2 FILLER_4_854 ();
 sg13g2_decap_4 FILLER_4_864 ();
 sg13g2_fill_1 FILLER_4_882 ();
 sg13g2_fill_1 FILLER_4_909 ();
 sg13g2_decap_8 FILLER_4_914 ();
 sg13g2_fill_2 FILLER_4_921 ();
 sg13g2_fill_1 FILLER_4_932 ();
 sg13g2_fill_1 FILLER_4_950 ();
 sg13g2_fill_2 FILLER_4_963 ();
 sg13g2_fill_1 FILLER_4_965 ();
 sg13g2_fill_2 FILLER_4_1004 ();
 sg13g2_decap_4 FILLER_4_1019 ();
 sg13g2_fill_1 FILLER_4_1023 ();
 sg13g2_decap_4 FILLER_4_1028 ();
 sg13g2_fill_1 FILLER_4_1032 ();
 sg13g2_fill_1 FILLER_4_1063 ();
 sg13g2_decap_8 FILLER_4_1072 ();
 sg13g2_decap_4 FILLER_4_1079 ();
 sg13g2_fill_1 FILLER_4_1083 ();
 sg13g2_fill_2 FILLER_4_1126 ();
 sg13g2_fill_1 FILLER_4_1128 ();
 sg13g2_decap_8 FILLER_4_1211 ();
 sg13g2_fill_2 FILLER_4_1218 ();
 sg13g2_fill_1 FILLER_4_1220 ();
 sg13g2_fill_2 FILLER_4_1225 ();
 sg13g2_fill_1 FILLER_4_1227 ();
 sg13g2_decap_8 FILLER_4_1249 ();
 sg13g2_decap_8 FILLER_4_1256 ();
 sg13g2_fill_2 FILLER_4_1263 ();
 sg13g2_fill_1 FILLER_4_1265 ();
 sg13g2_fill_2 FILLER_4_1302 ();
 sg13g2_fill_1 FILLER_4_1304 ();
 sg13g2_decap_8 FILLER_4_1341 ();
 sg13g2_decap_8 FILLER_4_1348 ();
 sg13g2_decap_8 FILLER_4_1355 ();
 sg13g2_fill_1 FILLER_4_1366 ();
 sg13g2_decap_8 FILLER_4_1371 ();
 sg13g2_decap_8 FILLER_4_1378 ();
 sg13g2_decap_8 FILLER_4_1385 ();
 sg13g2_fill_2 FILLER_4_1392 ();
 sg13g2_fill_2 FILLER_4_1398 ();
 sg13g2_fill_1 FILLER_4_1400 ();
 sg13g2_decap_8 FILLER_4_1405 ();
 sg13g2_decap_8 FILLER_4_1412 ();
 sg13g2_decap_4 FILLER_4_1429 ();
 sg13g2_fill_1 FILLER_4_1433 ();
 sg13g2_fill_2 FILLER_4_1438 ();
 sg13g2_fill_2 FILLER_4_1450 ();
 sg13g2_fill_1 FILLER_4_1452 ();
 sg13g2_fill_1 FILLER_4_1457 ();
 sg13g2_fill_1 FILLER_4_1462 ();
 sg13g2_fill_2 FILLER_4_1489 ();
 sg13g2_decap_8 FILLER_4_1503 ();
 sg13g2_fill_1 FILLER_4_1510 ();
 sg13g2_decap_4 FILLER_4_1519 ();
 sg13g2_fill_1 FILLER_4_1543 ();
 sg13g2_fill_2 FILLER_4_1593 ();
 sg13g2_fill_2 FILLER_4_1614 ();
 sg13g2_fill_1 FILLER_4_1619 ();
 sg13g2_decap_8 FILLER_4_1650 ();
 sg13g2_decap_8 FILLER_4_1657 ();
 sg13g2_fill_2 FILLER_4_1664 ();
 sg13g2_fill_1 FILLER_4_1666 ();
 sg13g2_fill_2 FILLER_4_1703 ();
 sg13g2_fill_1 FILLER_4_1705 ();
 sg13g2_fill_1 FILLER_4_1710 ();
 sg13g2_fill_1 FILLER_4_1789 ();
 sg13g2_fill_1 FILLER_4_1795 ();
 sg13g2_fill_1 FILLER_4_1802 ();
 sg13g2_fill_1 FILLER_4_1813 ();
 sg13g2_fill_2 FILLER_4_1819 ();
 sg13g2_fill_1 FILLER_4_1821 ();
 sg13g2_fill_2 FILLER_4_1831 ();
 sg13g2_fill_1 FILLER_4_1833 ();
 sg13g2_decap_4 FILLER_4_1839 ();
 sg13g2_fill_1 FILLER_4_1843 ();
 sg13g2_fill_1 FILLER_4_1887 ();
 sg13g2_decap_8 FILLER_4_1901 ();
 sg13g2_fill_1 FILLER_4_1908 ();
 sg13g2_decap_4 FILLER_4_1936 ();
 sg13g2_decap_4 FILLER_4_1950 ();
 sg13g2_decap_8 FILLER_4_1958 ();
 sg13g2_decap_8 FILLER_4_1969 ();
 sg13g2_fill_2 FILLER_4_1976 ();
 sg13g2_decap_8 FILLER_4_1988 ();
 sg13g2_decap_8 FILLER_4_1995 ();
 sg13g2_decap_8 FILLER_4_2032 ();
 sg13g2_fill_2 FILLER_4_2039 ();
 sg13g2_fill_1 FILLER_4_2041 ();
 sg13g2_decap_8 FILLER_4_2063 ();
 sg13g2_fill_1 FILLER_4_2070 ();
 sg13g2_decap_8 FILLER_4_2097 ();
 sg13g2_fill_2 FILLER_4_2104 ();
 sg13g2_fill_1 FILLER_4_2106 ();
 sg13g2_fill_1 FILLER_4_2205 ();
 sg13g2_fill_2 FILLER_4_2214 ();
 sg13g2_fill_1 FILLER_4_2216 ();
 sg13g2_fill_2 FILLER_4_2225 ();
 sg13g2_fill_2 FILLER_4_2266 ();
 sg13g2_fill_2 FILLER_4_2297 ();
 sg13g2_fill_1 FILLER_4_2309 ();
 sg13g2_fill_2 FILLER_4_2331 ();
 sg13g2_fill_1 FILLER_4_2333 ();
 sg13g2_decap_8 FILLER_4_2347 ();
 sg13g2_fill_1 FILLER_4_2354 ();
 sg13g2_fill_2 FILLER_4_2365 ();
 sg13g2_decap_8 FILLER_4_2388 ();
 sg13g2_decap_4 FILLER_4_2395 ();
 sg13g2_decap_4 FILLER_4_2409 ();
 sg13g2_decap_4 FILLER_4_2423 ();
 sg13g2_fill_1 FILLER_4_2427 ();
 sg13g2_decap_8 FILLER_4_2432 ();
 sg13g2_decap_4 FILLER_4_2439 ();
 sg13g2_fill_1 FILLER_4_2443 ();
 sg13g2_decap_8 FILLER_4_2488 ();
 sg13g2_fill_1 FILLER_4_2495 ();
 sg13g2_fill_1 FILLER_4_2506 ();
 sg13g2_decap_4 FILLER_4_2532 ();
 sg13g2_fill_1 FILLER_4_2536 ();
 sg13g2_fill_1 FILLER_4_2547 ();
 sg13g2_decap_8 FILLER_4_2574 ();
 sg13g2_decap_8 FILLER_4_2581 ();
 sg13g2_decap_8 FILLER_4_2588 ();
 sg13g2_decap_8 FILLER_4_2595 ();
 sg13g2_decap_8 FILLER_4_2602 ();
 sg13g2_decap_8 FILLER_4_2609 ();
 sg13g2_decap_8 FILLER_4_2616 ();
 sg13g2_decap_8 FILLER_4_2623 ();
 sg13g2_decap_8 FILLER_4_2630 ();
 sg13g2_decap_8 FILLER_4_2637 ();
 sg13g2_decap_8 FILLER_4_2644 ();
 sg13g2_decap_8 FILLER_4_2651 ();
 sg13g2_decap_8 FILLER_4_2658 ();
 sg13g2_decap_4 FILLER_4_2665 ();
 sg13g2_fill_1 FILLER_4_2669 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_7 ();
 sg13g2_fill_1 FILLER_5_13 ();
 sg13g2_fill_2 FILLER_5_39 ();
 sg13g2_fill_1 FILLER_5_41 ();
 sg13g2_decap_8 FILLER_5_86 ();
 sg13g2_decap_8 FILLER_5_93 ();
 sg13g2_fill_2 FILLER_5_100 ();
 sg13g2_fill_1 FILLER_5_106 ();
 sg13g2_fill_1 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_fill_1 FILLER_5_135 ();
 sg13g2_fill_1 FILLER_5_140 ();
 sg13g2_decap_4 FILLER_5_175 ();
 sg13g2_fill_1 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_255 ();
 sg13g2_decap_8 FILLER_5_262 ();
 sg13g2_decap_4 FILLER_5_269 ();
 sg13g2_fill_1 FILLER_5_282 ();
 sg13g2_fill_2 FILLER_5_288 ();
 sg13g2_fill_2 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_307 ();
 sg13g2_fill_2 FILLER_5_314 ();
 sg13g2_fill_1 FILLER_5_330 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_359 ();
 sg13g2_fill_2 FILLER_5_391 ();
 sg13g2_fill_2 FILLER_5_409 ();
 sg13g2_fill_2 FILLER_5_421 ();
 sg13g2_fill_1 FILLER_5_423 ();
 sg13g2_fill_2 FILLER_5_433 ();
 sg13g2_fill_2 FILLER_5_448 ();
 sg13g2_decap_4 FILLER_5_460 ();
 sg13g2_fill_1 FILLER_5_464 ();
 sg13g2_fill_1 FILLER_5_470 ();
 sg13g2_fill_1 FILLER_5_489 ();
 sg13g2_decap_8 FILLER_5_505 ();
 sg13g2_fill_2 FILLER_5_512 ();
 sg13g2_decap_4 FILLER_5_522 ();
 sg13g2_fill_1 FILLER_5_535 ();
 sg13g2_decap_8 FILLER_5_556 ();
 sg13g2_decap_8 FILLER_5_563 ();
 sg13g2_fill_2 FILLER_5_570 ();
 sg13g2_fill_1 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_583 ();
 sg13g2_fill_2 FILLER_5_589 ();
 sg13g2_fill_1 FILLER_5_591 ();
 sg13g2_fill_1 FILLER_5_602 ();
 sg13g2_fill_1 FILLER_5_641 ();
 sg13g2_fill_2 FILLER_5_647 ();
 sg13g2_fill_2 FILLER_5_659 ();
 sg13g2_decap_8 FILLER_5_674 ();
 sg13g2_decap_8 FILLER_5_681 ();
 sg13g2_decap_4 FILLER_5_693 ();
 sg13g2_fill_1 FILLER_5_728 ();
 sg13g2_fill_2 FILLER_5_737 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_4 FILLER_5_809 ();
 sg13g2_fill_2 FILLER_5_813 ();
 sg13g2_decap_4 FILLER_5_825 ();
 sg13g2_decap_8 FILLER_5_833 ();
 sg13g2_decap_8 FILLER_5_840 ();
 sg13g2_fill_1 FILLER_5_847 ();
 sg13g2_decap_4 FILLER_5_852 ();
 sg13g2_fill_1 FILLER_5_856 ();
 sg13g2_decap_8 FILLER_5_867 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_fill_1 FILLER_5_911 ();
 sg13g2_decap_8 FILLER_5_926 ();
 sg13g2_decap_8 FILLER_5_933 ();
 sg13g2_fill_2 FILLER_5_940 ();
 sg13g2_fill_2 FILLER_5_947 ();
 sg13g2_fill_1 FILLER_5_957 ();
 sg13g2_decap_4 FILLER_5_962 ();
 sg13g2_fill_1 FILLER_5_976 ();
 sg13g2_fill_2 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1080 ();
 sg13g2_fill_2 FILLER_5_1087 ();
 sg13g2_fill_2 FILLER_5_1118 ();
 sg13g2_fill_1 FILLER_5_1120 ();
 sg13g2_decap_8 FILLER_5_1142 ();
 sg13g2_decap_4 FILLER_5_1149 ();
 sg13g2_fill_1 FILLER_5_1153 ();
 sg13g2_decap_8 FILLER_5_1158 ();
 sg13g2_decap_8 FILLER_5_1165 ();
 sg13g2_decap_8 FILLER_5_1172 ();
 sg13g2_decap_4 FILLER_5_1179 ();
 sg13g2_decap_4 FILLER_5_1187 ();
 sg13g2_fill_1 FILLER_5_1191 ();
 sg13g2_decap_8 FILLER_5_1196 ();
 sg13g2_decap_8 FILLER_5_1203 ();
 sg13g2_decap_8 FILLER_5_1210 ();
 sg13g2_decap_8 FILLER_5_1217 ();
 sg13g2_decap_4 FILLER_5_1224 ();
 sg13g2_decap_4 FILLER_5_1249 ();
 sg13g2_fill_1 FILLER_5_1253 ();
 sg13g2_decap_8 FILLER_5_1294 ();
 sg13g2_fill_1 FILLER_5_1301 ();
 sg13g2_decap_8 FILLER_5_1306 ();
 sg13g2_fill_2 FILLER_5_1313 ();
 sg13g2_fill_1 FILLER_5_1315 ();
 sg13g2_fill_2 FILLER_5_1320 ();
 sg13g2_decap_8 FILLER_5_1326 ();
 sg13g2_decap_8 FILLER_5_1333 ();
 sg13g2_decap_4 FILLER_5_1340 ();
 sg13g2_fill_1 FILLER_5_1344 ();
 sg13g2_fill_2 FILLER_5_1385 ();
 sg13g2_fill_2 FILLER_5_1423 ();
 sg13g2_fill_2 FILLER_5_1435 ();
 sg13g2_fill_1 FILLER_5_1437 ();
 sg13g2_decap_4 FILLER_5_1442 ();
 sg13g2_decap_4 FILLER_5_1456 ();
 sg13g2_fill_2 FILLER_5_1474 ();
 sg13g2_decap_8 FILLER_5_1484 ();
 sg13g2_decap_4 FILLER_5_1501 ();
 sg13g2_fill_1 FILLER_5_1505 ();
 sg13g2_decap_4 FILLER_5_1519 ();
 sg13g2_fill_1 FILLER_5_1523 ();
 sg13g2_fill_2 FILLER_5_1528 ();
 sg13g2_decap_8 FILLER_5_1539 ();
 sg13g2_decap_8 FILLER_5_1546 ();
 sg13g2_fill_1 FILLER_5_1557 ();
 sg13g2_fill_1 FILLER_5_1568 ();
 sg13g2_fill_2 FILLER_5_1599 ();
 sg13g2_fill_1 FILLER_5_1601 ();
 sg13g2_decap_8 FILLER_5_1653 ();
 sg13g2_fill_2 FILLER_5_1660 ();
 sg13g2_fill_1 FILLER_5_1662 ();
 sg13g2_decap_8 FILLER_5_1677 ();
 sg13g2_decap_4 FILLER_5_1684 ();
 sg13g2_fill_2 FILLER_5_1688 ();
 sg13g2_decap_8 FILLER_5_1694 ();
 sg13g2_decap_4 FILLER_5_1701 ();
 sg13g2_fill_2 FILLER_5_1741 ();
 sg13g2_fill_1 FILLER_5_1756 ();
 sg13g2_decap_4 FILLER_5_1763 ();
 sg13g2_decap_8 FILLER_5_1772 ();
 sg13g2_decap_8 FILLER_5_1779 ();
 sg13g2_decap_8 FILLER_5_1821 ();
 sg13g2_decap_8 FILLER_5_1828 ();
 sg13g2_fill_2 FILLER_5_1835 ();
 sg13g2_fill_2 FILLER_5_1857 ();
 sg13g2_fill_2 FILLER_5_1889 ();
 sg13g2_fill_1 FILLER_5_1891 ();
 sg13g2_decap_4 FILLER_5_1897 ();
 sg13g2_decap_8 FILLER_5_1905 ();
 sg13g2_decap_8 FILLER_5_1912 ();
 sg13g2_fill_2 FILLER_5_1919 ();
 sg13g2_fill_1 FILLER_5_1921 ();
 sg13g2_decap_8 FILLER_5_1926 ();
 sg13g2_decap_4 FILLER_5_1933 ();
 sg13g2_fill_2 FILLER_5_1937 ();
 sg13g2_decap_8 FILLER_5_1985 ();
 sg13g2_decap_4 FILLER_5_1992 ();
 sg13g2_fill_2 FILLER_5_1996 ();
 sg13g2_decap_8 FILLER_5_2096 ();
 sg13g2_decap_8 FILLER_5_2103 ();
 sg13g2_fill_1 FILLER_5_2110 ();
 sg13g2_fill_2 FILLER_5_2119 ();
 sg13g2_fill_1 FILLER_5_2121 ();
 sg13g2_fill_1 FILLER_5_2126 ();
 sg13g2_fill_2 FILLER_5_2150 ();
 sg13g2_fill_1 FILLER_5_2156 ();
 sg13g2_decap_4 FILLER_5_2199 ();
 sg13g2_fill_1 FILLER_5_2221 ();
 sg13g2_fill_1 FILLER_5_2230 ();
 sg13g2_decap_8 FILLER_5_2284 ();
 sg13g2_decap_8 FILLER_5_2291 ();
 sg13g2_decap_8 FILLER_5_2298 ();
 sg13g2_fill_2 FILLER_5_2305 ();
 sg13g2_decap_8 FILLER_5_2343 ();
 sg13g2_decap_8 FILLER_5_2350 ();
 sg13g2_decap_4 FILLER_5_2357 ();
 sg13g2_fill_2 FILLER_5_2361 ();
 sg13g2_decap_8 FILLER_5_2397 ();
 sg13g2_decap_8 FILLER_5_2404 ();
 sg13g2_decap_4 FILLER_5_2411 ();
 sg13g2_decap_4 FILLER_5_2425 ();
 sg13g2_fill_2 FILLER_5_2450 ();
 sg13g2_fill_2 FILLER_5_2476 ();
 sg13g2_fill_2 FILLER_5_2496 ();
 sg13g2_fill_1 FILLER_5_2498 ();
 sg13g2_fill_2 FILLER_5_2535 ();
 sg13g2_fill_1 FILLER_5_2537 ();
 sg13g2_decap_4 FILLER_5_2561 ();
 sg13g2_fill_1 FILLER_5_2565 ();
 sg13g2_decap_8 FILLER_5_2570 ();
 sg13g2_decap_8 FILLER_5_2577 ();
 sg13g2_decap_8 FILLER_5_2584 ();
 sg13g2_decap_8 FILLER_5_2591 ();
 sg13g2_decap_8 FILLER_5_2598 ();
 sg13g2_decap_8 FILLER_5_2605 ();
 sg13g2_decap_8 FILLER_5_2612 ();
 sg13g2_decap_8 FILLER_5_2619 ();
 sg13g2_decap_8 FILLER_5_2626 ();
 sg13g2_decap_8 FILLER_5_2633 ();
 sg13g2_decap_8 FILLER_5_2640 ();
 sg13g2_decap_8 FILLER_5_2647 ();
 sg13g2_decap_8 FILLER_5_2654 ();
 sg13g2_decap_8 FILLER_5_2661 ();
 sg13g2_fill_2 FILLER_5_2668 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_1 FILLER_6_4 ();
 sg13g2_decap_8 FILLER_6_31 ();
 sg13g2_decap_8 FILLER_6_38 ();
 sg13g2_decap_8 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_decap_4 FILLER_6_58 ();
 sg13g2_fill_1 FILLER_6_62 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_96 ();
 sg13g2_fill_2 FILLER_6_103 ();
 sg13g2_fill_1 FILLER_6_125 ();
 sg13g2_fill_2 FILLER_6_140 ();
 sg13g2_fill_1 FILLER_6_142 ();
 sg13g2_fill_1 FILLER_6_147 ();
 sg13g2_fill_1 FILLER_6_158 ();
 sg13g2_fill_2 FILLER_6_167 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_fill_1 FILLER_6_236 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_fill_1 FILLER_6_247 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_decap_4 FILLER_6_257 ();
 sg13g2_fill_1 FILLER_6_300 ();
 sg13g2_fill_2 FILLER_6_305 ();
 sg13g2_fill_1 FILLER_6_337 ();
 sg13g2_fill_2 FILLER_6_348 ();
 sg13g2_fill_1 FILLER_6_350 ();
 sg13g2_fill_2 FILLER_6_360 ();
 sg13g2_fill_2 FILLER_6_376 ();
 sg13g2_fill_2 FILLER_6_382 ();
 sg13g2_fill_1 FILLER_6_384 ();
 sg13g2_fill_2 FILLER_6_400 ();
 sg13g2_fill_1 FILLER_6_406 ();
 sg13g2_fill_2 FILLER_6_412 ();
 sg13g2_fill_1 FILLER_6_459 ();
 sg13g2_fill_2 FILLER_6_480 ();
 sg13g2_fill_2 FILLER_6_497 ();
 sg13g2_fill_1 FILLER_6_499 ();
 sg13g2_decap_8 FILLER_6_508 ();
 sg13g2_fill_2 FILLER_6_515 ();
 sg13g2_fill_1 FILLER_6_517 ();
 sg13g2_decap_4 FILLER_6_522 ();
 sg13g2_decap_8 FILLER_6_557 ();
 sg13g2_decap_8 FILLER_6_564 ();
 sg13g2_decap_4 FILLER_6_571 ();
 sg13g2_fill_1 FILLER_6_575 ();
 sg13g2_fill_2 FILLER_6_590 ();
 sg13g2_fill_1 FILLER_6_597 ();
 sg13g2_fill_1 FILLER_6_608 ();
 sg13g2_fill_1 FILLER_6_615 ();
 sg13g2_decap_8 FILLER_6_622 ();
 sg13g2_decap_8 FILLER_6_635 ();
 sg13g2_fill_1 FILLER_6_642 ();
 sg13g2_fill_1 FILLER_6_692 ();
 sg13g2_fill_1 FILLER_6_697 ();
 sg13g2_fill_2 FILLER_6_703 ();
 sg13g2_fill_1 FILLER_6_705 ();
 sg13g2_fill_1 FILLER_6_715 ();
 sg13g2_fill_2 FILLER_6_726 ();
 sg13g2_fill_2 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_778 ();
 sg13g2_fill_2 FILLER_6_785 ();
 sg13g2_fill_1 FILLER_6_787 ();
 sg13g2_decap_4 FILLER_6_814 ();
 sg13g2_fill_1 FILLER_6_818 ();
 sg13g2_fill_1 FILLER_6_827 ();
 sg13g2_decap_8 FILLER_6_878 ();
 sg13g2_decap_4 FILLER_6_885 ();
 sg13g2_fill_1 FILLER_6_889 ();
 sg13g2_decap_8 FILLER_6_921 ();
 sg13g2_decap_8 FILLER_6_928 ();
 sg13g2_decap_8 FILLER_6_935 ();
 sg13g2_decap_8 FILLER_6_942 ();
 sg13g2_fill_2 FILLER_6_949 ();
 sg13g2_fill_2 FILLER_6_977 ();
 sg13g2_fill_1 FILLER_6_979 ();
 sg13g2_decap_4 FILLER_6_989 ();
 sg13g2_fill_1 FILLER_6_993 ();
 sg13g2_fill_1 FILLER_6_1051 ();
 sg13g2_fill_1 FILLER_6_1078 ();
 sg13g2_fill_1 FILLER_6_1087 ();
 sg13g2_fill_2 FILLER_6_1093 ();
 sg13g2_fill_2 FILLER_6_1121 ();
 sg13g2_fill_2 FILLER_6_1149 ();
 sg13g2_decap_4 FILLER_6_1155 ();
 sg13g2_fill_2 FILLER_6_1159 ();
 sg13g2_decap_8 FILLER_6_1197 ();
 sg13g2_fill_2 FILLER_6_1204 ();
 sg13g2_fill_2 FILLER_6_1242 ();
 sg13g2_decap_4 FILLER_6_1265 ();
 sg13g2_fill_1 FILLER_6_1269 ();
 sg13g2_decap_4 FILLER_6_1274 ();
 sg13g2_fill_2 FILLER_6_1299 ();
 sg13g2_fill_1 FILLER_6_1311 ();
 sg13g2_decap_8 FILLER_6_1338 ();
 sg13g2_decap_8 FILLER_6_1345 ();
 sg13g2_fill_2 FILLER_6_1352 ();
 sg13g2_decap_8 FILLER_6_1390 ();
 sg13g2_fill_2 FILLER_6_1427 ();
 sg13g2_fill_1 FILLER_6_1429 ();
 sg13g2_decap_8 FILLER_6_1491 ();
 sg13g2_decap_8 FILLER_6_1498 ();
 sg13g2_fill_2 FILLER_6_1505 ();
 sg13g2_decap_4 FILLER_6_1543 ();
 sg13g2_fill_2 FILLER_6_1547 ();
 sg13g2_fill_2 FILLER_6_1608 ();
 sg13g2_fill_2 FILLER_6_1632 ();
 sg13g2_decap_8 FILLER_6_1644 ();
 sg13g2_fill_2 FILLER_6_1651 ();
 sg13g2_fill_1 FILLER_6_1653 ();
 sg13g2_fill_1 FILLER_6_1690 ();
 sg13g2_fill_2 FILLER_6_1717 ();
 sg13g2_fill_1 FILLER_6_1719 ();
 sg13g2_fill_2 FILLER_6_1749 ();
 sg13g2_fill_1 FILLER_6_1764 ();
 sg13g2_decap_8 FILLER_6_1775 ();
 sg13g2_fill_2 FILLER_6_1796 ();
 sg13g2_decap_8 FILLER_6_1832 ();
 sg13g2_decap_4 FILLER_6_1839 ();
 sg13g2_fill_2 FILLER_6_1904 ();
 sg13g2_decap_8 FILLER_6_1916 ();
 sg13g2_fill_2 FILLER_6_1923 ();
 sg13g2_decap_4 FILLER_6_1946 ();
 sg13g2_fill_2 FILLER_6_1950 ();
 sg13g2_decap_8 FILLER_6_1956 ();
 sg13g2_decap_4 FILLER_6_1963 ();
 sg13g2_fill_2 FILLER_6_1967 ();
 sg13g2_decap_4 FILLER_6_1977 ();
 sg13g2_fill_2 FILLER_6_1981 ();
 sg13g2_decap_8 FILLER_6_1987 ();
 sg13g2_decap_8 FILLER_6_1994 ();
 sg13g2_fill_2 FILLER_6_2001 ();
 sg13g2_fill_1 FILLER_6_2003 ();
 sg13g2_fill_2 FILLER_6_2008 ();
 sg13g2_fill_1 FILLER_6_2010 ();
 sg13g2_decap_4 FILLER_6_2016 ();
 sg13g2_fill_1 FILLER_6_2020 ();
 sg13g2_decap_4 FILLER_6_2031 ();
 sg13g2_fill_1 FILLER_6_2035 ();
 sg13g2_decap_4 FILLER_6_2040 ();
 sg13g2_fill_1 FILLER_6_2044 ();
 sg13g2_fill_2 FILLER_6_2062 ();
 sg13g2_fill_1 FILLER_6_2078 ();
 sg13g2_fill_2 FILLER_6_2083 ();
 sg13g2_fill_1 FILLER_6_2085 ();
 sg13g2_decap_8 FILLER_6_2107 ();
 sg13g2_decap_8 FILLER_6_2114 ();
 sg13g2_decap_4 FILLER_6_2121 ();
 sg13g2_fill_2 FILLER_6_2125 ();
 sg13g2_fill_2 FILLER_6_2182 ();
 sg13g2_decap_8 FILLER_6_2205 ();
 sg13g2_fill_2 FILLER_6_2238 ();
 sg13g2_fill_1 FILLER_6_2271 ();
 sg13g2_decap_4 FILLER_6_2311 ();
 sg13g2_fill_1 FILLER_6_2344 ();
 sg13g2_decap_8 FILLER_6_2378 ();
 sg13g2_decap_8 FILLER_6_2446 ();
 sg13g2_fill_2 FILLER_6_2453 ();
 sg13g2_decap_8 FILLER_6_2511 ();
 sg13g2_decap_4 FILLER_6_2518 ();
 sg13g2_fill_2 FILLER_6_2522 ();
 sg13g2_decap_8 FILLER_6_2586 ();
 sg13g2_decap_8 FILLER_6_2593 ();
 sg13g2_decap_8 FILLER_6_2600 ();
 sg13g2_decap_8 FILLER_6_2607 ();
 sg13g2_decap_8 FILLER_6_2614 ();
 sg13g2_decap_8 FILLER_6_2621 ();
 sg13g2_decap_8 FILLER_6_2628 ();
 sg13g2_decap_8 FILLER_6_2635 ();
 sg13g2_decap_8 FILLER_6_2642 ();
 sg13g2_decap_8 FILLER_6_2649 ();
 sg13g2_decap_8 FILLER_6_2656 ();
 sg13g2_decap_8 FILLER_6_2663 ();
 sg13g2_fill_2 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_45 ();
 sg13g2_decap_4 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_60 ();
 sg13g2_fill_2 FILLER_7_71 ();
 sg13g2_fill_2 FILLER_7_78 ();
 sg13g2_decap_4 FILLER_7_85 ();
 sg13g2_decap_8 FILLER_7_93 ();
 sg13g2_fill_2 FILLER_7_100 ();
 sg13g2_fill_1 FILLER_7_102 ();
 sg13g2_fill_1 FILLER_7_205 ();
 sg13g2_fill_2 FILLER_7_225 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_fill_2 FILLER_7_265 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_fill_1 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_283 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_4 FILLER_7_297 ();
 sg13g2_decap_4 FILLER_7_305 ();
 sg13g2_decap_4 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_decap_4 FILLER_7_326 ();
 sg13g2_fill_2 FILLER_7_330 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_fill_2 FILLER_7_393 ();
 sg13g2_decap_8 FILLER_7_447 ();
 sg13g2_decap_4 FILLER_7_454 ();
 sg13g2_fill_1 FILLER_7_458 ();
 sg13g2_fill_1 FILLER_7_515 ();
 sg13g2_decap_8 FILLER_7_520 ();
 sg13g2_fill_1 FILLER_7_527 ();
 sg13g2_fill_2 FILLER_7_532 ();
 sg13g2_fill_1 FILLER_7_538 ();
 sg13g2_decap_8 FILLER_7_544 ();
 sg13g2_decap_8 FILLER_7_551 ();
 sg13g2_decap_8 FILLER_7_558 ();
 sg13g2_decap_8 FILLER_7_565 ();
 sg13g2_fill_2 FILLER_7_572 ();
 sg13g2_fill_1 FILLER_7_574 ();
 sg13g2_fill_2 FILLER_7_615 ();
 sg13g2_fill_1 FILLER_7_632 ();
 sg13g2_decap_4 FILLER_7_639 ();
 sg13g2_decap_4 FILLER_7_658 ();
 sg13g2_fill_1 FILLER_7_662 ();
 sg13g2_fill_2 FILLER_7_693 ();
 sg13g2_fill_1 FILLER_7_695 ();
 sg13g2_fill_2 FILLER_7_704 ();
 sg13g2_fill_2 FILLER_7_715 ();
 sg13g2_fill_2 FILLER_7_722 ();
 sg13g2_fill_1 FILLER_7_724 ();
 sg13g2_fill_2 FILLER_7_730 ();
 sg13g2_fill_1 FILLER_7_732 ();
 sg13g2_fill_2 FILLER_7_738 ();
 sg13g2_decap_8 FILLER_7_778 ();
 sg13g2_fill_2 FILLER_7_785 ();
 sg13g2_fill_2 FILLER_7_879 ();
 sg13g2_fill_2 FILLER_7_924 ();
 sg13g2_decap_8 FILLER_7_987 ();
 sg13g2_decap_4 FILLER_7_994 ();
 sg13g2_fill_2 FILLER_7_998 ();
 sg13g2_decap_4 FILLER_7_1004 ();
 sg13g2_fill_2 FILLER_7_1008 ();
 sg13g2_fill_2 FILLER_7_1014 ();
 sg13g2_fill_1 FILLER_7_1016 ();
 sg13g2_fill_2 FILLER_7_1022 ();
 sg13g2_fill_1 FILLER_7_1024 ();
 sg13g2_fill_2 FILLER_7_1029 ();
 sg13g2_fill_1 FILLER_7_1057 ();
 sg13g2_fill_1 FILLER_7_1063 ();
 sg13g2_fill_1 FILLER_7_1095 ();
 sg13g2_fill_1 FILLER_7_1122 ();
 sg13g2_fill_1 FILLER_7_1131 ();
 sg13g2_fill_1 FILLER_7_1158 ();
 sg13g2_fill_2 FILLER_7_1169 ();
 sg13g2_fill_2 FILLER_7_1192 ();
 sg13g2_fill_2 FILLER_7_1198 ();
 sg13g2_decap_8 FILLER_7_1238 ();
 sg13g2_decap_8 FILLER_7_1245 ();
 sg13g2_decap_4 FILLER_7_1321 ();
 sg13g2_fill_1 FILLER_7_1325 ();
 sg13g2_fill_2 FILLER_7_1336 ();
 sg13g2_decap_8 FILLER_7_1346 ();
 sg13g2_decap_8 FILLER_7_1353 ();
 sg13g2_decap_8 FILLER_7_1360 ();
 sg13g2_fill_1 FILLER_7_1367 ();
 sg13g2_decap_4 FILLER_7_1398 ();
 sg13g2_decap_8 FILLER_7_1428 ();
 sg13g2_decap_8 FILLER_7_1435 ();
 sg13g2_decap_4 FILLER_7_1442 ();
 sg13g2_decap_8 FILLER_7_1454 ();
 sg13g2_fill_1 FILLER_7_1461 ();
 sg13g2_fill_1 FILLER_7_1488 ();
 sg13g2_decap_8 FILLER_7_1493 ();
 sg13g2_fill_2 FILLER_7_1500 ();
 sg13g2_decap_4 FILLER_7_1512 ();
 sg13g2_fill_1 FILLER_7_1516 ();
 sg13g2_decap_4 FILLER_7_1589 ();
 sg13g2_fill_1 FILLER_7_1593 ();
 sg13g2_decap_4 FILLER_7_1601 ();
 sg13g2_fill_2 FILLER_7_1605 ();
 sg13g2_fill_1 FILLER_7_1611 ();
 sg13g2_fill_1 FILLER_7_1615 ();
 sg13g2_fill_1 FILLER_7_1656 ();
 sg13g2_decap_4 FILLER_7_1661 ();
 sg13g2_fill_1 FILLER_7_1755 ();
 sg13g2_fill_2 FILLER_7_1762 ();
 sg13g2_fill_2 FILLER_7_1769 ();
 sg13g2_fill_2 FILLER_7_1776 ();
 sg13g2_fill_1 FILLER_7_1778 ();
 sg13g2_fill_1 FILLER_7_1804 ();
 sg13g2_fill_1 FILLER_7_1809 ();
 sg13g2_fill_2 FILLER_7_1824 ();
 sg13g2_fill_1 FILLER_7_1826 ();
 sg13g2_fill_1 FILLER_7_1832 ();
 sg13g2_fill_1 FILLER_7_1839 ();
 sg13g2_fill_1 FILLER_7_1860 ();
 sg13g2_fill_1 FILLER_7_1865 ();
 sg13g2_fill_1 FILLER_7_1872 ();
 sg13g2_fill_1 FILLER_7_1879 ();
 sg13g2_fill_1 FILLER_7_1884 ();
 sg13g2_fill_2 FILLER_7_1916 ();
 sg13g2_fill_1 FILLER_7_1918 ();
 sg13g2_decap_8 FILLER_7_1923 ();
 sg13g2_decap_4 FILLER_7_1930 ();
 sg13g2_fill_2 FILLER_7_1943 ();
 sg13g2_fill_1 FILLER_7_1945 ();
 sg13g2_fill_1 FILLER_7_2002 ();
 sg13g2_decap_4 FILLER_7_2055 ();
 sg13g2_fill_2 FILLER_7_2059 ();
 sg13g2_decap_4 FILLER_7_2113 ();
 sg13g2_fill_2 FILLER_7_2160 ();
 sg13g2_decap_8 FILLER_7_2238 ();
 sg13g2_decap_8 FILLER_7_2245 ();
 sg13g2_fill_2 FILLER_7_2252 ();
 sg13g2_fill_1 FILLER_7_2254 ();
 sg13g2_fill_2 FILLER_7_2305 ();
 sg13g2_fill_1 FILLER_7_2317 ();
 sg13g2_fill_2 FILLER_7_2364 ();
 sg13g2_fill_2 FILLER_7_2370 ();
 sg13g2_fill_1 FILLER_7_2372 ();
 sg13g2_fill_1 FILLER_7_2399 ();
 sg13g2_fill_2 FILLER_7_2426 ();
 sg13g2_fill_1 FILLER_7_2454 ();
 sg13g2_fill_2 FILLER_7_2481 ();
 sg13g2_decap_8 FILLER_7_2509 ();
 sg13g2_decap_8 FILLER_7_2516 ();
 sg13g2_decap_8 FILLER_7_2523 ();
 sg13g2_fill_1 FILLER_7_2530 ();
 sg13g2_decap_4 FILLER_7_2556 ();
 sg13g2_fill_1 FILLER_7_2560 ();
 sg13g2_decap_8 FILLER_7_2565 ();
 sg13g2_decap_8 FILLER_7_2572 ();
 sg13g2_decap_8 FILLER_7_2579 ();
 sg13g2_decap_8 FILLER_7_2586 ();
 sg13g2_decap_8 FILLER_7_2593 ();
 sg13g2_decap_8 FILLER_7_2600 ();
 sg13g2_decap_8 FILLER_7_2607 ();
 sg13g2_decap_8 FILLER_7_2614 ();
 sg13g2_decap_8 FILLER_7_2621 ();
 sg13g2_decap_8 FILLER_7_2628 ();
 sg13g2_decap_8 FILLER_7_2635 ();
 sg13g2_decap_8 FILLER_7_2642 ();
 sg13g2_decap_8 FILLER_7_2649 ();
 sg13g2_decap_8 FILLER_7_2656 ();
 sg13g2_decap_8 FILLER_7_2663 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_34 ();
 sg13g2_fill_1 FILLER_8_53 ();
 sg13g2_decap_4 FILLER_8_78 ();
 sg13g2_fill_1 FILLER_8_82 ();
 sg13g2_fill_1 FILLER_8_91 ();
 sg13g2_fill_1 FILLER_8_127 ();
 sg13g2_fill_1 FILLER_8_133 ();
 sg13g2_fill_2 FILLER_8_139 ();
 sg13g2_fill_2 FILLER_8_145 ();
 sg13g2_fill_2 FILLER_8_151 ();
 sg13g2_decap_4 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_222 ();
 sg13g2_fill_2 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_272 ();
 sg13g2_decap_8 FILLER_8_277 ();
 sg13g2_decap_8 FILLER_8_284 ();
 sg13g2_fill_2 FILLER_8_291 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_1 FILLER_8_330 ();
 sg13g2_fill_1 FILLER_8_367 ();
 sg13g2_decap_4 FILLER_8_409 ();
 sg13g2_fill_1 FILLER_8_413 ();
 sg13g2_decap_4 FILLER_8_422 ();
 sg13g2_fill_2 FILLER_8_426 ();
 sg13g2_fill_1 FILLER_8_436 ();
 sg13g2_fill_2 FILLER_8_447 ();
 sg13g2_decap_8 FILLER_8_454 ();
 sg13g2_fill_2 FILLER_8_461 ();
 sg13g2_fill_1 FILLER_8_463 ();
 sg13g2_fill_2 FILLER_8_490 ();
 sg13g2_fill_1 FILLER_8_492 ();
 sg13g2_decap_8 FILLER_8_499 ();
 sg13g2_decap_4 FILLER_8_511 ();
 sg13g2_fill_2 FILLER_8_545 ();
 sg13g2_decap_8 FILLER_8_551 ();
 sg13g2_decap_8 FILLER_8_558 ();
 sg13g2_fill_2 FILLER_8_565 ();
 sg13g2_fill_1 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_573 ();
 sg13g2_fill_1 FILLER_8_580 ();
 sg13g2_fill_2 FILLER_8_617 ();
 sg13g2_fill_1 FILLER_8_629 ();
 sg13g2_fill_1 FILLER_8_666 ();
 sg13g2_fill_2 FILLER_8_672 ();
 sg13g2_fill_1 FILLER_8_674 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_fill_1 FILLER_8_747 ();
 sg13g2_fill_2 FILLER_8_766 ();
 sg13g2_decap_8 FILLER_8_772 ();
 sg13g2_decap_4 FILLER_8_779 ();
 sg13g2_fill_1 FILLER_8_783 ();
 sg13g2_fill_2 FILLER_8_788 ();
 sg13g2_fill_1 FILLER_8_790 ();
 sg13g2_fill_1 FILLER_8_795 ();
 sg13g2_fill_1 FILLER_8_822 ();
 sg13g2_fill_2 FILLER_8_849 ();
 sg13g2_decap_8 FILLER_8_872 ();
 sg13g2_fill_2 FILLER_8_966 ();
 sg13g2_fill_1 FILLER_8_998 ();
 sg13g2_decap_4 FILLER_8_1034 ();
 sg13g2_fill_1 FILLER_8_1042 ();
 sg13g2_decap_8 FILLER_8_1081 ();
 sg13g2_fill_2 FILLER_8_1088 ();
 sg13g2_fill_1 FILLER_8_1090 ();
 sg13g2_fill_2 FILLER_8_1100 ();
 sg13g2_fill_1 FILLER_8_1102 ();
 sg13g2_decap_8 FILLER_8_1145 ();
 sg13g2_fill_1 FILLER_8_1182 ();
 sg13g2_fill_2 FILLER_8_1209 ();
 sg13g2_decap_8 FILLER_8_1237 ();
 sg13g2_fill_2 FILLER_8_1244 ();
 sg13g2_decap_4 FILLER_8_1272 ();
 sg13g2_fill_2 FILLER_8_1276 ();
 sg13g2_fill_1 FILLER_8_1283 ();
 sg13g2_decap_8 FILLER_8_1325 ();
 sg13g2_fill_2 FILLER_8_1332 ();
 sg13g2_fill_1 FILLER_8_1334 ();
 sg13g2_decap_4 FILLER_8_1375 ();
 sg13g2_fill_1 FILLER_8_1379 ();
 sg13g2_fill_2 FILLER_8_1384 ();
 sg13g2_fill_2 FILLER_8_1413 ();
 sg13g2_fill_1 FILLER_8_1441 ();
 sg13g2_decap_8 FILLER_8_1446 ();
 sg13g2_decap_4 FILLER_8_1453 ();
 sg13g2_fill_2 FILLER_8_1457 ();
 sg13g2_fill_1 FILLER_8_1473 ();
 sg13g2_fill_1 FILLER_8_1478 ();
 sg13g2_decap_4 FILLER_8_1505 ();
 sg13g2_decap_4 FILLER_8_1513 ();
 sg13g2_fill_2 FILLER_8_1517 ();
 sg13g2_fill_2 FILLER_8_1546 ();
 sg13g2_fill_1 FILLER_8_1548 ();
 sg13g2_fill_2 FILLER_8_1552 ();
 sg13g2_fill_1 FILLER_8_1584 ();
 sg13g2_fill_1 FILLER_8_1611 ();
 sg13g2_fill_2 FILLER_8_1622 ();
 sg13g2_fill_1 FILLER_8_1624 ();
 sg13g2_fill_2 FILLER_8_1629 ();
 sg13g2_fill_2 FILLER_8_1656 ();
 sg13g2_fill_1 FILLER_8_1658 ();
 sg13g2_fill_2 FILLER_8_1695 ();
 sg13g2_fill_1 FILLER_8_1697 ();
 sg13g2_decap_8 FILLER_8_1702 ();
 sg13g2_decap_8 FILLER_8_1709 ();
 sg13g2_fill_1 FILLER_8_1716 ();
 sg13g2_fill_1 FILLER_8_1788 ();
 sg13g2_fill_1 FILLER_8_1793 ();
 sg13g2_fill_2 FILLER_8_1799 ();
 sg13g2_fill_1 FILLER_8_1822 ();
 sg13g2_fill_2 FILLER_8_1880 ();
 sg13g2_fill_1 FILLER_8_1882 ();
 sg13g2_fill_2 FILLER_8_1893 ();
 sg13g2_fill_1 FILLER_8_1895 ();
 sg13g2_fill_1 FILLER_8_1922 ();
 sg13g2_fill_1 FILLER_8_1928 ();
 sg13g2_fill_1 FILLER_8_1934 ();
 sg13g2_fill_2 FILLER_8_1945 ();
 sg13g2_fill_1 FILLER_8_1951 ();
 sg13g2_fill_1 FILLER_8_1962 ();
 sg13g2_decap_4 FILLER_8_1999 ();
 sg13g2_fill_1 FILLER_8_2003 ();
 sg13g2_decap_8 FILLER_8_2018 ();
 sg13g2_decap_8 FILLER_8_2025 ();
 sg13g2_fill_2 FILLER_8_2068 ();
 sg13g2_fill_1 FILLER_8_2070 ();
 sg13g2_decap_8 FILLER_8_2075 ();
 sg13g2_fill_1 FILLER_8_2082 ();
 sg13g2_decap_8 FILLER_8_2122 ();
 sg13g2_fill_2 FILLER_8_2129 ();
 sg13g2_decap_4 FILLER_8_2139 ();
 sg13g2_decap_4 FILLER_8_2167 ();
 sg13g2_fill_1 FILLER_8_2196 ();
 sg13g2_fill_1 FILLER_8_2201 ();
 sg13g2_fill_1 FILLER_8_2212 ();
 sg13g2_fill_1 FILLER_8_2217 ();
 sg13g2_fill_2 FILLER_8_2249 ();
 sg13g2_fill_1 FILLER_8_2251 ();
 sg13g2_fill_2 FILLER_8_2307 ();
 sg13g2_fill_1 FILLER_8_2309 ();
 sg13g2_fill_2 FILLER_8_2362 ();
 sg13g2_fill_1 FILLER_8_2400 ();
 sg13g2_decap_4 FILLER_8_2405 ();
 sg13g2_decap_8 FILLER_8_2436 ();
 sg13g2_decap_8 FILLER_8_2443 ();
 sg13g2_decap_8 FILLER_8_2450 ();
 sg13g2_decap_4 FILLER_8_2457 ();
 sg13g2_fill_1 FILLER_8_2461 ();
 sg13g2_fill_1 FILLER_8_2466 ();
 sg13g2_fill_2 FILLER_8_2488 ();
 sg13g2_fill_1 FILLER_8_2490 ();
 sg13g2_fill_2 FILLER_8_2521 ();
 sg13g2_decap_8 FILLER_8_2580 ();
 sg13g2_decap_8 FILLER_8_2587 ();
 sg13g2_decap_8 FILLER_8_2594 ();
 sg13g2_decap_8 FILLER_8_2601 ();
 sg13g2_decap_8 FILLER_8_2608 ();
 sg13g2_decap_8 FILLER_8_2615 ();
 sg13g2_decap_8 FILLER_8_2622 ();
 sg13g2_decap_8 FILLER_8_2629 ();
 sg13g2_decap_8 FILLER_8_2636 ();
 sg13g2_decap_8 FILLER_8_2643 ();
 sg13g2_decap_8 FILLER_8_2650 ();
 sg13g2_decap_8 FILLER_8_2657 ();
 sg13g2_decap_4 FILLER_8_2664 ();
 sg13g2_fill_2 FILLER_8_2668 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_11 ();
 sg13g2_fill_1 FILLER_9_13 ();
 sg13g2_decap_8 FILLER_9_92 ();
 sg13g2_decap_4 FILLER_9_99 ();
 sg13g2_fill_2 FILLER_9_103 ();
 sg13g2_fill_2 FILLER_9_115 ();
 sg13g2_fill_1 FILLER_9_117 ();
 sg13g2_fill_2 FILLER_9_166 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_193 ();
 sg13g2_fill_2 FILLER_9_239 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_4 FILLER_9_262 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_2 FILLER_9_307 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_fill_2 FILLER_9_336 ();
 sg13g2_fill_1 FILLER_9_338 ();
 sg13g2_fill_2 FILLER_9_343 ();
 sg13g2_decap_4 FILLER_9_375 ();
 sg13g2_fill_2 FILLER_9_379 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_fill_1 FILLER_9_392 ();
 sg13g2_fill_2 FILLER_9_399 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_decap_4 FILLER_9_411 ();
 sg13g2_fill_2 FILLER_9_415 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_fill_2 FILLER_9_434 ();
 sg13g2_fill_1 FILLER_9_436 ();
 sg13g2_fill_1 FILLER_9_459 ();
 sg13g2_decap_4 FILLER_9_511 ();
 sg13g2_fill_2 FILLER_9_525 ();
 sg13g2_fill_1 FILLER_9_527 ();
 sg13g2_decap_8 FILLER_9_568 ();
 sg13g2_decap_8 FILLER_9_670 ();
 sg13g2_decap_8 FILLER_9_677 ();
 sg13g2_decap_4 FILLER_9_684 ();
 sg13g2_fill_2 FILLER_9_688 ();
 sg13g2_fill_1 FILLER_9_704 ();
 sg13g2_fill_1 FILLER_9_722 ();
 sg13g2_fill_2 FILLER_9_733 ();
 sg13g2_decap_4 FILLER_9_779 ();
 sg13g2_fill_1 FILLER_9_803 ();
 sg13g2_fill_2 FILLER_9_814 ();
 sg13g2_fill_2 FILLER_9_837 ();
 sg13g2_fill_2 FILLER_9_843 ();
 sg13g2_fill_1 FILLER_9_855 ();
 sg13g2_fill_2 FILLER_9_869 ();
 sg13g2_fill_2 FILLER_9_906 ();
 sg13g2_fill_2 FILLER_9_916 ();
 sg13g2_fill_1 FILLER_9_918 ();
 sg13g2_decap_4 FILLER_9_954 ();
 sg13g2_fill_1 FILLER_9_958 ();
 sg13g2_fill_2 FILLER_9_976 ();
 sg13g2_decap_4 FILLER_9_987 ();
 sg13g2_decap_4 FILLER_9_1021 ();
 sg13g2_fill_2 FILLER_9_1025 ();
 sg13g2_fill_2 FILLER_9_1032 ();
 sg13g2_decap_4 FILLER_9_1039 ();
 sg13g2_fill_2 FILLER_9_1043 ();
 sg13g2_decap_4 FILLER_9_1050 ();
 sg13g2_fill_1 FILLER_9_1054 ();
 sg13g2_decap_4 FILLER_9_1059 ();
 sg13g2_fill_1 FILLER_9_1063 ();
 sg13g2_decap_4 FILLER_9_1068 ();
 sg13g2_fill_2 FILLER_9_1080 ();
 sg13g2_decap_4 FILLER_9_1087 ();
 sg13g2_decap_4 FILLER_9_1095 ();
 sg13g2_fill_2 FILLER_9_1134 ();
 sg13g2_fill_1 FILLER_9_1198 ();
 sg13g2_fill_2 FILLER_9_1232 ();
 sg13g2_decap_4 FILLER_9_1244 ();
 sg13g2_fill_2 FILLER_9_1248 ();
 sg13g2_fill_2 FILLER_9_1271 ();
 sg13g2_fill_1 FILLER_9_1273 ();
 sg13g2_decap_4 FILLER_9_1298 ();
 sg13g2_fill_1 FILLER_9_1302 ();
 sg13g2_decap_8 FILLER_9_1307 ();
 sg13g2_decap_4 FILLER_9_1314 ();
 sg13g2_fill_1 FILLER_9_1318 ();
 sg13g2_decap_8 FILLER_9_1365 ();
 sg13g2_decap_8 FILLER_9_1372 ();
 sg13g2_decap_8 FILLER_9_1379 ();
 sg13g2_decap_8 FILLER_9_1386 ();
 sg13g2_fill_2 FILLER_9_1393 ();
 sg13g2_fill_2 FILLER_9_1409 ();
 sg13g2_fill_1 FILLER_9_1411 ();
 sg13g2_fill_1 FILLER_9_1435 ();
 sg13g2_decap_8 FILLER_9_1472 ();
 sg13g2_fill_2 FILLER_9_1479 ();
 sg13g2_fill_1 FILLER_9_1481 ();
 sg13g2_fill_2 FILLER_9_1490 ();
 sg13g2_fill_1 FILLER_9_1495 ();
 sg13g2_fill_2 FILLER_9_1501 ();
 sg13g2_fill_2 FILLER_9_1532 ();
 sg13g2_fill_2 FILLER_9_1544 ();
 sg13g2_fill_1 FILLER_9_1567 ();
 sg13g2_fill_2 FILLER_9_1572 ();
 sg13g2_fill_1 FILLER_9_1586 ();
 sg13g2_fill_1 FILLER_9_1617 ();
 sg13g2_fill_2 FILLER_9_1644 ();
 sg13g2_fill_2 FILLER_9_1676 ();
 sg13g2_decap_8 FILLER_9_1686 ();
 sg13g2_decap_8 FILLER_9_1693 ();
 sg13g2_decap_8 FILLER_9_1700 ();
 sg13g2_decap_8 FILLER_9_1707 ();
 sg13g2_decap_8 FILLER_9_1714 ();
 sg13g2_decap_8 FILLER_9_1721 ();
 sg13g2_fill_1 FILLER_9_1728 ();
 sg13g2_decap_4 FILLER_9_1737 ();
 sg13g2_fill_1 FILLER_9_1780 ();
 sg13g2_fill_1 FILLER_9_1786 ();
 sg13g2_decap_8 FILLER_9_1813 ();
 sg13g2_fill_1 FILLER_9_1820 ();
 sg13g2_fill_2 FILLER_9_1830 ();
 sg13g2_fill_1 FILLER_9_1832 ();
 sg13g2_fill_2 FILLER_9_1837 ();
 sg13g2_fill_1 FILLER_9_1850 ();
 sg13g2_fill_1 FILLER_9_1877 ();
 sg13g2_fill_2 FILLER_9_1899 ();
 sg13g2_fill_1 FILLER_9_1901 ();
 sg13g2_decap_8 FILLER_9_1912 ();
 sg13g2_decap_4 FILLER_9_1919 ();
 sg13g2_fill_1 FILLER_9_1937 ();
 sg13g2_fill_1 FILLER_9_1948 ();
 sg13g2_fill_1 FILLER_9_1953 ();
 sg13g2_fill_1 FILLER_9_1958 ();
 sg13g2_fill_1 FILLER_9_1963 ();
 sg13g2_decap_4 FILLER_9_1989 ();
 sg13g2_fill_2 FILLER_9_1993 ();
 sg13g2_fill_1 FILLER_9_2021 ();
 sg13g2_decap_8 FILLER_9_2096 ();
 sg13g2_decap_4 FILLER_9_2103 ();
 sg13g2_fill_2 FILLER_9_2147 ();
 sg13g2_fill_1 FILLER_9_2149 ();
 sg13g2_fill_1 FILLER_9_2202 ();
 sg13g2_decap_8 FILLER_9_2220 ();
 sg13g2_decap_4 FILLER_9_2227 ();
 sg13g2_fill_2 FILLER_9_2235 ();
 sg13g2_fill_1 FILLER_9_2237 ();
 sg13g2_fill_1 FILLER_9_2273 ();
 sg13g2_fill_1 FILLER_9_2287 ();
 sg13g2_fill_1 FILLER_9_2292 ();
 sg13g2_fill_1 FILLER_9_2297 ();
 sg13g2_fill_1 FILLER_9_2319 ();
 sg13g2_decap_4 FILLER_9_2324 ();
 sg13g2_decap_4 FILLER_9_2338 ();
 sg13g2_decap_4 FILLER_9_2359 ();
 sg13g2_fill_1 FILLER_9_2363 ();
 sg13g2_decap_8 FILLER_9_2394 ();
 sg13g2_decap_8 FILLER_9_2401 ();
 sg13g2_decap_4 FILLER_9_2408 ();
 sg13g2_fill_1 FILLER_9_2412 ();
 sg13g2_fill_2 FILLER_9_2416 ();
 sg13g2_fill_1 FILLER_9_2418 ();
 sg13g2_fill_2 FILLER_9_2470 ();
 sg13g2_fill_1 FILLER_9_2472 ();
 sg13g2_decap_8 FILLER_9_2483 ();
 sg13g2_fill_1 FILLER_9_2490 ();
 sg13g2_decap_4 FILLER_9_2560 ();
 sg13g2_fill_2 FILLER_9_2564 ();
 sg13g2_decap_8 FILLER_9_2576 ();
 sg13g2_decap_8 FILLER_9_2583 ();
 sg13g2_decap_8 FILLER_9_2590 ();
 sg13g2_decap_8 FILLER_9_2597 ();
 sg13g2_decap_8 FILLER_9_2604 ();
 sg13g2_decap_8 FILLER_9_2611 ();
 sg13g2_decap_8 FILLER_9_2618 ();
 sg13g2_decap_8 FILLER_9_2625 ();
 sg13g2_decap_8 FILLER_9_2632 ();
 sg13g2_decap_8 FILLER_9_2639 ();
 sg13g2_decap_8 FILLER_9_2646 ();
 sg13g2_decap_8 FILLER_9_2653 ();
 sg13g2_decap_8 FILLER_9_2660 ();
 sg13g2_fill_2 FILLER_9_2667 ();
 sg13g2_fill_1 FILLER_9_2669 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_4 FILLER_10_7 ();
 sg13g2_fill_1 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_16 ();
 sg13g2_decap_4 FILLER_10_23 ();
 sg13g2_fill_1 FILLER_10_27 ();
 sg13g2_decap_4 FILLER_10_33 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_47 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_85 ();
 sg13g2_decap_8 FILLER_10_92 ();
 sg13g2_decap_4 FILLER_10_99 ();
 sg13g2_fill_2 FILLER_10_107 ();
 sg13g2_fill_1 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_4 FILLER_10_125 ();
 sg13g2_fill_2 FILLER_10_129 ();
 sg13g2_decap_8 FILLER_10_136 ();
 sg13g2_fill_2 FILLER_10_153 ();
 sg13g2_fill_1 FILLER_10_174 ();
 sg13g2_fill_2 FILLER_10_180 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_219 ();
 sg13g2_decap_4 FILLER_10_226 ();
 sg13g2_fill_2 FILLER_10_230 ();
 sg13g2_decap_8 FILLER_10_245 ();
 sg13g2_decap_8 FILLER_10_252 ();
 sg13g2_decap_4 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_decap_4 FILLER_10_300 ();
 sg13g2_fill_2 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_316 ();
 sg13g2_fill_1 FILLER_10_362 ();
 sg13g2_fill_2 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_379 ();
 sg13g2_decap_8 FILLER_10_386 ();
 sg13g2_decap_4 FILLER_10_428 ();
 sg13g2_fill_2 FILLER_10_467 ();
 sg13g2_decap_8 FILLER_10_478 ();
 sg13g2_fill_2 FILLER_10_485 ();
 sg13g2_fill_1 FILLER_10_487 ();
 sg13g2_fill_1 FILLER_10_493 ();
 sg13g2_fill_2 FILLER_10_498 ();
 sg13g2_decap_8 FILLER_10_504 ();
 sg13g2_decap_4 FILLER_10_511 ();
 sg13g2_fill_1 FILLER_10_515 ();
 sg13g2_decap_4 FILLER_10_534 ();
 sg13g2_fill_1 FILLER_10_552 ();
 sg13g2_decap_4 FILLER_10_579 ();
 sg13g2_fill_1 FILLER_10_583 ();
 sg13g2_decap_4 FILLER_10_620 ();
 sg13g2_fill_1 FILLER_10_624 ();
 sg13g2_decap_8 FILLER_10_629 ();
 sg13g2_fill_2 FILLER_10_636 ();
 sg13g2_decap_8 FILLER_10_649 ();
 sg13g2_decap_8 FILLER_10_656 ();
 sg13g2_decap_8 FILLER_10_663 ();
 sg13g2_decap_8 FILLER_10_670 ();
 sg13g2_decap_8 FILLER_10_677 ();
 sg13g2_fill_1 FILLER_10_688 ();
 sg13g2_fill_1 FILLER_10_710 ();
 sg13g2_fill_2 FILLER_10_745 ();
 sg13g2_decap_8 FILLER_10_773 ();
 sg13g2_decap_8 FILLER_10_780 ();
 sg13g2_decap_8 FILLER_10_787 ();
 sg13g2_fill_1 FILLER_10_794 ();
 sg13g2_fill_2 FILLER_10_821 ();
 sg13g2_fill_1 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_834 ();
 sg13g2_decap_8 FILLER_10_841 ();
 sg13g2_decap_4 FILLER_10_848 ();
 sg13g2_decap_8 FILLER_10_911 ();
 sg13g2_decap_4 FILLER_10_918 ();
 sg13g2_fill_1 FILLER_10_922 ();
 sg13g2_decap_4 FILLER_10_937 ();
 sg13g2_fill_1 FILLER_10_941 ();
 sg13g2_fill_2 FILLER_10_946 ();
 sg13g2_decap_8 FILLER_10_973 ();
 sg13g2_fill_2 FILLER_10_980 ();
 sg13g2_fill_2 FILLER_10_1007 ();
 sg13g2_fill_2 FILLER_10_1014 ();
 sg13g2_decap_8 FILLER_10_1024 ();
 sg13g2_decap_8 FILLER_10_1031 ();
 sg13g2_decap_8 FILLER_10_1038 ();
 sg13g2_decap_8 FILLER_10_1045 ();
 sg13g2_decap_8 FILLER_10_1052 ();
 sg13g2_decap_8 FILLER_10_1059 ();
 sg13g2_decap_8 FILLER_10_1066 ();
 sg13g2_decap_8 FILLER_10_1073 ();
 sg13g2_fill_2 FILLER_10_1080 ();
 sg13g2_fill_2 FILLER_10_1125 ();
 sg13g2_fill_1 FILLER_10_1127 ();
 sg13g2_decap_8 FILLER_10_1158 ();
 sg13g2_decap_8 FILLER_10_1165 ();
 sg13g2_decap_4 FILLER_10_1172 ();
 sg13g2_fill_1 FILLER_10_1176 ();
 sg13g2_fill_2 FILLER_10_1181 ();
 sg13g2_decap_4 FILLER_10_1215 ();
 sg13g2_fill_1 FILLER_10_1219 ();
 sg13g2_fill_2 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1274 ();
 sg13g2_decap_4 FILLER_10_1315 ();
 sg13g2_decap_4 FILLER_10_1324 ();
 sg13g2_fill_1 FILLER_10_1328 ();
 sg13g2_fill_2 FILLER_10_1337 ();
 sg13g2_fill_2 FILLER_10_1343 ();
 sg13g2_fill_1 FILLER_10_1371 ();
 sg13g2_decap_8 FILLER_10_1398 ();
 sg13g2_decap_4 FILLER_10_1405 ();
 sg13g2_fill_1 FILLER_10_1409 ();
 sg13g2_decap_4 FILLER_10_1428 ();
 sg13g2_fill_2 FILLER_10_1432 ();
 sg13g2_fill_2 FILLER_10_1456 ();
 sg13g2_decap_4 FILLER_10_1461 ();
 sg13g2_fill_1 FILLER_10_1465 ();
 sg13g2_decap_8 FILLER_10_1479 ();
 sg13g2_fill_1 FILLER_10_1486 ();
 sg13g2_fill_2 FILLER_10_1492 ();
 sg13g2_fill_1 FILLER_10_1494 ();
 sg13g2_fill_2 FILLER_10_1505 ();
 sg13g2_fill_1 FILLER_10_1516 ();
 sg13g2_fill_2 FILLER_10_1550 ();
 sg13g2_fill_1 FILLER_10_1552 ();
 sg13g2_decap_4 FILLER_10_1566 ();
 sg13g2_fill_1 FILLER_10_1599 ();
 sg13g2_fill_1 FILLER_10_1655 ();
 sg13g2_decap_8 FILLER_10_1674 ();
 sg13g2_fill_2 FILLER_10_1681 ();
 sg13g2_fill_1 FILLER_10_1683 ();
 sg13g2_decap_8 FILLER_10_1688 ();
 sg13g2_decap_4 FILLER_10_1712 ();
 sg13g2_fill_2 FILLER_10_1716 ();
 sg13g2_fill_2 FILLER_10_1722 ();
 sg13g2_decap_4 FILLER_10_1729 ();
 sg13g2_fill_1 FILLER_10_1741 ();
 sg13g2_fill_2 FILLER_10_1754 ();
 sg13g2_fill_2 FILLER_10_1764 ();
 sg13g2_fill_2 FILLER_10_1778 ();
 sg13g2_decap_4 FILLER_10_1785 ();
 sg13g2_decap_8 FILLER_10_1793 ();
 sg13g2_fill_2 FILLER_10_1800 ();
 sg13g2_decap_4 FILLER_10_1826 ();
 sg13g2_fill_2 FILLER_10_1830 ();
 sg13g2_fill_2 FILLER_10_1837 ();
 sg13g2_fill_2 FILLER_10_1843 ();
 sg13g2_fill_1 FILLER_10_1851 ();
 sg13g2_fill_2 FILLER_10_1860 ();
 sg13g2_fill_2 FILLER_10_1882 ();
 sg13g2_decap_4 FILLER_10_1909 ();
 sg13g2_fill_2 FILLER_10_1913 ();
 sg13g2_fill_2 FILLER_10_1919 ();
 sg13g2_fill_1 FILLER_10_1921 ();
 sg13g2_fill_1 FILLER_10_1927 ();
 sg13g2_decap_4 FILLER_10_1954 ();
 sg13g2_fill_2 FILLER_10_1958 ();
 sg13g2_decap_8 FILLER_10_1970 ();
 sg13g2_decap_8 FILLER_10_1977 ();
 sg13g2_decap_8 FILLER_10_1984 ();
 sg13g2_decap_4 FILLER_10_1991 ();
 sg13g2_fill_2 FILLER_10_1995 ();
 sg13g2_fill_2 FILLER_10_2069 ();
 sg13g2_fill_1 FILLER_10_2071 ();
 sg13g2_decap_4 FILLER_10_2108 ();
 sg13g2_fill_2 FILLER_10_2112 ();
 sg13g2_decap_8 FILLER_10_2128 ();
 sg13g2_fill_2 FILLER_10_2135 ();
 sg13g2_fill_1 FILLER_10_2137 ();
 sg13g2_decap_4 FILLER_10_2154 ();
 sg13g2_fill_2 FILLER_10_2188 ();
 sg13g2_fill_1 FILLER_10_2190 ();
 sg13g2_decap_4 FILLER_10_2201 ();
 sg13g2_decap_8 FILLER_10_2278 ();
 sg13g2_fill_2 FILLER_10_2285 ();
 sg13g2_decap_8 FILLER_10_2297 ();
 sg13g2_decap_8 FILLER_10_2304 ();
 sg13g2_decap_8 FILLER_10_2311 ();
 sg13g2_decap_8 FILLER_10_2318 ();
 sg13g2_decap_8 FILLER_10_2325 ();
 sg13g2_decap_8 FILLER_10_2332 ();
 sg13g2_fill_2 FILLER_10_2339 ();
 sg13g2_decap_8 FILLER_10_2398 ();
 sg13g2_fill_2 FILLER_10_2410 ();
 sg13g2_decap_8 FILLER_10_2463 ();
 sg13g2_decap_8 FILLER_10_2470 ();
 sg13g2_decap_8 FILLER_10_2477 ();
 sg13g2_decap_8 FILLER_10_2484 ();
 sg13g2_decap_8 FILLER_10_2491 ();
 sg13g2_decap_4 FILLER_10_2498 ();
 sg13g2_fill_2 FILLER_10_2502 ();
 sg13g2_fill_2 FILLER_10_2508 ();
 sg13g2_fill_2 FILLER_10_2560 ();
 sg13g2_decap_8 FILLER_10_2588 ();
 sg13g2_decap_8 FILLER_10_2595 ();
 sg13g2_decap_8 FILLER_10_2602 ();
 sg13g2_decap_8 FILLER_10_2609 ();
 sg13g2_decap_8 FILLER_10_2616 ();
 sg13g2_decap_8 FILLER_10_2623 ();
 sg13g2_decap_8 FILLER_10_2630 ();
 sg13g2_decap_8 FILLER_10_2637 ();
 sg13g2_decap_8 FILLER_10_2644 ();
 sg13g2_decap_8 FILLER_10_2651 ();
 sg13g2_decap_8 FILLER_10_2658 ();
 sg13g2_decap_4 FILLER_10_2665 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_2 FILLER_11_29 ();
 sg13g2_decap_8 FILLER_11_45 ();
 sg13g2_decap_4 FILLER_11_56 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_1 FILLER_11_101 ();
 sg13g2_fill_1 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_142 ();
 sg13g2_fill_2 FILLER_11_148 ();
 sg13g2_fill_1 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_205 ();
 sg13g2_fill_1 FILLER_11_212 ();
 sg13g2_fill_1 FILLER_11_218 ();
 sg13g2_fill_1 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_240 ();
 sg13g2_decap_8 FILLER_11_247 ();
 sg13g2_decap_8 FILLER_11_254 ();
 sg13g2_decap_4 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_265 ();
 sg13g2_decap_8 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_296 ();
 sg13g2_fill_1 FILLER_11_321 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_fill_2 FILLER_11_364 ();
 sg13g2_fill_2 FILLER_11_370 ();
 sg13g2_fill_1 FILLER_11_372 ();
 sg13g2_fill_2 FILLER_11_387 ();
 sg13g2_fill_1 FILLER_11_389 ();
 sg13g2_decap_4 FILLER_11_434 ();
 sg13g2_fill_1 FILLER_11_477 ();
 sg13g2_decap_8 FILLER_11_487 ();
 sg13g2_fill_1 FILLER_11_494 ();
 sg13g2_decap_4 FILLER_11_499 ();
 sg13g2_fill_2 FILLER_11_503 ();
 sg13g2_fill_1 FILLER_11_528 ();
 sg13g2_fill_1 FILLER_11_547 ();
 sg13g2_fill_2 FILLER_11_556 ();
 sg13g2_fill_1 FILLER_11_558 ();
 sg13g2_decap_8 FILLER_11_563 ();
 sg13g2_fill_1 FILLER_11_570 ();
 sg13g2_decap_4 FILLER_11_585 ();
 sg13g2_fill_1 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_615 ();
 sg13g2_decap_8 FILLER_11_622 ();
 sg13g2_decap_4 FILLER_11_629 ();
 sg13g2_decap_8 FILLER_11_652 ();
 sg13g2_fill_2 FILLER_11_659 ();
 sg13g2_fill_2 FILLER_11_671 ();
 sg13g2_fill_2 FILLER_11_677 ();
 sg13g2_fill_1 FILLER_11_679 ();
 sg13g2_fill_2 FILLER_11_715 ();
 sg13g2_fill_1 FILLER_11_736 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_fill_2 FILLER_11_798 ();
 sg13g2_fill_1 FILLER_11_800 ();
 sg13g2_fill_1 FILLER_11_831 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_fill_1 FILLER_11_875 ();
 sg13g2_decap_4 FILLER_11_907 ();
 sg13g2_fill_2 FILLER_11_915 ();
 sg13g2_decap_8 FILLER_11_951 ();
 sg13g2_decap_8 FILLER_11_958 ();
 sg13g2_decap_8 FILLER_11_965 ();
 sg13g2_fill_2 FILLER_11_972 ();
 sg13g2_fill_1 FILLER_11_974 ();
 sg13g2_fill_2 FILLER_11_980 ();
 sg13g2_fill_1 FILLER_11_1034 ();
 sg13g2_fill_1 FILLER_11_1061 ();
 sg13g2_fill_1 FILLER_11_1066 ();
 sg13g2_decap_8 FILLER_11_1071 ();
 sg13g2_fill_2 FILLER_11_1078 ();
 sg13g2_decap_8 FILLER_11_1084 ();
 sg13g2_decap_4 FILLER_11_1091 ();
 sg13g2_fill_1 FILLER_11_1095 ();
 sg13g2_decap_8 FILLER_11_1160 ();
 sg13g2_decap_8 FILLER_11_1167 ();
 sg13g2_decap_4 FILLER_11_1174 ();
 sg13g2_fill_2 FILLER_11_1178 ();
 sg13g2_decap_8 FILLER_11_1190 ();
 sg13g2_fill_2 FILLER_11_1202 ();
 sg13g2_decap_4 FILLER_11_1208 ();
 sg13g2_fill_2 FILLER_11_1212 ();
 sg13g2_decap_8 FILLER_11_1229 ();
 sg13g2_decap_8 FILLER_11_1236 ();
 sg13g2_decap_4 FILLER_11_1243 ();
 sg13g2_fill_1 FILLER_11_1251 ();
 sg13g2_fill_2 FILLER_11_1288 ();
 sg13g2_fill_2 FILLER_11_1294 ();
 sg13g2_fill_2 FILLER_11_1301 ();
 sg13g2_fill_1 FILLER_11_1303 ();
 sg13g2_decap_8 FILLER_11_1310 ();
 sg13g2_decap_8 FILLER_11_1317 ();
 sg13g2_decap_8 FILLER_11_1324 ();
 sg13g2_decap_8 FILLER_11_1331 ();
 sg13g2_decap_4 FILLER_11_1338 ();
 sg13g2_fill_2 FILLER_11_1342 ();
 sg13g2_fill_2 FILLER_11_1392 ();
 sg13g2_fill_2 FILLER_11_1434 ();
 sg13g2_fill_1 FILLER_11_1436 ();
 sg13g2_decap_8 FILLER_11_1442 ();
 sg13g2_decap_4 FILLER_11_1449 ();
 sg13g2_fill_2 FILLER_11_1453 ();
 sg13g2_decap_4 FILLER_11_1464 ();
 sg13g2_fill_2 FILLER_11_1468 ();
 sg13g2_fill_2 FILLER_11_1487 ();
 sg13g2_fill_2 FILLER_11_1504 ();
 sg13g2_fill_2 FILLER_11_1513 ();
 sg13g2_fill_2 FILLER_11_1548 ();
 sg13g2_decap_8 FILLER_11_1558 ();
 sg13g2_fill_1 FILLER_11_1565 ();
 sg13g2_fill_2 FILLER_11_1616 ();
 sg13g2_fill_1 FILLER_11_1622 ();
 sg13g2_fill_1 FILLER_11_1636 ();
 sg13g2_fill_1 FILLER_11_1702 ();
 sg13g2_fill_1 FILLER_11_1706 ();
 sg13g2_fill_2 FILLER_11_1732 ();
 sg13g2_fill_1 FILLER_11_1734 ();
 sg13g2_fill_1 FILLER_11_1752 ();
 sg13g2_fill_2 FILLER_11_1766 ();
 sg13g2_fill_1 FILLER_11_1830 ();
 sg13g2_fill_2 FILLER_11_1836 ();
 sg13g2_fill_2 FILLER_11_1878 ();
 sg13g2_fill_1 FILLER_11_1880 ();
 sg13g2_decap_8 FILLER_11_1911 ();
 sg13g2_fill_2 FILLER_11_1918 ();
 sg13g2_fill_1 FILLER_11_1920 ();
 sg13g2_fill_2 FILLER_11_1926 ();
 sg13g2_fill_1 FILLER_11_1928 ();
 sg13g2_decap_8 FILLER_11_1955 ();
 sg13g2_decap_4 FILLER_11_1962 ();
 sg13g2_fill_2 FILLER_11_1966 ();
 sg13g2_fill_2 FILLER_11_1998 ();
 sg13g2_decap_4 FILLER_11_2026 ();
 sg13g2_decap_4 FILLER_11_2034 ();
 sg13g2_fill_2 FILLER_11_2038 ();
 sg13g2_decap_8 FILLER_11_2080 ();
 sg13g2_fill_2 FILLER_11_2087 ();
 sg13g2_decap_8 FILLER_11_2093 ();
 sg13g2_fill_2 FILLER_11_2100 ();
 sg13g2_decap_8 FILLER_11_2106 ();
 sg13g2_fill_2 FILLER_11_2113 ();
 sg13g2_fill_1 FILLER_11_2115 ();
 sg13g2_decap_8 FILLER_11_2141 ();
 sg13g2_decap_4 FILLER_11_2148 ();
 sg13g2_decap_4 FILLER_11_2160 ();
 sg13g2_fill_2 FILLER_11_2178 ();
 sg13g2_fill_1 FILLER_11_2180 ();
 sg13g2_fill_1 FILLER_11_2191 ();
 sg13g2_decap_8 FILLER_11_2222 ();
 sg13g2_decap_8 FILLER_11_2229 ();
 sg13g2_fill_1 FILLER_11_2236 ();
 sg13g2_decap_4 FILLER_11_2273 ();
 sg13g2_fill_1 FILLER_11_2281 ();
 sg13g2_fill_1 FILLER_11_2318 ();
 sg13g2_decap_8 FILLER_11_2332 ();
 sg13g2_decap_8 FILLER_11_2339 ();
 sg13g2_decap_8 FILLER_11_2346 ();
 sg13g2_decap_4 FILLER_11_2353 ();
 sg13g2_fill_2 FILLER_11_2357 ();
 sg13g2_decap_8 FILLER_11_2363 ();
 sg13g2_fill_2 FILLER_11_2370 ();
 sg13g2_fill_1 FILLER_11_2372 ();
 sg13g2_decap_4 FILLER_11_2377 ();
 sg13g2_fill_2 FILLER_11_2385 ();
 sg13g2_decap_4 FILLER_11_2452 ();
 sg13g2_fill_2 FILLER_11_2512 ();
 sg13g2_fill_1 FILLER_11_2518 ();
 sg13g2_fill_1 FILLER_11_2523 ();
 sg13g2_decap_8 FILLER_11_2550 ();
 sg13g2_decap_8 FILLER_11_2597 ();
 sg13g2_decap_8 FILLER_11_2604 ();
 sg13g2_decap_8 FILLER_11_2611 ();
 sg13g2_decap_8 FILLER_11_2618 ();
 sg13g2_decap_8 FILLER_11_2625 ();
 sg13g2_decap_8 FILLER_11_2632 ();
 sg13g2_decap_8 FILLER_11_2639 ();
 sg13g2_decap_8 FILLER_11_2646 ();
 sg13g2_decap_8 FILLER_11_2653 ();
 sg13g2_decap_8 FILLER_11_2660 ();
 sg13g2_fill_2 FILLER_11_2667 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_fill_2 FILLER_12_0 ();
 sg13g2_fill_1 FILLER_12_2 ();
 sg13g2_fill_2 FILLER_12_34 ();
 sg13g2_fill_2 FILLER_12_46 ();
 sg13g2_fill_1 FILLER_12_48 ();
 sg13g2_fill_1 FILLER_12_72 ();
 sg13g2_fill_1 FILLER_12_77 ();
 sg13g2_fill_1 FILLER_12_83 ();
 sg13g2_fill_2 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_191 ();
 sg13g2_decap_8 FILLER_12_248 ();
 sg13g2_decap_8 FILLER_12_255 ();
 sg13g2_decap_4 FILLER_12_262 ();
 sg13g2_fill_1 FILLER_12_266 ();
 sg13g2_decap_8 FILLER_12_272 ();
 sg13g2_decap_4 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_283 ();
 sg13g2_fill_1 FILLER_12_294 ();
 sg13g2_decap_4 FILLER_12_304 ();
 sg13g2_fill_1 FILLER_12_317 ();
 sg13g2_fill_2 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_fill_2 FILLER_12_387 ();
 sg13g2_fill_2 FILLER_12_411 ();
 sg13g2_fill_1 FILLER_12_434 ();
 sg13g2_fill_2 FILLER_12_449 ();
 sg13g2_fill_1 FILLER_12_460 ();
 sg13g2_fill_1 FILLER_12_489 ();
 sg13g2_fill_1 FILLER_12_530 ();
 sg13g2_fill_2 FILLER_12_541 ();
 sg13g2_decap_4 FILLER_12_548 ();
 sg13g2_fill_1 FILLER_12_552 ();
 sg13g2_decap_8 FILLER_12_691 ();
 sg13g2_fill_2 FILLER_12_698 ();
 sg13g2_decap_4 FILLER_12_709 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_fill_1 FILLER_12_732 ();
 sg13g2_fill_2 FILLER_12_801 ();
 sg13g2_fill_1 FILLER_12_889 ();
 sg13g2_fill_1 FILLER_12_916 ();
 sg13g2_fill_1 FILLER_12_943 ();
 sg13g2_fill_1 FILLER_12_970 ();
 sg13g2_fill_1 FILLER_12_1040 ();
 sg13g2_fill_2 FILLER_12_1091 ();
 sg13g2_fill_1 FILLER_12_1093 ();
 sg13g2_decap_4 FILLER_12_1098 ();
 sg13g2_fill_1 FILLER_12_1107 ();
 sg13g2_fill_1 FILLER_12_1112 ();
 sg13g2_fill_2 FILLER_12_1117 ();
 sg13g2_fill_2 FILLER_12_1144 ();
 sg13g2_fill_2 FILLER_12_1150 ();
 sg13g2_fill_1 FILLER_12_1152 ();
 sg13g2_fill_1 FILLER_12_1179 ();
 sg13g2_fill_2 FILLER_12_1219 ();
 sg13g2_decap_8 FILLER_12_1275 ();
 sg13g2_fill_1 FILLER_12_1282 ();
 sg13g2_fill_2 FILLER_12_1288 ();
 sg13g2_decap_4 FILLER_12_1306 ();
 sg13g2_fill_1 FILLER_12_1310 ();
 sg13g2_decap_8 FILLER_12_1321 ();
 sg13g2_decap_8 FILLER_12_1328 ();
 sg13g2_decap_8 FILLER_12_1335 ();
 sg13g2_fill_1 FILLER_12_1342 ();
 sg13g2_decap_8 FILLER_12_1353 ();
 sg13g2_fill_2 FILLER_12_1360 ();
 sg13g2_fill_1 FILLER_12_1362 ();
 sg13g2_fill_2 FILLER_12_1373 ();
 sg13g2_fill_2 FILLER_12_1379 ();
 sg13g2_decap_8 FILLER_12_1385 ();
 sg13g2_decap_8 FILLER_12_1392 ();
 sg13g2_fill_2 FILLER_12_1399 ();
 sg13g2_fill_1 FILLER_12_1401 ();
 sg13g2_fill_2 FILLER_12_1405 ();
 sg13g2_fill_2 FILLER_12_1417 ();
 sg13g2_fill_1 FILLER_12_1419 ();
 sg13g2_decap_8 FILLER_12_1426 ();
 sg13g2_fill_2 FILLER_12_1433 ();
 sg13g2_fill_1 FILLER_12_1435 ();
 sg13g2_decap_8 FILLER_12_1441 ();
 sg13g2_fill_2 FILLER_12_1454 ();
 sg13g2_fill_1 FILLER_12_1472 ();
 sg13g2_fill_1 FILLER_12_1486 ();
 sg13g2_fill_1 FILLER_12_1499 ();
 sg13g2_fill_2 FILLER_12_1505 ();
 sg13g2_fill_1 FILLER_12_1512 ();
 sg13g2_fill_2 FILLER_12_1525 ();
 sg13g2_fill_2 FILLER_12_1550 ();
 sg13g2_fill_1 FILLER_12_1562 ();
 sg13g2_fill_2 FILLER_12_1591 ();
 sg13g2_decap_4 FILLER_12_1617 ();
 sg13g2_fill_2 FILLER_12_1642 ();
 sg13g2_decap_8 FILLER_12_1661 ();
 sg13g2_decap_8 FILLER_12_1668 ();
 sg13g2_decap_8 FILLER_12_1675 ();
 sg13g2_decap_8 FILLER_12_1682 ();
 sg13g2_fill_2 FILLER_12_1693 ();
 sg13g2_decap_4 FILLER_12_1699 ();
 sg13g2_fill_1 FILLER_12_1703 ();
 sg13g2_fill_2 FILLER_12_1717 ();
 sg13g2_fill_1 FILLER_12_1724 ();
 sg13g2_fill_1 FILLER_12_1732 ();
 sg13g2_fill_2 FILLER_12_1746 ();
 sg13g2_fill_1 FILLER_12_1832 ();
 sg13g2_decap_8 FILLER_12_1840 ();
 sg13g2_fill_2 FILLER_12_1847 ();
 sg13g2_decap_4 FILLER_12_1858 ();
 sg13g2_fill_1 FILLER_12_1862 ();
 sg13g2_decap_8 FILLER_12_1867 ();
 sg13g2_fill_1 FILLER_12_1874 ();
 sg13g2_decap_8 FILLER_12_1905 ();
 sg13g2_decap_8 FILLER_12_1912 ();
 sg13g2_fill_2 FILLER_12_1919 ();
 sg13g2_fill_1 FILLER_12_1921 ();
 sg13g2_fill_2 FILLER_12_1949 ();
 sg13g2_fill_2 FILLER_12_1962 ();
 sg13g2_decap_8 FILLER_12_1982 ();
 sg13g2_decap_8 FILLER_12_1989 ();
 sg13g2_decap_8 FILLER_12_1996 ();
 sg13g2_fill_2 FILLER_12_2003 ();
 sg13g2_fill_2 FILLER_12_2009 ();
 sg13g2_decap_8 FILLER_12_2015 ();
 sg13g2_decap_8 FILLER_12_2022 ();
 sg13g2_decap_8 FILLER_12_2029 ();
 sg13g2_fill_2 FILLER_12_2080 ();
 sg13g2_fill_1 FILLER_12_2082 ();
 sg13g2_decap_4 FILLER_12_2087 ();
 sg13g2_fill_2 FILLER_12_2091 ();
 sg13g2_fill_2 FILLER_12_2097 ();
 sg13g2_fill_2 FILLER_12_2109 ();
 sg13g2_fill_1 FILLER_12_2111 ();
 sg13g2_fill_1 FILLER_12_2160 ();
 sg13g2_decap_4 FILLER_12_2195 ();
 sg13g2_decap_8 FILLER_12_2209 ();
 sg13g2_decap_8 FILLER_12_2216 ();
 sg13g2_fill_1 FILLER_12_2223 ();
 sg13g2_decap_8 FILLER_12_2253 ();
 sg13g2_decap_4 FILLER_12_2260 ();
 sg13g2_fill_1 FILLER_12_2268 ();
 sg13g2_decap_4 FILLER_12_2295 ();
 sg13g2_fill_2 FILLER_12_2303 ();
 sg13g2_fill_1 FILLER_12_2305 ();
 sg13g2_decap_8 FILLER_12_2357 ();
 sg13g2_decap_4 FILLER_12_2364 ();
 sg13g2_fill_2 FILLER_12_2368 ();
 sg13g2_fill_2 FILLER_12_2400 ();
 sg13g2_fill_1 FILLER_12_2408 ();
 sg13g2_fill_2 FILLER_12_2452 ();
 sg13g2_decap_8 FILLER_12_2480 ();
 sg13g2_fill_1 FILLER_12_2487 ();
 sg13g2_decap_4 FILLER_12_2502 ();
 sg13g2_decap_8 FILLER_12_2543 ();
 sg13g2_decap_4 FILLER_12_2550 ();
 sg13g2_fill_1 FILLER_12_2554 ();
 sg13g2_decap_4 FILLER_12_2559 ();
 sg13g2_fill_1 FILLER_12_2563 ();
 sg13g2_decap_8 FILLER_12_2589 ();
 sg13g2_decap_8 FILLER_12_2596 ();
 sg13g2_decap_8 FILLER_12_2603 ();
 sg13g2_decap_8 FILLER_12_2610 ();
 sg13g2_decap_8 FILLER_12_2617 ();
 sg13g2_decap_8 FILLER_12_2624 ();
 sg13g2_decap_8 FILLER_12_2631 ();
 sg13g2_decap_8 FILLER_12_2638 ();
 sg13g2_decap_8 FILLER_12_2645 ();
 sg13g2_decap_8 FILLER_12_2652 ();
 sg13g2_decap_8 FILLER_12_2659 ();
 sg13g2_decap_4 FILLER_12_2666 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_17 ();
 sg13g2_fill_1 FILLER_13_24 ();
 sg13g2_decap_4 FILLER_13_41 ();
 sg13g2_fill_1 FILLER_13_45 ();
 sg13g2_fill_2 FILLER_13_86 ();
 sg13g2_decap_8 FILLER_13_93 ();
 sg13g2_fill_2 FILLER_13_120 ();
 sg13g2_fill_2 FILLER_13_137 ();
 sg13g2_fill_1 FILLER_13_139 ();
 sg13g2_decap_4 FILLER_13_155 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_1 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_200 ();
 sg13g2_fill_1 FILLER_13_205 ();
 sg13g2_fill_1 FILLER_13_212 ();
 sg13g2_fill_1 FILLER_13_217 ();
 sg13g2_decap_4 FILLER_13_223 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_255 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_decap_8 FILLER_13_297 ();
 sg13g2_decap_4 FILLER_13_304 ();
 sg13g2_fill_2 FILLER_13_308 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_411 ();
 sg13g2_fill_1 FILLER_13_419 ();
 sg13g2_fill_2 FILLER_13_463 ();
 sg13g2_decap_4 FILLER_13_499 ();
 sg13g2_fill_1 FILLER_13_503 ();
 sg13g2_decap_8 FILLER_13_508 ();
 sg13g2_fill_2 FILLER_13_515 ();
 sg13g2_fill_1 FILLER_13_517 ();
 sg13g2_decap_4 FILLER_13_548 ();
 sg13g2_fill_1 FILLER_13_552 ();
 sg13g2_fill_2 FILLER_13_558 ();
 sg13g2_fill_1 FILLER_13_560 ();
 sg13g2_fill_2 FILLER_13_584 ();
 sg13g2_fill_1 FILLER_13_586 ();
 sg13g2_fill_2 FILLER_13_624 ();
 sg13g2_fill_2 FILLER_13_630 ();
 sg13g2_fill_1 FILLER_13_636 ();
 sg13g2_fill_1 FILLER_13_668 ();
 sg13g2_fill_2 FILLER_13_673 ();
 sg13g2_fill_2 FILLER_13_680 ();
 sg13g2_fill_1 FILLER_13_686 ();
 sg13g2_fill_2 FILLER_13_691 ();
 sg13g2_fill_1 FILLER_13_693 ();
 sg13g2_fill_2 FILLER_13_699 ();
 sg13g2_fill_1 FILLER_13_701 ();
 sg13g2_decap_4 FILLER_13_732 ();
 sg13g2_fill_2 FILLER_13_736 ();
 sg13g2_fill_2 FILLER_13_809 ();
 sg13g2_fill_2 FILLER_13_815 ();
 sg13g2_fill_1 FILLER_13_817 ();
 sg13g2_fill_1 FILLER_13_828 ();
 sg13g2_fill_2 FILLER_13_850 ();
 sg13g2_fill_1 FILLER_13_852 ();
 sg13g2_decap_8 FILLER_13_857 ();
 sg13g2_decap_4 FILLER_13_864 ();
 sg13g2_fill_2 FILLER_13_868 ();
 sg13g2_fill_1 FILLER_13_900 ();
 sg13g2_decap_8 FILLER_13_905 ();
 sg13g2_decap_4 FILLER_13_912 ();
 sg13g2_fill_2 FILLER_13_916 ();
 sg13g2_decap_8 FILLER_13_937 ();
 sg13g2_fill_1 FILLER_13_944 ();
 sg13g2_fill_1 FILLER_13_954 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_fill_2 FILLER_13_1001 ();
 sg13g2_fill_1 FILLER_13_1038 ();
 sg13g2_fill_1 FILLER_13_1074 ();
 sg13g2_fill_2 FILLER_13_1079 ();
 sg13g2_decap_8 FILLER_13_1134 ();
 sg13g2_decap_4 FILLER_13_1141 ();
 sg13g2_decap_8 FILLER_13_1153 ();
 sg13g2_fill_1 FILLER_13_1204 ();
 sg13g2_fill_2 FILLER_13_1250 ();
 sg13g2_fill_1 FILLER_13_1252 ();
 sg13g2_decap_8 FILLER_13_1263 ();
 sg13g2_decap_8 FILLER_13_1270 ();
 sg13g2_fill_2 FILLER_13_1277 ();
 sg13g2_fill_1 FILLER_13_1284 ();
 sg13g2_fill_1 FILLER_13_1300 ();
 sg13g2_decap_4 FILLER_13_1316 ();
 sg13g2_fill_2 FILLER_13_1320 ();
 sg13g2_decap_8 FILLER_13_1351 ();
 sg13g2_decap_4 FILLER_13_1358 ();
 sg13g2_fill_1 FILLER_13_1362 ();
 sg13g2_fill_2 FILLER_13_1367 ();
 sg13g2_fill_1 FILLER_13_1369 ();
 sg13g2_decap_4 FILLER_13_1406 ();
 sg13g2_fill_2 FILLER_13_1442 ();
 sg13g2_fill_1 FILLER_13_1469 ();
 sg13g2_fill_1 FILLER_13_1477 ();
 sg13g2_fill_1 FILLER_13_1491 ();
 sg13g2_fill_2 FILLER_13_1514 ();
 sg13g2_fill_2 FILLER_13_1556 ();
 sg13g2_decap_8 FILLER_13_1573 ();
 sg13g2_fill_1 FILLER_13_1585 ();
 sg13g2_decap_8 FILLER_13_1612 ();
 sg13g2_fill_1 FILLER_13_1619 ();
 sg13g2_decap_8 FILLER_13_1630 ();
 sg13g2_decap_8 FILLER_13_1637 ();
 sg13g2_fill_2 FILLER_13_1644 ();
 sg13g2_fill_1 FILLER_13_1646 ();
 sg13g2_decap_8 FILLER_13_1653 ();
 sg13g2_decap_8 FILLER_13_1660 ();
 sg13g2_fill_2 FILLER_13_1667 ();
 sg13g2_fill_2 FILLER_13_1699 ();
 sg13g2_fill_1 FILLER_13_1701 ();
 sg13g2_fill_2 FILLER_13_1747 ();
 sg13g2_fill_1 FILLER_13_1772 ();
 sg13g2_fill_2 FILLER_13_1781 ();
 sg13g2_fill_1 FILLER_13_1802 ();
 sg13g2_fill_2 FILLER_13_1842 ();
 sg13g2_fill_1 FILLER_13_1844 ();
 sg13g2_fill_1 FILLER_13_1849 ();
 sg13g2_fill_2 FILLER_13_1856 ();
 sg13g2_fill_1 FILLER_13_1863 ();
 sg13g2_fill_2 FILLER_13_1890 ();
 sg13g2_fill_1 FILLER_13_1968 ();
 sg13g2_decap_4 FILLER_13_1995 ();
 sg13g2_fill_2 FILLER_13_2013 ();
 sg13g2_fill_1 FILLER_13_2015 ();
 sg13g2_decap_8 FILLER_13_2020 ();
 sg13g2_decap_8 FILLER_13_2027 ();
 sg13g2_decap_4 FILLER_13_2034 ();
 sg13g2_fill_1 FILLER_13_2074 ();
 sg13g2_fill_1 FILLER_13_2080 ();
 sg13g2_fill_2 FILLER_13_2138 ();
 sg13g2_decap_8 FILLER_13_2169 ();
 sg13g2_fill_1 FILLER_13_2245 ();
 sg13g2_fill_2 FILLER_13_2256 ();
 sg13g2_decap_4 FILLER_13_2354 ();
 sg13g2_decap_4 FILLER_13_2363 ();
 sg13g2_fill_2 FILLER_13_2367 ();
 sg13g2_fill_1 FILLER_13_2442 ();
 sg13g2_fill_1 FILLER_13_2500 ();
 sg13g2_decap_8 FILLER_13_2527 ();
 sg13g2_decap_4 FILLER_13_2534 ();
 sg13g2_fill_1 FILLER_13_2538 ();
 sg13g2_decap_4 FILLER_13_2575 ();
 sg13g2_fill_1 FILLER_13_2589 ();
 sg13g2_decap_8 FILLER_13_2616 ();
 sg13g2_decap_8 FILLER_13_2623 ();
 sg13g2_decap_8 FILLER_13_2630 ();
 sg13g2_decap_8 FILLER_13_2637 ();
 sg13g2_decap_8 FILLER_13_2644 ();
 sg13g2_decap_8 FILLER_13_2651 ();
 sg13g2_decap_8 FILLER_13_2658 ();
 sg13g2_decap_4 FILLER_13_2665 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_fill_2 FILLER_14_0 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_decap_8 FILLER_14_93 ();
 sg13g2_decap_8 FILLER_14_100 ();
 sg13g2_decap_4 FILLER_14_107 ();
 sg13g2_fill_2 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_132 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_decap_8 FILLER_14_139 ();
 sg13g2_fill_2 FILLER_14_146 ();
 sg13g2_fill_1 FILLER_14_148 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_fill_2 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_172 ();
 sg13g2_fill_1 FILLER_14_179 ();
 sg13g2_fill_1 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_195 ();
 sg13g2_decap_8 FILLER_14_201 ();
 sg13g2_decap_8 FILLER_14_208 ();
 sg13g2_decap_4 FILLER_14_215 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_235 ();
 sg13g2_decap_8 FILLER_14_240 ();
 sg13g2_decap_8 FILLER_14_247 ();
 sg13g2_decap_4 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_337 ();
 sg13g2_decap_4 FILLER_14_344 ();
 sg13g2_fill_2 FILLER_14_348 ();
 sg13g2_fill_1 FILLER_14_367 ();
 sg13g2_fill_1 FILLER_14_403 ();
 sg13g2_fill_2 FILLER_14_448 ();
 sg13g2_fill_1 FILLER_14_467 ();
 sg13g2_fill_2 FILLER_14_472 ();
 sg13g2_fill_1 FILLER_14_484 ();
 sg13g2_decap_4 FILLER_14_537 ();
 sg13g2_fill_1 FILLER_14_541 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_fill_1 FILLER_14_560 ();
 sg13g2_fill_1 FILLER_14_573 ();
 sg13g2_fill_2 FILLER_14_579 ();
 sg13g2_fill_1 FILLER_14_581 ();
 sg13g2_fill_2 FILLER_14_591 ();
 sg13g2_fill_1 FILLER_14_593 ();
 sg13g2_fill_1 FILLER_14_598 ();
 sg13g2_decap_4 FILLER_14_662 ();
 sg13g2_fill_2 FILLER_14_666 ();
 sg13g2_fill_2 FILLER_14_673 ();
 sg13g2_fill_2 FILLER_14_680 ();
 sg13g2_fill_2 FILLER_14_691 ();
 sg13g2_fill_1 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_734 ();
 sg13g2_fill_2 FILLER_14_741 ();
 sg13g2_fill_1 FILLER_14_743 ();
 sg13g2_fill_1 FILLER_14_794 ();
 sg13g2_decap_8 FILLER_14_799 ();
 sg13g2_decap_8 FILLER_14_806 ();
 sg13g2_decap_8 FILLER_14_813 ();
 sg13g2_decap_8 FILLER_14_820 ();
 sg13g2_decap_8 FILLER_14_827 ();
 sg13g2_fill_2 FILLER_14_834 ();
 sg13g2_decap_8 FILLER_14_846 ();
 sg13g2_decap_8 FILLER_14_853 ();
 sg13g2_decap_8 FILLER_14_860 ();
 sg13g2_decap_8 FILLER_14_867 ();
 sg13g2_fill_1 FILLER_14_874 ();
 sg13g2_decap_4 FILLER_14_880 ();
 sg13g2_fill_1 FILLER_14_889 ();
 sg13g2_fill_1 FILLER_14_895 ();
 sg13g2_fill_1 FILLER_14_900 ();
 sg13g2_fill_1 FILLER_14_932 ();
 sg13g2_fill_1 FILLER_14_959 ();
 sg13g2_decap_4 FILLER_14_969 ();
 sg13g2_fill_2 FILLER_14_973 ();
 sg13g2_fill_1 FILLER_14_1001 ();
 sg13g2_decap_4 FILLER_14_1010 ();
 sg13g2_fill_1 FILLER_14_1014 ();
 sg13g2_decap_4 FILLER_14_1040 ();
 sg13g2_fill_1 FILLER_14_1052 ();
 sg13g2_decap_4 FILLER_14_1079 ();
 sg13g2_fill_1 FILLER_14_1083 ();
 sg13g2_fill_2 FILLER_14_1115 ();
 sg13g2_fill_1 FILLER_14_1117 ();
 sg13g2_fill_2 FILLER_14_1144 ();
 sg13g2_fill_1 FILLER_14_1146 ();
 sg13g2_decap_8 FILLER_14_1177 ();
 sg13g2_fill_2 FILLER_14_1184 ();
 sg13g2_decap_4 FILLER_14_1199 ();
 sg13g2_fill_2 FILLER_14_1203 ();
 sg13g2_fill_1 FILLER_14_1236 ();
 sg13g2_decap_4 FILLER_14_1273 ();
 sg13g2_decap_4 FILLER_14_1315 ();
 sg13g2_fill_2 FILLER_14_1345 ();
 sg13g2_fill_1 FILLER_14_1347 ();
 sg13g2_fill_2 FILLER_14_1358 ();
 sg13g2_fill_2 FILLER_14_1386 ();
 sg13g2_decap_4 FILLER_14_1392 ();
 sg13g2_decap_8 FILLER_14_1401 ();
 sg13g2_decap_8 FILLER_14_1408 ();
 sg13g2_decap_4 FILLER_14_1415 ();
 sg13g2_decap_8 FILLER_14_1424 ();
 sg13g2_decap_4 FILLER_14_1431 ();
 sg13g2_decap_4 FILLER_14_1450 ();
 sg13g2_fill_1 FILLER_14_1454 ();
 sg13g2_fill_1 FILLER_14_1492 ();
 sg13g2_fill_1 FILLER_14_1506 ();
 sg13g2_fill_1 FILLER_14_1570 ();
 sg13g2_fill_2 FILLER_14_1578 ();
 sg13g2_fill_1 FILLER_14_1580 ();
 sg13g2_decap_8 FILLER_14_1589 ();
 sg13g2_decap_4 FILLER_14_1596 ();
 sg13g2_fill_2 FILLER_14_1618 ();
 sg13g2_decap_8 FILLER_14_1636 ();
 sg13g2_fill_2 FILLER_14_1643 ();
 sg13g2_fill_2 FILLER_14_1739 ();
 sg13g2_fill_2 FILLER_14_1764 ();
 sg13g2_fill_1 FILLER_14_1771 ();
 sg13g2_fill_1 FILLER_14_1948 ();
 sg13g2_decap_8 FILLER_14_1993 ();
 sg13g2_decap_8 FILLER_14_2000 ();
 sg13g2_decap_8 FILLER_14_2033 ();
 sg13g2_fill_1 FILLER_14_2053 ();
 sg13g2_decap_8 FILLER_14_2058 ();
 sg13g2_decap_8 FILLER_14_2065 ();
 sg13g2_decap_8 FILLER_14_2072 ();
 sg13g2_decap_8 FILLER_14_2105 ();
 sg13g2_decap_8 FILLER_14_2112 ();
 sg13g2_decap_4 FILLER_14_2133 ();
 sg13g2_fill_1 FILLER_14_2137 ();
 sg13g2_decap_8 FILLER_14_2174 ();
 sg13g2_decap_8 FILLER_14_2181 ();
 sg13g2_fill_2 FILLER_14_2188 ();
 sg13g2_fill_1 FILLER_14_2190 ();
 sg13g2_decap_8 FILLER_14_2201 ();
 sg13g2_decap_8 FILLER_14_2208 ();
 sg13g2_fill_2 FILLER_14_2219 ();
 sg13g2_fill_1 FILLER_14_2221 ();
 sg13g2_fill_1 FILLER_14_2230 ();
 sg13g2_fill_1 FILLER_14_2245 ();
 sg13g2_decap_8 FILLER_14_2273 ();
 sg13g2_decap_8 FILLER_14_2280 ();
 sg13g2_fill_2 FILLER_14_2287 ();
 sg13g2_fill_1 FILLER_14_2289 ();
 sg13g2_fill_2 FILLER_14_2300 ();
 sg13g2_fill_1 FILLER_14_2302 ();
 sg13g2_fill_1 FILLER_14_2311 ();
 sg13g2_fill_1 FILLER_14_2316 ();
 sg13g2_fill_2 FILLER_14_2330 ();
 sg13g2_fill_1 FILLER_14_2358 ();
 sg13g2_decap_4 FILLER_14_2363 ();
 sg13g2_fill_1 FILLER_14_2431 ();
 sg13g2_fill_1 FILLER_14_2489 ();
 sg13g2_decap_8 FILLER_14_2520 ();
 sg13g2_decap_8 FILLER_14_2527 ();
 sg13g2_decap_4 FILLER_14_2544 ();
 sg13g2_decap_4 FILLER_14_2574 ();
 sg13g2_decap_8 FILLER_14_2614 ();
 sg13g2_decap_8 FILLER_14_2621 ();
 sg13g2_decap_8 FILLER_14_2628 ();
 sg13g2_decap_8 FILLER_14_2635 ();
 sg13g2_decap_8 FILLER_14_2642 ();
 sg13g2_decap_8 FILLER_14_2649 ();
 sg13g2_decap_8 FILLER_14_2656 ();
 sg13g2_decap_8 FILLER_14_2663 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_13 ();
 sg13g2_decap_8 FILLER_15_20 ();
 sg13g2_decap_8 FILLER_15_31 ();
 sg13g2_fill_2 FILLER_15_71 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_1 FILLER_15_82 ();
 sg13g2_decap_4 FILLER_15_93 ();
 sg13g2_fill_1 FILLER_15_97 ();
 sg13g2_fill_2 FILLER_15_129 ();
 sg13g2_fill_1 FILLER_15_131 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_decap_4 FILLER_15_210 ();
 sg13g2_decap_4 FILLER_15_250 ();
 sg13g2_decap_4 FILLER_15_331 ();
 sg13g2_decap_8 FILLER_15_345 ();
 sg13g2_decap_4 FILLER_15_352 ();
 sg13g2_fill_1 FILLER_15_356 ();
 sg13g2_decap_8 FILLER_15_366 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_decap_4 FILLER_15_388 ();
 sg13g2_fill_2 FILLER_15_392 ();
 sg13g2_fill_1 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_15_419 ();
 sg13g2_fill_2 FILLER_15_444 ();
 sg13g2_decap_8 FILLER_15_485 ();
 sg13g2_fill_1 FILLER_15_492 ();
 sg13g2_fill_1 FILLER_15_498 ();
 sg13g2_decap_4 FILLER_15_512 ();
 sg13g2_fill_1 FILLER_15_530 ();
 sg13g2_decap_8 FILLER_15_535 ();
 sg13g2_fill_2 FILLER_15_542 ();
 sg13g2_fill_2 FILLER_15_582 ();
 sg13g2_decap_4 FILLER_15_594 ();
 sg13g2_fill_1 FILLER_15_598 ();
 sg13g2_fill_2 FILLER_15_604 ();
 sg13g2_fill_1 FILLER_15_606 ();
 sg13g2_fill_2 FILLER_15_619 ();
 sg13g2_fill_1 FILLER_15_621 ();
 sg13g2_decap_8 FILLER_15_661 ();
 sg13g2_decap_8 FILLER_15_668 ();
 sg13g2_decap_8 FILLER_15_675 ();
 sg13g2_decap_4 FILLER_15_682 ();
 sg13g2_fill_1 FILLER_15_695 ();
 sg13g2_fill_1 FILLER_15_701 ();
 sg13g2_fill_2 FILLER_15_737 ();
 sg13g2_fill_1 FILLER_15_739 ();
 sg13g2_fill_1 FILLER_15_750 ();
 sg13g2_fill_2 FILLER_15_771 ();
 sg13g2_decap_8 FILLER_15_778 ();
 sg13g2_decap_8 FILLER_15_785 ();
 sg13g2_decap_8 FILLER_15_792 ();
 sg13g2_decap_8 FILLER_15_799 ();
 sg13g2_decap_8 FILLER_15_806 ();
 sg13g2_decap_8 FILLER_15_813 ();
 sg13g2_decap_8 FILLER_15_860 ();
 sg13g2_decap_4 FILLER_15_867 ();
 sg13g2_fill_2 FILLER_15_871 ();
 sg13g2_decap_8 FILLER_15_899 ();
 sg13g2_decap_8 FILLER_15_906 ();
 sg13g2_decap_8 FILLER_15_913 ();
 sg13g2_fill_2 FILLER_15_937 ();
 sg13g2_decap_8 FILLER_15_943 ();
 sg13g2_fill_2 FILLER_15_950 ();
 sg13g2_fill_1 FILLER_15_996 ();
 sg13g2_decap_4 FILLER_15_1040 ();
 sg13g2_fill_2 FILLER_15_1044 ();
 sg13g2_decap_4 FILLER_15_1054 ();
 sg13g2_fill_1 FILLER_15_1058 ();
 sg13g2_decap_8 FILLER_15_1080 ();
 sg13g2_decap_8 FILLER_15_1087 ();
 sg13g2_fill_2 FILLER_15_1094 ();
 sg13g2_fill_2 FILLER_15_1100 ();
 sg13g2_decap_8 FILLER_15_1106 ();
 sg13g2_decap_4 FILLER_15_1113 ();
 sg13g2_decap_8 FILLER_15_1147 ();
 sg13g2_fill_2 FILLER_15_1198 ();
 sg13g2_fill_2 FILLER_15_1204 ();
 sg13g2_decap_4 FILLER_15_1280 ();
 sg13g2_fill_2 FILLER_15_1284 ();
 sg13g2_fill_2 FILLER_15_1290 ();
 sg13g2_fill_1 FILLER_15_1328 ();
 sg13g2_decap_8 FILLER_15_1337 ();
 sg13g2_decap_4 FILLER_15_1344 ();
 sg13g2_fill_2 FILLER_15_1348 ();
 sg13g2_fill_2 FILLER_15_1412 ();
 sg13g2_fill_2 FILLER_15_1436 ();
 sg13g2_fill_1 FILLER_15_1461 ();
 sg13g2_fill_1 FILLER_15_1467 ();
 sg13g2_fill_1 FILLER_15_1519 ();
 sg13g2_decap_8 FILLER_15_1531 ();
 sg13g2_decap_4 FILLER_15_1538 ();
 sg13g2_fill_2 FILLER_15_1542 ();
 sg13g2_decap_4 FILLER_15_1548 ();
 sg13g2_decap_8 FILLER_15_1589 ();
 sg13g2_decap_4 FILLER_15_1596 ();
 sg13g2_fill_1 FILLER_15_1600 ();
 sg13g2_fill_1 FILLER_15_1606 ();
 sg13g2_fill_1 FILLER_15_1617 ();
 sg13g2_decap_4 FILLER_15_1654 ();
 sg13g2_fill_2 FILLER_15_1658 ();
 sg13g2_fill_1 FILLER_15_1673 ();
 sg13g2_fill_1 FILLER_15_1696 ();
 sg13g2_fill_1 FILLER_15_1700 ();
 sg13g2_fill_2 FILLER_15_1704 ();
 sg13g2_fill_1 FILLER_15_1706 ();
 sg13g2_fill_2 FILLER_15_1715 ();
 sg13g2_fill_1 FILLER_15_1735 ();
 sg13g2_fill_2 FILLER_15_1741 ();
 sg13g2_fill_2 FILLER_15_1758 ();
 sg13g2_fill_1 FILLER_15_1765 ();
 sg13g2_fill_2 FILLER_15_1798 ();
 sg13g2_fill_2 FILLER_15_1842 ();
 sg13g2_fill_1 FILLER_15_1876 ();
 sg13g2_fill_1 FILLER_15_1911 ();
 sg13g2_decap_8 FILLER_15_1962 ();
 sg13g2_decap_8 FILLER_15_1969 ();
 sg13g2_decap_8 FILLER_15_1980 ();
 sg13g2_fill_2 FILLER_15_1987 ();
 sg13g2_fill_1 FILLER_15_1989 ();
 sg13g2_fill_1 FILLER_15_2000 ();
 sg13g2_decap_4 FILLER_15_2031 ();
 sg13g2_fill_2 FILLER_15_2035 ();
 sg13g2_decap_4 FILLER_15_2073 ();
 sg13g2_decap_8 FILLER_15_2107 ();
 sg13g2_decap_8 FILLER_15_2114 ();
 sg13g2_decap_4 FILLER_15_2121 ();
 sg13g2_fill_1 FILLER_15_2125 ();
 sg13g2_decap_8 FILLER_15_2130 ();
 sg13g2_decap_4 FILLER_15_2137 ();
 sg13g2_fill_1 FILLER_15_2141 ();
 sg13g2_decap_4 FILLER_15_2168 ();
 sg13g2_fill_2 FILLER_15_2172 ();
 sg13g2_decap_4 FILLER_15_2188 ();
 sg13g2_decap_8 FILLER_15_2222 ();
 sg13g2_decap_8 FILLER_15_2229 ();
 sg13g2_decap_4 FILLER_15_2236 ();
 sg13g2_decap_8 FILLER_15_2260 ();
 sg13g2_decap_8 FILLER_15_2267 ();
 sg13g2_fill_1 FILLER_15_2274 ();
 sg13g2_fill_1 FILLER_15_2322 ();
 sg13g2_fill_1 FILLER_15_2336 ();
 sg13g2_fill_2 FILLER_15_2379 ();
 sg13g2_fill_1 FILLER_15_2381 ();
 sg13g2_fill_2 FILLER_15_2418 ();
 sg13g2_fill_1 FILLER_15_2483 ();
 sg13g2_decap_8 FILLER_15_2508 ();
 sg13g2_fill_1 FILLER_15_2515 ();
 sg13g2_decap_4 FILLER_15_2546 ();
 sg13g2_fill_2 FILLER_15_2593 ();
 sg13g2_decap_8 FILLER_15_2603 ();
 sg13g2_decap_8 FILLER_15_2610 ();
 sg13g2_decap_8 FILLER_15_2617 ();
 sg13g2_decap_8 FILLER_15_2624 ();
 sg13g2_decap_8 FILLER_15_2631 ();
 sg13g2_decap_8 FILLER_15_2638 ();
 sg13g2_decap_8 FILLER_15_2645 ();
 sg13g2_decap_8 FILLER_15_2652 ();
 sg13g2_decap_8 FILLER_15_2659 ();
 sg13g2_decap_4 FILLER_15_2666 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_59 ();
 sg13g2_fill_1 FILLER_16_66 ();
 sg13g2_fill_2 FILLER_16_76 ();
 sg13g2_fill_1 FILLER_16_78 ();
 sg13g2_decap_4 FILLER_16_90 ();
 sg13g2_fill_2 FILLER_16_94 ();
 sg13g2_fill_2 FILLER_16_145 ();
 sg13g2_fill_1 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_2 FILLER_16_212 ();
 sg13g2_fill_1 FILLER_16_214 ();
 sg13g2_decap_8 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_fill_1 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_decap_4 FILLER_16_281 ();
 sg13g2_fill_2 FILLER_16_285 ();
 sg13g2_fill_1 FILLER_16_292 ();
 sg13g2_fill_1 FILLER_16_297 ();
 sg13g2_fill_1 FILLER_16_303 ();
 sg13g2_fill_2 FILLER_16_313 ();
 sg13g2_fill_1 FILLER_16_320 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_decap_4 FILLER_16_359 ();
 sg13g2_fill_2 FILLER_16_367 ();
 sg13g2_fill_2 FILLER_16_420 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_fill_1 FILLER_16_441 ();
 sg13g2_decap_4 FILLER_16_459 ();
 sg13g2_fill_1 FILLER_16_463 ();
 sg13g2_fill_2 FILLER_16_470 ();
 sg13g2_decap_4 FILLER_16_476 ();
 sg13g2_fill_2 FILLER_16_480 ();
 sg13g2_fill_1 FILLER_16_504 ();
 sg13g2_fill_2 FILLER_16_509 ();
 sg13g2_fill_2 FILLER_16_542 ();
 sg13g2_fill_2 FILLER_16_588 ();
 sg13g2_fill_1 FILLER_16_590 ();
 sg13g2_decap_4 FILLER_16_597 ();
 sg13g2_fill_2 FILLER_16_620 ();
 sg13g2_fill_1 FILLER_16_622 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_fill_2 FILLER_16_672 ();
 sg13g2_fill_1 FILLER_16_674 ();
 sg13g2_fill_1 FILLER_16_706 ();
 sg13g2_fill_2 FILLER_16_711 ();
 sg13g2_fill_1 FILLER_16_713 ();
 sg13g2_fill_1 FILLER_16_718 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_fill_1 FILLER_16_772 ();
 sg13g2_fill_1 FILLER_16_782 ();
 sg13g2_decap_8 FILLER_16_792 ();
 sg13g2_decap_8 FILLER_16_799 ();
 sg13g2_fill_2 FILLER_16_842 ();
 sg13g2_fill_1 FILLER_16_844 ();
 sg13g2_fill_1 FILLER_16_871 ();
 sg13g2_fill_1 FILLER_16_882 ();
 sg13g2_fill_1 FILLER_16_930 ();
 sg13g2_fill_2 FILLER_16_957 ();
 sg13g2_decap_8 FILLER_16_967 ();
 sg13g2_decap_8 FILLER_16_974 ();
 sg13g2_fill_2 FILLER_16_981 ();
 sg13g2_fill_1 FILLER_16_983 ();
 sg13g2_decap_8 FILLER_16_989 ();
 sg13g2_decap_8 FILLER_16_996 ();
 sg13g2_fill_1 FILLER_16_1003 ();
 sg13g2_fill_2 FILLER_16_1008 ();
 sg13g2_fill_1 FILLER_16_1010 ();
 sg13g2_fill_1 FILLER_16_1016 ();
 sg13g2_decap_4 FILLER_16_1085 ();
 sg13g2_fill_1 FILLER_16_1098 ();
 sg13g2_fill_2 FILLER_16_1129 ();
 sg13g2_fill_1 FILLER_16_1131 ();
 sg13g2_decap_8 FILLER_16_1136 ();
 sg13g2_decap_8 FILLER_16_1143 ();
 sg13g2_fill_2 FILLER_16_1191 ();
 sg13g2_fill_2 FILLER_16_1276 ();
 sg13g2_decap_4 FILLER_16_1282 ();
 sg13g2_fill_1 FILLER_16_1286 ();
 sg13g2_fill_2 FILLER_16_1292 ();
 sg13g2_decap_8 FILLER_16_1299 ();
 sg13g2_fill_2 FILLER_16_1306 ();
 sg13g2_decap_8 FILLER_16_1312 ();
 sg13g2_decap_8 FILLER_16_1319 ();
 sg13g2_decap_8 FILLER_16_1326 ();
 sg13g2_decap_8 FILLER_16_1333 ();
 sg13g2_decap_8 FILLER_16_1340 ();
 sg13g2_decap_8 FILLER_16_1347 ();
 sg13g2_decap_4 FILLER_16_1354 ();
 sg13g2_fill_1 FILLER_16_1358 ();
 sg13g2_decap_8 FILLER_16_1393 ();
 sg13g2_fill_2 FILLER_16_1400 ();
 sg13g2_fill_1 FILLER_16_1402 ();
 sg13g2_fill_2 FILLER_16_1438 ();
 sg13g2_decap_4 FILLER_16_1446 ();
 sg13g2_fill_2 FILLER_16_1455 ();
 sg13g2_fill_1 FILLER_16_1472 ();
 sg13g2_fill_2 FILLER_16_1487 ();
 sg13g2_fill_1 FILLER_16_1494 ();
 sg13g2_fill_1 FILLER_16_1500 ();
 sg13g2_fill_2 FILLER_16_1512 ();
 sg13g2_fill_2 FILLER_16_1519 ();
 sg13g2_fill_2 FILLER_16_1539 ();
 sg13g2_fill_2 FILLER_16_1565 ();
 sg13g2_fill_1 FILLER_16_1567 ();
 sg13g2_fill_1 FILLER_16_1573 ();
 sg13g2_fill_2 FILLER_16_1595 ();
 sg13g2_decap_8 FILLER_16_1605 ();
 sg13g2_fill_2 FILLER_16_1616 ();
 sg13g2_fill_2 FILLER_16_1632 ();
 sg13g2_decap_8 FILLER_16_1666 ();
 sg13g2_fill_2 FILLER_16_1722 ();
 sg13g2_fill_1 FILLER_16_1766 ();
 sg13g2_fill_1 FILLER_16_1776 ();
 sg13g2_fill_2 FILLER_16_1782 ();
 sg13g2_fill_1 FILLER_16_1841 ();
 sg13g2_fill_2 FILLER_16_1852 ();
 sg13g2_fill_1 FILLER_16_1858 ();
 sg13g2_fill_2 FILLER_16_1885 ();
 sg13g2_fill_2 FILLER_16_1948 ();
 sg13g2_fill_1 FILLER_16_1954 ();
 sg13g2_fill_1 FILLER_16_1996 ();
 sg13g2_fill_1 FILLER_16_2011 ();
 sg13g2_fill_2 FILLER_16_2017 ();
 sg13g2_fill_1 FILLER_16_2019 ();
 sg13g2_decap_4 FILLER_16_2030 ();
 sg13g2_fill_1 FILLER_16_2034 ();
 sg13g2_fill_2 FILLER_16_2095 ();
 sg13g2_decap_8 FILLER_16_2123 ();
 sg13g2_decap_8 FILLER_16_2130 ();
 sg13g2_decap_4 FILLER_16_2147 ();
 sg13g2_decap_4 FILLER_16_2155 ();
 sg13g2_fill_1 FILLER_16_2193 ();
 sg13g2_fill_1 FILLER_16_2204 ();
 sg13g2_decap_4 FILLER_16_2362 ();
 sg13g2_fill_2 FILLER_16_2387 ();
 sg13g2_fill_1 FILLER_16_2415 ();
 sg13g2_fill_1 FILLER_16_2456 ();
 sg13g2_fill_2 FILLER_16_2488 ();
 sg13g2_fill_1 FILLER_16_2516 ();
 sg13g2_decap_8 FILLER_16_2547 ();
 sg13g2_fill_2 FILLER_16_2554 ();
 sg13g2_fill_1 FILLER_16_2556 ();
 sg13g2_decap_8 FILLER_16_2567 ();
 sg13g2_fill_2 FILLER_16_2574 ();
 sg13g2_fill_1 FILLER_16_2576 ();
 sg13g2_fill_1 FILLER_16_2581 ();
 sg13g2_decap_8 FILLER_16_2603 ();
 sg13g2_decap_8 FILLER_16_2636 ();
 sg13g2_decap_8 FILLER_16_2643 ();
 sg13g2_decap_8 FILLER_16_2650 ();
 sg13g2_decap_8 FILLER_16_2657 ();
 sg13g2_decap_4 FILLER_16_2664 ();
 sg13g2_fill_2 FILLER_16_2668 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_fill_1 FILLER_17_33 ();
 sg13g2_fill_1 FILLER_17_57 ();
 sg13g2_fill_1 FILLER_17_63 ();
 sg13g2_fill_2 FILLER_17_72 ();
 sg13g2_fill_1 FILLER_17_87 ();
 sg13g2_fill_2 FILLER_17_94 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_2 FILLER_17_111 ();
 sg13g2_fill_1 FILLER_17_113 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_1 FILLER_17_120 ();
 sg13g2_fill_2 FILLER_17_131 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_162 ();
 sg13g2_fill_1 FILLER_17_164 ();
 sg13g2_fill_1 FILLER_17_170 ();
 sg13g2_fill_1 FILLER_17_175 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_206 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_fill_1 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_233 ();
 sg13g2_fill_2 FILLER_17_240 ();
 sg13g2_fill_1 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_247 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_265 ();
 sg13g2_decap_4 FILLER_17_272 ();
 sg13g2_fill_2 FILLER_17_276 ();
 sg13g2_decap_8 FILLER_17_283 ();
 sg13g2_fill_1 FILLER_17_290 ();
 sg13g2_decap_8 FILLER_17_303 ();
 sg13g2_decap_4 FILLER_17_310 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_327 ();
 sg13g2_decap_4 FILLER_17_339 ();
 sg13g2_fill_1 FILLER_17_374 ();
 sg13g2_fill_2 FILLER_17_395 ();
 sg13g2_fill_1 FILLER_17_403 ();
 sg13g2_fill_1 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_470 ();
 sg13g2_fill_2 FILLER_17_477 ();
 sg13g2_fill_2 FILLER_17_484 ();
 sg13g2_decap_8 FILLER_17_491 ();
 sg13g2_fill_1 FILLER_17_498 ();
 sg13g2_fill_2 FILLER_17_538 ();
 sg13g2_fill_2 FILLER_17_586 ();
 sg13g2_fill_1 FILLER_17_588 ();
 sg13g2_decap_4 FILLER_17_630 ();
 sg13g2_fill_1 FILLER_17_634 ();
 sg13g2_fill_1 FILLER_17_649 ();
 sg13g2_fill_2 FILLER_17_676 ();
 sg13g2_fill_2 FILLER_17_733 ();
 sg13g2_fill_2 FILLER_17_739 ();
 sg13g2_decap_4 FILLER_17_772 ();
 sg13g2_fill_2 FILLER_17_776 ();
 sg13g2_decap_8 FILLER_17_808 ();
 sg13g2_fill_1 FILLER_17_819 ();
 sg13g2_fill_2 FILLER_17_866 ();
 sg13g2_decap_4 FILLER_17_878 ();
 sg13g2_fill_1 FILLER_17_882 ();
 sg13g2_decap_8 FILLER_17_893 ();
 sg13g2_fill_2 FILLER_17_900 ();
 sg13g2_decap_4 FILLER_17_928 ();
 sg13g2_decap_8 FILLER_17_958 ();
 sg13g2_fill_2 FILLER_17_965 ();
 sg13g2_decap_8 FILLER_17_988 ();
 sg13g2_decap_8 FILLER_17_995 ();
 sg13g2_decap_8 FILLER_17_1002 ();
 sg13g2_decap_4 FILLER_17_1009 ();
 sg13g2_decap_8 FILLER_17_1124 ();
 sg13g2_decap_8 FILLER_17_1131 ();
 sg13g2_decap_8 FILLER_17_1138 ();
 sg13g2_decap_8 FILLER_17_1145 ();
 sg13g2_fill_2 FILLER_17_1152 ();
 sg13g2_decap_8 FILLER_17_1158 ();
 sg13g2_decap_8 FILLER_17_1165 ();
 sg13g2_fill_1 FILLER_17_1172 ();
 sg13g2_decap_8 FILLER_17_1177 ();
 sg13g2_decap_8 FILLER_17_1184 ();
 sg13g2_fill_2 FILLER_17_1196 ();
 sg13g2_fill_1 FILLER_17_1198 ();
 sg13g2_fill_1 FILLER_17_1203 ();
 sg13g2_fill_2 FILLER_17_1214 ();
 sg13g2_fill_2 FILLER_17_1231 ();
 sg13g2_fill_1 FILLER_17_1233 ();
 sg13g2_decap_4 FILLER_17_1246 ();
 sg13g2_fill_2 FILLER_17_1250 ();
 sg13g2_fill_1 FILLER_17_1262 ();
 sg13g2_fill_2 FILLER_17_1297 ();
 sg13g2_decap_4 FILLER_17_1335 ();
 sg13g2_decap_8 FILLER_17_1349 ();
 sg13g2_decap_8 FILLER_17_1356 ();
 sg13g2_decap_4 FILLER_17_1363 ();
 sg13g2_fill_2 FILLER_17_1367 ();
 sg13g2_decap_8 FILLER_17_1409 ();
 sg13g2_fill_1 FILLER_17_1431 ();
 sg13g2_decap_4 FILLER_17_1449 ();
 sg13g2_fill_2 FILLER_17_1453 ();
 sg13g2_fill_2 FILLER_17_1461 ();
 sg13g2_fill_1 FILLER_17_1463 ();
 sg13g2_fill_2 FILLER_17_1471 ();
 sg13g2_fill_1 FILLER_17_1473 ();
 sg13g2_decap_8 FILLER_17_1485 ();
 sg13g2_decap_8 FILLER_17_1499 ();
 sg13g2_decap_4 FILLER_17_1506 ();
 sg13g2_fill_2 FILLER_17_1510 ();
 sg13g2_fill_2 FILLER_17_1539 ();
 sg13g2_fill_1 FILLER_17_1541 ();
 sg13g2_decap_8 FILLER_17_1589 ();
 sg13g2_decap_8 FILLER_17_1606 ();
 sg13g2_decap_4 FILLER_17_1613 ();
 sg13g2_decap_8 FILLER_17_1679 ();
 sg13g2_decap_8 FILLER_17_1686 ();
 sg13g2_decap_8 FILLER_17_1693 ();
 sg13g2_fill_1 FILLER_17_1700 ();
 sg13g2_fill_2 FILLER_17_1709 ();
 sg13g2_fill_1 FILLER_17_1753 ();
 sg13g2_fill_1 FILLER_17_1777 ();
 sg13g2_fill_1 FILLER_17_1807 ();
 sg13g2_fill_2 FILLER_17_1818 ();
 sg13g2_fill_2 FILLER_17_1829 ();
 sg13g2_fill_1 FILLER_17_1841 ();
 sg13g2_fill_2 FILLER_17_1847 ();
 sg13g2_fill_2 FILLER_17_1863 ();
 sg13g2_decap_8 FILLER_17_1869 ();
 sg13g2_fill_2 FILLER_17_1880 ();
 sg13g2_fill_1 FILLER_17_1887 ();
 sg13g2_fill_1 FILLER_17_1894 ();
 sg13g2_decap_4 FILLER_17_1899 ();
 sg13g2_fill_2 FILLER_17_1903 ();
 sg13g2_fill_1 FILLER_17_1926 ();
 sg13g2_fill_1 FILLER_17_1954 ();
 sg13g2_fill_2 FILLER_17_2057 ();
 sg13g2_fill_1 FILLER_17_2059 ();
 sg13g2_fill_1 FILLER_17_2068 ();
 sg13g2_decap_4 FILLER_17_2083 ();
 sg13g2_fill_2 FILLER_17_2117 ();
 sg13g2_decap_4 FILLER_17_2145 ();
 sg13g2_decap_8 FILLER_17_2159 ();
 sg13g2_fill_2 FILLER_17_2166 ();
 sg13g2_fill_2 FILLER_17_2194 ();
 sg13g2_fill_1 FILLER_17_2217 ();
 sg13g2_fill_1 FILLER_17_2223 ();
 sg13g2_fill_1 FILLER_17_2250 ();
 sg13g2_fill_2 FILLER_17_2404 ();
 sg13g2_fill_2 FILLER_17_2442 ();
 sg13g2_fill_1 FILLER_17_2493 ();
 sg13g2_fill_2 FILLER_17_2530 ();
 sg13g2_decap_8 FILLER_17_2576 ();
 sg13g2_decap_8 FILLER_17_2583 ();
 sg13g2_decap_8 FILLER_17_2590 ();
 sg13g2_decap_4 FILLER_17_2597 ();
 sg13g2_fill_2 FILLER_17_2601 ();
 sg13g2_decap_8 FILLER_17_2621 ();
 sg13g2_decap_8 FILLER_17_2628 ();
 sg13g2_decap_8 FILLER_17_2635 ();
 sg13g2_decap_8 FILLER_17_2642 ();
 sg13g2_decap_8 FILLER_17_2649 ();
 sg13g2_decap_8 FILLER_17_2656 ();
 sg13g2_decap_8 FILLER_17_2663 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_7 ();
 sg13g2_decap_4 FILLER_18_17 ();
 sg13g2_fill_2 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_82 ();
 sg13g2_decap_8 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_107 ();
 sg13g2_decap_8 FILLER_18_114 ();
 sg13g2_decap_8 FILLER_18_121 ();
 sg13g2_decap_8 FILLER_18_128 ();
 sg13g2_decap_4 FILLER_18_135 ();
 sg13g2_fill_1 FILLER_18_139 ();
 sg13g2_fill_2 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_155 ();
 sg13g2_fill_1 FILLER_18_187 ();
 sg13g2_decap_4 FILLER_18_206 ();
 sg13g2_fill_1 FILLER_18_210 ();
 sg13g2_fill_1 FILLER_18_237 ();
 sg13g2_fill_2 FILLER_18_243 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_310 ();
 sg13g2_fill_1 FILLER_18_316 ();
 sg13g2_fill_2 FILLER_18_343 ();
 sg13g2_fill_1 FILLER_18_371 ();
 sg13g2_fill_1 FILLER_18_382 ();
 sg13g2_fill_2 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_402 ();
 sg13g2_decap_4 FILLER_18_409 ();
 sg13g2_fill_1 FILLER_18_446 ();
 sg13g2_fill_2 FILLER_18_479 ();
 sg13g2_fill_2 FILLER_18_524 ();
 sg13g2_fill_1 FILLER_18_526 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_fill_1 FILLER_18_539 ();
 sg13g2_decap_4 FILLER_18_544 ();
 sg13g2_fill_2 FILLER_18_562 ();
 sg13g2_fill_1 FILLER_18_564 ();
 sg13g2_fill_1 FILLER_18_569 ();
 sg13g2_fill_1 FILLER_18_580 ();
 sg13g2_fill_1 FILLER_18_591 ();
 sg13g2_fill_1 FILLER_18_598 ();
 sg13g2_fill_1 FILLER_18_603 ();
 sg13g2_decap_4 FILLER_18_633 ();
 sg13g2_fill_1 FILLER_18_637 ();
 sg13g2_fill_2 FILLER_18_647 ();
 sg13g2_fill_1 FILLER_18_649 ();
 sg13g2_fill_2 FILLER_18_655 ();
 sg13g2_fill_2 FILLER_18_661 ();
 sg13g2_fill_2 FILLER_18_675 ();
 sg13g2_fill_1 FILLER_18_686 ();
 sg13g2_fill_2 FILLER_18_696 ();
 sg13g2_fill_1 FILLER_18_698 ();
 sg13g2_decap_4 FILLER_18_709 ();
 sg13g2_fill_1 FILLER_18_713 ();
 sg13g2_fill_1 FILLER_18_722 ();
 sg13g2_fill_2 FILLER_18_737 ();
 sg13g2_decap_4 FILLER_18_748 ();
 sg13g2_fill_1 FILLER_18_752 ();
 sg13g2_fill_1 FILLER_18_776 ();
 sg13g2_decap_8 FILLER_18_808 ();
 sg13g2_decap_8 FILLER_18_815 ();
 sg13g2_fill_2 FILLER_18_822 ();
 sg13g2_fill_1 FILLER_18_824 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_4 FILLER_18_840 ();
 sg13g2_decap_4 FILLER_18_865 ();
 sg13g2_fill_1 FILLER_18_869 ();
 sg13g2_fill_1 FILLER_18_896 ();
 sg13g2_fill_1 FILLER_18_911 ();
 sg13g2_decap_8 FILLER_18_963 ();
 sg13g2_decap_4 FILLER_18_1006 ();
 sg13g2_decap_8 FILLER_18_1044 ();
 sg13g2_decap_4 FILLER_18_1051 ();
 sg13g2_fill_1 FILLER_18_1055 ();
 sg13g2_fill_2 FILLER_18_1061 ();
 sg13g2_decap_4 FILLER_18_1067 ();
 sg13g2_fill_2 FILLER_18_1071 ();
 sg13g2_fill_1 FILLER_18_1116 ();
 sg13g2_decap_4 FILLER_18_1183 ();
 sg13g2_fill_2 FILLER_18_1187 ();
 sg13g2_decap_8 FILLER_18_1194 ();
 sg13g2_fill_2 FILLER_18_1201 ();
 sg13g2_fill_2 FILLER_18_1211 ();
 sg13g2_fill_2 FILLER_18_1240 ();
 sg13g2_fill_1 FILLER_18_1242 ();
 sg13g2_fill_2 FILLER_18_1289 ();
 sg13g2_fill_1 FILLER_18_1291 ();
 sg13g2_fill_2 FILLER_18_1296 ();
 sg13g2_fill_1 FILLER_18_1312 ();
 sg13g2_fill_1 FILLER_18_1339 ();
 sg13g2_decap_4 FILLER_18_1366 ();
 sg13g2_fill_1 FILLER_18_1370 ();
 sg13g2_decap_8 FILLER_18_1381 ();
 sg13g2_decap_8 FILLER_18_1388 ();
 sg13g2_decap_8 FILLER_18_1395 ();
 sg13g2_decap_8 FILLER_18_1402 ();
 sg13g2_decap_8 FILLER_18_1409 ();
 sg13g2_decap_8 FILLER_18_1416 ();
 sg13g2_decap_8 FILLER_18_1423 ();
 sg13g2_decap_4 FILLER_18_1430 ();
 sg13g2_fill_1 FILLER_18_1434 ();
 sg13g2_fill_2 FILLER_18_1445 ();
 sg13g2_fill_1 FILLER_18_1453 ();
 sg13g2_decap_8 FILLER_18_1510 ();
 sg13g2_fill_1 FILLER_18_1517 ();
 sg13g2_fill_1 FILLER_18_1546 ();
 sg13g2_decap_4 FILLER_18_1551 ();
 sg13g2_decap_8 FILLER_18_1561 ();
 sg13g2_decap_8 FILLER_18_1568 ();
 sg13g2_decap_4 FILLER_18_1575 ();
 sg13g2_fill_1 FILLER_18_1579 ();
 sg13g2_decap_8 FILLER_18_1595 ();
 sg13g2_fill_2 FILLER_18_1602 ();
 sg13g2_fill_2 FILLER_18_1637 ();
 sg13g2_fill_1 FILLER_18_1639 ();
 sg13g2_fill_2 FILLER_18_1660 ();
 sg13g2_fill_1 FILLER_18_1672 ();
 sg13g2_fill_1 FILLER_18_1679 ();
 sg13g2_decap_8 FILLER_18_1684 ();
 sg13g2_decap_8 FILLER_18_1691 ();
 sg13g2_decap_4 FILLER_18_1702 ();
 sg13g2_fill_2 FILLER_18_1706 ();
 sg13g2_fill_1 FILLER_18_1713 ();
 sg13g2_fill_2 FILLER_18_1717 ();
 sg13g2_fill_2 FILLER_18_1730 ();
 sg13g2_decap_4 FILLER_18_1803 ();
 sg13g2_fill_1 FILLER_18_1814 ();
 sg13g2_decap_4 FILLER_18_1832 ();
 sg13g2_fill_2 FILLER_18_1836 ();
 sg13g2_decap_8 FILLER_18_1852 ();
 sg13g2_decap_8 FILLER_18_1859 ();
 sg13g2_decap_8 FILLER_18_1866 ();
 sg13g2_decap_8 FILLER_18_1873 ();
 sg13g2_decap_4 FILLER_18_1880 ();
 sg13g2_decap_8 FILLER_18_1894 ();
 sg13g2_decap_8 FILLER_18_1901 ();
 sg13g2_decap_8 FILLER_18_1908 ();
 sg13g2_decap_4 FILLER_18_1915 ();
 sg13g2_fill_1 FILLER_18_1934 ();
 sg13g2_fill_1 FILLER_18_1961 ();
 sg13g2_fill_2 FILLER_18_1983 ();
 sg13g2_decap_8 FILLER_18_2010 ();
 sg13g2_decap_4 FILLER_18_2017 ();
 sg13g2_fill_1 FILLER_18_2021 ();
 sg13g2_decap_4 FILLER_18_2043 ();
 sg13g2_fill_1 FILLER_18_2047 ();
 sg13g2_decap_8 FILLER_18_2052 ();
 sg13g2_fill_1 FILLER_18_2059 ();
 sg13g2_fill_2 FILLER_18_2111 ();
 sg13g2_fill_1 FILLER_18_2113 ();
 sg13g2_decap_4 FILLER_18_2140 ();
 sg13g2_fill_1 FILLER_18_2227 ();
 sg13g2_decap_8 FILLER_18_2267 ();
 sg13g2_fill_2 FILLER_18_2274 ();
 sg13g2_decap_8 FILLER_18_2304 ();
 sg13g2_fill_2 FILLER_18_2311 ();
 sg13g2_fill_1 FILLER_18_2313 ();
 sg13g2_decap_4 FILLER_18_2318 ();
 sg13g2_fill_2 FILLER_18_2361 ();
 sg13g2_decap_4 FILLER_18_2380 ();
 sg13g2_fill_1 FILLER_18_2443 ();
 sg13g2_fill_2 FILLER_18_2471 ();
 sg13g2_fill_2 FILLER_18_2504 ();
 sg13g2_fill_1 FILLER_18_2561 ();
 sg13g2_decap_8 FILLER_18_2588 ();
 sg13g2_fill_1 FILLER_18_2595 ();
 sg13g2_decap_8 FILLER_18_2632 ();
 sg13g2_decap_8 FILLER_18_2639 ();
 sg13g2_decap_8 FILLER_18_2646 ();
 sg13g2_decap_8 FILLER_18_2653 ();
 sg13g2_decap_8 FILLER_18_2660 ();
 sg13g2_fill_2 FILLER_18_2667 ();
 sg13g2_fill_1 FILLER_18_2669 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_decap_4 FILLER_19_37 ();
 sg13g2_fill_1 FILLER_19_41 ();
 sg13g2_fill_2 FILLER_19_51 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_74 ();
 sg13g2_fill_2 FILLER_19_93 ();
 sg13g2_fill_1 FILLER_19_116 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_1 FILLER_19_140 ();
 sg13g2_decap_4 FILLER_19_177 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_decap_8 FILLER_19_187 ();
 sg13g2_decap_4 FILLER_19_194 ();
 sg13g2_fill_1 FILLER_19_198 ();
 sg13g2_fill_2 FILLER_19_203 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_fill_1 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_247 ();
 sg13g2_fill_1 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_286 ();
 sg13g2_fill_1 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_323 ();
 sg13g2_decap_8 FILLER_19_328 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_4 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_19_401 ();
 sg13g2_fill_2 FILLER_19_438 ();
 sg13g2_fill_1 FILLER_19_448 ();
 sg13g2_fill_2 FILLER_19_464 ();
 sg13g2_decap_4 FILLER_19_482 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_4 FILLER_19_525 ();
 sg13g2_fill_2 FILLER_19_529 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_fill_1 FILLER_19_542 ();
 sg13g2_fill_2 FILLER_19_552 ();
 sg13g2_decap_4 FILLER_19_588 ();
 sg13g2_decap_4 FILLER_19_597 ();
 sg13g2_fill_1 FILLER_19_610 ();
 sg13g2_decap_4 FILLER_19_655 ();
 sg13g2_fill_1 FILLER_19_659 ();
 sg13g2_fill_1 FILLER_19_667 ();
 sg13g2_fill_1 FILLER_19_698 ();
 sg13g2_fill_2 FILLER_19_704 ();
 sg13g2_fill_1 FILLER_19_712 ();
 sg13g2_fill_1 FILLER_19_719 ();
 sg13g2_fill_1 FILLER_19_726 ();
 sg13g2_fill_1 FILLER_19_732 ();
 sg13g2_fill_2 FILLER_19_769 ();
 sg13g2_fill_1 FILLER_19_771 ();
 sg13g2_fill_2 FILLER_19_790 ();
 sg13g2_fill_1 FILLER_19_792 ();
 sg13g2_decap_4 FILLER_19_797 ();
 sg13g2_fill_1 FILLER_19_801 ();
 sg13g2_decap_8 FILLER_19_838 ();
 sg13g2_decap_8 FILLER_19_845 ();
 sg13g2_decap_8 FILLER_19_852 ();
 sg13g2_decap_8 FILLER_19_859 ();
 sg13g2_decap_8 FILLER_19_866 ();
 sg13g2_fill_2 FILLER_19_873 ();
 sg13g2_decap_8 FILLER_19_883 ();
 sg13g2_fill_2 FILLER_19_890 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_4 FILLER_19_903 ();
 sg13g2_fill_1 FILLER_19_907 ();
 sg13g2_decap_4 FILLER_19_935 ();
 sg13g2_decap_4 FILLER_19_943 ();
 sg13g2_fill_1 FILLER_19_947 ();
 sg13g2_fill_2 FILLER_19_999 ();
 sg13g2_fill_1 FILLER_19_1001 ();
 sg13g2_decap_4 FILLER_19_1007 ();
 sg13g2_fill_1 FILLER_19_1011 ();
 sg13g2_decap_4 FILLER_19_1016 ();
 sg13g2_fill_1 FILLER_19_1020 ();
 sg13g2_decap_4 FILLER_19_1034 ();
 sg13g2_fill_1 FILLER_19_1038 ();
 sg13g2_decap_4 FILLER_19_1064 ();
 sg13g2_fill_1 FILLER_19_1072 ();
 sg13g2_fill_1 FILLER_19_1103 ();
 sg13g2_decap_4 FILLER_19_1125 ();
 sg13g2_fill_1 FILLER_19_1129 ();
 sg13g2_decap_8 FILLER_19_1134 ();
 sg13g2_decap_4 FILLER_19_1141 ();
 sg13g2_fill_1 FILLER_19_1202 ();
 sg13g2_fill_2 FILLER_19_1208 ();
 sg13g2_decap_8 FILLER_19_1220 ();
 sg13g2_decap_4 FILLER_19_1227 ();
 sg13g2_fill_1 FILLER_19_1241 ();
 sg13g2_decap_8 FILLER_19_1281 ();
 sg13g2_decap_4 FILLER_19_1288 ();
 sg13g2_fill_1 FILLER_19_1305 ();
 sg13g2_fill_1 FILLER_19_1325 ();
 sg13g2_fill_2 FILLER_19_1330 ();
 sg13g2_decap_8 FILLER_19_1373 ();
 sg13g2_decap_8 FILLER_19_1380 ();
 sg13g2_decap_8 FILLER_19_1387 ();
 sg13g2_decap_8 FILLER_19_1394 ();
 sg13g2_decap_8 FILLER_19_1401 ();
 sg13g2_decap_8 FILLER_19_1408 ();
 sg13g2_decap_8 FILLER_19_1415 ();
 sg13g2_decap_8 FILLER_19_1422 ();
 sg13g2_decap_4 FILLER_19_1429 ();
 sg13g2_fill_1 FILLER_19_1433 ();
 sg13g2_decap_4 FILLER_19_1448 ();
 sg13g2_fill_2 FILLER_19_1452 ();
 sg13g2_decap_4 FILLER_19_1464 ();
 sg13g2_fill_1 FILLER_19_1489 ();
 sg13g2_decap_4 FILLER_19_1498 ();
 sg13g2_fill_2 FILLER_19_1527 ();
 sg13g2_fill_2 FILLER_19_1546 ();
 sg13g2_fill_1 FILLER_19_1548 ();
 sg13g2_fill_1 FILLER_19_1571 ();
 sg13g2_fill_1 FILLER_19_1577 ();
 sg13g2_fill_1 FILLER_19_1583 ();
 sg13g2_decap_8 FILLER_19_1589 ();
 sg13g2_fill_1 FILLER_19_1606 ();
 sg13g2_fill_2 FILLER_19_1616 ();
 sg13g2_fill_1 FILLER_19_1618 ();
 sg13g2_fill_2 FILLER_19_1706 ();
 sg13g2_fill_1 FILLER_19_1708 ();
 sg13g2_fill_2 FILLER_19_1730 ();
 sg13g2_fill_2 FILLER_19_1764 ();
 sg13g2_fill_2 FILLER_19_1773 ();
 sg13g2_fill_2 FILLER_19_1779 ();
 sg13g2_fill_1 FILLER_19_1781 ();
 sg13g2_fill_1 FILLER_19_1789 ();
 sg13g2_decap_4 FILLER_19_1806 ();
 sg13g2_fill_2 FILLER_19_1810 ();
 sg13g2_decap_8 FILLER_19_1872 ();
 sg13g2_fill_2 FILLER_19_1879 ();
 sg13g2_fill_2 FILLER_19_1890 ();
 sg13g2_fill_2 FILLER_19_1901 ();
 sg13g2_fill_2 FILLER_19_1922 ();
 sg13g2_fill_1 FILLER_19_1929 ();
 sg13g2_fill_2 FILLER_19_1949 ();
 sg13g2_decap_8 FILLER_19_1956 ();
 sg13g2_fill_1 FILLER_19_1963 ();
 sg13g2_fill_2 FILLER_19_1974 ();
 sg13g2_fill_1 FILLER_19_1990 ();
 sg13g2_decap_4 FILLER_19_2017 ();
 sg13g2_fill_2 FILLER_19_2021 ();
 sg13g2_decap_8 FILLER_19_2027 ();
 sg13g2_decap_4 FILLER_19_2034 ();
 sg13g2_decap_8 FILLER_19_2094 ();
 sg13g2_fill_2 FILLER_19_2101 ();
 sg13g2_fill_1 FILLER_19_2103 ();
 sg13g2_fill_2 FILLER_19_2112 ();
 sg13g2_decap_4 FILLER_19_2118 ();
 sg13g2_fill_2 FILLER_19_2158 ();
 sg13g2_fill_2 FILLER_19_2177 ();
 sg13g2_fill_2 FILLER_19_2256 ();
 sg13g2_decap_4 FILLER_19_2265 ();
 sg13g2_fill_2 FILLER_19_2269 ();
 sg13g2_decap_8 FILLER_19_2275 ();
 sg13g2_fill_2 FILLER_19_2282 ();
 sg13g2_decap_8 FILLER_19_2289 ();
 sg13g2_decap_4 FILLER_19_2296 ();
 sg13g2_fill_1 FILLER_19_2300 ();
 sg13g2_fill_1 FILLER_19_2359 ();
 sg13g2_decap_8 FILLER_19_2370 ();
 sg13g2_fill_2 FILLER_19_2384 ();
 sg13g2_fill_2 FILLER_19_2395 ();
 sg13g2_fill_2 FILLER_19_2436 ();
 sg13g2_fill_2 FILLER_19_2448 ();
 sg13g2_fill_1 FILLER_19_2460 ();
 sg13g2_decap_8 FILLER_19_2508 ();
 sg13g2_decap_8 FILLER_19_2515 ();
 sg13g2_fill_1 FILLER_19_2522 ();
 sg13g2_decap_8 FILLER_19_2532 ();
 sg13g2_decap_8 FILLER_19_2539 ();
 sg13g2_decap_8 FILLER_19_2620 ();
 sg13g2_decap_8 FILLER_19_2627 ();
 sg13g2_decap_8 FILLER_19_2634 ();
 sg13g2_decap_8 FILLER_19_2641 ();
 sg13g2_decap_8 FILLER_19_2648 ();
 sg13g2_decap_8 FILLER_19_2655 ();
 sg13g2_decap_8 FILLER_19_2662 ();
 sg13g2_fill_1 FILLER_19_2669 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_28 ();
 sg13g2_fill_1 FILLER_20_30 ();
 sg13g2_fill_2 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_fill_1 FILLER_20_70 ();
 sg13g2_decap_4 FILLER_20_115 ();
 sg13g2_fill_2 FILLER_20_119 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_189 ();
 sg13g2_fill_1 FILLER_20_202 ();
 sg13g2_fill_2 FILLER_20_238 ();
 sg13g2_decap_4 FILLER_20_303 ();
 sg13g2_decap_4 FILLER_20_312 ();
 sg13g2_fill_2 FILLER_20_316 ();
 sg13g2_fill_1 FILLER_20_322 ();
 sg13g2_decap_8 FILLER_20_331 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_344 ();
 sg13g2_fill_1 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_355 ();
 sg13g2_fill_2 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_366 ();
 sg13g2_decap_4 FILLER_20_404 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_fill_2 FILLER_20_442 ();
 sg13g2_decap_8 FILLER_20_478 ();
 sg13g2_fill_1 FILLER_20_485 ();
 sg13g2_fill_2 FILLER_20_491 ();
 sg13g2_decap_8 FILLER_20_498 ();
 sg13g2_decap_8 FILLER_20_505 ();
 sg13g2_decap_4 FILLER_20_516 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_fill_2 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_570 ();
 sg13g2_decap_8 FILLER_20_577 ();
 sg13g2_fill_2 FILLER_20_584 ();
 sg13g2_fill_1 FILLER_20_591 ();
 sg13g2_fill_2 FILLER_20_597 ();
 sg13g2_fill_2 FILLER_20_612 ();
 sg13g2_fill_1 FILLER_20_637 ();
 sg13g2_decap_8 FILLER_20_651 ();
 sg13g2_decap_8 FILLER_20_658 ();
 sg13g2_decap_8 FILLER_20_665 ();
 sg13g2_fill_1 FILLER_20_672 ();
 sg13g2_fill_1 FILLER_20_708 ();
 sg13g2_fill_2 FILLER_20_743 ();
 sg13g2_fill_2 FILLER_20_776 ();
 sg13g2_fill_1 FILLER_20_778 ();
 sg13g2_fill_2 FILLER_20_820 ();
 sg13g2_fill_1 FILLER_20_822 ();
 sg13g2_decap_8 FILLER_20_827 ();
 sg13g2_decap_8 FILLER_20_834 ();
 sg13g2_decap_8 FILLER_20_841 ();
 sg13g2_decap_4 FILLER_20_848 ();
 sg13g2_fill_2 FILLER_20_852 ();
 sg13g2_decap_8 FILLER_20_880 ();
 sg13g2_decap_8 FILLER_20_887 ();
 sg13g2_fill_2 FILLER_20_894 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_fill_1 FILLER_20_914 ();
 sg13g2_decap_4 FILLER_20_930 ();
 sg13g2_fill_2 FILLER_20_934 ();
 sg13g2_fill_2 FILLER_20_972 ();
 sg13g2_fill_1 FILLER_20_974 ();
 sg13g2_fill_2 FILLER_20_1001 ();
 sg13g2_fill_1 FILLER_20_1003 ();
 sg13g2_fill_2 FILLER_20_1030 ();
 sg13g2_fill_2 FILLER_20_1084 ();
 sg13g2_fill_2 FILLER_20_1095 ();
 sg13g2_fill_1 FILLER_20_1097 ();
 sg13g2_decap_8 FILLER_20_1106 ();
 sg13g2_fill_1 FILLER_20_1113 ();
 sg13g2_decap_4 FILLER_20_1127 ();
 sg13g2_fill_2 FILLER_20_1131 ();
 sg13g2_decap_4 FILLER_20_1143 ();
 sg13g2_fill_1 FILLER_20_1147 ();
 sg13g2_fill_2 FILLER_20_1178 ();
 sg13g2_fill_1 FILLER_20_1180 ();
 sg13g2_decap_8 FILLER_20_1195 ();
 sg13g2_decap_8 FILLER_20_1202 ();
 sg13g2_decap_4 FILLER_20_1209 ();
 sg13g2_fill_1 FILLER_20_1213 ();
 sg13g2_decap_8 FILLER_20_1250 ();
 sg13g2_decap_8 FILLER_20_1257 ();
 sg13g2_decap_4 FILLER_20_1264 ();
 sg13g2_decap_4 FILLER_20_1273 ();
 sg13g2_fill_1 FILLER_20_1277 ();
 sg13g2_fill_1 FILLER_20_1288 ();
 sg13g2_fill_2 FILLER_20_1303 ();
 sg13g2_decap_4 FILLER_20_1313 ();
 sg13g2_decap_8 FILLER_20_1321 ();
 sg13g2_decap_8 FILLER_20_1332 ();
 sg13g2_decap_4 FILLER_20_1343 ();
 sg13g2_fill_2 FILLER_20_1351 ();
 sg13g2_fill_1 FILLER_20_1353 ();
 sg13g2_decap_4 FILLER_20_1384 ();
 sg13g2_fill_1 FILLER_20_1388 ();
 sg13g2_decap_8 FILLER_20_1393 ();
 sg13g2_fill_1 FILLER_20_1400 ();
 sg13g2_decap_4 FILLER_20_1427 ();
 sg13g2_fill_2 FILLER_20_1431 ();
 sg13g2_decap_4 FILLER_20_1465 ();
 sg13g2_fill_2 FILLER_20_1469 ();
 sg13g2_fill_1 FILLER_20_1481 ();
 sg13g2_fill_1 FILLER_20_1490 ();
 sg13g2_decap_8 FILLER_20_1508 ();
 sg13g2_fill_2 FILLER_20_1523 ();
 sg13g2_fill_1 FILLER_20_1525 ();
 sg13g2_fill_2 FILLER_20_1531 ();
 sg13g2_decap_4 FILLER_20_1541 ();
 sg13g2_fill_2 FILLER_20_1545 ();
 sg13g2_fill_2 FILLER_20_1556 ();
 sg13g2_fill_1 FILLER_20_1558 ();
 sg13g2_decap_4 FILLER_20_1566 ();
 sg13g2_fill_1 FILLER_20_1570 ();
 sg13g2_fill_1 FILLER_20_1576 ();
 sg13g2_fill_2 FILLER_20_1636 ();
 sg13g2_decap_8 FILLER_20_1642 ();
 sg13g2_fill_1 FILLER_20_1649 ();
 sg13g2_fill_2 FILLER_20_1734 ();
 sg13g2_fill_1 FILLER_20_1749 ();
 sg13g2_fill_1 FILLER_20_1770 ();
 sg13g2_decap_8 FILLER_20_1807 ();
 sg13g2_decap_8 FILLER_20_1814 ();
 sg13g2_fill_2 FILLER_20_1821 ();
 sg13g2_fill_1 FILLER_20_1823 ();
 sg13g2_fill_1 FILLER_20_1828 ();
 sg13g2_fill_1 FILLER_20_1834 ();
 sg13g2_decap_4 FILLER_20_1882 ();
 sg13g2_decap_8 FILLER_20_1895 ();
 sg13g2_decap_4 FILLER_20_1902 ();
 sg13g2_fill_1 FILLER_20_1918 ();
 sg13g2_fill_2 FILLER_20_1924 ();
 sg13g2_fill_2 FILLER_20_1935 ();
 sg13g2_fill_2 FILLER_20_1951 ();
 sg13g2_decap_8 FILLER_20_1974 ();
 sg13g2_decap_8 FILLER_20_1981 ();
 sg13g2_decap_8 FILLER_20_1988 ();
 sg13g2_fill_1 FILLER_20_2005 ();
 sg13g2_decap_8 FILLER_20_2042 ();
 sg13g2_decap_8 FILLER_20_2049 ();
 sg13g2_fill_1 FILLER_20_2072 ();
 sg13g2_decap_8 FILLER_20_2109 ();
 sg13g2_decap_8 FILLER_20_2116 ();
 sg13g2_fill_2 FILLER_20_2123 ();
 sg13g2_fill_1 FILLER_20_2125 ();
 sg13g2_decap_4 FILLER_20_2134 ();
 sg13g2_fill_2 FILLER_20_2159 ();
 sg13g2_fill_1 FILLER_20_2161 ();
 sg13g2_fill_1 FILLER_20_2171 ();
 sg13g2_fill_2 FILLER_20_2219 ();
 sg13g2_decap_4 FILLER_20_2231 ();
 sg13g2_fill_2 FILLER_20_2235 ();
 sg13g2_fill_1 FILLER_20_2241 ();
 sg13g2_decap_8 FILLER_20_2263 ();
 sg13g2_decap_4 FILLER_20_2306 ();
 sg13g2_fill_1 FILLER_20_2320 ();
 sg13g2_fill_2 FILLER_20_2350 ();
 sg13g2_fill_2 FILLER_20_2355 ();
 sg13g2_fill_1 FILLER_20_2357 ();
 sg13g2_fill_1 FILLER_20_2402 ();
 sg13g2_fill_2 FILLER_20_2420 ();
 sg13g2_fill_1 FILLER_20_2457 ();
 sg13g2_fill_1 FILLER_20_2465 ();
 sg13g2_decap_4 FILLER_20_2511 ();
 sg13g2_decap_8 FILLER_20_2541 ();
 sg13g2_fill_1 FILLER_20_2548 ();
 sg13g2_decap_4 FILLER_20_2559 ();
 sg13g2_decap_8 FILLER_20_2629 ();
 sg13g2_decap_8 FILLER_20_2636 ();
 sg13g2_decap_8 FILLER_20_2643 ();
 sg13g2_decap_8 FILLER_20_2650 ();
 sg13g2_decap_8 FILLER_20_2657 ();
 sg13g2_decap_4 FILLER_20_2664 ();
 sg13g2_fill_2 FILLER_20_2668 ();
 sg13g2_fill_1 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_11 ();
 sg13g2_fill_1 FILLER_21_16 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_2 FILLER_21_98 ();
 sg13g2_fill_1 FILLER_21_108 ();
 sg13g2_decap_8 FILLER_21_114 ();
 sg13g2_decap_4 FILLER_21_121 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_decap_8 FILLER_21_152 ();
 sg13g2_fill_2 FILLER_21_159 ();
 sg13g2_fill_1 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_4 FILLER_21_189 ();
 sg13g2_fill_1 FILLER_21_193 ();
 sg13g2_fill_2 FILLER_21_254 ();
 sg13g2_decap_4 FILLER_21_260 ();
 sg13g2_fill_1 FILLER_21_269 ();
 sg13g2_decap_4 FILLER_21_278 ();
 sg13g2_fill_2 FILLER_21_297 ();
 sg13g2_fill_1 FILLER_21_299 ();
 sg13g2_decap_8 FILLER_21_305 ();
 sg13g2_decap_4 FILLER_21_322 ();
 sg13g2_fill_1 FILLER_21_326 ();
 sg13g2_fill_1 FILLER_21_331 ();
 sg13g2_fill_2 FILLER_21_336 ();
 sg13g2_fill_2 FILLER_21_343 ();
 sg13g2_fill_2 FILLER_21_349 ();
 sg13g2_fill_1 FILLER_21_351 ();
 sg13g2_decap_8 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_369 ();
 sg13g2_decap_8 FILLER_21_376 ();
 sg13g2_fill_1 FILLER_21_383 ();
 sg13g2_decap_4 FILLER_21_393 ();
 sg13g2_fill_2 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_433 ();
 sg13g2_fill_2 FILLER_21_437 ();
 sg13g2_fill_2 FILLER_21_449 ();
 sg13g2_decap_8 FILLER_21_477 ();
 sg13g2_fill_2 FILLER_21_484 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_fill_2 FILLER_21_497 ();
 sg13g2_fill_1 FILLER_21_507 ();
 sg13g2_fill_1 FILLER_21_512 ();
 sg13g2_fill_2 FILLER_21_521 ();
 sg13g2_fill_1 FILLER_21_555 ();
 sg13g2_decap_4 FILLER_21_561 ();
 sg13g2_fill_2 FILLER_21_565 ();
 sg13g2_decap_8 FILLER_21_573 ();
 sg13g2_fill_2 FILLER_21_580 ();
 sg13g2_fill_2 FILLER_21_586 ();
 sg13g2_fill_1 FILLER_21_588 ();
 sg13g2_fill_1 FILLER_21_602 ();
 sg13g2_fill_1 FILLER_21_608 ();
 sg13g2_decap_4 FILLER_21_624 ();
 sg13g2_fill_1 FILLER_21_628 ();
 sg13g2_decap_8 FILLER_21_670 ();
 sg13g2_fill_2 FILLER_21_677 ();
 sg13g2_fill_1 FILLER_21_683 ();
 sg13g2_fill_1 FILLER_21_692 ();
 sg13g2_fill_2 FILLER_21_726 ();
 sg13g2_fill_2 FILLER_21_757 ();
 sg13g2_decap_8 FILLER_21_835 ();
 sg13g2_fill_2 FILLER_21_842 ();
 sg13g2_fill_1 FILLER_21_844 ();
 sg13g2_decap_8 FILLER_21_931 ();
 sg13g2_decap_8 FILLER_21_938 ();
 sg13g2_fill_2 FILLER_21_945 ();
 sg13g2_fill_2 FILLER_21_956 ();
 sg13g2_fill_1 FILLER_21_958 ();
 sg13g2_fill_2 FILLER_21_979 ();
 sg13g2_decap_8 FILLER_21_985 ();
 sg13g2_fill_2 FILLER_21_992 ();
 sg13g2_fill_1 FILLER_21_994 ();
 sg13g2_fill_2 FILLER_21_1068 ();
 sg13g2_fill_1 FILLER_21_1070 ();
 sg13g2_fill_1 FILLER_21_1110 ();
 sg13g2_fill_2 FILLER_21_1115 ();
 sg13g2_decap_4 FILLER_21_1162 ();
 sg13g2_decap_4 FILLER_21_1170 ();
 sg13g2_decap_4 FILLER_21_1200 ();
 sg13g2_decap_8 FILLER_21_1208 ();
 sg13g2_fill_2 FILLER_21_1215 ();
 sg13g2_fill_2 FILLER_21_1235 ();
 sg13g2_decap_4 FILLER_21_1263 ();
 sg13g2_fill_2 FILLER_21_1267 ();
 sg13g2_decap_8 FILLER_21_1283 ();
 sg13g2_decap_8 FILLER_21_1290 ();
 sg13g2_decap_4 FILLER_21_1297 ();
 sg13g2_fill_2 FILLER_21_1301 ();
 sg13g2_decap_8 FILLER_21_1333 ();
 sg13g2_decap_8 FILLER_21_1340 ();
 sg13g2_decap_8 FILLER_21_1347 ();
 sg13g2_fill_2 FILLER_21_1354 ();
 sg13g2_fill_1 FILLER_21_1356 ();
 sg13g2_fill_2 FILLER_21_1367 ();
 sg13g2_fill_1 FILLER_21_1395 ();
 sg13g2_fill_2 FILLER_21_1411 ();
 sg13g2_fill_1 FILLER_21_1413 ();
 sg13g2_fill_2 FILLER_21_1423 ();
 sg13g2_fill_2 FILLER_21_1451 ();
 sg13g2_decap_4 FILLER_21_1458 ();
 sg13g2_fill_2 FILLER_21_1488 ();
 sg13g2_fill_1 FILLER_21_1490 ();
 sg13g2_decap_4 FILLER_21_1496 ();
 sg13g2_fill_1 FILLER_21_1500 ();
 sg13g2_decap_4 FILLER_21_1506 ();
 sg13g2_fill_2 FILLER_21_1510 ();
 sg13g2_decap_4 FILLER_21_1522 ();
 sg13g2_fill_2 FILLER_21_1526 ();
 sg13g2_fill_1 FILLER_21_1541 ();
 sg13g2_fill_2 FILLER_21_1561 ();
 sg13g2_fill_1 FILLER_21_1563 ();
 sg13g2_decap_4 FILLER_21_1579 ();
 sg13g2_fill_1 FILLER_21_1593 ();
 sg13g2_fill_2 FILLER_21_1605 ();
 sg13g2_fill_1 FILLER_21_1607 ();
 sg13g2_fill_1 FILLER_21_1621 ();
 sg13g2_decap_8 FILLER_21_1653 ();
 sg13g2_decap_8 FILLER_21_1660 ();
 sg13g2_fill_2 FILLER_21_1667 ();
 sg13g2_fill_2 FILLER_21_1683 ();
 sg13g2_fill_1 FILLER_21_1702 ();
 sg13g2_fill_1 FILLER_21_1707 ();
 sg13g2_decap_4 FILLER_21_1727 ();
 sg13g2_fill_1 FILLER_21_1731 ();
 sg13g2_fill_1 FILLER_21_1744 ();
 sg13g2_fill_1 FILLER_21_1785 ();
 sg13g2_fill_1 FILLER_21_1812 ();
 sg13g2_decap_8 FILLER_21_1818 ();
 sg13g2_decap_4 FILLER_21_1825 ();
 sg13g2_fill_1 FILLER_21_1829 ();
 sg13g2_fill_1 FILLER_21_1864 ();
 sg13g2_fill_1 FILLER_21_1870 ();
 sg13g2_decap_4 FILLER_21_1897 ();
 sg13g2_fill_1 FILLER_21_1901 ();
 sg13g2_fill_2 FILLER_21_1911 ();
 sg13g2_fill_1 FILLER_21_1913 ();
 sg13g2_fill_2 FILLER_21_1961 ();
 sg13g2_fill_1 FILLER_21_1963 ();
 sg13g2_decap_8 FILLER_21_1974 ();
 sg13g2_decap_8 FILLER_21_1981 ();
 sg13g2_decap_8 FILLER_21_1988 ();
 sg13g2_fill_2 FILLER_21_1995 ();
 sg13g2_fill_1 FILLER_21_2001 ();
 sg13g2_fill_1 FILLER_21_2048 ();
 sg13g2_fill_1 FILLER_21_2083 ();
 sg13g2_decap_8 FILLER_21_2109 ();
 sg13g2_decap_8 FILLER_21_2116 ();
 sg13g2_fill_2 FILLER_21_2123 ();
 sg13g2_fill_1 FILLER_21_2125 ();
 sg13g2_decap_8 FILLER_21_2130 ();
 sg13g2_decap_4 FILLER_21_2137 ();
 sg13g2_decap_4 FILLER_21_2151 ();
 sg13g2_fill_2 FILLER_21_2155 ();
 sg13g2_fill_1 FILLER_21_2174 ();
 sg13g2_fill_1 FILLER_21_2198 ();
 sg13g2_fill_2 FILLER_21_2212 ();
 sg13g2_decap_4 FILLER_21_2240 ();
 sg13g2_fill_2 FILLER_21_2244 ();
 sg13g2_decap_8 FILLER_21_2255 ();
 sg13g2_decap_8 FILLER_21_2262 ();
 sg13g2_fill_2 FILLER_21_2269 ();
 sg13g2_fill_1 FILLER_21_2271 ();
 sg13g2_decap_8 FILLER_21_2319 ();
 sg13g2_decap_8 FILLER_21_2330 ();
 sg13g2_decap_8 FILLER_21_2337 ();
 sg13g2_decap_4 FILLER_21_2344 ();
 sg13g2_fill_1 FILLER_21_2348 ();
 sg13g2_fill_1 FILLER_21_2390 ();
 sg13g2_fill_2 FILLER_21_2498 ();
 sg13g2_fill_1 FILLER_21_2500 ();
 sg13g2_decap_8 FILLER_21_2541 ();
 sg13g2_decap_8 FILLER_21_2548 ();
 sg13g2_decap_8 FILLER_21_2555 ();
 sg13g2_fill_2 FILLER_21_2562 ();
 sg13g2_fill_1 FILLER_21_2564 ();
 sg13g2_fill_2 FILLER_21_2592 ();
 sg13g2_fill_2 FILLER_21_2615 ();
 sg13g2_fill_1 FILLER_21_2617 ();
 sg13g2_decap_8 FILLER_21_2644 ();
 sg13g2_decap_8 FILLER_21_2651 ();
 sg13g2_decap_8 FILLER_21_2658 ();
 sg13g2_decap_4 FILLER_21_2665 ();
 sg13g2_fill_1 FILLER_21_2669 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_1 FILLER_22_2 ();
 sg13g2_decap_4 FILLER_22_7 ();
 sg13g2_fill_1 FILLER_22_25 ();
 sg13g2_fill_1 FILLER_22_86 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_4 FILLER_22_130 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_decap_4 FILLER_22_144 ();
 sg13g2_fill_2 FILLER_22_156 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_197 ();
 sg13g2_fill_1 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_223 ();
 sg13g2_decap_8 FILLER_22_275 ();
 sg13g2_decap_8 FILLER_22_282 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_fill_1 FILLER_22_291 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_fill_1 FILLER_22_332 ();
 sg13g2_fill_1 FILLER_22_337 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_fill_1 FILLER_22_375 ();
 sg13g2_fill_2 FILLER_22_390 ();
 sg13g2_fill_2 FILLER_22_452 ();
 sg13g2_fill_2 FILLER_22_459 ();
 sg13g2_fill_2 FILLER_22_491 ();
 sg13g2_fill_2 FILLER_22_503 ();
 sg13g2_fill_1 FILLER_22_505 ();
 sg13g2_fill_1 FILLER_22_559 ();
 sg13g2_fill_2 FILLER_22_590 ();
 sg13g2_fill_1 FILLER_22_592 ();
 sg13g2_fill_1 FILLER_22_603 ();
 sg13g2_fill_2 FILLER_22_618 ();
 sg13g2_fill_1 FILLER_22_620 ();
 sg13g2_fill_2 FILLER_22_625 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_fill_2 FILLER_22_648 ();
 sg13g2_fill_1 FILLER_22_650 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_fill_1 FILLER_22_736 ();
 sg13g2_fill_2 FILLER_22_778 ();
 sg13g2_fill_1 FILLER_22_780 ();
 sg13g2_fill_1 FILLER_22_815 ();
 sg13g2_fill_1 FILLER_22_837 ();
 sg13g2_fill_1 FILLER_22_868 ();
 sg13g2_fill_1 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_942 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_956 ();
 sg13g2_decap_8 FILLER_22_963 ();
 sg13g2_decap_8 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_fill_2 FILLER_22_991 ();
 sg13g2_fill_2 FILLER_22_1062 ();
 sg13g2_fill_1 FILLER_22_1064 ();
 sg13g2_decap_4 FILLER_22_1174 ();
 sg13g2_decap_4 FILLER_22_1218 ();
 sg13g2_fill_1 FILLER_22_1256 ();
 sg13g2_decap_4 FILLER_22_1261 ();
 sg13g2_fill_2 FILLER_22_1265 ();
 sg13g2_decap_4 FILLER_22_1272 ();
 sg13g2_fill_2 FILLER_22_1302 ();
 sg13g2_fill_1 FILLER_22_1309 ();
 sg13g2_fill_2 FILLER_22_1336 ();
 sg13g2_fill_2 FILLER_22_1364 ();
 sg13g2_fill_1 FILLER_22_1366 ();
 sg13g2_fill_2 FILLER_22_1371 ();
 sg13g2_fill_1 FILLER_22_1373 ();
 sg13g2_fill_2 FILLER_22_1378 ();
 sg13g2_fill_1 FILLER_22_1380 ();
 sg13g2_fill_2 FILLER_22_1391 ();
 sg13g2_fill_1 FILLER_22_1393 ();
 sg13g2_fill_2 FILLER_22_1412 ();
 sg13g2_decap_4 FILLER_22_1427 ();
 sg13g2_decap_8 FILLER_22_1457 ();
 sg13g2_fill_1 FILLER_22_1464 ();
 sg13g2_decap_4 FILLER_22_1481 ();
 sg13g2_fill_2 FILLER_22_1490 ();
 sg13g2_decap_8 FILLER_22_1500 ();
 sg13g2_fill_2 FILLER_22_1507 ();
 sg13g2_fill_1 FILLER_22_1509 ();
 sg13g2_fill_2 FILLER_22_1520 ();
 sg13g2_decap_8 FILLER_22_1527 ();
 sg13g2_fill_1 FILLER_22_1551 ();
 sg13g2_decap_8 FILLER_22_1571 ();
 sg13g2_decap_8 FILLER_22_1592 ();
 sg13g2_fill_2 FILLER_22_1616 ();
 sg13g2_fill_1 FILLER_22_1623 ();
 sg13g2_decap_4 FILLER_22_1632 ();
 sg13g2_fill_2 FILLER_22_1640 ();
 sg13g2_fill_2 FILLER_22_1692 ();
 sg13g2_fill_1 FILLER_22_1694 ();
 sg13g2_fill_2 FILLER_22_1717 ();
 sg13g2_fill_1 FILLER_22_1719 ();
 sg13g2_decap_8 FILLER_22_1726 ();
 sg13g2_decap_4 FILLER_22_1733 ();
 sg13g2_fill_2 FILLER_22_1780 ();
 sg13g2_fill_2 FILLER_22_1795 ();
 sg13g2_fill_1 FILLER_22_1797 ();
 sg13g2_fill_2 FILLER_22_1808 ();
 sg13g2_fill_1 FILLER_22_1810 ();
 sg13g2_fill_2 FILLER_22_1816 ();
 sg13g2_fill_1 FILLER_22_1818 ();
 sg13g2_fill_1 FILLER_22_1854 ();
 sg13g2_fill_2 FILLER_22_1884 ();
 sg13g2_fill_1 FILLER_22_1886 ();
 sg13g2_decap_8 FILLER_22_1892 ();
 sg13g2_decap_8 FILLER_22_1899 ();
 sg13g2_fill_1 FILLER_22_1906 ();
 sg13g2_fill_2 FILLER_22_1912 ();
 sg13g2_fill_1 FILLER_22_1941 ();
 sg13g2_fill_1 FILLER_22_1973 ();
 sg13g2_decap_4 FILLER_22_2000 ();
 sg13g2_fill_2 FILLER_22_2004 ();
 sg13g2_fill_1 FILLER_22_2010 ();
 sg13g2_fill_1 FILLER_22_2059 ();
 sg13g2_decap_8 FILLER_22_2064 ();
 sg13g2_fill_2 FILLER_22_2071 ();
 sg13g2_fill_1 FILLER_22_2073 ();
 sg13g2_fill_1 FILLER_22_2084 ();
 sg13g2_fill_1 FILLER_22_2110 ();
 sg13g2_decap_4 FILLER_22_2187 ();
 sg13g2_fill_1 FILLER_22_2191 ();
 sg13g2_decap_8 FILLER_22_2223 ();
 sg13g2_decap_8 FILLER_22_2230 ();
 sg13g2_decap_4 FILLER_22_2237 ();
 sg13g2_fill_1 FILLER_22_2241 ();
 sg13g2_decap_4 FILLER_22_2250 ();
 sg13g2_fill_1 FILLER_22_2254 ();
 sg13g2_fill_2 FILLER_22_2351 ();
 sg13g2_fill_2 FILLER_22_2383 ();
 sg13g2_fill_1 FILLER_22_2411 ();
 sg13g2_fill_2 FILLER_22_2429 ();
 sg13g2_fill_2 FILLER_22_2525 ();
 sg13g2_fill_1 FILLER_22_2527 ();
 sg13g2_fill_2 FILLER_22_2538 ();
 sg13g2_fill_1 FILLER_22_2540 ();
 sg13g2_decap_8 FILLER_22_2567 ();
 sg13g2_decap_4 FILLER_22_2574 ();
 sg13g2_fill_1 FILLER_22_2578 ();
 sg13g2_decap_8 FILLER_22_2605 ();
 sg13g2_decap_8 FILLER_22_2612 ();
 sg13g2_decap_4 FILLER_22_2619 ();
 sg13g2_fill_2 FILLER_22_2623 ();
 sg13g2_decap_8 FILLER_22_2629 ();
 sg13g2_decap_4 FILLER_22_2636 ();
 sg13g2_decap_8 FILLER_22_2644 ();
 sg13g2_decap_8 FILLER_22_2651 ();
 sg13g2_decap_8 FILLER_22_2658 ();
 sg13g2_decap_4 FILLER_22_2665 ();
 sg13g2_fill_1 FILLER_22_2669 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_2 ();
 sg13g2_fill_1 FILLER_23_29 ();
 sg13g2_fill_1 FILLER_23_61 ();
 sg13g2_fill_1 FILLER_23_87 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_decap_4 FILLER_23_181 ();
 sg13g2_fill_2 FILLER_23_190 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_fill_1 FILLER_23_243 ();
 sg13g2_fill_2 FILLER_23_342 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_358 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_fill_1 FILLER_23_365 ();
 sg13g2_fill_2 FILLER_23_371 ();
 sg13g2_fill_2 FILLER_23_378 ();
 sg13g2_fill_2 FILLER_23_406 ();
 sg13g2_fill_2 FILLER_23_426 ();
 sg13g2_fill_1 FILLER_23_468 ();
 sg13g2_fill_1 FILLER_23_526 ();
 sg13g2_fill_1 FILLER_23_531 ();
 sg13g2_decap_8 FILLER_23_596 ();
 sg13g2_decap_8 FILLER_23_603 ();
 sg13g2_fill_1 FILLER_23_610 ();
 sg13g2_decap_4 FILLER_23_637 ();
 sg13g2_decap_4 FILLER_23_647 ();
 sg13g2_fill_1 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_656 ();
 sg13g2_decap_8 FILLER_23_663 ();
 sg13g2_fill_1 FILLER_23_670 ();
 sg13g2_fill_2 FILLER_23_718 ();
 sg13g2_fill_2 FILLER_23_724 ();
 sg13g2_decap_8 FILLER_23_778 ();
 sg13g2_decap_8 FILLER_23_785 ();
 sg13g2_decap_8 FILLER_23_792 ();
 sg13g2_fill_2 FILLER_23_799 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_4 FILLER_23_812 ();
 sg13g2_fill_2 FILLER_23_816 ();
 sg13g2_fill_2 FILLER_23_875 ();
 sg13g2_fill_2 FILLER_23_881 ();
 sg13g2_fill_1 FILLER_23_883 ();
 sg13g2_decap_8 FILLER_23_935 ();
 sg13g2_decap_4 FILLER_23_942 ();
 sg13g2_fill_1 FILLER_23_946 ();
 sg13g2_fill_2 FILLER_23_973 ();
 sg13g2_fill_1 FILLER_23_975 ();
 sg13g2_fill_2 FILLER_23_981 ();
 sg13g2_fill_2 FILLER_23_996 ();
 sg13g2_fill_1 FILLER_23_1039 ();
 sg13g2_fill_2 FILLER_23_1049 ();
 sg13g2_decap_4 FILLER_23_1121 ();
 sg13g2_fill_1 FILLER_23_1125 ();
 sg13g2_fill_2 FILLER_23_1130 ();
 sg13g2_fill_2 FILLER_23_1142 ();
 sg13g2_fill_1 FILLER_23_1144 ();
 sg13g2_fill_1 FILLER_23_1171 ();
 sg13g2_decap_8 FILLER_23_1182 ();
 sg13g2_fill_1 FILLER_23_1189 ();
 sg13g2_fill_2 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1289 ();
 sg13g2_decap_4 FILLER_23_1296 ();
 sg13g2_decap_4 FILLER_23_1304 ();
 sg13g2_decap_4 FILLER_23_1313 ();
 sg13g2_fill_1 FILLER_23_1317 ();
 sg13g2_decap_4 FILLER_23_1322 ();
 sg13g2_fill_1 FILLER_23_1334 ();
 sg13g2_fill_2 FILLER_23_1345 ();
 sg13g2_decap_4 FILLER_23_1377 ();
 sg13g2_fill_2 FILLER_23_1385 ();
 sg13g2_fill_1 FILLER_23_1387 ();
 sg13g2_fill_1 FILLER_23_1417 ();
 sg13g2_fill_1 FILLER_23_1448 ();
 sg13g2_fill_1 FILLER_23_1469 ();
 sg13g2_decap_8 FILLER_23_1495 ();
 sg13g2_fill_2 FILLER_23_1502 ();
 sg13g2_fill_1 FILLER_23_1504 ();
 sg13g2_decap_8 FILLER_23_1515 ();
 sg13g2_decap_8 FILLER_23_1522 ();
 sg13g2_fill_2 FILLER_23_1529 ();
 sg13g2_fill_1 FILLER_23_1531 ();
 sg13g2_decap_8 FILLER_23_1538 ();
 sg13g2_fill_2 FILLER_23_1545 ();
 sg13g2_fill_1 FILLER_23_1559 ();
 sg13g2_fill_1 FILLER_23_1569 ();
 sg13g2_fill_2 FILLER_23_1581 ();
 sg13g2_fill_1 FILLER_23_1583 ();
 sg13g2_fill_1 FILLER_23_1590 ();
 sg13g2_fill_2 FILLER_23_1656 ();
 sg13g2_fill_1 FILLER_23_1677 ();
 sg13g2_fill_2 FILLER_23_1683 ();
 sg13g2_fill_1 FILLER_23_1729 ();
 sg13g2_fill_2 FILLER_23_1737 ();
 sg13g2_fill_1 FILLER_23_1739 ();
 sg13g2_decap_8 FILLER_23_1766 ();
 sg13g2_decap_8 FILLER_23_1773 ();
 sg13g2_decap_4 FILLER_23_1780 ();
 sg13g2_fill_1 FILLER_23_1784 ();
 sg13g2_fill_2 FILLER_23_1790 ();
 sg13g2_fill_1 FILLER_23_1792 ();
 sg13g2_fill_2 FILLER_23_1797 ();
 sg13g2_decap_8 FILLER_23_1815 ();
 sg13g2_fill_1 FILLER_23_1822 ();
 sg13g2_fill_2 FILLER_23_1857 ();
 sg13g2_decap_8 FILLER_23_1897 ();
 sg13g2_fill_2 FILLER_23_1959 ();
 sg13g2_decap_8 FILLER_23_1971 ();
 sg13g2_fill_2 FILLER_23_1978 ();
 sg13g2_decap_4 FILLER_23_1984 ();
 sg13g2_fill_1 FILLER_23_1988 ();
 sg13g2_fill_1 FILLER_23_2076 ();
 sg13g2_decap_4 FILLER_23_2107 ();
 sg13g2_fill_1 FILLER_23_2111 ();
 sg13g2_fill_1 FILLER_23_2138 ();
 sg13g2_fill_2 FILLER_23_2149 ();
 sg13g2_decap_4 FILLER_23_2177 ();
 sg13g2_decap_8 FILLER_23_2220 ();
 sg13g2_fill_2 FILLER_23_2227 ();
 sg13g2_fill_1 FILLER_23_2285 ();
 sg13g2_fill_1 FILLER_23_2358 ();
 sg13g2_fill_1 FILLER_23_2402 ();
 sg13g2_fill_1 FILLER_23_2433 ();
 sg13g2_fill_1 FILLER_23_2455 ();
 sg13g2_fill_1 FILLER_23_2481 ();
 sg13g2_decap_4 FILLER_23_2492 ();
 sg13g2_fill_1 FILLER_23_2496 ();
 sg13g2_fill_1 FILLER_23_2523 ();
 sg13g2_decap_4 FILLER_23_2538 ();
 sg13g2_fill_2 FILLER_23_2542 ();
 sg13g2_decap_8 FILLER_23_2570 ();
 sg13g2_decap_4 FILLER_23_2577 ();
 sg13g2_fill_1 FILLER_23_2581 ();
 sg13g2_decap_4 FILLER_23_2603 ();
 sg13g2_fill_1 FILLER_23_2607 ();
 sg13g2_decap_8 FILLER_23_2628 ();
 sg13g2_fill_1 FILLER_23_2635 ();
 sg13g2_decap_8 FILLER_23_2662 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_fill_2 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_13 ();
 sg13g2_decap_8 FILLER_24_20 ();
 sg13g2_decap_8 FILLER_24_27 ();
 sg13g2_fill_2 FILLER_24_34 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_2 FILLER_24_60 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_114 ();
 sg13g2_decap_4 FILLER_24_134 ();
 sg13g2_decap_4 FILLER_24_167 ();
 sg13g2_fill_1 FILLER_24_171 ();
 sg13g2_fill_2 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_209 ();
 sg13g2_fill_1 FILLER_24_215 ();
 sg13g2_fill_1 FILLER_24_224 ();
 sg13g2_fill_2 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_253 ();
 sg13g2_fill_1 FILLER_24_288 ();
 sg13g2_fill_1 FILLER_24_293 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_1 FILLER_24_304 ();
 sg13g2_fill_1 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_364 ();
 sg13g2_fill_1 FILLER_24_366 ();
 sg13g2_fill_1 FILLER_24_474 ();
 sg13g2_fill_1 FILLER_24_479 ();
 sg13g2_fill_1 FILLER_24_490 ();
 sg13g2_fill_2 FILLER_24_505 ();
 sg13g2_fill_1 FILLER_24_511 ();
 sg13g2_fill_1 FILLER_24_517 ();
 sg13g2_fill_2 FILLER_24_523 ();
 sg13g2_fill_1 FILLER_24_525 ();
 sg13g2_fill_2 FILLER_24_537 ();
 sg13g2_fill_1 FILLER_24_539 ();
 sg13g2_fill_2 FILLER_24_544 ();
 sg13g2_fill_1 FILLER_24_552 ();
 sg13g2_fill_2 FILLER_24_558 ();
 sg13g2_fill_2 FILLER_24_611 ();
 sg13g2_fill_1 FILLER_24_616 ();
 sg13g2_fill_2 FILLER_24_621 ();
 sg13g2_fill_1 FILLER_24_623 ();
 sg13g2_decap_8 FILLER_24_629 ();
 sg13g2_decap_4 FILLER_24_636 ();
 sg13g2_decap_4 FILLER_24_646 ();
 sg13g2_fill_2 FILLER_24_650 ();
 sg13g2_fill_2 FILLER_24_709 ();
 sg13g2_fill_2 FILLER_24_714 ();
 sg13g2_fill_1 FILLER_24_736 ();
 sg13g2_decap_8 FILLER_24_787 ();
 sg13g2_decap_8 FILLER_24_794 ();
 sg13g2_decap_8 FILLER_24_801 ();
 sg13g2_fill_2 FILLER_24_808 ();
 sg13g2_decap_8 FILLER_24_820 ();
 sg13g2_decap_8 FILLER_24_827 ();
 sg13g2_fill_2 FILLER_24_834 ();
 sg13g2_fill_2 FILLER_24_840 ();
 sg13g2_decap_4 FILLER_24_852 ();
 sg13g2_decap_4 FILLER_24_877 ();
 sg13g2_decap_4 FILLER_24_891 ();
 sg13g2_fill_2 FILLER_24_905 ();
 sg13g2_fill_1 FILLER_24_907 ();
 sg13g2_decap_4 FILLER_24_931 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_fill_1 FILLER_24_956 ();
 sg13g2_fill_2 FILLER_24_1009 ();
 sg13g2_decap_4 FILLER_24_1020 ();
 sg13g2_fill_1 FILLER_24_1024 ();
 sg13g2_fill_2 FILLER_24_1056 ();
 sg13g2_fill_1 FILLER_24_1058 ();
 sg13g2_fill_1 FILLER_24_1063 ();
 sg13g2_fill_2 FILLER_24_1085 ();
 sg13g2_decap_4 FILLER_24_1096 ();
 sg13g2_fill_2 FILLER_24_1100 ();
 sg13g2_fill_2 FILLER_24_1106 ();
 sg13g2_decap_8 FILLER_24_1120 ();
 sg13g2_decap_4 FILLER_24_1127 ();
 sg13g2_fill_1 FILLER_24_1131 ();
 sg13g2_fill_1 FILLER_24_1140 ();
 sg13g2_fill_2 FILLER_24_1151 ();
 sg13g2_fill_1 FILLER_24_1153 ();
 sg13g2_fill_2 FILLER_24_1196 ();
 sg13g2_fill_1 FILLER_24_1198 ();
 sg13g2_fill_1 FILLER_24_1225 ();
 sg13g2_fill_2 FILLER_24_1230 ();
 sg13g2_fill_2 FILLER_24_1263 ();
 sg13g2_fill_1 FILLER_24_1265 ();
 sg13g2_fill_2 FILLER_24_1301 ();
 sg13g2_decap_8 FILLER_24_1329 ();
 sg13g2_decap_4 FILLER_24_1336 ();
 sg13g2_fill_1 FILLER_24_1350 ();
 sg13g2_decap_4 FILLER_24_1365 ();
 sg13g2_fill_2 FILLER_24_1379 ();
 sg13g2_fill_1 FILLER_24_1381 ();
 sg13g2_decap_8 FILLER_24_1385 ();
 sg13g2_fill_1 FILLER_24_1420 ();
 sg13g2_decap_8 FILLER_24_1427 ();
 sg13g2_fill_2 FILLER_24_1434 ();
 sg13g2_fill_1 FILLER_24_1436 ();
 sg13g2_decap_4 FILLER_24_1446 ();
 sg13g2_fill_2 FILLER_24_1450 ();
 sg13g2_fill_1 FILLER_24_1471 ();
 sg13g2_fill_2 FILLER_24_1485 ();
 sg13g2_fill_1 FILLER_24_1487 ();
 sg13g2_fill_2 FILLER_24_1493 ();
 sg13g2_fill_1 FILLER_24_1511 ();
 sg13g2_decap_8 FILLER_24_1517 ();
 sg13g2_decap_4 FILLER_24_1524 ();
 sg13g2_fill_2 FILLER_24_1543 ();
 sg13g2_fill_1 FILLER_24_1545 ();
 sg13g2_decap_8 FILLER_24_1555 ();
 sg13g2_decap_8 FILLER_24_1573 ();
 sg13g2_fill_1 FILLER_24_1580 ();
 sg13g2_decap_4 FILLER_24_1594 ();
 sg13g2_decap_8 FILLER_24_1608 ();
 sg13g2_fill_1 FILLER_24_1615 ();
 sg13g2_decap_4 FILLER_24_1621 ();
 sg13g2_fill_1 FILLER_24_1625 ();
 sg13g2_decap_8 FILLER_24_1645 ();
 sg13g2_decap_8 FILLER_24_1652 ();
 sg13g2_fill_2 FILLER_24_1662 ();
 sg13g2_decap_4 FILLER_24_1684 ();
 sg13g2_fill_1 FILLER_24_1688 ();
 sg13g2_decap_8 FILLER_24_1728 ();
 sg13g2_fill_2 FILLER_24_1735 ();
 sg13g2_fill_1 FILLER_24_1737 ();
 sg13g2_fill_2 FILLER_24_1742 ();
 sg13g2_fill_1 FILLER_24_1744 ();
 sg13g2_fill_1 FILLER_24_1750 ();
 sg13g2_fill_1 FILLER_24_1756 ();
 sg13g2_fill_1 FILLER_24_1762 ();
 sg13g2_fill_2 FILLER_24_1788 ();
 sg13g2_fill_2 FILLER_24_1794 ();
 sg13g2_fill_1 FILLER_24_1796 ();
 sg13g2_decap_4 FILLER_24_1827 ();
 sg13g2_fill_2 FILLER_24_1855 ();
 sg13g2_decap_8 FILLER_24_1883 ();
 sg13g2_fill_2 FILLER_24_1890 ();
 sg13g2_decap_4 FILLER_24_1897 ();
 sg13g2_fill_1 FILLER_24_1901 ();
 sg13g2_decap_4 FILLER_24_1909 ();
 sg13g2_fill_2 FILLER_24_1913 ();
 sg13g2_fill_1 FILLER_24_1953 ();
 sg13g2_decap_8 FILLER_24_1958 ();
 sg13g2_decap_8 FILLER_24_1965 ();
 sg13g2_decap_8 FILLER_24_1972 ();
 sg13g2_decap_8 FILLER_24_1979 ();
 sg13g2_decap_8 FILLER_24_1996 ();
 sg13g2_decap_4 FILLER_24_2003 ();
 sg13g2_fill_2 FILLER_24_2007 ();
 sg13g2_fill_1 FILLER_24_2035 ();
 sg13g2_fill_1 FILLER_24_2049 ();
 sg13g2_fill_2 FILLER_24_2076 ();
 sg13g2_fill_1 FILLER_24_2082 ();
 sg13g2_fill_2 FILLER_24_2091 ();
 sg13g2_fill_1 FILLER_24_2103 ();
 sg13g2_fill_2 FILLER_24_2138 ();
 sg13g2_decap_4 FILLER_24_2164 ();
 sg13g2_fill_2 FILLER_24_2168 ();
 sg13g2_decap_8 FILLER_24_2200 ();
 sg13g2_fill_2 FILLER_24_2207 ();
 sg13g2_fill_1 FILLER_24_2209 ();
 sg13g2_decap_8 FILLER_24_2214 ();
 sg13g2_decap_8 FILLER_24_2221 ();
 sg13g2_decap_4 FILLER_24_2228 ();
 sg13g2_fill_2 FILLER_24_2232 ();
 sg13g2_decap_8 FILLER_24_2326 ();
 sg13g2_decap_8 FILLER_24_2333 ();
 sg13g2_decap_8 FILLER_24_2340 ();
 sg13g2_fill_2 FILLER_24_2463 ();
 sg13g2_decap_8 FILLER_24_2470 ();
 sg13g2_fill_2 FILLER_24_2477 ();
 sg13g2_decap_4 FILLER_24_2483 ();
 sg13g2_decap_8 FILLER_24_2491 ();
 sg13g2_decap_4 FILLER_24_2498 ();
 sg13g2_fill_1 FILLER_24_2502 ();
 sg13g2_decap_8 FILLER_24_2507 ();
 sg13g2_decap_8 FILLER_24_2514 ();
 sg13g2_decap_4 FILLER_24_2521 ();
 sg13g2_fill_1 FILLER_24_2525 ();
 sg13g2_decap_8 FILLER_24_2597 ();
 sg13g2_fill_2 FILLER_24_2604 ();
 sg13g2_fill_1 FILLER_24_2616 ();
 sg13g2_decap_8 FILLER_24_2647 ();
 sg13g2_decap_8 FILLER_24_2654 ();
 sg13g2_decap_8 FILLER_24_2661 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_28 ();
 sg13g2_fill_1 FILLER_25_30 ();
 sg13g2_fill_1 FILLER_25_36 ();
 sg13g2_fill_1 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_60 ();
 sg13g2_fill_1 FILLER_25_72 ();
 sg13g2_fill_1 FILLER_25_81 ();
 sg13g2_fill_2 FILLER_25_87 ();
 sg13g2_fill_2 FILLER_25_93 ();
 sg13g2_fill_2 FILLER_25_105 ();
 sg13g2_decap_4 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_151 ();
 sg13g2_fill_1 FILLER_25_171 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_200 ();
 sg13g2_fill_2 FILLER_25_235 ();
 sg13g2_fill_1 FILLER_25_246 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_312 ();
 sg13g2_fill_1 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_fill_2 FILLER_25_424 ();
 sg13g2_fill_1 FILLER_25_431 ();
 sg13g2_fill_1 FILLER_25_456 ();
 sg13g2_fill_2 FILLER_25_477 ();
 sg13g2_fill_1 FILLER_25_493 ();
 sg13g2_decap_8 FILLER_25_524 ();
 sg13g2_fill_2 FILLER_25_531 ();
 sg13g2_fill_1 FILLER_25_533 ();
 sg13g2_decap_4 FILLER_25_539 ();
 sg13g2_fill_2 FILLER_25_561 ();
 sg13g2_fill_1 FILLER_25_563 ();
 sg13g2_fill_1 FILLER_25_568 ();
 sg13g2_decap_4 FILLER_25_631 ();
 sg13g2_fill_2 FILLER_25_697 ();
 sg13g2_fill_2 FILLER_25_737 ();
 sg13g2_fill_1 FILLER_25_743 ();
 sg13g2_fill_2 FILLER_25_769 ();
 sg13g2_fill_1 FILLER_25_780 ();
 sg13g2_fill_2 FILLER_25_791 ();
 sg13g2_fill_1 FILLER_25_793 ();
 sg13g2_fill_1 FILLER_25_820 ();
 sg13g2_decap_8 FILLER_25_842 ();
 sg13g2_decap_8 FILLER_25_849 ();
 sg13g2_decap_8 FILLER_25_856 ();
 sg13g2_fill_1 FILLER_25_873 ();
 sg13g2_fill_1 FILLER_25_910 ();
 sg13g2_fill_1 FILLER_25_951 ();
 sg13g2_fill_2 FILLER_25_1015 ();
 sg13g2_fill_2 FILLER_25_1038 ();
 sg13g2_decap_4 FILLER_25_1048 ();
 sg13g2_fill_1 FILLER_25_1052 ();
 sg13g2_fill_2 FILLER_25_1082 ();
 sg13g2_fill_1 FILLER_25_1084 ();
 sg13g2_decap_4 FILLER_25_1116 ();
 sg13g2_fill_1 FILLER_25_1120 ();
 sg13g2_decap_8 FILLER_25_1129 ();
 sg13g2_decap_8 FILLER_25_1140 ();
 sg13g2_fill_2 FILLER_25_1147 ();
 sg13g2_fill_1 FILLER_25_1149 ();
 sg13g2_fill_1 FILLER_25_1154 ();
 sg13g2_fill_1 FILLER_25_1165 ();
 sg13g2_decap_8 FILLER_25_1170 ();
 sg13g2_fill_1 FILLER_25_1203 ();
 sg13g2_decap_8 FILLER_25_1208 ();
 sg13g2_decap_8 FILLER_25_1215 ();
 sg13g2_decap_8 FILLER_25_1222 ();
 sg13g2_fill_2 FILLER_25_1229 ();
 sg13g2_fill_1 FILLER_25_1231 ();
 sg13g2_fill_1 FILLER_25_1237 ();
 sg13g2_fill_1 FILLER_25_1269 ();
 sg13g2_decap_4 FILLER_25_1275 ();
 sg13g2_fill_1 FILLER_25_1279 ();
 sg13g2_decap_4 FILLER_25_1284 ();
 sg13g2_fill_2 FILLER_25_1288 ();
 sg13g2_decap_8 FILLER_25_1294 ();
 sg13g2_decap_8 FILLER_25_1301 ();
 sg13g2_decap_4 FILLER_25_1308 ();
 sg13g2_decap_8 FILLER_25_1316 ();
 sg13g2_fill_2 FILLER_25_1357 ();
 sg13g2_fill_2 FILLER_25_1389 ();
 sg13g2_fill_2 FILLER_25_1424 ();
 sg13g2_decap_8 FILLER_25_1456 ();
 sg13g2_decap_4 FILLER_25_1463 ();
 sg13g2_fill_1 FILLER_25_1467 ();
 sg13g2_decap_4 FILLER_25_1480 ();
 sg13g2_fill_1 FILLER_25_1484 ();
 sg13g2_fill_2 FILLER_25_1490 ();
 sg13g2_fill_1 FILLER_25_1492 ();
 sg13g2_decap_8 FILLER_25_1500 ();
 sg13g2_fill_1 FILLER_25_1507 ();
 sg13g2_decap_4 FILLER_25_1528 ();
 sg13g2_fill_2 FILLER_25_1537 ();
 sg13g2_fill_1 FILLER_25_1539 ();
 sg13g2_decap_4 FILLER_25_1556 ();
 sg13g2_fill_2 FILLER_25_1560 ();
 sg13g2_fill_1 FILLER_25_1584 ();
 sg13g2_fill_2 FILLER_25_1590 ();
 sg13g2_fill_1 FILLER_25_1592 ();
 sg13g2_decap_4 FILLER_25_1608 ();
 sg13g2_decap_8 FILLER_25_1616 ();
 sg13g2_decap_8 FILLER_25_1623 ();
 sg13g2_decap_4 FILLER_25_1630 ();
 sg13g2_decap_8 FILLER_25_1647 ();
 sg13g2_fill_2 FILLER_25_1654 ();
 sg13g2_fill_2 FILLER_25_1698 ();
 sg13g2_fill_1 FILLER_25_1713 ();
 sg13g2_decap_4 FILLER_25_1740 ();
 sg13g2_fill_2 FILLER_25_1744 ();
 sg13g2_fill_1 FILLER_25_1756 ();
 sg13g2_fill_2 FILLER_25_1797 ();
 sg13g2_decap_8 FILLER_25_1819 ();
 sg13g2_decap_8 FILLER_25_1877 ();
 sg13g2_fill_1 FILLER_25_1884 ();
 sg13g2_fill_1 FILLER_25_1900 ();
 sg13g2_fill_1 FILLER_25_1906 ();
 sg13g2_fill_2 FILLER_25_1929 ();
 sg13g2_decap_8 FILLER_25_1957 ();
 sg13g2_decap_4 FILLER_25_1964 ();
 sg13g2_fill_2 FILLER_25_1968 ();
 sg13g2_decap_8 FILLER_25_2022 ();
 sg13g2_fill_1 FILLER_25_2029 ();
 sg13g2_fill_2 FILLER_25_2060 ();
 sg13g2_fill_1 FILLER_25_2062 ();
 sg13g2_fill_2 FILLER_25_2073 ();
 sg13g2_fill_1 FILLER_25_2075 ();
 sg13g2_decap_4 FILLER_25_2102 ();
 sg13g2_fill_1 FILLER_25_2106 ();
 sg13g2_fill_2 FILLER_25_2132 ();
 sg13g2_decap_4 FILLER_25_2142 ();
 sg13g2_fill_2 FILLER_25_2146 ();
 sg13g2_decap_8 FILLER_25_2157 ();
 sg13g2_fill_1 FILLER_25_2168 ();
 sg13g2_decap_8 FILLER_25_2183 ();
 sg13g2_fill_2 FILLER_25_2190 ();
 sg13g2_fill_1 FILLER_25_2192 ();
 sg13g2_fill_2 FILLER_25_2229 ();
 sg13g2_decap_4 FILLER_25_2252 ();
 sg13g2_fill_2 FILLER_25_2256 ();
 sg13g2_decap_8 FILLER_25_2341 ();
 sg13g2_decap_4 FILLER_25_2348 ();
 sg13g2_fill_2 FILLER_25_2352 ();
 sg13g2_decap_4 FILLER_25_2358 ();
 sg13g2_fill_1 FILLER_25_2362 ();
 sg13g2_fill_2 FILLER_25_2434 ();
 sg13g2_fill_1 FILLER_25_2459 ();
 sg13g2_decap_8 FILLER_25_2506 ();
 sg13g2_decap_8 FILLER_25_2513 ();
 sg13g2_decap_8 FILLER_25_2526 ();
 sg13g2_decap_8 FILLER_25_2533 ();
 sg13g2_decap_4 FILLER_25_2540 ();
 sg13g2_fill_1 FILLER_25_2544 ();
 sg13g2_decap_4 FILLER_25_2553 ();
 sg13g2_fill_2 FILLER_25_2557 ();
 sg13g2_decap_4 FILLER_25_2611 ();
 sg13g2_fill_2 FILLER_25_2615 ();
 sg13g2_decap_8 FILLER_25_2643 ();
 sg13g2_decap_8 FILLER_25_2650 ();
 sg13g2_decap_8 FILLER_25_2657 ();
 sg13g2_decap_4 FILLER_25_2664 ();
 sg13g2_fill_2 FILLER_25_2668 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_33 ();
 sg13g2_fill_2 FILLER_26_81 ();
 sg13g2_fill_2 FILLER_26_107 ();
 sg13g2_fill_2 FILLER_26_113 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_129 ();
 sg13g2_fill_2 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_154 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_fill_2 FILLER_26_229 ();
 sg13g2_fill_2 FILLER_26_252 ();
 sg13g2_fill_1 FILLER_26_254 ();
 sg13g2_decap_4 FILLER_26_260 ();
 sg13g2_fill_2 FILLER_26_286 ();
 sg13g2_fill_1 FILLER_26_288 ();
 sg13g2_fill_1 FILLER_26_299 ();
 sg13g2_decap_8 FILLER_26_309 ();
 sg13g2_decap_8 FILLER_26_316 ();
 sg13g2_decap_4 FILLER_26_323 ();
 sg13g2_decap_4 FILLER_26_336 ();
 sg13g2_fill_2 FILLER_26_340 ();
 sg13g2_decap_4 FILLER_26_347 ();
 sg13g2_fill_1 FILLER_26_351 ();
 sg13g2_decap_8 FILLER_26_360 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_369 ();
 sg13g2_fill_2 FILLER_26_380 ();
 sg13g2_decap_4 FILLER_26_388 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_fill_1 FILLER_26_414 ();
 sg13g2_fill_1 FILLER_26_427 ();
 sg13g2_fill_1 FILLER_26_499 ();
 sg13g2_decap_8 FILLER_26_505 ();
 sg13g2_decap_8 FILLER_26_512 ();
 sg13g2_decap_4 FILLER_26_519 ();
 sg13g2_fill_2 FILLER_26_523 ();
 sg13g2_fill_1 FILLER_26_534 ();
 sg13g2_decap_8 FILLER_26_561 ();
 sg13g2_decap_4 FILLER_26_568 ();
 sg13g2_fill_1 FILLER_26_572 ();
 sg13g2_fill_1 FILLER_26_577 ();
 sg13g2_fill_1 FILLER_26_582 ();
 sg13g2_fill_2 FILLER_26_587 ();
 sg13g2_fill_2 FILLER_26_594 ();
 sg13g2_fill_2 FILLER_26_600 ();
 sg13g2_fill_1 FILLER_26_606 ();
 sg13g2_fill_2 FILLER_26_612 ();
 sg13g2_fill_1 FILLER_26_614 ();
 sg13g2_fill_2 FILLER_26_624 ();
 sg13g2_fill_1 FILLER_26_626 ();
 sg13g2_fill_1 FILLER_26_657 ();
 sg13g2_fill_1 FILLER_26_668 ();
 sg13g2_fill_1 FILLER_26_695 ();
 sg13g2_fill_1 FILLER_26_706 ();
 sg13g2_fill_1 FILLER_26_711 ();
 sg13g2_fill_2 FILLER_26_750 ();
 sg13g2_fill_1 FILLER_26_793 ();
 sg13g2_fill_2 FILLER_26_871 ();
 sg13g2_fill_1 FILLER_26_873 ();
 sg13g2_fill_2 FILLER_26_900 ();
 sg13g2_fill_2 FILLER_26_928 ();
 sg13g2_decap_4 FILLER_26_934 ();
 sg13g2_decap_8 FILLER_26_974 ();
 sg13g2_fill_2 FILLER_26_981 ();
 sg13g2_fill_1 FILLER_26_988 ();
 sg13g2_fill_1 FILLER_26_994 ();
 sg13g2_fill_2 FILLER_26_1033 ();
 sg13g2_decap_8 FILLER_26_1039 ();
 sg13g2_fill_2 FILLER_26_1046 ();
 sg13g2_fill_1 FILLER_26_1053 ();
 sg13g2_fill_2 FILLER_26_1080 ();
 sg13g2_fill_1 FILLER_26_1082 ();
 sg13g2_fill_1 FILLER_26_1109 ();
 sg13g2_fill_2 FILLER_26_1136 ();
 sg13g2_decap_8 FILLER_26_1150 ();
 sg13g2_decap_8 FILLER_26_1157 ();
 sg13g2_fill_1 FILLER_26_1164 ();
 sg13g2_decap_8 FILLER_26_1182 ();
 sg13g2_fill_2 FILLER_26_1189 ();
 sg13g2_decap_4 FILLER_26_1209 ();
 sg13g2_fill_1 FILLER_26_1213 ();
 sg13g2_decap_4 FILLER_26_1254 ();
 sg13g2_fill_2 FILLER_26_1258 ();
 sg13g2_fill_2 FILLER_26_1270 ();
 sg13g2_decap_4 FILLER_26_1298 ();
 sg13g2_decap_8 FILLER_26_1332 ();
 sg13g2_decap_8 FILLER_26_1339 ();
 sg13g2_decap_8 FILLER_26_1346 ();
 sg13g2_fill_2 FILLER_26_1353 ();
 sg13g2_fill_1 FILLER_26_1372 ();
 sg13g2_fill_1 FILLER_26_1384 ();
 sg13g2_fill_2 FILLER_26_1396 ();
 sg13g2_fill_2 FILLER_26_1410 ();
 sg13g2_fill_1 FILLER_26_1447 ();
 sg13g2_decap_8 FILLER_26_1459 ();
 sg13g2_decap_4 FILLER_26_1466 ();
 sg13g2_decap_8 FILLER_26_1482 ();
 sg13g2_fill_2 FILLER_26_1489 ();
 sg13g2_fill_1 FILLER_26_1491 ();
 sg13g2_fill_1 FILLER_26_1496 ();
 sg13g2_fill_2 FILLER_26_1505 ();
 sg13g2_fill_1 FILLER_26_1515 ();
 sg13g2_fill_1 FILLER_26_1522 ();
 sg13g2_fill_1 FILLER_26_1528 ();
 sg13g2_fill_1 FILLER_26_1533 ();
 sg13g2_fill_1 FILLER_26_1539 ();
 sg13g2_decap_8 FILLER_26_1549 ();
 sg13g2_decap_8 FILLER_26_1556 ();
 sg13g2_decap_8 FILLER_26_1563 ();
 sg13g2_decap_8 FILLER_26_1570 ();
 sg13g2_fill_2 FILLER_26_1577 ();
 sg13g2_fill_1 FILLER_26_1579 ();
 sg13g2_decap_4 FILLER_26_1592 ();
 sg13g2_fill_1 FILLER_26_1596 ();
 sg13g2_fill_1 FILLER_26_1603 ();
 sg13g2_fill_2 FILLER_26_1609 ();
 sg13g2_fill_2 FILLER_26_1615 ();
 sg13g2_fill_2 FILLER_26_1622 ();
 sg13g2_fill_1 FILLER_26_1633 ();
 sg13g2_decap_8 FILLER_26_1638 ();
 sg13g2_decap_8 FILLER_26_1645 ();
 sg13g2_decap_8 FILLER_26_1652 ();
 sg13g2_decap_8 FILLER_26_1659 ();
 sg13g2_decap_8 FILLER_26_1666 ();
 sg13g2_fill_2 FILLER_26_1673 ();
 sg13g2_fill_1 FILLER_26_1675 ();
 sg13g2_fill_1 FILLER_26_1697 ();
 sg13g2_decap_8 FILLER_26_1728 ();
 sg13g2_fill_2 FILLER_26_1735 ();
 sg13g2_fill_1 FILLER_26_1737 ();
 sg13g2_fill_2 FILLER_26_1748 ();
 sg13g2_fill_2 FILLER_26_1754 ();
 sg13g2_fill_1 FILLER_26_1756 ();
 sg13g2_fill_2 FILLER_26_1763 ();
 sg13g2_fill_1 FILLER_26_1796 ();
 sg13g2_fill_2 FILLER_26_1801 ();
 sg13g2_fill_2 FILLER_26_1862 ();
 sg13g2_fill_1 FILLER_26_1864 ();
 sg13g2_fill_2 FILLER_26_1869 ();
 sg13g2_fill_1 FILLER_26_1871 ();
 sg13g2_decap_4 FILLER_26_1898 ();
 sg13g2_fill_1 FILLER_26_1902 ();
 sg13g2_fill_1 FILLER_26_1933 ();
 sg13g2_fill_2 FILLER_26_1943 ();
 sg13g2_fill_1 FILLER_26_1945 ();
 sg13g2_decap_4 FILLER_26_1950 ();
 sg13g2_fill_1 FILLER_26_1990 ();
 sg13g2_decap_4 FILLER_26_2001 ();
 sg13g2_fill_1 FILLER_26_2005 ();
 sg13g2_decap_4 FILLER_26_2027 ();
 sg13g2_fill_1 FILLER_26_2070 ();
 sg13g2_decap_8 FILLER_26_2076 ();
 sg13g2_fill_2 FILLER_26_2087 ();
 sg13g2_decap_8 FILLER_26_2125 ();
 sg13g2_decap_8 FILLER_26_2132 ();
 sg13g2_decap_8 FILLER_26_2139 ();
 sg13g2_fill_1 FILLER_26_2146 ();
 sg13g2_fill_1 FILLER_26_2151 ();
 sg13g2_fill_2 FILLER_26_2173 ();
 sg13g2_fill_1 FILLER_26_2175 ();
 sg13g2_decap_4 FILLER_26_2202 ();
 sg13g2_fill_2 FILLER_26_2206 ();
 sg13g2_fill_2 FILLER_26_2234 ();
 sg13g2_fill_1 FILLER_26_2236 ();
 sg13g2_decap_8 FILLER_26_2247 ();
 sg13g2_fill_1 FILLER_26_2254 ();
 sg13g2_fill_1 FILLER_26_2291 ();
 sg13g2_fill_2 FILLER_26_2302 ();
 sg13g2_decap_8 FILLER_26_2356 ();
 sg13g2_decap_8 FILLER_26_2363 ();
 sg13g2_decap_8 FILLER_26_2396 ();
 sg13g2_fill_1 FILLER_26_2403 ();
 sg13g2_fill_2 FILLER_26_2413 ();
 sg13g2_fill_1 FILLER_26_2436 ();
 sg13g2_fill_1 FILLER_26_2453 ();
 sg13g2_decap_8 FILLER_26_2490 ();
 sg13g2_decap_4 FILLER_26_2497 ();
 sg13g2_decap_8 FILLER_26_2505 ();
 sg13g2_fill_2 FILLER_26_2512 ();
 sg13g2_decap_8 FILLER_26_2533 ();
 sg13g2_decap_8 FILLER_26_2540 ();
 sg13g2_decap_8 FILLER_26_2547 ();
 sg13g2_fill_2 FILLER_26_2554 ();
 sg13g2_fill_1 FILLER_26_2556 ();
 sg13g2_decap_4 FILLER_26_2584 ();
 sg13g2_fill_1 FILLER_26_2588 ();
 sg13g2_decap_8 FILLER_26_2593 ();
 sg13g2_decap_4 FILLER_26_2600 ();
 sg13g2_fill_2 FILLER_26_2604 ();
 sg13g2_fill_1 FILLER_26_2616 ();
 sg13g2_decap_8 FILLER_26_2643 ();
 sg13g2_decap_8 FILLER_26_2650 ();
 sg13g2_decap_8 FILLER_26_2657 ();
 sg13g2_decap_4 FILLER_26_2664 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_43 ();
 sg13g2_decap_8 FILLER_27_85 ();
 sg13g2_decap_4 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_134 ();
 sg13g2_decap_4 FILLER_27_141 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_decap_4 FILLER_27_196 ();
 sg13g2_fill_2 FILLER_27_200 ();
 sg13g2_fill_1 FILLER_27_210 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_fill_1 FILLER_27_226 ();
 sg13g2_fill_1 FILLER_27_250 ();
 sg13g2_decap_4 FILLER_27_266 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_decap_4 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_279 ();
 sg13g2_fill_2 FILLER_27_291 ();
 sg13g2_fill_2 FILLER_27_297 ();
 sg13g2_decap_4 FILLER_27_304 ();
 sg13g2_fill_1 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_314 ();
 sg13g2_fill_2 FILLER_27_325 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_fill_2 FILLER_27_354 ();
 sg13g2_fill_2 FILLER_27_382 ();
 sg13g2_fill_1 FILLER_27_466 ();
 sg13g2_fill_2 FILLER_27_472 ();
 sg13g2_decap_4 FILLER_27_479 ();
 sg13g2_fill_1 FILLER_27_483 ();
 sg13g2_decap_8 FILLER_27_488 ();
 sg13g2_fill_2 FILLER_27_495 ();
 sg13g2_decap_4 FILLER_27_501 ();
 sg13g2_fill_1 FILLER_27_505 ();
 sg13g2_decap_8 FILLER_27_511 ();
 sg13g2_decap_4 FILLER_27_529 ();
 sg13g2_fill_2 FILLER_27_547 ();
 sg13g2_decap_4 FILLER_27_563 ();
 sg13g2_fill_2 FILLER_27_567 ();
 sg13g2_decap_4 FILLER_27_632 ();
 sg13g2_fill_2 FILLER_27_645 ();
 sg13g2_fill_2 FILLER_27_674 ();
 sg13g2_fill_2 FILLER_27_680 ();
 sg13g2_fill_2 FILLER_27_692 ();
 sg13g2_fill_1 FILLER_27_710 ();
 sg13g2_fill_1 FILLER_27_724 ();
 sg13g2_fill_1 FILLER_27_735 ();
 sg13g2_fill_2 FILLER_27_753 ();
 sg13g2_fill_1 FILLER_27_775 ();
 sg13g2_fill_1 FILLER_27_810 ();
 sg13g2_fill_2 FILLER_27_844 ();
 sg13g2_decap_4 FILLER_27_915 ();
 sg13g2_fill_2 FILLER_27_919 ();
 sg13g2_decap_8 FILLER_27_929 ();
 sg13g2_decap_4 FILLER_27_940 ();
 sg13g2_fill_1 FILLER_27_944 ();
 sg13g2_fill_2 FILLER_27_955 ();
 sg13g2_fill_1 FILLER_27_1004 ();
 sg13g2_fill_2 FILLER_27_1031 ();
 sg13g2_fill_1 FILLER_27_1033 ();
 sg13g2_decap_8 FILLER_27_1039 ();
 sg13g2_fill_1 FILLER_27_1046 ();
 sg13g2_fill_2 FILLER_27_1051 ();
 sg13g2_fill_1 FILLER_27_1053 ();
 sg13g2_fill_1 FILLER_27_1085 ();
 sg13g2_fill_2 FILLER_27_1107 ();
 sg13g2_fill_1 FILLER_27_1114 ();
 sg13g2_fill_2 FILLER_27_1123 ();
 sg13g2_decap_4 FILLER_27_1155 ();
 sg13g2_fill_2 FILLER_27_1182 ();
 sg13g2_fill_1 FILLER_27_1246 ();
 sg13g2_fill_2 FILLER_27_1268 ();
 sg13g2_fill_2 FILLER_27_1274 ();
 sg13g2_fill_2 FILLER_27_1302 ();
 sg13g2_fill_1 FILLER_27_1309 ();
 sg13g2_fill_2 FILLER_27_1314 ();
 sg13g2_fill_1 FILLER_27_1316 ();
 sg13g2_decap_4 FILLER_27_1353 ();
 sg13g2_fill_2 FILLER_27_1357 ();
 sg13g2_fill_2 FILLER_27_1373 ();
 sg13g2_fill_1 FILLER_27_1415 ();
 sg13g2_fill_2 FILLER_27_1422 ();
 sg13g2_fill_2 FILLER_27_1429 ();
 sg13g2_fill_2 FILLER_27_1436 ();
 sg13g2_fill_1 FILLER_27_1438 ();
 sg13g2_fill_2 FILLER_27_1443 ();
 sg13g2_fill_1 FILLER_27_1445 ();
 sg13g2_fill_2 FILLER_27_1454 ();
 sg13g2_decap_8 FILLER_27_1466 ();
 sg13g2_fill_2 FILLER_27_1473 ();
 sg13g2_decap_8 FILLER_27_1482 ();
 sg13g2_decap_4 FILLER_27_1489 ();
 sg13g2_decap_4 FILLER_27_1498 ();
 sg13g2_fill_2 FILLER_27_1507 ();
 sg13g2_fill_1 FILLER_27_1509 ();
 sg13g2_fill_1 FILLER_27_1515 ();
 sg13g2_fill_2 FILLER_27_1521 ();
 sg13g2_fill_1 FILLER_27_1523 ();
 sg13g2_fill_2 FILLER_27_1534 ();
 sg13g2_fill_2 FILLER_27_1550 ();
 sg13g2_fill_1 FILLER_27_1552 ();
 sg13g2_decap_4 FILLER_27_1569 ();
 sg13g2_fill_2 FILLER_27_1573 ();
 sg13g2_decap_4 FILLER_27_1607 ();
 sg13g2_fill_1 FILLER_27_1611 ();
 sg13g2_decap_4 FILLER_27_1657 ();
 sg13g2_decap_4 FILLER_27_1674 ();
 sg13g2_decap_8 FILLER_27_1734 ();
 sg13g2_decap_8 FILLER_27_1741 ();
 sg13g2_fill_2 FILLER_27_1748 ();
 sg13g2_fill_1 FILLER_27_1750 ();
 sg13g2_fill_2 FILLER_27_1797 ();
 sg13g2_decap_8 FILLER_27_1825 ();
 sg13g2_fill_2 FILLER_27_1841 ();
 sg13g2_fill_1 FILLER_27_1843 ();
 sg13g2_fill_2 FILLER_27_1860 ();
 sg13g2_decap_8 FILLER_27_1887 ();
 sg13g2_decap_8 FILLER_27_1894 ();
 sg13g2_decap_8 FILLER_27_1901 ();
 sg13g2_decap_4 FILLER_27_1908 ();
 sg13g2_fill_1 FILLER_27_1912 ();
 sg13g2_fill_2 FILLER_27_1927 ();
 sg13g2_fill_2 FILLER_27_1948 ();
 sg13g2_fill_1 FILLER_27_1950 ();
 sg13g2_decap_8 FILLER_27_1961 ();
 sg13g2_fill_2 FILLER_27_1968 ();
 sg13g2_fill_1 FILLER_27_1970 ();
 sg13g2_fill_1 FILLER_27_1975 ();
 sg13g2_decap_8 FILLER_27_1980 ();
 sg13g2_fill_2 FILLER_27_1987 ();
 sg13g2_fill_2 FILLER_27_2027 ();
 sg13g2_decap_8 FILLER_27_2033 ();
 sg13g2_decap_8 FILLER_27_2080 ();
 sg13g2_fill_2 FILLER_27_2087 ();
 sg13g2_fill_1 FILLER_27_2089 ();
 sg13g2_fill_2 FILLER_27_2094 ();
 sg13g2_fill_1 FILLER_27_2096 ();
 sg13g2_fill_2 FILLER_27_2139 ();
 sg13g2_fill_1 FILLER_27_2211 ();
 sg13g2_fill_2 FILLER_27_2329 ();
 sg13g2_decap_8 FILLER_27_2357 ();
 sg13g2_decap_4 FILLER_27_2364 ();
 sg13g2_decap_4 FILLER_27_2411 ();
 sg13g2_fill_1 FILLER_27_2441 ();
 sg13g2_fill_1 FILLER_27_2566 ();
 sg13g2_decap_4 FILLER_27_2577 ();
 sg13g2_fill_2 FILLER_27_2581 ();
 sg13g2_decap_8 FILLER_27_2587 ();
 sg13g2_decap_8 FILLER_27_2594 ();
 sg13g2_fill_1 FILLER_27_2601 ();
 sg13g2_decap_8 FILLER_27_2631 ();
 sg13g2_decap_8 FILLER_27_2638 ();
 sg13g2_decap_8 FILLER_27_2645 ();
 sg13g2_decap_8 FILLER_27_2652 ();
 sg13g2_decap_8 FILLER_27_2659 ();
 sg13g2_decap_4 FILLER_27_2666 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_38 ();
 sg13g2_fill_1 FILLER_28_43 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_decap_8 FILLER_28_132 ();
 sg13g2_decap_4 FILLER_28_139 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_4 FILLER_28_173 ();
 sg13g2_fill_1 FILLER_28_177 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_fill_1 FILLER_28_286 ();
 sg13g2_fill_1 FILLER_28_292 ();
 sg13g2_fill_2 FILLER_28_323 ();
 sg13g2_decap_4 FILLER_28_344 ();
 sg13g2_fill_2 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_fill_2 FILLER_28_360 ();
 sg13g2_decap_4 FILLER_28_381 ();
 sg13g2_decap_4 FILLER_28_394 ();
 sg13g2_decap_4 FILLER_28_402 ();
 sg13g2_fill_1 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_4 FILLER_28_420 ();
 sg13g2_fill_2 FILLER_28_453 ();
 sg13g2_fill_2 FILLER_28_458 ();
 sg13g2_fill_2 FILLER_28_474 ();
 sg13g2_fill_1 FILLER_28_476 ();
 sg13g2_fill_1 FILLER_28_492 ();
 sg13g2_fill_1 FILLER_28_612 ();
 sg13g2_fill_2 FILLER_28_661 ();
 sg13g2_decap_4 FILLER_28_690 ();
 sg13g2_fill_2 FILLER_28_763 ();
 sg13g2_fill_2 FILLER_28_832 ();
 sg13g2_fill_2 FILLER_28_855 ();
 sg13g2_fill_1 FILLER_28_857 ();
 sg13g2_fill_2 FILLER_28_868 ();
 sg13g2_fill_1 FILLER_28_870 ();
 sg13g2_fill_2 FILLER_28_875 ();
 sg13g2_fill_1 FILLER_28_877 ();
 sg13g2_fill_2 FILLER_28_892 ();
 sg13g2_fill_1 FILLER_28_894 ();
 sg13g2_decap_8 FILLER_28_899 ();
 sg13g2_decap_8 FILLER_28_906 ();
 sg13g2_decap_4 FILLER_28_913 ();
 sg13g2_fill_2 FILLER_28_917 ();
 sg13g2_decap_8 FILLER_28_955 ();
 sg13g2_decap_4 FILLER_28_962 ();
 sg13g2_decap_8 FILLER_28_974 ();
 sg13g2_fill_2 FILLER_28_981 ();
 sg13g2_fill_2 FILLER_28_987 ();
 sg13g2_fill_1 FILLER_28_989 ();
 sg13g2_decap_4 FILLER_28_994 ();
 sg13g2_fill_2 FILLER_28_998 ();
 sg13g2_decap_8 FILLER_28_1004 ();
 sg13g2_fill_2 FILLER_28_1011 ();
 sg13g2_fill_1 FILLER_28_1013 ();
 sg13g2_decap_8 FILLER_28_1018 ();
 sg13g2_fill_1 FILLER_28_1025 ();
 sg13g2_decap_4 FILLER_28_1030 ();
 sg13g2_decap_4 FILLER_28_1064 ();
 sg13g2_decap_8 FILLER_28_1072 ();
 sg13g2_decap_8 FILLER_28_1083 ();
 sg13g2_fill_2 FILLER_28_1098 ();
 sg13g2_fill_1 FILLER_28_1105 ();
 sg13g2_fill_1 FILLER_28_1112 ();
 sg13g2_decap_4 FILLER_28_1127 ();
 sg13g2_fill_2 FILLER_28_1191 ();
 sg13g2_fill_1 FILLER_28_1197 ();
 sg13g2_fill_1 FILLER_28_1202 ();
 sg13g2_fill_1 FILLER_28_1239 ();
 sg13g2_decap_4 FILLER_28_1266 ();
 sg13g2_fill_2 FILLER_28_1278 ();
 sg13g2_decap_8 FILLER_28_1310 ();
 sg13g2_decap_4 FILLER_28_1317 ();
 sg13g2_fill_1 FILLER_28_1321 ();
 sg13g2_decap_8 FILLER_28_1336 ();
 sg13g2_decap_4 FILLER_28_1343 ();
 sg13g2_fill_1 FILLER_28_1378 ();
 sg13g2_fill_2 FILLER_28_1409 ();
 sg13g2_fill_1 FILLER_28_1411 ();
 sg13g2_fill_2 FILLER_28_1423 ();
 sg13g2_decap_8 FILLER_28_1430 ();
 sg13g2_decap_8 FILLER_28_1437 ();
 sg13g2_decap_4 FILLER_28_1464 ();
 sg13g2_fill_1 FILLER_28_1475 ();
 sg13g2_decap_4 FILLER_28_1494 ();
 sg13g2_fill_2 FILLER_28_1518 ();
 sg13g2_fill_1 FILLER_28_1525 ();
 sg13g2_fill_2 FILLER_28_1547 ();
 sg13g2_fill_1 FILLER_28_1549 ();
 sg13g2_fill_2 FILLER_28_1555 ();
 sg13g2_fill_2 FILLER_28_1564 ();
 sg13g2_fill_2 FILLER_28_1570 ();
 sg13g2_fill_1 FILLER_28_1579 ();
 sg13g2_decap_4 FILLER_28_1599 ();
 sg13g2_fill_2 FILLER_28_1603 ();
 sg13g2_fill_1 FILLER_28_1610 ();
 sg13g2_fill_1 FILLER_28_1680 ();
 sg13g2_fill_1 FILLER_28_1684 ();
 sg13g2_fill_1 FILLER_28_1697 ();
 sg13g2_decap_8 FILLER_28_1730 ();
 sg13g2_decap_8 FILLER_28_1737 ();
 sg13g2_fill_2 FILLER_28_1744 ();
 sg13g2_decap_4 FILLER_28_1749 ();
 sg13g2_fill_1 FILLER_28_1753 ();
 sg13g2_decap_8 FILLER_28_1796 ();
 sg13g2_fill_2 FILLER_28_1803 ();
 sg13g2_fill_1 FILLER_28_1805 ();
 sg13g2_decap_8 FILLER_28_1820 ();
 sg13g2_decap_8 FILLER_28_1827 ();
 sg13g2_decap_8 FILLER_28_1834 ();
 sg13g2_decap_4 FILLER_28_1841 ();
 sg13g2_decap_4 FILLER_28_1879 ();
 sg13g2_fill_2 FILLER_28_1883 ();
 sg13g2_decap_4 FILLER_28_1898 ();
 sg13g2_fill_2 FILLER_28_1958 ();
 sg13g2_fill_1 FILLER_28_1960 ();
 sg13g2_decap_8 FILLER_28_1971 ();
 sg13g2_decap_8 FILLER_28_1978 ();
 sg13g2_decap_4 FILLER_28_1999 ();
 sg13g2_fill_1 FILLER_28_2007 ();
 sg13g2_fill_1 FILLER_28_2047 ();
 sg13g2_decap_4 FILLER_28_2058 ();
 sg13g2_decap_8 FILLER_28_2070 ();
 sg13g2_decap_4 FILLER_28_2077 ();
 sg13g2_fill_2 FILLER_28_2081 ();
 sg13g2_fill_2 FILLER_28_2088 ();
 sg13g2_fill_1 FILLER_28_2090 ();
 sg13g2_decap_8 FILLER_28_2099 ();
 sg13g2_decap_4 FILLER_28_2106 ();
 sg13g2_fill_1 FILLER_28_2110 ();
 sg13g2_decap_4 FILLER_28_2141 ();
 sg13g2_fill_1 FILLER_28_2145 ();
 sg13g2_decap_4 FILLER_28_2169 ();
 sg13g2_fill_1 FILLER_28_2173 ();
 sg13g2_fill_2 FILLER_28_2200 ();
 sg13g2_decap_4 FILLER_28_2225 ();
 sg13g2_decap_8 FILLER_28_2239 ();
 sg13g2_fill_1 FILLER_28_2250 ();
 sg13g2_fill_2 FILLER_28_2274 ();
 sg13g2_fill_2 FILLER_28_2286 ();
 sg13g2_fill_2 FILLER_28_2307 ();
 sg13g2_fill_2 FILLER_28_2322 ();
 sg13g2_fill_1 FILLER_28_2342 ();
 sg13g2_fill_1 FILLER_28_2373 ();
 sg13g2_fill_2 FILLER_28_2396 ();
 sg13g2_fill_1 FILLER_28_2431 ();
 sg13g2_fill_1 FILLER_28_2458 ();
 sg13g2_fill_1 FILLER_28_2480 ();
 sg13g2_fill_1 FILLER_28_2485 ();
 sg13g2_decap_8 FILLER_28_2542 ();
 sg13g2_decap_8 FILLER_28_2622 ();
 sg13g2_decap_8 FILLER_28_2629 ();
 sg13g2_decap_8 FILLER_28_2636 ();
 sg13g2_decap_8 FILLER_28_2643 ();
 sg13g2_decap_8 FILLER_28_2650 ();
 sg13g2_decap_8 FILLER_28_2657 ();
 sg13g2_decap_4 FILLER_28_2664 ();
 sg13g2_fill_2 FILLER_28_2668 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_24 ();
 sg13g2_decap_4 FILLER_29_35 ();
 sg13g2_fill_1 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_44 ();
 sg13g2_decap_4 FILLER_29_51 ();
 sg13g2_fill_1 FILLER_29_59 ();
 sg13g2_decap_8 FILLER_29_86 ();
 sg13g2_fill_1 FILLER_29_93 ();
 sg13g2_fill_2 FILLER_29_99 ();
 sg13g2_fill_1 FILLER_29_101 ();
 sg13g2_fill_2 FILLER_29_154 ();
 sg13g2_decap_4 FILLER_29_187 ();
 sg13g2_fill_2 FILLER_29_209 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_fill_1 FILLER_29_283 ();
 sg13g2_fill_1 FILLER_29_289 ();
 sg13g2_decap_8 FILLER_29_351 ();
 sg13g2_decap_4 FILLER_29_358 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_411 ();
 sg13g2_decap_8 FILLER_29_439 ();
 sg13g2_fill_1 FILLER_29_463 ();
 sg13g2_decap_4 FILLER_29_478 ();
 sg13g2_fill_1 FILLER_29_508 ();
 sg13g2_fill_1 FILLER_29_518 ();
 sg13g2_decap_8 FILLER_29_560 ();
 sg13g2_decap_8 FILLER_29_567 ();
 sg13g2_fill_2 FILLER_29_630 ();
 sg13g2_fill_1 FILLER_29_632 ();
 sg13g2_fill_2 FILLER_29_664 ();
 sg13g2_fill_1 FILLER_29_696 ();
 sg13g2_fill_1 FILLER_29_741 ();
 sg13g2_fill_1 FILLER_29_825 ();
 sg13g2_fill_1 FILLER_29_852 ();
 sg13g2_fill_2 FILLER_29_879 ();
 sg13g2_fill_1 FILLER_29_902 ();
 sg13g2_decap_4 FILLER_29_924 ();
 sg13g2_fill_2 FILLER_29_928 ();
 sg13g2_decap_4 FILLER_29_970 ();
 sg13g2_fill_1 FILLER_29_974 ();
 sg13g2_fill_1 FILLER_29_1015 ();
 sg13g2_decap_8 FILLER_29_1020 ();
 sg13g2_decap_8 FILLER_29_1027 ();
 sg13g2_decap_8 FILLER_29_1034 ();
 sg13g2_fill_1 FILLER_29_1041 ();
 sg13g2_decap_8 FILLER_29_1046 ();
 sg13g2_fill_2 FILLER_29_1053 ();
 sg13g2_fill_1 FILLER_29_1068 ();
 sg13g2_fill_2 FILLER_29_1086 ();
 sg13g2_fill_1 FILLER_29_1088 ();
 sg13g2_fill_1 FILLER_29_1164 ();
 sg13g2_fill_1 FILLER_29_1169 ();
 sg13g2_decap_8 FILLER_29_1196 ();
 sg13g2_decap_8 FILLER_29_1203 ();
 sg13g2_decap_8 FILLER_29_1210 ();
 sg13g2_fill_1 FILLER_29_1217 ();
 sg13g2_fill_2 FILLER_29_1222 ();
 sg13g2_fill_1 FILLER_29_1224 ();
 sg13g2_decap_8 FILLER_29_1229 ();
 sg13g2_decap_8 FILLER_29_1236 ();
 sg13g2_decap_4 FILLER_29_1243 ();
 sg13g2_fill_1 FILLER_29_1247 ();
 sg13g2_decap_8 FILLER_29_1252 ();
 sg13g2_decap_8 FILLER_29_1259 ();
 sg13g2_fill_2 FILLER_29_1266 ();
 sg13g2_fill_1 FILLER_29_1268 ();
 sg13g2_fill_2 FILLER_29_1335 ();
 sg13g2_fill_1 FILLER_29_1337 ();
 sg13g2_fill_2 FILLER_29_1347 ();
 sg13g2_fill_2 FILLER_29_1416 ();
 sg13g2_decap_8 FILLER_29_1429 ();
 sg13g2_fill_1 FILLER_29_1445 ();
 sg13g2_fill_1 FILLER_29_1451 ();
 sg13g2_fill_2 FILLER_29_1476 ();
 sg13g2_fill_1 FILLER_29_1488 ();
 sg13g2_fill_1 FILLER_29_1553 ();
 sg13g2_fill_1 FILLER_29_1569 ();
 sg13g2_fill_2 FILLER_29_1581 ();
 sg13g2_fill_1 FILLER_29_1590 ();
 sg13g2_fill_2 FILLER_29_1644 ();
 sg13g2_fill_1 FILLER_29_1680 ();
 sg13g2_decap_4 FILLER_29_1734 ();
 sg13g2_fill_1 FILLER_29_1746 ();
 sg13g2_fill_2 FILLER_29_1754 ();
 sg13g2_fill_2 FILLER_29_1769 ();
 sg13g2_decap_4 FILLER_29_1793 ();
 sg13g2_fill_1 FILLER_29_1797 ();
 sg13g2_fill_1 FILLER_29_1838 ();
 sg13g2_fill_1 FILLER_29_1870 ();
 sg13g2_fill_2 FILLER_29_1875 ();
 sg13g2_fill_2 FILLER_29_1932 ();
 sg13g2_fill_2 FILLER_29_1974 ();
 sg13g2_fill_1 FILLER_29_1976 ();
 sg13g2_fill_2 FILLER_29_1987 ();
 sg13g2_fill_1 FILLER_29_1989 ();
 sg13g2_fill_2 FILLER_29_1994 ();
 sg13g2_fill_1 FILLER_29_2006 ();
 sg13g2_decap_4 FILLER_29_2052 ();
 sg13g2_fill_2 FILLER_29_2056 ();
 sg13g2_decap_8 FILLER_29_2088 ();
 sg13g2_decap_4 FILLER_29_2095 ();
 sg13g2_fill_2 FILLER_29_2109 ();
 sg13g2_fill_2 FILLER_29_2147 ();
 sg13g2_fill_1 FILLER_29_2149 ();
 sg13g2_fill_1 FILLER_29_2171 ();
 sg13g2_fill_2 FILLER_29_2176 ();
 sg13g2_fill_1 FILLER_29_2192 ();
 sg13g2_decap_8 FILLER_29_2227 ();
 sg13g2_decap_8 FILLER_29_2234 ();
 sg13g2_decap_8 FILLER_29_2241 ();
 sg13g2_fill_2 FILLER_29_2248 ();
 sg13g2_fill_1 FILLER_29_2250 ();
 sg13g2_decap_4 FILLER_29_2263 ();
 sg13g2_fill_1 FILLER_29_2267 ();
 sg13g2_fill_2 FILLER_29_2271 ();
 sg13g2_decap_4 FILLER_29_2318 ();
 sg13g2_fill_1 FILLER_29_2322 ();
 sg13g2_decap_8 FILLER_29_2333 ();
 sg13g2_decap_8 FILLER_29_2340 ();
 sg13g2_fill_2 FILLER_29_2347 ();
 sg13g2_fill_1 FILLER_29_2349 ();
 sg13g2_decap_4 FILLER_29_2354 ();
 sg13g2_fill_2 FILLER_29_2358 ();
 sg13g2_decap_8 FILLER_29_2363 ();
 sg13g2_decap_4 FILLER_29_2370 ();
 sg13g2_fill_1 FILLER_29_2428 ();
 sg13g2_decap_4 FILLER_29_2446 ();
 sg13g2_fill_1 FILLER_29_2454 ();
 sg13g2_fill_1 FILLER_29_2459 ();
 sg13g2_decap_4 FILLER_29_2469 ();
 sg13g2_fill_1 FILLER_29_2477 ();
 sg13g2_fill_2 FILLER_29_2491 ();
 sg13g2_fill_1 FILLER_29_2493 ();
 sg13g2_fill_2 FILLER_29_2498 ();
 sg13g2_fill_2 FILLER_29_2510 ();
 sg13g2_fill_1 FILLER_29_2512 ();
 sg13g2_fill_1 FILLER_29_2523 ();
 sg13g2_decap_8 FILLER_29_2598 ();
 sg13g2_fill_2 FILLER_29_2605 ();
 sg13g2_fill_1 FILLER_29_2607 ();
 sg13g2_decap_8 FILLER_29_2618 ();
 sg13g2_decap_8 FILLER_29_2625 ();
 sg13g2_decap_8 FILLER_29_2632 ();
 sg13g2_decap_8 FILLER_29_2639 ();
 sg13g2_decap_8 FILLER_29_2646 ();
 sg13g2_decap_8 FILLER_29_2653 ();
 sg13g2_decap_8 FILLER_29_2660 ();
 sg13g2_fill_2 FILLER_29_2667 ();
 sg13g2_fill_1 FILLER_29_2669 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_fill_2 FILLER_30_56 ();
 sg13g2_fill_1 FILLER_30_58 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_104 ();
 sg13g2_fill_2 FILLER_30_122 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_fill_2 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_141 ();
 sg13g2_fill_1 FILLER_30_143 ();
 sg13g2_decap_4 FILLER_30_148 ();
 sg13g2_fill_2 FILLER_30_152 ();
 sg13g2_decap_8 FILLER_30_158 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_191 ();
 sg13g2_fill_1 FILLER_30_218 ();
 sg13g2_fill_1 FILLER_30_249 ();
 sg13g2_fill_1 FILLER_30_256 ();
 sg13g2_fill_1 FILLER_30_266 ();
 sg13g2_decap_4 FILLER_30_302 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_1 FILLER_30_317 ();
 sg13g2_fill_2 FILLER_30_344 ();
 sg13g2_fill_1 FILLER_30_346 ();
 sg13g2_fill_2 FILLER_30_373 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_30_428 ();
 sg13g2_fill_1 FILLER_30_447 ();
 sg13g2_fill_2 FILLER_30_456 ();
 sg13g2_fill_1 FILLER_30_481 ();
 sg13g2_fill_1 FILLER_30_508 ();
 sg13g2_fill_2 FILLER_30_513 ();
 sg13g2_fill_2 FILLER_30_521 ();
 sg13g2_fill_2 FILLER_30_529 ();
 sg13g2_fill_1 FILLER_30_531 ();
 sg13g2_fill_2 FILLER_30_548 ();
 sg13g2_decap_4 FILLER_30_554 ();
 sg13g2_decap_4 FILLER_30_566 ();
 sg13g2_fill_1 FILLER_30_570 ();
 sg13g2_fill_1 FILLER_30_586 ();
 sg13g2_fill_2 FILLER_30_605 ();
 sg13g2_decap_8 FILLER_30_611 ();
 sg13g2_decap_8 FILLER_30_618 ();
 sg13g2_fill_1 FILLER_30_625 ();
 sg13g2_fill_2 FILLER_30_638 ();
 sg13g2_decap_4 FILLER_30_662 ();
 sg13g2_decap_8 FILLER_30_685 ();
 sg13g2_fill_1 FILLER_30_758 ();
 sg13g2_fill_2 FILLER_30_799 ();
 sg13g2_fill_2 FILLER_30_804 ();
 sg13g2_fill_2 FILLER_30_810 ();
 sg13g2_fill_1 FILLER_30_866 ();
 sg13g2_fill_1 FILLER_30_872 ();
 sg13g2_decap_8 FILLER_30_899 ();
 sg13g2_decap_8 FILLER_30_906 ();
 sg13g2_fill_1 FILLER_30_956 ();
 sg13g2_fill_2 FILLER_30_987 ();
 sg13g2_decap_4 FILLER_30_993 ();
 sg13g2_fill_2 FILLER_30_1023 ();
 sg13g2_fill_1 FILLER_30_1025 ();
 sg13g2_fill_1 FILLER_30_1082 ();
 sg13g2_fill_2 FILLER_30_1139 ();
 sg13g2_fill_1 FILLER_30_1141 ();
 sg13g2_fill_2 FILLER_30_1155 ();
 sg13g2_fill_1 FILLER_30_1178 ();
 sg13g2_fill_1 FILLER_30_1184 ();
 sg13g2_decap_8 FILLER_30_1210 ();
 sg13g2_decap_8 FILLER_30_1217 ();
 sg13g2_decap_8 FILLER_30_1224 ();
 sg13g2_decap_8 FILLER_30_1231 ();
 sg13g2_fill_1 FILLER_30_1238 ();
 sg13g2_fill_2 FILLER_30_1263 ();
 sg13g2_fill_1 FILLER_30_1265 ();
 sg13g2_decap_8 FILLER_30_1327 ();
 sg13g2_fill_2 FILLER_30_1334 ();
 sg13g2_fill_1 FILLER_30_1336 ();
 sg13g2_fill_1 FILLER_30_1373 ();
 sg13g2_fill_1 FILLER_30_1390 ();
 sg13g2_fill_2 FILLER_30_1400 ();
 sg13g2_fill_1 FILLER_30_1415 ();
 sg13g2_fill_2 FILLER_30_1424 ();
 sg13g2_fill_2 FILLER_30_1441 ();
 sg13g2_fill_1 FILLER_30_1449 ();
 sg13g2_fill_2 FILLER_30_1479 ();
 sg13g2_fill_1 FILLER_30_1505 ();
 sg13g2_fill_2 FILLER_30_1510 ();
 sg13g2_fill_1 FILLER_30_1512 ();
 sg13g2_fill_1 FILLER_30_1518 ();
 sg13g2_fill_1 FILLER_30_1529 ();
 sg13g2_decap_8 FILLER_30_1535 ();
 sg13g2_decap_4 FILLER_30_1542 ();
 sg13g2_fill_2 FILLER_30_1546 ();
 sg13g2_fill_2 FILLER_30_1553 ();
 sg13g2_fill_1 FILLER_30_1567 ();
 sg13g2_fill_1 FILLER_30_1573 ();
 sg13g2_fill_2 FILLER_30_1587 ();
 sg13g2_fill_2 FILLER_30_1638 ();
 sg13g2_fill_1 FILLER_30_1694 ();
 sg13g2_fill_1 FILLER_30_1731 ();
 sg13g2_fill_1 FILLER_30_1741 ();
 sg13g2_fill_2 FILLER_30_1778 ();
 sg13g2_decap_8 FILLER_30_1802 ();
 sg13g2_decap_4 FILLER_30_1809 ();
 sg13g2_fill_2 FILLER_30_1813 ();
 sg13g2_fill_2 FILLER_30_1823 ();
 sg13g2_fill_2 FILLER_30_1839 ();
 sg13g2_fill_1 FILLER_30_1841 ();
 sg13g2_fill_1 FILLER_30_1855 ();
 sg13g2_decap_8 FILLER_30_1882 ();
 sg13g2_fill_2 FILLER_30_1900 ();
 sg13g2_fill_2 FILLER_30_1938 ();
 sg13g2_fill_1 FILLER_30_1948 ();
 sg13g2_fill_2 FILLER_30_1953 ();
 sg13g2_fill_2 FILLER_30_1976 ();
 sg13g2_fill_1 FILLER_30_1978 ();
 sg13g2_decap_4 FILLER_30_2005 ();
 sg13g2_fill_2 FILLER_30_2009 ();
 sg13g2_fill_1 FILLER_30_2032 ();
 sg13g2_fill_2 FILLER_30_2066 ();
 sg13g2_fill_1 FILLER_30_2127 ();
 sg13g2_decap_4 FILLER_30_2154 ();
 sg13g2_decap_8 FILLER_30_2184 ();
 sg13g2_fill_2 FILLER_30_2201 ();
 sg13g2_fill_2 FILLER_30_2229 ();
 sg13g2_fill_1 FILLER_30_2231 ();
 sg13g2_decap_4 FILLER_30_2246 ();
 sg13g2_fill_1 FILLER_30_2250 ();
 sg13g2_fill_1 FILLER_30_2261 ();
 sg13g2_fill_2 FILLER_30_2302 ();
 sg13g2_decap_4 FILLER_30_2312 ();
 sg13g2_decap_8 FILLER_30_2320 ();
 sg13g2_decap_8 FILLER_30_2327 ();
 sg13g2_decap_8 FILLER_30_2334 ();
 sg13g2_fill_1 FILLER_30_2341 ();
 sg13g2_decap_8 FILLER_30_2352 ();
 sg13g2_fill_1 FILLER_30_2359 ();
 sg13g2_decap_8 FILLER_30_2370 ();
 sg13g2_fill_1 FILLER_30_2377 ();
 sg13g2_decap_8 FILLER_30_2381 ();
 sg13g2_fill_2 FILLER_30_2388 ();
 sg13g2_fill_1 FILLER_30_2390 ();
 sg13g2_fill_2 FILLER_30_2444 ();
 sg13g2_fill_1 FILLER_30_2446 ();
 sg13g2_decap_8 FILLER_30_2451 ();
 sg13g2_decap_4 FILLER_30_2458 ();
 sg13g2_decap_8 FILLER_30_2482 ();
 sg13g2_decap_8 FILLER_30_2489 ();
 sg13g2_decap_8 FILLER_30_2496 ();
 sg13g2_decap_8 FILLER_30_2503 ();
 sg13g2_decap_8 FILLER_30_2510 ();
 sg13g2_fill_1 FILLER_30_2553 ();
 sg13g2_fill_1 FILLER_30_2584 ();
 sg13g2_decap_4 FILLER_30_2589 ();
 sg13g2_decap_8 FILLER_30_2644 ();
 sg13g2_decap_8 FILLER_30_2651 ();
 sg13g2_decap_8 FILLER_30_2658 ();
 sg13g2_decap_4 FILLER_30_2665 ();
 sg13g2_fill_1 FILLER_30_2669 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_2 FILLER_31_46 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_82 ();
 sg13g2_fill_1 FILLER_31_87 ();
 sg13g2_decap_8 FILLER_31_92 ();
 sg13g2_fill_1 FILLER_31_99 ();
 sg13g2_decap_8 FILLER_31_135 ();
 sg13g2_decap_8 FILLER_31_142 ();
 sg13g2_decap_8 FILLER_31_149 ();
 sg13g2_decap_8 FILLER_31_156 ();
 sg13g2_decap_8 FILLER_31_163 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_fill_1 FILLER_31_177 ();
 sg13g2_fill_2 FILLER_31_208 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_fill_2 FILLER_31_232 ();
 sg13g2_fill_1 FILLER_31_234 ();
 sg13g2_fill_1 FILLER_31_239 ();
 sg13g2_fill_1 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_288 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_1 FILLER_31_297 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_4 FILLER_31_309 ();
 sg13g2_decap_4 FILLER_31_318 ();
 sg13g2_fill_1 FILLER_31_322 ();
 sg13g2_fill_1 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_352 ();
 sg13g2_fill_2 FILLER_31_399 ();
 sg13g2_fill_1 FILLER_31_411 ();
 sg13g2_fill_2 FILLER_31_499 ();
 sg13g2_fill_1 FILLER_31_501 ();
 sg13g2_decap_8 FILLER_31_537 ();
 sg13g2_decap_4 FILLER_31_544 ();
 sg13g2_fill_2 FILLER_31_548 ();
 sg13g2_decap_4 FILLER_31_553 ();
 sg13g2_fill_2 FILLER_31_557 ();
 sg13g2_fill_1 FILLER_31_594 ();
 sg13g2_decap_4 FILLER_31_615 ();
 sg13g2_fill_2 FILLER_31_619 ();
 sg13g2_decap_8 FILLER_31_633 ();
 sg13g2_fill_1 FILLER_31_640 ();
 sg13g2_fill_2 FILLER_31_649 ();
 sg13g2_fill_2 FILLER_31_661 ();
 sg13g2_fill_2 FILLER_31_689 ();
 sg13g2_fill_2 FILLER_31_700 ();
 sg13g2_fill_2 FILLER_31_710 ();
 sg13g2_fill_2 FILLER_31_742 ();
 sg13g2_fill_2 FILLER_31_812 ();
 sg13g2_fill_2 FILLER_31_842 ();
 sg13g2_decap_8 FILLER_31_848 ();
 sg13g2_decap_4 FILLER_31_855 ();
 sg13g2_fill_1 FILLER_31_859 ();
 sg13g2_decap_8 FILLER_31_906 ();
 sg13g2_fill_2 FILLER_31_913 ();
 sg13g2_fill_1 FILLER_31_925 ();
 sg13g2_fill_2 FILLER_31_930 ();
 sg13g2_decap_8 FILLER_31_937 ();
 sg13g2_fill_2 FILLER_31_1069 ();
 sg13g2_fill_1 FILLER_31_1110 ();
 sg13g2_fill_1 FILLER_31_1138 ();
 sg13g2_fill_1 FILLER_31_1149 ();
 sg13g2_fill_2 FILLER_31_1154 ();
 sg13g2_decap_4 FILLER_31_1169 ();
 sg13g2_fill_1 FILLER_31_1173 ();
 sg13g2_fill_1 FILLER_31_1179 ();
 sg13g2_fill_1 FILLER_31_1184 ();
 sg13g2_fill_2 FILLER_31_1189 ();
 sg13g2_fill_1 FILLER_31_1191 ();
 sg13g2_decap_4 FILLER_31_1231 ();
 sg13g2_fill_1 FILLER_31_1248 ();
 sg13g2_decap_4 FILLER_31_1288 ();
 sg13g2_fill_1 FILLER_31_1292 ();
 sg13g2_decap_8 FILLER_31_1297 ();
 sg13g2_decap_8 FILLER_31_1304 ();
 sg13g2_fill_2 FILLER_31_1311 ();
 sg13g2_fill_1 FILLER_31_1313 ();
 sg13g2_decap_8 FILLER_31_1328 ();
 sg13g2_decap_4 FILLER_31_1335 ();
 sg13g2_fill_2 FILLER_31_1353 ();
 sg13g2_decap_4 FILLER_31_1429 ();
 sg13g2_fill_1 FILLER_31_1433 ();
 sg13g2_fill_2 FILLER_31_1447 ();
 sg13g2_fill_1 FILLER_31_1449 ();
 sg13g2_fill_2 FILLER_31_1473 ();
 sg13g2_fill_1 FILLER_31_1475 ();
 sg13g2_fill_1 FILLER_31_1517 ();
 sg13g2_fill_1 FILLER_31_1523 ();
 sg13g2_decap_4 FILLER_31_1530 ();
 sg13g2_fill_2 FILLER_31_1534 ();
 sg13g2_decap_4 FILLER_31_1541 ();
 sg13g2_decap_8 FILLER_31_1551 ();
 sg13g2_fill_2 FILLER_31_1558 ();
 sg13g2_fill_1 FILLER_31_1560 ();
 sg13g2_fill_1 FILLER_31_1566 ();
 sg13g2_fill_1 FILLER_31_1572 ();
 sg13g2_fill_1 FILLER_31_1583 ();
 sg13g2_fill_1 FILLER_31_1589 ();
 sg13g2_fill_1 FILLER_31_1597 ();
 sg13g2_fill_1 FILLER_31_1646 ();
 sg13g2_fill_1 FILLER_31_1707 ();
 sg13g2_fill_2 FILLER_31_1756 ();
 sg13g2_decap_4 FILLER_31_1808 ();
 sg13g2_fill_1 FILLER_31_1812 ();
 sg13g2_decap_4 FILLER_31_1818 ();
 sg13g2_fill_1 FILLER_31_1822 ();
 sg13g2_fill_2 FILLER_31_1863 ();
 sg13g2_decap_8 FILLER_31_1903 ();
 sg13g2_fill_2 FILLER_31_1910 ();
 sg13g2_fill_1 FILLER_31_1941 ();
 sg13g2_fill_1 FILLER_31_1968 ();
 sg13g2_fill_1 FILLER_31_1979 ();
 sg13g2_fill_2 FILLER_31_2032 ();
 sg13g2_decap_4 FILLER_31_2077 ();
 sg13g2_decap_8 FILLER_31_2111 ();
 sg13g2_decap_4 FILLER_31_2130 ();
 sg13g2_fill_2 FILLER_31_2148 ();
 sg13g2_fill_1 FILLER_31_2150 ();
 sg13g2_decap_4 FILLER_31_2161 ();
 sg13g2_fill_2 FILLER_31_2165 ();
 sg13g2_decap_8 FILLER_31_2171 ();
 sg13g2_decap_8 FILLER_31_2178 ();
 sg13g2_fill_2 FILLER_31_2185 ();
 sg13g2_fill_1 FILLER_31_2187 ();
 sg13g2_fill_1 FILLER_31_2192 ();
 sg13g2_fill_2 FILLER_31_2219 ();
 sg13g2_fill_2 FILLER_31_2298 ();
 sg13g2_fill_1 FILLER_31_2340 ();
 sg13g2_fill_2 FILLER_31_2367 ();
 sg13g2_fill_2 FILLER_31_2395 ();
 sg13g2_fill_1 FILLER_31_2397 ();
 sg13g2_fill_2 FILLER_31_2435 ();
 sg13g2_fill_1 FILLER_31_2437 ();
 sg13g2_fill_2 FILLER_31_2468 ();
 sg13g2_fill_1 FILLER_31_2470 ();
 sg13g2_decap_4 FILLER_31_2501 ();
 sg13g2_fill_2 FILLER_31_2509 ();
 sg13g2_decap_4 FILLER_31_2536 ();
 sg13g2_fill_1 FILLER_31_2540 ();
 sg13g2_decap_8 FILLER_31_2551 ();
 sg13g2_decap_8 FILLER_31_2558 ();
 sg13g2_fill_1 FILLER_31_2565 ();
 sg13g2_decap_8 FILLER_31_2570 ();
 sg13g2_decap_4 FILLER_31_2577 ();
 sg13g2_decap_8 FILLER_31_2651 ();
 sg13g2_decap_8 FILLER_31_2658 ();
 sg13g2_decap_4 FILLER_31_2665 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_decap_4 FILLER_32_32 ();
 sg13g2_decap_4 FILLER_32_40 ();
 sg13g2_decap_8 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_76 ();
 sg13g2_decap_8 FILLER_32_83 ();
 sg13g2_decap_8 FILLER_32_90 ();
 sg13g2_decap_8 FILLER_32_97 ();
 sg13g2_fill_2 FILLER_32_104 ();
 sg13g2_fill_1 FILLER_32_106 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_4 FILLER_32_144 ();
 sg13g2_fill_1 FILLER_32_148 ();
 sg13g2_fill_2 FILLER_32_175 ();
 sg13g2_decap_4 FILLER_32_203 ();
 sg13g2_fill_2 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_1 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_242 ();
 sg13g2_decap_4 FILLER_32_247 ();
 sg13g2_fill_2 FILLER_32_251 ();
 sg13g2_fill_1 FILLER_32_261 ();
 sg13g2_fill_1 FILLER_32_269 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_decap_4 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_fill_2 FILLER_32_300 ();
 sg13g2_fill_2 FILLER_32_307 ();
 sg13g2_fill_2 FILLER_32_313 ();
 sg13g2_fill_1 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_fill_2 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_349 ();
 sg13g2_fill_2 FILLER_32_359 ();
 sg13g2_fill_1 FILLER_32_361 ();
 sg13g2_fill_2 FILLER_32_400 ();
 sg13g2_fill_1 FILLER_32_402 ();
 sg13g2_fill_1 FILLER_32_501 ();
 sg13g2_fill_2 FILLER_32_517 ();
 sg13g2_decap_4 FILLER_32_525 ();
 sg13g2_fill_1 FILLER_32_529 ();
 sg13g2_decap_4 FILLER_32_535 ();
 sg13g2_fill_1 FILLER_32_539 ();
 sg13g2_decap_4 FILLER_32_545 ();
 sg13g2_fill_1 FILLER_32_549 ();
 sg13g2_fill_2 FILLER_32_668 ();
 sg13g2_fill_2 FILLER_32_674 ();
 sg13g2_fill_1 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_681 ();
 sg13g2_decap_8 FILLER_32_688 ();
 sg13g2_fill_1 FILLER_32_699 ();
 sg13g2_fill_2 FILLER_32_737 ();
 sg13g2_fill_1 FILLER_32_758 ();
 sg13g2_fill_1 FILLER_32_767 ();
 sg13g2_fill_2 FILLER_32_776 ();
 sg13g2_fill_2 FILLER_32_788 ();
 sg13g2_fill_1 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_843 ();
 sg13g2_decap_8 FILLER_32_850 ();
 sg13g2_decap_8 FILLER_32_857 ();
 sg13g2_fill_2 FILLER_32_864 ();
 sg13g2_fill_1 FILLER_32_866 ();
 sg13g2_decap_8 FILLER_32_897 ();
 sg13g2_decap_8 FILLER_32_904 ();
 sg13g2_decap_8 FILLER_32_911 ();
 sg13g2_fill_2 FILLER_32_918 ();
 sg13g2_fill_1 FILLER_32_920 ();
 sg13g2_fill_2 FILLER_32_947 ();
 sg13g2_fill_1 FILLER_32_949 ();
 sg13g2_fill_1 FILLER_32_967 ();
 sg13g2_decap_8 FILLER_32_977 ();
 sg13g2_decap_8 FILLER_32_984 ();
 sg13g2_fill_1 FILLER_32_991 ();
 sg13g2_fill_2 FILLER_32_1070 ();
 sg13g2_decap_4 FILLER_32_1098 ();
 sg13g2_fill_1 FILLER_32_1102 ();
 sg13g2_fill_1 FILLER_32_1107 ();
 sg13g2_fill_2 FILLER_32_1137 ();
 sg13g2_fill_1 FILLER_32_1139 ();
 sg13g2_fill_2 FILLER_32_1148 ();
 sg13g2_fill_2 FILLER_32_1197 ();
 sg13g2_fill_2 FILLER_32_1204 ();
 sg13g2_fill_2 FILLER_32_1232 ();
 sg13g2_fill_1 FILLER_32_1234 ();
 sg13g2_fill_1 FILLER_32_1261 ();
 sg13g2_decap_8 FILLER_32_1288 ();
 sg13g2_decap_8 FILLER_32_1295 ();
 sg13g2_decap_8 FILLER_32_1328 ();
 sg13g2_fill_2 FILLER_32_1335 ();
 sg13g2_fill_2 FILLER_32_1344 ();
 sg13g2_fill_1 FILLER_32_1346 ();
 sg13g2_fill_2 FILLER_32_1383 ();
 sg13g2_decap_4 FILLER_32_1391 ();
 sg13g2_fill_1 FILLER_32_1395 ();
 sg13g2_fill_2 FILLER_32_1418 ();
 sg13g2_fill_2 FILLER_32_1435 ();
 sg13g2_fill_1 FILLER_32_1442 ();
 sg13g2_fill_1 FILLER_32_1450 ();
 sg13g2_fill_1 FILLER_32_1461 ();
 sg13g2_fill_2 FILLER_32_1472 ();
 sg13g2_fill_1 FILLER_32_1474 ();
 sg13g2_fill_1 FILLER_32_1491 ();
 sg13g2_decap_8 FILLER_32_1498 ();
 sg13g2_decap_4 FILLER_32_1505 ();
 sg13g2_fill_2 FILLER_32_1509 ();
 sg13g2_decap_4 FILLER_32_1528 ();
 sg13g2_fill_1 FILLER_32_1532 ();
 sg13g2_fill_2 FILLER_32_1543 ();
 sg13g2_fill_2 FILLER_32_1553 ();
 sg13g2_fill_1 FILLER_32_1555 ();
 sg13g2_fill_1 FILLER_32_1585 ();
 sg13g2_fill_2 FILLER_32_1602 ();
 sg13g2_fill_1 FILLER_32_1635 ();
 sg13g2_fill_1 FILLER_32_1702 ();
 sg13g2_fill_2 FILLER_32_1707 ();
 sg13g2_fill_1 FILLER_32_1752 ();
 sg13g2_decap_8 FILLER_32_1798 ();
 sg13g2_decap_8 FILLER_32_1805 ();
 sg13g2_fill_1 FILLER_32_1812 ();
 sg13g2_fill_2 FILLER_32_1817 ();
 sg13g2_decap_8 FILLER_32_1824 ();
 sg13g2_decap_8 FILLER_32_1831 ();
 sg13g2_decap_4 FILLER_32_1838 ();
 sg13g2_fill_1 FILLER_32_1842 ();
 sg13g2_fill_2 FILLER_32_1856 ();
 sg13g2_decap_8 FILLER_32_1876 ();
 sg13g2_decap_8 FILLER_32_1883 ();
 sg13g2_decap_8 FILLER_32_1890 ();
 sg13g2_decap_4 FILLER_32_1897 ();
 sg13g2_fill_1 FILLER_32_1950 ();
 sg13g2_fill_2 FILLER_32_1991 ();
 sg13g2_decap_8 FILLER_32_1998 ();
 sg13g2_fill_2 FILLER_32_2005 ();
 sg13g2_fill_2 FILLER_32_2012 ();
 sg13g2_decap_8 FILLER_32_2018 ();
 sg13g2_fill_2 FILLER_32_2025 ();
 sg13g2_fill_1 FILLER_32_2039 ();
 sg13g2_fill_2 FILLER_32_2121 ();
 sg13g2_decap_4 FILLER_32_2159 ();
 sg13g2_fill_1 FILLER_32_2163 ();
 sg13g2_decap_4 FILLER_32_2190 ();
 sg13g2_fill_1 FILLER_32_2219 ();
 sg13g2_decap_8 FILLER_32_2252 ();
 sg13g2_decap_8 FILLER_32_2289 ();
 sg13g2_decap_8 FILLER_32_2296 ();
 sg13g2_decap_8 FILLER_32_2303 ();
 sg13g2_fill_2 FILLER_32_2310 ();
 sg13g2_fill_1 FILLER_32_2312 ();
 sg13g2_fill_2 FILLER_32_2317 ();
 sg13g2_decap_4 FILLER_32_2340 ();
 sg13g2_fill_2 FILLER_32_2344 ();
 sg13g2_fill_1 FILLER_32_2350 ();
 sg13g2_fill_1 FILLER_32_2361 ();
 sg13g2_fill_2 FILLER_32_2396 ();
 sg13g2_fill_1 FILLER_32_2398 ();
 sg13g2_decap_8 FILLER_32_2403 ();
 sg13g2_fill_2 FILLER_32_2410 ();
 sg13g2_fill_2 FILLER_32_2427 ();
 sg13g2_decap_8 FILLER_32_2463 ();
 sg13g2_fill_2 FILLER_32_2470 ();
 sg13g2_decap_8 FILLER_32_2534 ();
 sg13g2_decap_8 FILLER_32_2541 ();
 sg13g2_decap_4 FILLER_32_2548 ();
 sg13g2_fill_1 FILLER_32_2552 ();
 sg13g2_decap_8 FILLER_32_2563 ();
 sg13g2_fill_2 FILLER_32_2570 ();
 sg13g2_fill_1 FILLER_32_2572 ();
 sg13g2_fill_2 FILLER_32_2583 ();
 sg13g2_decap_8 FILLER_32_2644 ();
 sg13g2_decap_8 FILLER_32_2651 ();
 sg13g2_decap_8 FILLER_32_2658 ();
 sg13g2_decap_4 FILLER_32_2665 ();
 sg13g2_fill_1 FILLER_32_2669 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_22 ();
 sg13g2_fill_2 FILLER_33_53 ();
 sg13g2_fill_1 FILLER_33_55 ();
 sg13g2_fill_2 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_128 ();
 sg13g2_fill_1 FILLER_33_155 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_decap_4 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_222 ();
 sg13g2_fill_2 FILLER_33_250 ();
 sg13g2_fill_1 FILLER_33_252 ();
 sg13g2_fill_2 FILLER_33_282 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_8 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_360 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_419 ();
 sg13g2_fill_2 FILLER_33_430 ();
 sg13g2_fill_1 FILLER_33_441 ();
 sg13g2_fill_2 FILLER_33_455 ();
 sg13g2_fill_2 FILLER_33_502 ();
 sg13g2_fill_2 FILLER_33_516 ();
 sg13g2_fill_1 FILLER_33_530 ();
 sg13g2_fill_1 FILLER_33_562 ();
 sg13g2_fill_2 FILLER_33_591 ();
 sg13g2_fill_1 FILLER_33_593 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_1 FILLER_33_610 ();
 sg13g2_decap_8 FILLER_33_619 ();
 sg13g2_fill_2 FILLER_33_626 ();
 sg13g2_decap_4 FILLER_33_634 ();
 sg13g2_fill_1 FILLER_33_638 ();
 sg13g2_fill_1 FILLER_33_643 ();
 sg13g2_fill_2 FILLER_33_650 ();
 sg13g2_fill_1 FILLER_33_655 ();
 sg13g2_decap_4 FILLER_33_661 ();
 sg13g2_fill_1 FILLER_33_665 ();
 sg13g2_fill_2 FILLER_33_675 ();
 sg13g2_fill_1 FILLER_33_677 ();
 sg13g2_decap_8 FILLER_33_683 ();
 sg13g2_fill_1 FILLER_33_708 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_808 ();
 sg13g2_decap_8 FILLER_33_815 ();
 sg13g2_decap_8 FILLER_33_822 ();
 sg13g2_decap_8 FILLER_33_829 ();
 sg13g2_decap_8 FILLER_33_836 ();
 sg13g2_decap_8 FILLER_33_843 ();
 sg13g2_fill_1 FILLER_33_850 ();
 sg13g2_decap_8 FILLER_33_859 ();
 sg13g2_fill_2 FILLER_33_866 ();
 sg13g2_fill_1 FILLER_33_868 ();
 sg13g2_fill_2 FILLER_33_890 ();
 sg13g2_fill_1 FILLER_33_892 ();
 sg13g2_decap_8 FILLER_33_897 ();
 sg13g2_decap_4 FILLER_33_904 ();
 sg13g2_fill_2 FILLER_33_908 ();
 sg13g2_decap_4 FILLER_33_917 ();
 sg13g2_fill_2 FILLER_33_925 ();
 sg13g2_fill_1 FILLER_33_927 ();
 sg13g2_fill_2 FILLER_33_946 ();
 sg13g2_decap_8 FILLER_33_982 ();
 sg13g2_decap_8 FILLER_33_989 ();
 sg13g2_fill_2 FILLER_33_996 ();
 sg13g2_fill_1 FILLER_33_998 ();
 sg13g2_decap_4 FILLER_33_1007 ();
 sg13g2_fill_1 FILLER_33_1011 ();
 sg13g2_decap_8 FILLER_33_1025 ();
 sg13g2_decap_4 FILLER_33_1032 ();
 sg13g2_fill_1 FILLER_33_1046 ();
 sg13g2_fill_2 FILLER_33_1074 ();
 sg13g2_fill_1 FILLER_33_1076 ();
 sg13g2_fill_2 FILLER_33_1108 ();
 sg13g2_fill_1 FILLER_33_1118 ();
 sg13g2_fill_2 FILLER_33_1124 ();
 sg13g2_decap_8 FILLER_33_1140 ();
 sg13g2_fill_2 FILLER_33_1147 ();
 sg13g2_fill_1 FILLER_33_1149 ();
 sg13g2_fill_1 FILLER_33_1220 ();
 sg13g2_decap_8 FILLER_33_1225 ();
 sg13g2_decap_4 FILLER_33_1232 ();
 sg13g2_fill_2 FILLER_33_1236 ();
 sg13g2_fill_1 FILLER_33_1260 ();
 sg13g2_fill_1 FILLER_33_1294 ();
 sg13g2_fill_2 FILLER_33_1300 ();
 sg13g2_decap_8 FILLER_33_1310 ();
 sg13g2_decap_8 FILLER_33_1317 ();
 sg13g2_decap_8 FILLER_33_1324 ();
 sg13g2_fill_2 FILLER_33_1331 ();
 sg13g2_decap_4 FILLER_33_1398 ();
 sg13g2_fill_1 FILLER_33_1415 ();
 sg13g2_decap_8 FILLER_33_1426 ();
 sg13g2_fill_1 FILLER_33_1433 ();
 sg13g2_decap_4 FILLER_33_1445 ();
 sg13g2_fill_1 FILLER_33_1449 ();
 sg13g2_fill_2 FILLER_33_1455 ();
 sg13g2_fill_1 FILLER_33_1465 ();
 sg13g2_fill_2 FILLER_33_1476 ();
 sg13g2_fill_2 FILLER_33_1485 ();
 sg13g2_decap_8 FILLER_33_1496 ();
 sg13g2_decap_4 FILLER_33_1503 ();
 sg13g2_fill_2 FILLER_33_1524 ();
 sg13g2_decap_8 FILLER_33_1547 ();
 sg13g2_decap_8 FILLER_33_1554 ();
 sg13g2_decap_8 FILLER_33_1561 ();
 sg13g2_fill_2 FILLER_33_1577 ();
 sg13g2_fill_1 FILLER_33_1579 ();
 sg13g2_fill_2 FILLER_33_1585 ();
 sg13g2_fill_1 FILLER_33_1587 ();
 sg13g2_fill_1 FILLER_33_1593 ();
 sg13g2_fill_1 FILLER_33_1688 ();
 sg13g2_decap_8 FILLER_33_1787 ();
 sg13g2_decap_4 FILLER_33_1794 ();
 sg13g2_fill_1 FILLER_33_1798 ();
 sg13g2_decap_8 FILLER_33_1818 ();
 sg13g2_decap_8 FILLER_33_1825 ();
 sg13g2_decap_8 FILLER_33_1832 ();
 sg13g2_decap_8 FILLER_33_1839 ();
 sg13g2_fill_1 FILLER_33_1846 ();
 sg13g2_decap_4 FILLER_33_1860 ();
 sg13g2_decap_8 FILLER_33_1877 ();
 sg13g2_decap_8 FILLER_33_1884 ();
 sg13g2_decap_8 FILLER_33_1891 ();
 sg13g2_decap_8 FILLER_33_1898 ();
 sg13g2_decap_8 FILLER_33_1905 ();
 sg13g2_fill_1 FILLER_33_1912 ();
 sg13g2_decap_4 FILLER_33_1917 ();
 sg13g2_fill_2 FILLER_33_1921 ();
 sg13g2_fill_2 FILLER_33_1929 ();
 sg13g2_fill_1 FILLER_33_1964 ();
 sg13g2_decap_8 FILLER_33_1998 ();
 sg13g2_fill_1 FILLER_33_2005 ();
 sg13g2_decap_8 FILLER_33_2011 ();
 sg13g2_fill_1 FILLER_33_2018 ();
 sg13g2_decap_4 FILLER_33_2031 ();
 sg13g2_decap_4 FILLER_33_2061 ();
 sg13g2_fill_2 FILLER_33_2065 ();
 sg13g2_fill_2 FILLER_33_2096 ();
 sg13g2_fill_2 FILLER_33_2145 ();
 sg13g2_fill_1 FILLER_33_2147 ();
 sg13g2_decap_8 FILLER_33_2182 ();
 sg13g2_fill_1 FILLER_33_2189 ();
 sg13g2_fill_2 FILLER_33_2205 ();
 sg13g2_fill_1 FILLER_33_2221 ();
 sg13g2_fill_2 FILLER_33_2230 ();
 sg13g2_fill_2 FILLER_33_2235 ();
 sg13g2_fill_1 FILLER_33_2271 ();
 sg13g2_fill_2 FILLER_33_2276 ();
 sg13g2_fill_1 FILLER_33_2282 ();
 sg13g2_fill_2 FILLER_33_2291 ();
 sg13g2_fill_1 FILLER_33_2293 ();
 sg13g2_fill_1 FILLER_33_2330 ();
 sg13g2_fill_1 FILLER_33_2433 ();
 sg13g2_fill_2 FILLER_33_2444 ();
 sg13g2_fill_1 FILLER_33_2490 ();
 sg13g2_fill_1 FILLER_33_2553 ();
 sg13g2_fill_1 FILLER_33_2558 ();
 sg13g2_fill_2 FILLER_33_2569 ();
 sg13g2_decap_4 FILLER_33_2602 ();
 sg13g2_fill_1 FILLER_33_2606 ();
 sg13g2_decap_8 FILLER_33_2617 ();
 sg13g2_fill_2 FILLER_33_2624 ();
 sg13g2_fill_1 FILLER_33_2626 ();
 sg13g2_decap_8 FILLER_33_2631 ();
 sg13g2_decap_8 FILLER_33_2638 ();
 sg13g2_decap_8 FILLER_33_2645 ();
 sg13g2_decap_8 FILLER_33_2652 ();
 sg13g2_decap_8 FILLER_33_2659 ();
 sg13g2_decap_4 FILLER_33_2666 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_2 FILLER_34_33 ();
 sg13g2_fill_1 FILLER_34_65 ();
 sg13g2_decap_4 FILLER_34_106 ();
 sg13g2_fill_1 FILLER_34_110 ();
 sg13g2_fill_2 FILLER_34_119 ();
 sg13g2_decap_8 FILLER_34_131 ();
 sg13g2_fill_2 FILLER_34_138 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_4 FILLER_34_151 ();
 sg13g2_fill_1 FILLER_34_155 ();
 sg13g2_fill_1 FILLER_34_190 ();
 sg13g2_fill_1 FILLER_34_259 ();
 sg13g2_fill_2 FILLER_34_286 ();
 sg13g2_decap_4 FILLER_34_314 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_decap_4 FILLER_34_330 ();
 sg13g2_decap_4 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_372 ();
 sg13g2_decap_8 FILLER_34_377 ();
 sg13g2_decap_8 FILLER_34_384 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_fill_1 FILLER_34_397 ();
 sg13g2_fill_1 FILLER_34_428 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_478 ();
 sg13g2_fill_2 FILLER_34_493 ();
 sg13g2_fill_2 FILLER_34_512 ();
 sg13g2_fill_1 FILLER_34_519 ();
 sg13g2_decap_8 FILLER_34_537 ();
 sg13g2_fill_2 FILLER_34_544 ();
 sg13g2_decap_8 FILLER_34_550 ();
 sg13g2_decap_4 FILLER_34_557 ();
 sg13g2_fill_1 FILLER_34_561 ();
 sg13g2_fill_1 FILLER_34_566 ();
 sg13g2_decap_8 FILLER_34_571 ();
 sg13g2_fill_1 FILLER_34_578 ();
 sg13g2_decap_8 FILLER_34_592 ();
 sg13g2_decap_8 FILLER_34_599 ();
 sg13g2_decap_8 FILLER_34_606 ();
 sg13g2_fill_1 FILLER_34_613 ();
 sg13g2_fill_2 FILLER_34_629 ();
 sg13g2_fill_2 FILLER_34_635 ();
 sg13g2_fill_1 FILLER_34_637 ();
 sg13g2_fill_1 FILLER_34_648 ();
 sg13g2_fill_2 FILLER_34_654 ();
 sg13g2_fill_1 FILLER_34_656 ();
 sg13g2_decap_8 FILLER_34_661 ();
 sg13g2_decap_8 FILLER_34_668 ();
 sg13g2_decap_8 FILLER_34_675 ();
 sg13g2_decap_8 FILLER_34_682 ();
 sg13g2_fill_1 FILLER_34_689 ();
 sg13g2_fill_1 FILLER_34_722 ();
 sg13g2_fill_2 FILLER_34_758 ();
 sg13g2_decap_8 FILLER_34_794 ();
 sg13g2_fill_1 FILLER_34_801 ();
 sg13g2_fill_1 FILLER_34_818 ();
 sg13g2_decap_8 FILLER_34_866 ();
 sg13g2_fill_1 FILLER_34_873 ();
 sg13g2_fill_1 FILLER_34_900 ();
 sg13g2_fill_1 FILLER_34_911 ();
 sg13g2_fill_1 FILLER_34_938 ();
 sg13g2_fill_1 FILLER_34_943 ();
 sg13g2_fill_2 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_994 ();
 sg13g2_fill_1 FILLER_34_1001 ();
 sg13g2_decap_4 FILLER_34_1011 ();
 sg13g2_fill_1 FILLER_34_1019 ();
 sg13g2_decap_8 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_34_1035 ();
 sg13g2_decap_4 FILLER_34_1042 ();
 sg13g2_fill_2 FILLER_34_1054 ();
 sg13g2_fill_2 FILLER_34_1076 ();
 sg13g2_fill_1 FILLER_34_1078 ();
 sg13g2_decap_4 FILLER_34_1091 ();
 sg13g2_fill_1 FILLER_34_1100 ();
 sg13g2_fill_2 FILLER_34_1110 ();
 sg13g2_fill_1 FILLER_34_1117 ();
 sg13g2_decap_8 FILLER_34_1144 ();
 sg13g2_decap_4 FILLER_34_1151 ();
 sg13g2_decap_8 FILLER_34_1186 ();
 sg13g2_decap_4 FILLER_34_1193 ();
 sg13g2_decap_4 FILLER_34_1201 ();
 sg13g2_fill_1 FILLER_34_1205 ();
 sg13g2_decap_8 FILLER_34_1210 ();
 sg13g2_decap_8 FILLER_34_1217 ();
 sg13g2_decap_8 FILLER_34_1224 ();
 sg13g2_fill_2 FILLER_34_1231 ();
 sg13g2_fill_1 FILLER_34_1263 ();
 sg13g2_fill_1 FILLER_34_1274 ();
 sg13g2_fill_1 FILLER_34_1279 ();
 sg13g2_fill_1 FILLER_34_1284 ();
 sg13g2_fill_1 FILLER_34_1311 ();
 sg13g2_fill_1 FILLER_34_1322 ();
 sg13g2_decap_4 FILLER_34_1362 ();
 sg13g2_fill_1 FILLER_34_1366 ();
 sg13g2_decap_8 FILLER_34_1371 ();
 sg13g2_fill_2 FILLER_34_1378 ();
 sg13g2_fill_1 FILLER_34_1380 ();
 sg13g2_fill_2 FILLER_34_1411 ();
 sg13g2_fill_2 FILLER_34_1421 ();
 sg13g2_fill_1 FILLER_34_1430 ();
 sg13g2_fill_1 FILLER_34_1490 ();
 sg13g2_decap_8 FILLER_34_1511 ();
 sg13g2_fill_2 FILLER_34_1518 ();
 sg13g2_fill_1 FILLER_34_1520 ();
 sg13g2_fill_2 FILLER_34_1526 ();
 sg13g2_fill_1 FILLER_34_1568 ();
 sg13g2_fill_2 FILLER_34_1583 ();
 sg13g2_fill_2 FILLER_34_1589 ();
 sg13g2_fill_1 FILLER_34_1591 ();
 sg13g2_fill_2 FILLER_34_1603 ();
 sg13g2_fill_2 FILLER_34_1625 ();
 sg13g2_fill_1 FILLER_34_1666 ();
 sg13g2_fill_1 FILLER_34_1693 ();
 sg13g2_fill_2 FILLER_34_1709 ();
 sg13g2_decap_4 FILLER_34_1762 ();
 sg13g2_decap_4 FILLER_34_1770 ();
 sg13g2_fill_2 FILLER_34_1774 ();
 sg13g2_decap_8 FILLER_34_1786 ();
 sg13g2_decap_8 FILLER_34_1793 ();
 sg13g2_fill_2 FILLER_34_1800 ();
 sg13g2_decap_8 FILLER_34_1837 ();
 sg13g2_decap_8 FILLER_34_1844 ();
 sg13g2_fill_2 FILLER_34_1851 ();
 sg13g2_fill_1 FILLER_34_1853 ();
 sg13g2_decap_8 FILLER_34_1897 ();
 sg13g2_decap_4 FILLER_34_1908 ();
 sg13g2_fill_1 FILLER_34_1912 ();
 sg13g2_fill_2 FILLER_34_1949 ();
 sg13g2_fill_2 FILLER_34_1996 ();
 sg13g2_fill_1 FILLER_34_2048 ();
 sg13g2_fill_2 FILLER_34_2080 ();
 sg13g2_fill_1 FILLER_34_2082 ();
 sg13g2_fill_1 FILLER_34_2104 ();
 sg13g2_fill_1 FILLER_34_2112 ();
 sg13g2_decap_8 FILLER_34_2184 ();
 sg13g2_decap_8 FILLER_34_2191 ();
 sg13g2_decap_4 FILLER_34_2198 ();
 sg13g2_decap_8 FILLER_34_2206 ();
 sg13g2_fill_2 FILLER_34_2213 ();
 sg13g2_fill_1 FILLER_34_2215 ();
 sg13g2_fill_2 FILLER_34_2230 ();
 sg13g2_fill_2 FILLER_34_2297 ();
 sg13g2_decap_4 FILLER_34_2339 ();
 sg13g2_fill_2 FILLER_34_2360 ();
 sg13g2_fill_1 FILLER_34_2362 ();
 sg13g2_decap_8 FILLER_34_2376 ();
 sg13g2_decap_4 FILLER_34_2383 ();
 sg13g2_fill_2 FILLER_34_2387 ();
 sg13g2_decap_8 FILLER_34_2397 ();
 sg13g2_fill_1 FILLER_34_2404 ();
 sg13g2_decap_8 FILLER_34_2409 ();
 sg13g2_decap_8 FILLER_34_2416 ();
 sg13g2_fill_2 FILLER_34_2423 ();
 sg13g2_decap_4 FILLER_34_2433 ();
 sg13g2_fill_2 FILLER_34_2441 ();
 sg13g2_fill_1 FILLER_34_2447 ();
 sg13g2_fill_2 FILLER_34_2460 ();
 sg13g2_fill_1 FILLER_34_2536 ();
 sg13g2_fill_1 FILLER_34_2541 ();
 sg13g2_decap_4 FILLER_34_2597 ();
 sg13g2_fill_1 FILLER_34_2601 ();
 sg13g2_fill_2 FILLER_34_2612 ();
 sg13g2_decap_8 FILLER_34_2640 ();
 sg13g2_decap_8 FILLER_34_2647 ();
 sg13g2_decap_8 FILLER_34_2654 ();
 sg13g2_decap_8 FILLER_34_2661 ();
 sg13g2_fill_2 FILLER_34_2668 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_2 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_30 ();
 sg13g2_decap_4 FILLER_35_37 ();
 sg13g2_fill_1 FILLER_35_41 ();
 sg13g2_decap_8 FILLER_35_46 ();
 sg13g2_fill_1 FILLER_35_105 ();
 sg13g2_fill_2 FILLER_35_112 ();
 sg13g2_fill_2 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_138 ();
 sg13g2_decap_4 FILLER_35_145 ();
 sg13g2_fill_2 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_166 ();
 sg13g2_fill_2 FILLER_35_173 ();
 sg13g2_fill_2 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_191 ();
 sg13g2_decap_8 FILLER_35_198 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_fill_1 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_225 ();
 sg13g2_fill_2 FILLER_35_231 ();
 sg13g2_fill_2 FILLER_35_237 ();
 sg13g2_fill_2 FILLER_35_243 ();
 sg13g2_fill_2 FILLER_35_254 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_334 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_fill_2 FILLER_35_373 ();
 sg13g2_decap_4 FILLER_35_379 ();
 sg13g2_fill_1 FILLER_35_388 ();
 sg13g2_decap_8 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_400 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_fill_2 FILLER_35_429 ();
 sg13g2_fill_2 FILLER_35_440 ();
 sg13g2_fill_2 FILLER_35_486 ();
 sg13g2_fill_2 FILLER_35_519 ();
 sg13g2_fill_2 FILLER_35_525 ();
 sg13g2_fill_2 FILLER_35_537 ();
 sg13g2_fill_2 FILLER_35_544 ();
 sg13g2_decap_4 FILLER_35_550 ();
 sg13g2_fill_1 FILLER_35_554 ();
 sg13g2_decap_4 FILLER_35_569 ();
 sg13g2_fill_1 FILLER_35_583 ();
 sg13g2_fill_1 FILLER_35_592 ();
 sg13g2_fill_1 FILLER_35_635 ();
 sg13g2_fill_2 FILLER_35_642 ();
 sg13g2_fill_1 FILLER_35_648 ();
 sg13g2_decap_4 FILLER_35_675 ();
 sg13g2_fill_2 FILLER_35_679 ();
 sg13g2_fill_1 FILLER_35_721 ();
 sg13g2_fill_1 FILLER_35_727 ();
 sg13g2_fill_1 FILLER_35_737 ();
 sg13g2_fill_2 FILLER_35_748 ();
 sg13g2_fill_2 FILLER_35_760 ();
 sg13g2_fill_2 FILLER_35_774 ();
 sg13g2_fill_1 FILLER_35_788 ();
 sg13g2_decap_4 FILLER_35_799 ();
 sg13g2_fill_2 FILLER_35_803 ();
 sg13g2_decap_4 FILLER_35_808 ();
 sg13g2_fill_2 FILLER_35_812 ();
 sg13g2_fill_2 FILLER_35_860 ();
 sg13g2_fill_1 FILLER_35_872 ();
 sg13g2_fill_1 FILLER_35_883 ();
 sg13g2_fill_1 FILLER_35_910 ();
 sg13g2_fill_1 FILLER_35_937 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_4 FILLER_35_966 ();
 sg13g2_decap_4 FILLER_35_974 ();
 sg13g2_fill_2 FILLER_35_1010 ();
 sg13g2_fill_1 FILLER_35_1012 ();
 sg13g2_decap_8 FILLER_35_1043 ();
 sg13g2_fill_2 FILLER_35_1050 ();
 sg13g2_fill_1 FILLER_35_1052 ();
 sg13g2_decap_8 FILLER_35_1069 ();
 sg13g2_fill_2 FILLER_35_1076 ();
 sg13g2_fill_1 FILLER_35_1099 ();
 sg13g2_decap_8 FILLER_35_1104 ();
 sg13g2_decap_8 FILLER_35_1111 ();
 sg13g2_fill_2 FILLER_35_1118 ();
 sg13g2_fill_2 FILLER_35_1133 ();
 sg13g2_fill_2 FILLER_35_1144 ();
 sg13g2_decap_8 FILLER_35_1175 ();
 sg13g2_decap_4 FILLER_35_1182 ();
 sg13g2_fill_1 FILLER_35_1186 ();
 sg13g2_decap_4 FILLER_35_1191 ();
 sg13g2_fill_1 FILLER_35_1230 ();
 sg13g2_fill_1 FILLER_35_1250 ();
 sg13g2_decap_8 FILLER_35_1286 ();
 sg13g2_fill_2 FILLER_35_1293 ();
 sg13g2_fill_2 FILLER_35_1299 ();
 sg13g2_fill_1 FILLER_35_1331 ();
 sg13g2_fill_2 FILLER_35_1360 ();
 sg13g2_fill_1 FILLER_35_1428 ();
 sg13g2_fill_1 FILLER_35_1435 ();
 sg13g2_decap_8 FILLER_35_1440 ();
 sg13g2_fill_2 FILLER_35_1447 ();
 sg13g2_fill_1 FILLER_35_1449 ();
 sg13g2_decap_4 FILLER_35_1461 ();
 sg13g2_fill_1 FILLER_35_1465 ();
 sg13g2_fill_1 FILLER_35_1472 ();
 sg13g2_fill_1 FILLER_35_1481 ();
 sg13g2_decap_8 FILLER_35_1493 ();
 sg13g2_fill_1 FILLER_35_1500 ();
 sg13g2_decap_4 FILLER_35_1506 ();
 sg13g2_decap_4 FILLER_35_1515 ();
 sg13g2_decap_4 FILLER_35_1524 ();
 sg13g2_fill_2 FILLER_35_1532 ();
 sg13g2_fill_1 FILLER_35_1534 ();
 sg13g2_fill_1 FILLER_35_1550 ();
 sg13g2_fill_1 FILLER_35_1561 ();
 sg13g2_fill_2 FILLER_35_1568 ();
 sg13g2_fill_1 FILLER_35_1576 ();
 sg13g2_fill_1 FILLER_35_1583 ();
 sg13g2_fill_1 FILLER_35_1588 ();
 sg13g2_fill_1 FILLER_35_1594 ();
 sg13g2_fill_2 FILLER_35_1605 ();
 sg13g2_fill_1 FILLER_35_1612 ();
 sg13g2_fill_1 FILLER_35_1618 ();
 sg13g2_fill_2 FILLER_35_1624 ();
 sg13g2_fill_2 FILLER_35_1631 ();
 sg13g2_fill_1 FILLER_35_1674 ();
 sg13g2_fill_1 FILLER_35_1696 ();
 sg13g2_fill_2 FILLER_35_1709 ();
 sg13g2_fill_1 FILLER_35_1737 ();
 sg13g2_fill_2 FILLER_35_1754 ();
 sg13g2_fill_2 FILLER_35_1791 ();
 sg13g2_fill_2 FILLER_35_1836 ();
 sg13g2_fill_1 FILLER_35_1838 ();
 sg13g2_decap_8 FILLER_35_1844 ();
 sg13g2_decap_8 FILLER_35_1881 ();
 sg13g2_fill_2 FILLER_35_1888 ();
 sg13g2_fill_1 FILLER_35_1890 ();
 sg13g2_fill_1 FILLER_35_1896 ();
 sg13g2_fill_2 FILLER_35_1923 ();
 sg13g2_decap_8 FILLER_35_1938 ();
 sg13g2_fill_1 FILLER_35_1975 ();
 sg13g2_fill_2 FILLER_35_2057 ();
 sg13g2_fill_1 FILLER_35_2067 ();
 sg13g2_fill_2 FILLER_35_2084 ();
 sg13g2_decap_8 FILLER_35_2096 ();
 sg13g2_decap_4 FILLER_35_2103 ();
 sg13g2_fill_1 FILLER_35_2123 ();
 sg13g2_fill_2 FILLER_35_2128 ();
 sg13g2_decap_8 FILLER_35_2134 ();
 sg13g2_decap_8 FILLER_35_2141 ();
 sg13g2_decap_8 FILLER_35_2148 ();
 sg13g2_fill_1 FILLER_35_2155 ();
 sg13g2_fill_2 FILLER_35_2177 ();
 sg13g2_fill_1 FILLER_35_2179 ();
 sg13g2_decap_8 FILLER_35_2194 ();
 sg13g2_fill_2 FILLER_35_2201 ();
 sg13g2_fill_2 FILLER_35_2211 ();
 sg13g2_fill_1 FILLER_35_2213 ();
 sg13g2_fill_1 FILLER_35_2240 ();
 sg13g2_fill_2 FILLER_35_2295 ();
 sg13g2_fill_1 FILLER_35_2297 ();
 sg13g2_fill_2 FILLER_35_2302 ();
 sg13g2_fill_1 FILLER_35_2304 ();
 sg13g2_fill_2 FILLER_35_2309 ();
 sg13g2_fill_2 FILLER_35_2327 ();
 sg13g2_fill_1 FILLER_35_2329 ();
 sg13g2_fill_2 FILLER_35_2355 ();
 sg13g2_decap_4 FILLER_35_2393 ();
 sg13g2_decap_4 FILLER_35_2428 ();
 sg13g2_fill_2 FILLER_35_2482 ();
 sg13g2_fill_2 FILLER_35_2492 ();
 sg13g2_decap_8 FILLER_35_2529 ();
 sg13g2_decap_8 FILLER_35_2536 ();
 sg13g2_fill_2 FILLER_35_2543 ();
 sg13g2_fill_1 FILLER_35_2545 ();
 sg13g2_decap_4 FILLER_35_2556 ();
 sg13g2_fill_2 FILLER_35_2560 ();
 sg13g2_decap_4 FILLER_35_2593 ();
 sg13g2_decap_8 FILLER_35_2641 ();
 sg13g2_decap_8 FILLER_35_2648 ();
 sg13g2_decap_8 FILLER_35_2655 ();
 sg13g2_decap_8 FILLER_35_2662 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_28 ();
 sg13g2_decap_4 FILLER_36_34 ();
 sg13g2_fill_1 FILLER_36_38 ();
 sg13g2_decap_4 FILLER_36_44 ();
 sg13g2_fill_2 FILLER_36_48 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_2 FILLER_36_71 ();
 sg13g2_decap_4 FILLER_36_103 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_1 FILLER_36_124 ();
 sg13g2_fill_2 FILLER_36_151 ();
 sg13g2_fill_2 FILLER_36_209 ();
 sg13g2_decap_4 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_249 ();
 sg13g2_decap_4 FILLER_36_256 ();
 sg13g2_fill_2 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_281 ();
 sg13g2_fill_1 FILLER_36_288 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_390 ();
 sg13g2_decap_8 FILLER_36_401 ();
 sg13g2_decap_4 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_433 ();
 sg13g2_fill_1 FILLER_36_440 ();
 sg13g2_fill_1 FILLER_36_450 ();
 sg13g2_fill_2 FILLER_36_456 ();
 sg13g2_fill_1 FILLER_36_487 ();
 sg13g2_fill_1 FILLER_36_498 ();
 sg13g2_fill_2 FILLER_36_516 ();
 sg13g2_fill_1 FILLER_36_528 ();
 sg13g2_fill_2 FILLER_36_555 ();
 sg13g2_fill_1 FILLER_36_557 ();
 sg13g2_fill_1 FILLER_36_649 ();
 sg13g2_fill_2 FILLER_36_680 ();
 sg13g2_fill_1 FILLER_36_682 ();
 sg13g2_fill_2 FILLER_36_700 ();
 sg13g2_fill_1 FILLER_36_707 ();
 sg13g2_fill_2 FILLER_36_713 ();
 sg13g2_fill_2 FILLER_36_719 ();
 sg13g2_fill_1 FILLER_36_822 ();
 sg13g2_fill_1 FILLER_36_853 ();
 sg13g2_fill_1 FILLER_36_890 ();
 sg13g2_fill_1 FILLER_36_912 ();
 sg13g2_fill_1 FILLER_36_918 ();
 sg13g2_fill_1 FILLER_36_923 ();
 sg13g2_fill_2 FILLER_36_934 ();
 sg13g2_fill_1 FILLER_36_936 ();
 sg13g2_decap_8 FILLER_36_963 ();
 sg13g2_decap_8 FILLER_36_970 ();
 sg13g2_fill_2 FILLER_36_977 ();
 sg13g2_fill_1 FILLER_36_983 ();
 sg13g2_fill_2 FILLER_36_1015 ();
 sg13g2_fill_1 FILLER_36_1022 ();
 sg13g2_fill_1 FILLER_36_1053 ();
 sg13g2_decap_8 FILLER_36_1101 ();
 sg13g2_decap_8 FILLER_36_1108 ();
 sg13g2_decap_8 FILLER_36_1115 ();
 sg13g2_fill_2 FILLER_36_1122 ();
 sg13g2_fill_1 FILLER_36_1124 ();
 sg13g2_fill_2 FILLER_36_1130 ();
 sg13g2_fill_1 FILLER_36_1132 ();
 sg13g2_decap_4 FILLER_36_1159 ();
 sg13g2_fill_1 FILLER_36_1163 ();
 sg13g2_decap_4 FILLER_36_1169 ();
 sg13g2_fill_1 FILLER_36_1173 ();
 sg13g2_decap_8 FILLER_36_1178 ();
 sg13g2_fill_2 FILLER_36_1185 ();
 sg13g2_decap_8 FILLER_36_1223 ();
 sg13g2_decap_4 FILLER_36_1230 ();
 sg13g2_fill_1 FILLER_36_1234 ();
 sg13g2_decap_4 FILLER_36_1286 ();
 sg13g2_fill_2 FILLER_36_1290 ();
 sg13g2_decap_8 FILLER_36_1305 ();
 sg13g2_decap_8 FILLER_36_1312 ();
 sg13g2_fill_2 FILLER_36_1329 ();
 sg13g2_fill_1 FILLER_36_1331 ();
 sg13g2_fill_2 FILLER_36_1345 ();
 sg13g2_fill_1 FILLER_36_1347 ();
 sg13g2_fill_1 FILLER_36_1358 ();
 sg13g2_decap_8 FILLER_36_1395 ();
 sg13g2_fill_1 FILLER_36_1402 ();
 sg13g2_fill_2 FILLER_36_1436 ();
 sg13g2_fill_1 FILLER_36_1454 ();
 sg13g2_fill_1 FILLER_36_1462 ();
 sg13g2_decap_4 FILLER_36_1482 ();
 sg13g2_fill_2 FILLER_36_1486 ();
 sg13g2_decap_8 FILLER_36_1505 ();
 sg13g2_fill_2 FILLER_36_1512 ();
 sg13g2_fill_1 FILLER_36_1514 ();
 sg13g2_decap_4 FILLER_36_1520 ();
 sg13g2_fill_2 FILLER_36_1544 ();
 sg13g2_fill_2 FILLER_36_1551 ();
 sg13g2_fill_2 FILLER_36_1558 ();
 sg13g2_fill_2 FILLER_36_1565 ();
 sg13g2_fill_2 FILLER_36_1573 ();
 sg13g2_fill_1 FILLER_36_1575 ();
 sg13g2_fill_2 FILLER_36_1581 ();
 sg13g2_fill_1 FILLER_36_1592 ();
 sg13g2_fill_1 FILLER_36_1603 ();
 sg13g2_fill_2 FILLER_36_1683 ();
 sg13g2_fill_2 FILLER_36_1688 ();
 sg13g2_decap_4 FILLER_36_1731 ();
 sg13g2_fill_2 FILLER_36_1735 ();
 sg13g2_decap_8 FILLER_36_1757 ();
 sg13g2_decap_4 FILLER_36_1764 ();
 sg13g2_fill_1 FILLER_36_1768 ();
 sg13g2_fill_1 FILLER_36_1799 ();
 sg13g2_fill_2 FILLER_36_1843 ();
 sg13g2_fill_1 FILLER_36_1845 ();
 sg13g2_fill_1 FILLER_36_1859 ();
 sg13g2_decap_8 FILLER_36_1868 ();
 sg13g2_decap_8 FILLER_36_1875 ();
 sg13g2_decap_8 FILLER_36_1882 ();
 sg13g2_fill_1 FILLER_36_1889 ();
 sg13g2_fill_1 FILLER_36_1895 ();
 sg13g2_fill_1 FILLER_36_1900 ();
 sg13g2_decap_4 FILLER_36_1905 ();
 sg13g2_fill_2 FILLER_36_1909 ();
 sg13g2_decap_8 FILLER_36_1924 ();
 sg13g2_decap_8 FILLER_36_1931 ();
 sg13g2_fill_2 FILLER_36_1951 ();
 sg13g2_fill_1 FILLER_36_1953 ();
 sg13g2_fill_1 FILLER_36_2001 ();
 sg13g2_fill_1 FILLER_36_2011 ();
 sg13g2_fill_1 FILLER_36_2033 ();
 sg13g2_decap_8 FILLER_36_2060 ();
 sg13g2_fill_1 FILLER_36_2081 ();
 sg13g2_decap_4 FILLER_36_2116 ();
 sg13g2_fill_1 FILLER_36_2120 ();
 sg13g2_decap_8 FILLER_36_2131 ();
 sg13g2_fill_1 FILLER_36_2138 ();
 sg13g2_decap_4 FILLER_36_2160 ();
 sg13g2_fill_2 FILLER_36_2164 ();
 sg13g2_fill_2 FILLER_36_2180 ();
 sg13g2_fill_2 FILLER_36_2288 ();
 sg13g2_fill_1 FILLER_36_2290 ();
 sg13g2_fill_2 FILLER_36_2338 ();
 sg13g2_fill_2 FILLER_36_2409 ();
 sg13g2_fill_1 FILLER_36_2411 ();
 sg13g2_fill_2 FILLER_36_2422 ();
 sg13g2_fill_2 FILLER_36_2434 ();
 sg13g2_fill_1 FILLER_36_2446 ();
 sg13g2_fill_2 FILLER_36_2483 ();
 sg13g2_fill_2 FILLER_36_2516 ();
 sg13g2_fill_1 FILLER_36_2518 ();
 sg13g2_decap_4 FILLER_36_2540 ();
 sg13g2_fill_2 FILLER_36_2544 ();
 sg13g2_decap_4 FILLER_36_2556 ();
 sg13g2_fill_2 FILLER_36_2560 ();
 sg13g2_decap_4 FILLER_36_2588 ();
 sg13g2_decap_8 FILLER_36_2628 ();
 sg13g2_decap_8 FILLER_36_2635 ();
 sg13g2_decap_8 FILLER_36_2642 ();
 sg13g2_decap_8 FILLER_36_2649 ();
 sg13g2_decap_8 FILLER_36_2656 ();
 sg13g2_decap_8 FILLER_36_2663 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_7 ();
 sg13g2_fill_1 FILLER_37_39 ();
 sg13g2_fill_2 FILLER_37_58 ();
 sg13g2_fill_1 FILLER_37_60 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_fill_1 FILLER_37_91 ();
 sg13g2_fill_1 FILLER_37_102 ();
 sg13g2_fill_2 FILLER_37_107 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_2 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_159 ();
 sg13g2_decap_4 FILLER_37_174 ();
 sg13g2_fill_1 FILLER_37_178 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_decap_4 FILLER_37_194 ();
 sg13g2_decap_8 FILLER_37_212 ();
 sg13g2_decap_4 FILLER_37_219 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_fill_2 FILLER_37_235 ();
 sg13g2_fill_1 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_fill_2 FILLER_37_248 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_fill_2 FILLER_37_266 ();
 sg13g2_decap_4 FILLER_37_273 ();
 sg13g2_decap_4 FILLER_37_285 ();
 sg13g2_fill_1 FILLER_37_319 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_344 ();
 sg13g2_decap_4 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_461 ();
 sg13g2_fill_1 FILLER_37_469 ();
 sg13g2_fill_1 FILLER_37_475 ();
 sg13g2_fill_2 FILLER_37_486 ();
 sg13g2_fill_1 FILLER_37_494 ();
 sg13g2_fill_1 FILLER_37_499 ();
 sg13g2_fill_2 FILLER_37_504 ();
 sg13g2_decap_8 FILLER_37_530 ();
 sg13g2_fill_1 FILLER_37_537 ();
 sg13g2_decap_4 FILLER_37_547 ();
 sg13g2_fill_1 FILLER_37_587 ();
 sg13g2_fill_2 FILLER_37_602 ();
 sg13g2_fill_1 FILLER_37_604 ();
 sg13g2_fill_2 FILLER_37_618 ();
 sg13g2_fill_2 FILLER_37_655 ();
 sg13g2_decap_4 FILLER_37_661 ();
 sg13g2_fill_1 FILLER_37_665 ();
 sg13g2_decap_4 FILLER_37_671 ();
 sg13g2_fill_1 FILLER_37_675 ();
 sg13g2_fill_1 FILLER_37_739 ();
 sg13g2_fill_1 FILLER_37_799 ();
 sg13g2_fill_2 FILLER_37_804 ();
 sg13g2_fill_1 FILLER_37_806 ();
 sg13g2_decap_4 FILLER_37_843 ();
 sg13g2_fill_1 FILLER_37_883 ();
 sg13g2_decap_8 FILLER_37_888 ();
 sg13g2_fill_2 FILLER_37_895 ();
 sg13g2_fill_1 FILLER_37_907 ();
 sg13g2_decap_8 FILLER_37_952 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_fill_1 FILLER_37_973 ();
 sg13g2_fill_1 FILLER_37_995 ();
 sg13g2_fill_1 FILLER_37_1000 ();
 sg13g2_fill_1 FILLER_37_1006 ();
 sg13g2_fill_1 FILLER_37_1011 ();
 sg13g2_fill_2 FILLER_37_1022 ();
 sg13g2_fill_2 FILLER_37_1045 ();
 sg13g2_fill_1 FILLER_37_1135 ();
 sg13g2_fill_2 FILLER_37_1144 ();
 sg13g2_fill_2 FILLER_37_1182 ();
 sg13g2_fill_2 FILLER_37_1194 ();
 sg13g2_decap_4 FILLER_37_1226 ();
 sg13g2_fill_2 FILLER_37_1233 ();
 sg13g2_fill_2 FILLER_37_1300 ();
 sg13g2_decap_8 FILLER_37_1358 ();
 sg13g2_decap_8 FILLER_37_1365 ();
 sg13g2_decap_8 FILLER_37_1376 ();
 sg13g2_fill_2 FILLER_37_1383 ();
 sg13g2_fill_1 FILLER_37_1385 ();
 sg13g2_decap_4 FILLER_37_1406 ();
 sg13g2_fill_2 FILLER_37_1410 ();
 sg13g2_fill_1 FILLER_37_1417 ();
 sg13g2_fill_2 FILLER_37_1424 ();
 sg13g2_fill_1 FILLER_37_1433 ();
 sg13g2_fill_1 FILLER_37_1444 ();
 sg13g2_decap_4 FILLER_37_1474 ();
 sg13g2_fill_1 FILLER_37_1484 ();
 sg13g2_fill_2 FILLER_37_1498 ();
 sg13g2_fill_1 FILLER_37_1531 ();
 sg13g2_fill_1 FILLER_37_1537 ();
 sg13g2_fill_2 FILLER_37_1543 ();
 sg13g2_fill_2 FILLER_37_1560 ();
 sg13g2_fill_1 FILLER_37_1567 ();
 sg13g2_fill_2 FILLER_37_1578 ();
 sg13g2_fill_2 FILLER_37_1585 ();
 sg13g2_fill_1 FILLER_37_1614 ();
 sg13g2_decap_8 FILLER_37_1632 ();
 sg13g2_fill_2 FILLER_37_1710 ();
 sg13g2_decap_4 FILLER_37_1734 ();
 sg13g2_fill_1 FILLER_37_1738 ();
 sg13g2_decap_8 FILLER_37_1781 ();
 sg13g2_decap_4 FILLER_37_1788 ();
 sg13g2_fill_1 FILLER_37_1792 ();
 sg13g2_decap_8 FILLER_37_1797 ();
 sg13g2_fill_2 FILLER_37_1804 ();
 sg13g2_decap_8 FILLER_37_1817 ();
 sg13g2_decap_8 FILLER_37_1824 ();
 sg13g2_decap_8 FILLER_37_1831 ();
 sg13g2_decap_8 FILLER_37_1838 ();
 sg13g2_decap_8 FILLER_37_1845 ();
 sg13g2_decap_4 FILLER_37_1852 ();
 sg13g2_decap_8 FILLER_37_1861 ();
 sg13g2_decap_8 FILLER_37_1868 ();
 sg13g2_decap_8 FILLER_37_1875 ();
 sg13g2_fill_1 FILLER_37_1886 ();
 sg13g2_fill_1 FILLER_37_1915 ();
 sg13g2_fill_2 FILLER_37_1920 ();
 sg13g2_decap_8 FILLER_37_1930 ();
 sg13g2_decap_8 FILLER_37_1937 ();
 sg13g2_fill_2 FILLER_37_1944 ();
 sg13g2_fill_1 FILLER_37_1946 ();
 sg13g2_fill_2 FILLER_37_1973 ();
 sg13g2_fill_1 FILLER_37_1995 ();
 sg13g2_fill_2 FILLER_37_2032 ();
 sg13g2_fill_2 FILLER_37_2073 ();
 sg13g2_fill_1 FILLER_37_2075 ();
 sg13g2_fill_1 FILLER_37_2081 ();
 sg13g2_fill_1 FILLER_37_2115 ();
 sg13g2_decap_8 FILLER_37_2152 ();
 sg13g2_fill_2 FILLER_37_2159 ();
 sg13g2_fill_1 FILLER_37_2161 ();
 sg13g2_fill_2 FILLER_37_2209 ();
 sg13g2_fill_2 FILLER_37_2241 ();
 sg13g2_fill_1 FILLER_37_2276 ();
 sg13g2_decap_8 FILLER_37_2313 ();
 sg13g2_decap_8 FILLER_37_2320 ();
 sg13g2_fill_1 FILLER_37_2327 ();
 sg13g2_decap_4 FILLER_37_2379 ();
 sg13g2_fill_1 FILLER_37_2383 ();
 sg13g2_fill_2 FILLER_37_2414 ();
 sg13g2_fill_1 FILLER_37_2416 ();
 sg13g2_fill_2 FILLER_37_2443 ();
 sg13g2_fill_1 FILLER_37_2470 ();
 sg13g2_decap_8 FILLER_37_2501 ();
 sg13g2_decap_4 FILLER_37_2508 ();
 sg13g2_fill_1 FILLER_37_2512 ();
 sg13g2_decap_4 FILLER_37_2523 ();
 sg13g2_fill_1 FILLER_37_2527 ();
 sg13g2_decap_8 FILLER_37_2580 ();
 sg13g2_decap_4 FILLER_37_2587 ();
 sg13g2_fill_1 FILLER_37_2591 ();
 sg13g2_decap_8 FILLER_37_2617 ();
 sg13g2_decap_8 FILLER_37_2624 ();
 sg13g2_decap_8 FILLER_37_2631 ();
 sg13g2_decap_8 FILLER_37_2638 ();
 sg13g2_decap_8 FILLER_37_2645 ();
 sg13g2_decap_8 FILLER_37_2652 ();
 sg13g2_decap_8 FILLER_37_2659 ();
 sg13g2_decap_4 FILLER_37_2666 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_fill_2 FILLER_38_25 ();
 sg13g2_fill_1 FILLER_38_32 ();
 sg13g2_fill_1 FILLER_38_37 ();
 sg13g2_decap_4 FILLER_38_68 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_fill_2 FILLER_38_77 ();
 sg13g2_fill_1 FILLER_38_79 ();
 sg13g2_fill_2 FILLER_38_106 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_fill_2 FILLER_38_126 ();
 sg13g2_fill_1 FILLER_38_137 ();
 sg13g2_fill_1 FILLER_38_142 ();
 sg13g2_fill_1 FILLER_38_169 ();
 sg13g2_fill_1 FILLER_38_200 ();
 sg13g2_fill_2 FILLER_38_253 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_decap_4 FILLER_38_287 ();
 sg13g2_fill_2 FILLER_38_301 ();
 sg13g2_decap_4 FILLER_38_308 ();
 sg13g2_fill_2 FILLER_38_316 ();
 sg13g2_fill_1 FILLER_38_318 ();
 sg13g2_decap_4 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_337 ();
 sg13g2_fill_2 FILLER_38_344 ();
 sg13g2_fill_1 FILLER_38_346 ();
 sg13g2_decap_4 FILLER_38_351 ();
 sg13g2_fill_1 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_374 ();
 sg13g2_decap_8 FILLER_38_381 ();
 sg13g2_decap_8 FILLER_38_388 ();
 sg13g2_fill_1 FILLER_38_395 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_412 ();
 sg13g2_decap_4 FILLER_38_419 ();
 sg13g2_fill_2 FILLER_38_423 ();
 sg13g2_fill_2 FILLER_38_429 ();
 sg13g2_fill_2 FILLER_38_447 ();
 sg13g2_fill_1 FILLER_38_449 ();
 sg13g2_decap_8 FILLER_38_465 ();
 sg13g2_fill_1 FILLER_38_485 ();
 sg13g2_fill_1 FILLER_38_505 ();
 sg13g2_fill_1 FILLER_38_514 ();
 sg13g2_decap_4 FILLER_38_522 ();
 sg13g2_decap_4 FILLER_38_530 ();
 sg13g2_fill_1 FILLER_38_534 ();
 sg13g2_fill_2 FILLER_38_539 ();
 sg13g2_fill_1 FILLER_38_541 ();
 sg13g2_decap_4 FILLER_38_552 ();
 sg13g2_fill_1 FILLER_38_556 ();
 sg13g2_fill_2 FILLER_38_566 ();
 sg13g2_fill_1 FILLER_38_568 ();
 sg13g2_fill_2 FILLER_38_583 ();
 sg13g2_fill_2 FILLER_38_611 ();
 sg13g2_fill_1 FILLER_38_613 ();
 sg13g2_fill_1 FILLER_38_629 ();
 sg13g2_decap_4 FILLER_38_638 ();
 sg13g2_fill_1 FILLER_38_642 ();
 sg13g2_decap_4 FILLER_38_649 ();
 sg13g2_fill_2 FILLER_38_653 ();
 sg13g2_decap_8 FILLER_38_661 ();
 sg13g2_fill_1 FILLER_38_668 ();
 sg13g2_fill_1 FILLER_38_674 ();
 sg13g2_fill_2 FILLER_38_684 ();
 sg13g2_fill_1 FILLER_38_696 ();
 sg13g2_fill_1 FILLER_38_701 ();
 sg13g2_fill_1 FILLER_38_706 ();
 sg13g2_fill_1 FILLER_38_711 ();
 sg13g2_fill_1 FILLER_38_717 ();
 sg13g2_fill_1 FILLER_38_722 ();
 sg13g2_fill_2 FILLER_38_776 ();
 sg13g2_fill_2 FILLER_38_784 ();
 sg13g2_decap_4 FILLER_38_789 ();
 sg13g2_decap_4 FILLER_38_819 ();
 sg13g2_decap_4 FILLER_38_827 ();
 sg13g2_fill_1 FILLER_38_831 ();
 sg13g2_fill_2 FILLER_38_836 ();
 sg13g2_decap_8 FILLER_38_848 ();
 sg13g2_decap_8 FILLER_38_855 ();
 sg13g2_fill_1 FILLER_38_862 ();
 sg13g2_fill_2 FILLER_38_867 ();
 sg13g2_fill_1 FILLER_38_869 ();
 sg13g2_decap_8 FILLER_38_874 ();
 sg13g2_fill_2 FILLER_38_881 ();
 sg13g2_decap_4 FILLER_38_887 ();
 sg13g2_fill_1 FILLER_38_891 ();
 sg13g2_fill_1 FILLER_38_909 ();
 sg13g2_decap_4 FILLER_38_936 ();
 sg13g2_fill_1 FILLER_38_940 ();
 sg13g2_decap_8 FILLER_38_982 ();
 sg13g2_decap_8 FILLER_38_999 ();
 sg13g2_fill_2 FILLER_38_1010 ();
 sg13g2_fill_2 FILLER_38_1017 ();
 sg13g2_fill_2 FILLER_38_1023 ();
 sg13g2_fill_2 FILLER_38_1034 ();
 sg13g2_fill_1 FILLER_38_1086 ();
 sg13g2_decap_4 FILLER_38_1123 ();
 sg13g2_fill_1 FILLER_38_1153 ();
 sg13g2_fill_1 FILLER_38_1210 ();
 sg13g2_fill_2 FILLER_38_1215 ();
 sg13g2_fill_1 FILLER_38_1217 ();
 sg13g2_fill_2 FILLER_38_1242 ();
 sg13g2_fill_2 FILLER_38_1248 ();
 sg13g2_fill_1 FILLER_38_1270 ();
 sg13g2_decap_8 FILLER_38_1321 ();
 sg13g2_decap_8 FILLER_38_1328 ();
 sg13g2_decap_4 FILLER_38_1335 ();
 sg13g2_decap_4 FILLER_38_1343 ();
 sg13g2_fill_1 FILLER_38_1347 ();
 sg13g2_decap_4 FILLER_38_1388 ();
 sg13g2_fill_2 FILLER_38_1392 ();
 sg13g2_decap_4 FILLER_38_1404 ();
 sg13g2_fill_1 FILLER_38_1430 ();
 sg13g2_decap_4 FILLER_38_1449 ();
 sg13g2_fill_1 FILLER_38_1453 ();
 sg13g2_fill_2 FILLER_38_1468 ();
 sg13g2_decap_8 FILLER_38_1475 ();
 sg13g2_fill_1 FILLER_38_1482 ();
 sg13g2_decap_8 FILLER_38_1488 ();
 sg13g2_decap_4 FILLER_38_1495 ();
 sg13g2_fill_2 FILLER_38_1499 ();
 sg13g2_fill_1 FILLER_38_1512 ();
 sg13g2_fill_1 FILLER_38_1541 ();
 sg13g2_fill_1 FILLER_38_1563 ();
 sg13g2_decap_8 FILLER_38_1579 ();
 sg13g2_decap_8 FILLER_38_1586 ();
 sg13g2_decap_8 FILLER_38_1593 ();
 sg13g2_fill_1 FILLER_38_1600 ();
 sg13g2_decap_8 FILLER_38_1605 ();
 sg13g2_decap_4 FILLER_38_1612 ();
 sg13g2_fill_1 FILLER_38_1616 ();
 sg13g2_fill_1 FILLER_38_1649 ();
 sg13g2_fill_1 FILLER_38_1684 ();
 sg13g2_fill_2 FILLER_38_1738 ();
 sg13g2_fill_2 FILLER_38_1794 ();
 sg13g2_fill_2 FILLER_38_1800 ();
 sg13g2_decap_8 FILLER_38_1812 ();
 sg13g2_decap_8 FILLER_38_1819 ();
 sg13g2_decap_8 FILLER_38_1826 ();
 sg13g2_decap_8 FILLER_38_1833 ();
 sg13g2_decap_4 FILLER_38_1840 ();
 sg13g2_fill_1 FILLER_38_1844 ();
 sg13g2_fill_1 FILLER_38_1865 ();
 sg13g2_fill_1 FILLER_38_1871 ();
 sg13g2_fill_1 FILLER_38_1877 ();
 sg13g2_fill_2 FILLER_38_1893 ();
 sg13g2_fill_1 FILLER_38_1895 ();
 sg13g2_fill_2 FILLER_38_1928 ();
 sg13g2_fill_1 FILLER_38_1930 ();
 sg13g2_fill_2 FILLER_38_1936 ();
 sg13g2_fill_1 FILLER_38_1938 ();
 sg13g2_decap_4 FILLER_38_1949 ();
 sg13g2_decap_8 FILLER_38_1957 ();
 sg13g2_decap_8 FILLER_38_1964 ();
 sg13g2_decap_4 FILLER_38_1971 ();
 sg13g2_fill_2 FILLER_38_1975 ();
 sg13g2_decap_4 FILLER_38_2015 ();
 sg13g2_fill_2 FILLER_38_2027 ();
 sg13g2_fill_1 FILLER_38_2041 ();
 sg13g2_fill_1 FILLER_38_2064 ();
 sg13g2_fill_1 FILLER_38_2091 ();
 sg13g2_fill_1 FILLER_38_2135 ();
 sg13g2_decap_8 FILLER_38_2162 ();
 sg13g2_decap_8 FILLER_38_2169 ();
 sg13g2_decap_4 FILLER_38_2176 ();
 sg13g2_fill_1 FILLER_38_2180 ();
 sg13g2_decap_8 FILLER_38_2184 ();
 sg13g2_decap_4 FILLER_38_2191 ();
 sg13g2_fill_1 FILLER_38_2229 ();
 sg13g2_fill_2 FILLER_38_2245 ();
 sg13g2_fill_1 FILLER_38_2358 ();
 sg13g2_decap_4 FILLER_38_2466 ();
 sg13g2_fill_1 FILLER_38_2470 ();
 sg13g2_decap_4 FILLER_38_2543 ();
 sg13g2_fill_2 FILLER_38_2547 ();
 sg13g2_fill_2 FILLER_38_2575 ();
 sg13g2_fill_1 FILLER_38_2577 ();
 sg13g2_decap_8 FILLER_38_2591 ();
 sg13g2_decap_8 FILLER_38_2628 ();
 sg13g2_decap_8 FILLER_38_2635 ();
 sg13g2_decap_8 FILLER_38_2642 ();
 sg13g2_decap_8 FILLER_38_2649 ();
 sg13g2_decap_8 FILLER_38_2656 ();
 sg13g2_decap_8 FILLER_38_2663 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_51 ();
 sg13g2_decap_4 FILLER_39_62 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_fill_2 FILLER_39_77 ();
 sg13g2_fill_1 FILLER_39_131 ();
 sg13g2_decap_8 FILLER_39_137 ();
 sg13g2_decap_4 FILLER_39_144 ();
 sg13g2_decap_4 FILLER_39_174 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_decap_4 FILLER_39_183 ();
 sg13g2_decap_4 FILLER_39_213 ();
 sg13g2_fill_2 FILLER_39_221 ();
 sg13g2_fill_1 FILLER_39_233 ();
 sg13g2_fill_1 FILLER_39_238 ();
 sg13g2_fill_2 FILLER_39_265 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_277 ();
 sg13g2_fill_2 FILLER_39_284 ();
 sg13g2_fill_2 FILLER_39_295 ();
 sg13g2_fill_1 FILLER_39_297 ();
 sg13g2_fill_2 FILLER_39_310 ();
 sg13g2_fill_1 FILLER_39_312 ();
 sg13g2_decap_4 FILLER_39_318 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_328 ();
 sg13g2_decap_8 FILLER_39_333 ();
 sg13g2_decap_8 FILLER_39_340 ();
 sg13g2_fill_1 FILLER_39_347 ();
 sg13g2_fill_2 FILLER_39_384 ();
 sg13g2_decap_8 FILLER_39_397 ();
 sg13g2_fill_2 FILLER_39_404 ();
 sg13g2_decap_4 FILLER_39_442 ();
 sg13g2_fill_2 FILLER_39_446 ();
 sg13g2_fill_2 FILLER_39_461 ();
 sg13g2_fill_1 FILLER_39_463 ();
 sg13g2_decap_4 FILLER_39_490 ();
 sg13g2_fill_2 FILLER_39_494 ();
 sg13g2_decap_8 FILLER_39_526 ();
 sg13g2_decap_4 FILLER_39_533 ();
 sg13g2_fill_2 FILLER_39_537 ();
 sg13g2_decap_4 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_566 ();
 sg13g2_decap_4 FILLER_39_573 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_fill_1 FILLER_39_610 ();
 sg13g2_decap_8 FILLER_39_616 ();
 sg13g2_decap_8 FILLER_39_623 ();
 sg13g2_fill_2 FILLER_39_630 ();
 sg13g2_fill_2 FILLER_39_640 ();
 sg13g2_decap_8 FILLER_39_650 ();
 sg13g2_fill_1 FILLER_39_668 ();
 sg13g2_fill_2 FILLER_39_691 ();
 sg13g2_fill_1 FILLER_39_693 ();
 sg13g2_decap_4 FILLER_39_706 ();
 sg13g2_fill_1 FILLER_39_715 ();
 sg13g2_fill_1 FILLER_39_742 ();
 sg13g2_decap_8 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_820 ();
 sg13g2_decap_8 FILLER_39_827 ();
 sg13g2_decap_4 FILLER_39_834 ();
 sg13g2_fill_2 FILLER_39_838 ();
 sg13g2_decap_4 FILLER_39_844 ();
 sg13g2_fill_1 FILLER_39_848 ();
 sg13g2_decap_8 FILLER_39_852 ();
 sg13g2_decap_8 FILLER_39_859 ();
 sg13g2_decap_4 FILLER_39_870 ();
 sg13g2_fill_2 FILLER_39_874 ();
 sg13g2_fill_1 FILLER_39_880 ();
 sg13g2_fill_2 FILLER_39_941 ();
 sg13g2_decap_8 FILLER_39_979 ();
 sg13g2_decap_8 FILLER_39_986 ();
 sg13g2_fill_2 FILLER_39_993 ();
 sg13g2_decap_8 FILLER_39_1025 ();
 sg13g2_decap_8 FILLER_39_1058 ();
 sg13g2_fill_1 FILLER_39_1065 ();
 sg13g2_decap_4 FILLER_39_1070 ();
 sg13g2_fill_1 FILLER_39_1074 ();
 sg13g2_fill_2 FILLER_39_1079 ();
 sg13g2_fill_1 FILLER_39_1081 ();
 sg13g2_fill_1 FILLER_39_1107 ();
 sg13g2_decap_8 FILLER_39_1112 ();
 sg13g2_decap_4 FILLER_39_1119 ();
 sg13g2_fill_1 FILLER_39_1123 ();
 sg13g2_fill_2 FILLER_39_1138 ();
 sg13g2_decap_4 FILLER_39_1144 ();
 sg13g2_fill_2 FILLER_39_1148 ();
 sg13g2_fill_2 FILLER_39_1154 ();
 sg13g2_decap_4 FILLER_39_1166 ();
 sg13g2_fill_1 FILLER_39_1170 ();
 sg13g2_decap_4 FILLER_39_1175 ();
 sg13g2_fill_2 FILLER_39_1213 ();
 sg13g2_fill_1 FILLER_39_1232 ();
 sg13g2_fill_1 FILLER_39_1270 ();
 sg13g2_fill_2 FILLER_39_1293 ();
 sg13g2_decap_8 FILLER_39_1331 ();
 sg13g2_decap_8 FILLER_39_1338 ();
 sg13g2_decap_8 FILLER_39_1345 ();
 sg13g2_decap_8 FILLER_39_1352 ();
 sg13g2_decap_8 FILLER_39_1359 ();
 sg13g2_fill_1 FILLER_39_1370 ();
 sg13g2_decap_8 FILLER_39_1401 ();
 sg13g2_decap_8 FILLER_39_1408 ();
 sg13g2_decap_4 FILLER_39_1415 ();
 sg13g2_fill_2 FILLER_39_1425 ();
 sg13g2_fill_2 FILLER_39_1432 ();
 sg13g2_fill_1 FILLER_39_1434 ();
 sg13g2_fill_2 FILLER_39_1441 ();
 sg13g2_fill_1 FILLER_39_1443 ();
 sg13g2_fill_1 FILLER_39_1449 ();
 sg13g2_decap_8 FILLER_39_1460 ();
 sg13g2_decap_4 FILLER_39_1467 ();
 sg13g2_fill_1 FILLER_39_1471 ();
 sg13g2_fill_2 FILLER_39_1491 ();
 sg13g2_fill_2 FILLER_39_1498 ();
 sg13g2_fill_1 FILLER_39_1500 ();
 sg13g2_decap_4 FILLER_39_1504 ();
 sg13g2_fill_1 FILLER_39_1508 ();
 sg13g2_fill_2 FILLER_39_1523 ();
 sg13g2_fill_1 FILLER_39_1525 ();
 sg13g2_fill_1 FILLER_39_1589 ();
 sg13g2_decap_4 FILLER_39_1594 ();
 sg13g2_fill_2 FILLER_39_1610 ();
 sg13g2_fill_1 FILLER_39_1612 ();
 sg13g2_fill_2 FILLER_39_1627 ();
 sg13g2_fill_1 FILLER_39_1629 ();
 sg13g2_fill_2 FILLER_39_1640 ();
 sg13g2_fill_2 FILLER_39_1657 ();
 sg13g2_fill_2 FILLER_39_1663 ();
 sg13g2_decap_8 FILLER_39_1669 ();
 sg13g2_decap_8 FILLER_39_1676 ();
 sg13g2_fill_1 FILLER_39_1687 ();
 sg13g2_decap_8 FILLER_39_1737 ();
 sg13g2_fill_2 FILLER_39_1744 ();
 sg13g2_decap_8 FILLER_39_1759 ();
 sg13g2_fill_2 FILLER_39_1766 ();
 sg13g2_decap_8 FILLER_39_1812 ();
 sg13g2_decap_8 FILLER_39_1819 ();
 sg13g2_decap_4 FILLER_39_1826 ();
 sg13g2_fill_1 FILLER_39_1870 ();
 sg13g2_fill_1 FILLER_39_1876 ();
 sg13g2_fill_1 FILLER_39_1890 ();
 sg13g2_fill_1 FILLER_39_1896 ();
 sg13g2_fill_1 FILLER_39_1921 ();
 sg13g2_fill_2 FILLER_39_1932 ();
 sg13g2_fill_1 FILLER_39_1939 ();
 sg13g2_fill_1 FILLER_39_1944 ();
 sg13g2_fill_1 FILLER_39_1949 ();
 sg13g2_fill_2 FILLER_39_1958 ();
 sg13g2_decap_4 FILLER_39_1968 ();
 sg13g2_fill_1 FILLER_39_1972 ();
 sg13g2_decap_8 FILLER_39_1977 ();
 sg13g2_fill_1 FILLER_39_1991 ();
 sg13g2_fill_2 FILLER_39_1999 ();
 sg13g2_decap_8 FILLER_39_2008 ();
 sg13g2_decap_8 FILLER_39_2015 ();
 sg13g2_fill_2 FILLER_39_2056 ();
 sg13g2_fill_1 FILLER_39_2094 ();
 sg13g2_decap_8 FILLER_39_2137 ();
 sg13g2_fill_1 FILLER_39_2144 ();
 sg13g2_decap_4 FILLER_39_2149 ();
 sg13g2_fill_1 FILLER_39_2153 ();
 sg13g2_decap_4 FILLER_39_2158 ();
 sg13g2_fill_1 FILLER_39_2185 ();
 sg13g2_fill_2 FILLER_39_2212 ();
 sg13g2_fill_1 FILLER_39_2214 ();
 sg13g2_decap_8 FILLER_39_2241 ();
 sg13g2_decap_4 FILLER_39_2314 ();
 sg13g2_fill_1 FILLER_39_2323 ();
 sg13g2_fill_2 FILLER_39_2328 ();
 sg13g2_fill_1 FILLER_39_2330 ();
 sg13g2_fill_1 FILLER_39_2340 ();
 sg13g2_fill_2 FILLER_39_2364 ();
 sg13g2_fill_1 FILLER_39_2370 ();
 sg13g2_decap_8 FILLER_39_2401 ();
 sg13g2_fill_2 FILLER_39_2408 ();
 sg13g2_fill_2 FILLER_39_2422 ();
 sg13g2_fill_1 FILLER_39_2424 ();
 sg13g2_fill_1 FILLER_39_2441 ();
 sg13g2_decap_8 FILLER_39_2468 ();
 sg13g2_fill_2 FILLER_39_2475 ();
 sg13g2_fill_1 FILLER_39_2477 ();
 sg13g2_fill_2 FILLER_39_2495 ();
 sg13g2_fill_2 FILLER_39_2521 ();
 sg13g2_fill_1 FILLER_39_2523 ();
 sg13g2_decap_8 FILLER_39_2528 ();
 sg13g2_decap_4 FILLER_39_2539 ();
 sg13g2_fill_2 FILLER_39_2557 ();
 sg13g2_fill_1 FILLER_39_2559 ();
 sg13g2_decap_8 FILLER_39_2564 ();
 sg13g2_decap_8 FILLER_39_2571 ();
 sg13g2_decap_8 FILLER_39_2578 ();
 sg13g2_decap_8 FILLER_39_2585 ();
 sg13g2_decap_8 FILLER_39_2592 ();
 sg13g2_decap_8 FILLER_39_2599 ();
 sg13g2_decap_8 FILLER_39_2606 ();
 sg13g2_decap_8 FILLER_39_2613 ();
 sg13g2_decap_8 FILLER_39_2620 ();
 sg13g2_decap_8 FILLER_39_2627 ();
 sg13g2_decap_8 FILLER_39_2634 ();
 sg13g2_decap_8 FILLER_39_2641 ();
 sg13g2_decap_8 FILLER_39_2648 ();
 sg13g2_decap_8 FILLER_39_2655 ();
 sg13g2_decap_8 FILLER_39_2662 ();
 sg13g2_fill_1 FILLER_39_2669 ();
 sg13g2_fill_2 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_2 ();
 sg13g2_decap_8 FILLER_40_74 ();
 sg13g2_decap_4 FILLER_40_81 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_124 ();
 sg13g2_decap_8 FILLER_40_129 ();
 sg13g2_decap_4 FILLER_40_136 ();
 sg13g2_fill_1 FILLER_40_140 ();
 sg13g2_decap_4 FILLER_40_151 ();
 sg13g2_fill_1 FILLER_40_155 ();
 sg13g2_decap_8 FILLER_40_160 ();
 sg13g2_decap_8 FILLER_40_167 ();
 sg13g2_decap_8 FILLER_40_174 ();
 sg13g2_fill_1 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_187 ();
 sg13g2_fill_1 FILLER_40_191 ();
 sg13g2_decap_4 FILLER_40_206 ();
 sg13g2_fill_1 FILLER_40_210 ();
 sg13g2_fill_2 FILLER_40_260 ();
 sg13g2_fill_1 FILLER_40_262 ();
 sg13g2_fill_2 FILLER_40_275 ();
 sg13g2_fill_1 FILLER_40_277 ();
 sg13g2_fill_2 FILLER_40_283 ();
 sg13g2_fill_1 FILLER_40_300 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_2 FILLER_40_362 ();
 sg13g2_decap_4 FILLER_40_434 ();
 sg13g2_fill_2 FILLER_40_438 ();
 sg13g2_decap_4 FILLER_40_443 ();
 sg13g2_fill_1 FILLER_40_447 ();
 sg13g2_fill_1 FILLER_40_474 ();
 sg13g2_fill_2 FILLER_40_479 ();
 sg13g2_fill_2 FILLER_40_489 ();
 sg13g2_fill_2 FILLER_40_496 ();
 sg13g2_decap_4 FILLER_40_537 ();
 sg13g2_fill_1 FILLER_40_549 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_4 FILLER_40_574 ();
 sg13g2_fill_1 FILLER_40_597 ();
 sg13g2_decap_4 FILLER_40_603 ();
 sg13g2_fill_2 FILLER_40_607 ();
 sg13g2_fill_1 FILLER_40_618 ();
 sg13g2_decap_4 FILLER_40_640 ();
 sg13g2_fill_1 FILLER_40_644 ();
 sg13g2_fill_2 FILLER_40_650 ();
 sg13g2_decap_4 FILLER_40_668 ();
 sg13g2_fill_1 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_678 ();
 sg13g2_decap_8 FILLER_40_690 ();
 sg13g2_fill_2 FILLER_40_697 ();
 sg13g2_fill_1 FILLER_40_699 ();
 sg13g2_fill_2 FILLER_40_793 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_fill_2 FILLER_40_826 ();
 sg13g2_fill_1 FILLER_40_828 ();
 sg13g2_fill_1 FILLER_40_852 ();
 sg13g2_decap_8 FILLER_40_889 ();
 sg13g2_fill_1 FILLER_40_930 ();
 sg13g2_fill_2 FILLER_40_957 ();
 sg13g2_fill_2 FILLER_40_963 ();
 sg13g2_decap_8 FILLER_40_991 ();
 sg13g2_fill_1 FILLER_40_1012 ();
 sg13g2_decap_4 FILLER_40_1081 ();
 sg13g2_fill_1 FILLER_40_1085 ();
 sg13g2_decap_8 FILLER_40_1091 ();
 sg13g2_decap_8 FILLER_40_1098 ();
 sg13g2_decap_4 FILLER_40_1105 ();
 sg13g2_fill_1 FILLER_40_1109 ();
 sg13g2_decap_8 FILLER_40_1131 ();
 sg13g2_fill_1 FILLER_40_1138 ();
 sg13g2_fill_2 FILLER_40_1144 ();
 sg13g2_fill_1 FILLER_40_1146 ();
 sg13g2_decap_8 FILLER_40_1157 ();
 sg13g2_decap_8 FILLER_40_1164 ();
 sg13g2_decap_8 FILLER_40_1171 ();
 sg13g2_fill_2 FILLER_40_1178 ();
 sg13g2_fill_1 FILLER_40_1189 ();
 sg13g2_decap_4 FILLER_40_1194 ();
 sg13g2_fill_1 FILLER_40_1198 ();
 sg13g2_fill_1 FILLER_40_1204 ();
 sg13g2_fill_1 FILLER_40_1209 ();
 sg13g2_fill_2 FILLER_40_1248 ();
 sg13g2_decap_8 FILLER_40_1332 ();
 sg13g2_decap_8 FILLER_40_1339 ();
 sg13g2_decap_8 FILLER_40_1346 ();
 sg13g2_decap_8 FILLER_40_1353 ();
 sg13g2_fill_2 FILLER_40_1360 ();
 sg13g2_decap_8 FILLER_40_1398 ();
 sg13g2_decap_8 FILLER_40_1405 ();
 sg13g2_decap_8 FILLER_40_1412 ();
 sg13g2_decap_8 FILLER_40_1419 ();
 sg13g2_decap_8 FILLER_40_1426 ();
 sg13g2_fill_2 FILLER_40_1433 ();
 sg13g2_fill_1 FILLER_40_1435 ();
 sg13g2_fill_1 FILLER_40_1441 ();
 sg13g2_fill_1 FILLER_40_1447 ();
 sg13g2_fill_1 FILLER_40_1458 ();
 sg13g2_decap_8 FILLER_40_1471 ();
 sg13g2_decap_4 FILLER_40_1519 ();
 sg13g2_fill_1 FILLER_40_1536 ();
 sg13g2_decap_4 FILLER_40_1582 ();
 sg13g2_fill_1 FILLER_40_1586 ();
 sg13g2_decap_4 FILLER_40_1610 ();
 sg13g2_fill_1 FILLER_40_1614 ();
 sg13g2_fill_1 FILLER_40_1631 ();
 sg13g2_fill_2 FILLER_40_1636 ();
 sg13g2_fill_1 FILLER_40_1642 ();
 sg13g2_fill_2 FILLER_40_1648 ();
 sg13g2_fill_2 FILLER_40_1658 ();
 sg13g2_fill_2 FILLER_40_1668 ();
 sg13g2_fill_1 FILLER_40_1683 ();
 sg13g2_fill_2 FILLER_40_1728 ();
 sg13g2_decap_8 FILLER_40_1761 ();
 sg13g2_decap_8 FILLER_40_1768 ();
 sg13g2_decap_8 FILLER_40_1775 ();
 sg13g2_decap_8 FILLER_40_1782 ();
 sg13g2_fill_2 FILLER_40_1789 ();
 sg13g2_decap_8 FILLER_40_1795 ();
 sg13g2_fill_1 FILLER_40_1832 ();
 sg13g2_fill_1 FILLER_40_1837 ();
 sg13g2_fill_2 FILLER_40_1875 ();
 sg13g2_fill_1 FILLER_40_1890 ();
 sg13g2_fill_2 FILLER_40_1960 ();
 sg13g2_fill_1 FILLER_40_1962 ();
 sg13g2_fill_1 FILLER_40_1979 ();
 sg13g2_fill_2 FILLER_40_2010 ();
 sg13g2_fill_1 FILLER_40_2012 ();
 sg13g2_decap_8 FILLER_40_2048 ();
 sg13g2_decap_8 FILLER_40_2055 ();
 sg13g2_decap_8 FILLER_40_2062 ();
 sg13g2_fill_1 FILLER_40_2069 ();
 sg13g2_decap_8 FILLER_40_2082 ();
 sg13g2_fill_2 FILLER_40_2089 ();
 sg13g2_fill_1 FILLER_40_2091 ();
 sg13g2_decap_8 FILLER_40_2097 ();
 sg13g2_fill_2 FILLER_40_2104 ();
 sg13g2_fill_1 FILLER_40_2106 ();
 sg13g2_decap_8 FILLER_40_2111 ();
 sg13g2_decap_4 FILLER_40_2118 ();
 sg13g2_fill_1 FILLER_40_2122 ();
 sg13g2_fill_1 FILLER_40_2127 ();
 sg13g2_decap_8 FILLER_40_2154 ();
 sg13g2_decap_8 FILLER_40_2161 ();
 sg13g2_decap_8 FILLER_40_2168 ();
 sg13g2_decap_4 FILLER_40_2175 ();
 sg13g2_fill_1 FILLER_40_2179 ();
 sg13g2_decap_4 FILLER_40_2206 ();
 sg13g2_fill_1 FILLER_40_2210 ();
 sg13g2_fill_1 FILLER_40_2220 ();
 sg13g2_fill_1 FILLER_40_2228 ();
 sg13g2_fill_2 FILLER_40_2265 ();
 sg13g2_fill_1 FILLER_40_2267 ();
 sg13g2_decap_4 FILLER_40_2271 ();
 sg13g2_fill_2 FILLER_40_2275 ();
 sg13g2_fill_1 FILLER_40_2286 ();
 sg13g2_fill_1 FILLER_40_2297 ();
 sg13g2_decap_8 FILLER_40_2311 ();
 sg13g2_fill_1 FILLER_40_2318 ();
 sg13g2_fill_2 FILLER_40_2329 ();
 sg13g2_fill_1 FILLER_40_2334 ();
 sg13g2_fill_1 FILLER_40_2357 ();
 sg13g2_fill_2 FILLER_40_2374 ();
 sg13g2_fill_1 FILLER_40_2376 ();
 sg13g2_decap_8 FILLER_40_2381 ();
 sg13g2_decap_8 FILLER_40_2388 ();
 sg13g2_decap_8 FILLER_40_2395 ();
 sg13g2_decap_8 FILLER_40_2402 ();
 sg13g2_decap_8 FILLER_40_2409 ();
 sg13g2_decap_4 FILLER_40_2416 ();
 sg13g2_fill_2 FILLER_40_2420 ();
 sg13g2_fill_1 FILLER_40_2426 ();
 sg13g2_fill_1 FILLER_40_2444 ();
 sg13g2_fill_1 FILLER_40_2451 ();
 sg13g2_decap_8 FILLER_40_2459 ();
 sg13g2_decap_8 FILLER_40_2466 ();
 sg13g2_fill_1 FILLER_40_2473 ();
 sg13g2_fill_1 FILLER_40_2491 ();
 sg13g2_decap_8 FILLER_40_2496 ();
 sg13g2_decap_8 FILLER_40_2503 ();
 sg13g2_decap_8 FILLER_40_2536 ();
 sg13g2_decap_8 FILLER_40_2543 ();
 sg13g2_decap_8 FILLER_40_2550 ();
 sg13g2_decap_8 FILLER_40_2557 ();
 sg13g2_decap_8 FILLER_40_2564 ();
 sg13g2_decap_8 FILLER_40_2571 ();
 sg13g2_decap_8 FILLER_40_2578 ();
 sg13g2_decap_8 FILLER_40_2585 ();
 sg13g2_decap_8 FILLER_40_2592 ();
 sg13g2_decap_8 FILLER_40_2599 ();
 sg13g2_decap_8 FILLER_40_2606 ();
 sg13g2_decap_8 FILLER_40_2613 ();
 sg13g2_decap_8 FILLER_40_2620 ();
 sg13g2_decap_8 FILLER_40_2627 ();
 sg13g2_decap_8 FILLER_40_2634 ();
 sg13g2_decap_8 FILLER_40_2641 ();
 sg13g2_decap_8 FILLER_40_2648 ();
 sg13g2_decap_8 FILLER_40_2655 ();
 sg13g2_decap_8 FILLER_40_2662 ();
 sg13g2_fill_1 FILLER_40_2669 ();
 sg13g2_fill_1 FILLER_41_44 ();
 sg13g2_fill_2 FILLER_41_62 ();
 sg13g2_decap_8 FILLER_41_68 ();
 sg13g2_decap_8 FILLER_41_75 ();
 sg13g2_decap_8 FILLER_41_82 ();
 sg13g2_decap_4 FILLER_41_89 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_fill_1 FILLER_41_110 ();
 sg13g2_decap_4 FILLER_41_115 ();
 sg13g2_decap_4 FILLER_41_124 ();
 sg13g2_fill_1 FILLER_41_128 ();
 sg13g2_decap_8 FILLER_41_136 ();
 sg13g2_fill_2 FILLER_41_157 ();
 sg13g2_fill_1 FILLER_41_159 ();
 sg13g2_decap_4 FILLER_41_168 ();
 sg13g2_fill_2 FILLER_41_172 ();
 sg13g2_decap_4 FILLER_41_184 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_fill_2 FILLER_41_216 ();
 sg13g2_fill_1 FILLER_41_218 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_4 FILLER_41_252 ();
 sg13g2_fill_1 FILLER_41_287 ();
 sg13g2_fill_1 FILLER_41_314 ();
 sg13g2_decap_8 FILLER_41_325 ();
 sg13g2_decap_8 FILLER_41_332 ();
 sg13g2_fill_1 FILLER_41_339 ();
 sg13g2_decap_4 FILLER_41_344 ();
 sg13g2_fill_2 FILLER_41_348 ();
 sg13g2_fill_1 FILLER_41_363 ();
 sg13g2_fill_2 FILLER_41_378 ();
 sg13g2_fill_1 FILLER_41_380 ();
 sg13g2_fill_1 FILLER_41_385 ();
 sg13g2_fill_1 FILLER_41_394 ();
 sg13g2_fill_2 FILLER_41_400 ();
 sg13g2_fill_1 FILLER_41_407 ();
 sg13g2_fill_2 FILLER_41_421 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_4 FILLER_41_441 ();
 sg13g2_fill_2 FILLER_41_449 ();
 sg13g2_fill_1 FILLER_41_451 ();
 sg13g2_fill_2 FILLER_41_456 ();
 sg13g2_fill_2 FILLER_41_462 ();
 sg13g2_fill_1 FILLER_41_464 ();
 sg13g2_fill_1 FILLER_41_469 ();
 sg13g2_fill_2 FILLER_41_475 ();
 sg13g2_fill_1 FILLER_41_477 ();
 sg13g2_fill_2 FILLER_41_482 ();
 sg13g2_fill_1 FILLER_41_484 ();
 sg13g2_fill_2 FILLER_41_493 ();
 sg13g2_fill_1 FILLER_41_495 ();
 sg13g2_decap_8 FILLER_41_527 ();
 sg13g2_fill_1 FILLER_41_534 ();
 sg13g2_decap_8 FILLER_41_566 ();
 sg13g2_decap_4 FILLER_41_592 ();
 sg13g2_fill_1 FILLER_41_608 ();
 sg13g2_decap_8 FILLER_41_643 ();
 sg13g2_fill_2 FILLER_41_650 ();
 sg13g2_decap_8 FILLER_41_698 ();
 sg13g2_fill_2 FILLER_41_705 ();
 sg13g2_fill_1 FILLER_41_707 ();
 sg13g2_decap_4 FILLER_41_712 ();
 sg13g2_fill_1 FILLER_41_770 ();
 sg13g2_fill_1 FILLER_41_787 ();
 sg13g2_decap_4 FILLER_41_814 ();
 sg13g2_fill_1 FILLER_41_848 ();
 sg13g2_fill_2 FILLER_41_892 ();
 sg13g2_decap_8 FILLER_41_902 ();
 sg13g2_fill_2 FILLER_41_913 ();
 sg13g2_fill_1 FILLER_41_915 ();
 sg13g2_fill_1 FILLER_41_936 ();
 sg13g2_decap_8 FILLER_41_981 ();
 sg13g2_fill_1 FILLER_41_993 ();
 sg13g2_fill_2 FILLER_41_1020 ();
 sg13g2_fill_2 FILLER_41_1026 ();
 sg13g2_fill_2 FILLER_41_1032 ();
 sg13g2_fill_1 FILLER_41_1034 ();
 sg13g2_fill_2 FILLER_41_1061 ();
 sg13g2_decap_8 FILLER_41_1067 ();
 sg13g2_decap_4 FILLER_41_1074 ();
 sg13g2_fill_2 FILLER_41_1078 ();
 sg13g2_decap_8 FILLER_41_1101 ();
 sg13g2_fill_1 FILLER_41_1108 ();
 sg13g2_fill_1 FILLER_41_1161 ();
 sg13g2_fill_2 FILLER_41_1213 ();
 sg13g2_fill_1 FILLER_41_1215 ();
 sg13g2_decap_4 FILLER_41_1224 ();
 sg13g2_fill_1 FILLER_41_1261 ();
 sg13g2_fill_2 FILLER_41_1306 ();
 sg13g2_decap_4 FILLER_41_1344 ();
 sg13g2_decap_8 FILLER_41_1358 ();
 sg13g2_decap_4 FILLER_41_1383 ();
 sg13g2_fill_2 FILLER_41_1387 ();
 sg13g2_decap_8 FILLER_41_1425 ();
 sg13g2_decap_8 FILLER_41_1432 ();
 sg13g2_fill_1 FILLER_41_1457 ();
 sg13g2_fill_2 FILLER_41_1471 ();
 sg13g2_fill_1 FILLER_41_1473 ();
 sg13g2_fill_2 FILLER_41_1512 ();
 sg13g2_fill_2 FILLER_41_1552 ();
 sg13g2_fill_1 FILLER_41_1554 ();
 sg13g2_fill_2 FILLER_41_1559 ();
 sg13g2_decap_8 FILLER_41_1585 ();
 sg13g2_decap_8 FILLER_41_1592 ();
 sg13g2_fill_2 FILLER_41_1599 ();
 sg13g2_fill_1 FILLER_41_1601 ();
 sg13g2_fill_2 FILLER_41_1607 ();
 sg13g2_fill_1 FILLER_41_1614 ();
 sg13g2_fill_1 FILLER_41_1619 ();
 sg13g2_fill_1 FILLER_41_1632 ();
 sg13g2_fill_1 FILLER_41_1638 ();
 sg13g2_decap_4 FILLER_41_1666 ();
 sg13g2_fill_2 FILLER_41_1679 ();
 sg13g2_fill_1 FILLER_41_1681 ();
 sg13g2_fill_1 FILLER_41_1700 ();
 sg13g2_decap_8 FILLER_41_1704 ();
 sg13g2_decap_4 FILLER_41_1711 ();
 sg13g2_decap_8 FILLER_41_1763 ();
 sg13g2_decap_4 FILLER_41_1770 ();
 sg13g2_fill_2 FILLER_41_1774 ();
 sg13g2_fill_2 FILLER_41_1780 ();
 sg13g2_decap_8 FILLER_41_1818 ();
 sg13g2_decap_8 FILLER_41_1825 ();
 sg13g2_fill_1 FILLER_41_1837 ();
 sg13g2_fill_1 FILLER_41_1888 ();
 sg13g2_fill_1 FILLER_41_1901 ();
 sg13g2_fill_1 FILLER_41_1912 ();
 sg13g2_fill_1 FILLER_41_1934 ();
 sg13g2_fill_2 FILLER_41_1963 ();
 sg13g2_fill_1 FILLER_41_1965 ();
 sg13g2_fill_2 FILLER_41_1979 ();
 sg13g2_decap_4 FILLER_41_2011 ();
 sg13g2_decap_8 FILLER_41_2055 ();
 sg13g2_decap_4 FILLER_41_2062 ();
 sg13g2_fill_1 FILLER_41_2092 ();
 sg13g2_decap_8 FILLER_41_2097 ();
 sg13g2_decap_8 FILLER_41_2104 ();
 sg13g2_fill_2 FILLER_41_2111 ();
 sg13g2_fill_1 FILLER_41_2113 ();
 sg13g2_fill_2 FILLER_41_2119 ();
 sg13g2_decap_8 FILLER_41_2173 ();
 sg13g2_decap_8 FILLER_41_2180 ();
 sg13g2_fill_1 FILLER_41_2187 ();
 sg13g2_fill_2 FILLER_41_2192 ();
 sg13g2_fill_1 FILLER_41_2194 ();
 sg13g2_fill_2 FILLER_41_2231 ();
 sg13g2_fill_1 FILLER_41_2241 ();
 sg13g2_fill_1 FILLER_41_2308 ();
 sg13g2_fill_2 FILLER_41_2325 ();
 sg13g2_decap_8 FILLER_41_2379 ();
 sg13g2_decap_8 FILLER_41_2386 ();
 sg13g2_fill_2 FILLER_41_2393 ();
 sg13g2_decap_8 FILLER_41_2405 ();
 sg13g2_fill_1 FILLER_41_2412 ();
 sg13g2_decap_4 FILLER_41_2417 ();
 sg13g2_fill_2 FILLER_41_2421 ();
 sg13g2_fill_1 FILLER_41_2474 ();
 sg13g2_fill_2 FILLER_41_2488 ();
 sg13g2_decap_8 FILLER_41_2494 ();
 sg13g2_decap_8 FILLER_41_2501 ();
 sg13g2_decap_8 FILLER_41_2508 ();
 sg13g2_decap_8 FILLER_41_2515 ();
 sg13g2_decap_8 FILLER_41_2522 ();
 sg13g2_fill_2 FILLER_41_2529 ();
 sg13g2_decap_8 FILLER_41_2534 ();
 sg13g2_fill_2 FILLER_41_2541 ();
 sg13g2_fill_1 FILLER_41_2543 ();
 sg13g2_decap_8 FILLER_41_2548 ();
 sg13g2_decap_8 FILLER_41_2555 ();
 sg13g2_decap_8 FILLER_41_2562 ();
 sg13g2_decap_8 FILLER_41_2569 ();
 sg13g2_decap_8 FILLER_41_2576 ();
 sg13g2_decap_8 FILLER_41_2583 ();
 sg13g2_decap_8 FILLER_41_2590 ();
 sg13g2_decap_8 FILLER_41_2597 ();
 sg13g2_decap_8 FILLER_41_2604 ();
 sg13g2_decap_8 FILLER_41_2611 ();
 sg13g2_decap_8 FILLER_41_2618 ();
 sg13g2_decap_8 FILLER_41_2625 ();
 sg13g2_decap_8 FILLER_41_2632 ();
 sg13g2_decap_8 FILLER_41_2639 ();
 sg13g2_decap_8 FILLER_41_2646 ();
 sg13g2_decap_8 FILLER_41_2653 ();
 sg13g2_decap_8 FILLER_41_2660 ();
 sg13g2_fill_2 FILLER_41_2667 ();
 sg13g2_fill_1 FILLER_41_2669 ();
 sg13g2_decap_4 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_4 ();
 sg13g2_fill_1 FILLER_42_40 ();
 sg13g2_fill_1 FILLER_42_46 ();
 sg13g2_fill_1 FILLER_42_52 ();
 sg13g2_fill_1 FILLER_42_57 ();
 sg13g2_decap_8 FILLER_42_62 ();
 sg13g2_decap_8 FILLER_42_69 ();
 sg13g2_decap_8 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_83 ();
 sg13g2_decap_4 FILLER_42_89 ();
 sg13g2_fill_2 FILLER_42_93 ();
 sg13g2_fill_1 FILLER_42_99 ();
 sg13g2_fill_2 FILLER_42_113 ();
 sg13g2_fill_1 FILLER_42_123 ();
 sg13g2_fill_2 FILLER_42_129 ();
 sg13g2_fill_1 FILLER_42_136 ();
 sg13g2_fill_2 FILLER_42_163 ();
 sg13g2_fill_2 FILLER_42_170 ();
 sg13g2_decap_4 FILLER_42_177 ();
 sg13g2_fill_1 FILLER_42_181 ();
 sg13g2_decap_8 FILLER_42_208 ();
 sg13g2_fill_1 FILLER_42_215 ();
 sg13g2_fill_1 FILLER_42_219 ();
 sg13g2_fill_2 FILLER_42_224 ();
 sg13g2_fill_1 FILLER_42_226 ();
 sg13g2_decap_4 FILLER_42_231 ();
 sg13g2_fill_2 FILLER_42_235 ();
 sg13g2_fill_2 FILLER_42_241 ();
 sg13g2_fill_1 FILLER_42_243 ();
 sg13g2_fill_2 FILLER_42_267 ();
 sg13g2_fill_1 FILLER_42_269 ();
 sg13g2_decap_4 FILLER_42_274 ();
 sg13g2_fill_2 FILLER_42_282 ();
 sg13g2_fill_1 FILLER_42_284 ();
 sg13g2_fill_1 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_299 ();
 sg13g2_decap_8 FILLER_42_314 ();
 sg13g2_decap_8 FILLER_42_321 ();
 sg13g2_decap_8 FILLER_42_328 ();
 sg13g2_fill_1 FILLER_42_335 ();
 sg13g2_decap_4 FILLER_42_339 ();
 sg13g2_fill_2 FILLER_42_343 ();
 sg13g2_fill_2 FILLER_42_357 ();
 sg13g2_decap_8 FILLER_42_392 ();
 sg13g2_fill_2 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_409 ();
 sg13g2_fill_1 FILLER_42_411 ();
 sg13g2_decap_8 FILLER_42_418 ();
 sg13g2_fill_2 FILLER_42_425 ();
 sg13g2_fill_1 FILLER_42_427 ();
 sg13g2_fill_1 FILLER_42_443 ();
 sg13g2_fill_2 FILLER_42_470 ();
 sg13g2_fill_1 FILLER_42_482 ();
 sg13g2_fill_2 FILLER_42_509 ();
 sg13g2_decap_4 FILLER_42_516 ();
 sg13g2_decap_4 FILLER_42_524 ();
 sg13g2_fill_2 FILLER_42_538 ();
 sg13g2_fill_1 FILLER_42_540 ();
 sg13g2_decap_8 FILLER_42_545 ();
 sg13g2_decap_8 FILLER_42_552 ();
 sg13g2_decap_8 FILLER_42_559 ();
 sg13g2_decap_8 FILLER_42_566 ();
 sg13g2_decap_4 FILLER_42_578 ();
 sg13g2_fill_1 FILLER_42_587 ();
 sg13g2_fill_1 FILLER_42_609 ();
 sg13g2_decap_8 FILLER_42_657 ();
 sg13g2_decap_8 FILLER_42_664 ();
 sg13g2_fill_2 FILLER_42_671 ();
 sg13g2_fill_1 FILLER_42_693 ();
 sg13g2_fill_1 FILLER_42_699 ();
 sg13g2_decap_4 FILLER_42_705 ();
 sg13g2_fill_1 FILLER_42_713 ();
 sg13g2_decap_4 FILLER_42_723 ();
 sg13g2_fill_2 FILLER_42_731 ();
 sg13g2_fill_2 FILLER_42_746 ();
 sg13g2_decap_4 FILLER_42_810 ();
 sg13g2_fill_2 FILLER_42_884 ();
 sg13g2_fill_2 FILLER_42_912 ();
 sg13g2_decap_8 FILLER_42_924 ();
 sg13g2_decap_8 FILLER_42_931 ();
 sg13g2_decap_8 FILLER_42_938 ();
 sg13g2_fill_2 FILLER_42_945 ();
 sg13g2_fill_1 FILLER_42_947 ();
 sg13g2_decap_8 FILLER_42_952 ();
 sg13g2_decap_8 FILLER_42_959 ();
 sg13g2_decap_8 FILLER_42_966 ();
 sg13g2_decap_8 FILLER_42_973 ();
 sg13g2_decap_8 FILLER_42_980 ();
 sg13g2_fill_1 FILLER_42_987 ();
 sg13g2_fill_2 FILLER_42_1035 ();
 sg13g2_fill_2 FILLER_42_1072 ();
 sg13g2_fill_1 FILLER_42_1074 ();
 sg13g2_decap_8 FILLER_42_1079 ();
 sg13g2_fill_1 FILLER_42_1086 ();
 sg13g2_fill_2 FILLER_42_1095 ();
 sg13g2_fill_2 FILLER_42_1145 ();
 sg13g2_fill_1 FILLER_42_1147 ();
 sg13g2_fill_2 FILLER_42_1153 ();
 sg13g2_fill_1 FILLER_42_1155 ();
 sg13g2_fill_1 FILLER_42_1182 ();
 sg13g2_fill_1 FILLER_42_1222 ();
 sg13g2_fill_1 FILLER_42_1270 ();
 sg13g2_fill_2 FILLER_42_1304 ();
 sg13g2_decap_4 FILLER_42_1310 ();
 sg13g2_decap_4 FILLER_42_1322 ();
 sg13g2_fill_1 FILLER_42_1378 ();
 sg13g2_decap_8 FILLER_42_1419 ();
 sg13g2_decap_4 FILLER_42_1426 ();
 sg13g2_decap_4 FILLER_42_1461 ();
 sg13g2_decap_8 FILLER_42_1485 ();
 sg13g2_fill_2 FILLER_42_1492 ();
 sg13g2_fill_1 FILLER_42_1510 ();
 sg13g2_decap_4 FILLER_42_1521 ();
 sg13g2_fill_1 FILLER_42_1525 ();
 sg13g2_decap_8 FILLER_42_1534 ();
 sg13g2_decap_8 FILLER_42_1541 ();
 sg13g2_decap_4 FILLER_42_1548 ();
 sg13g2_decap_4 FILLER_42_1565 ();
 sg13g2_fill_1 FILLER_42_1586 ();
 sg13g2_fill_1 FILLER_42_1593 ();
 sg13g2_fill_2 FILLER_42_1609 ();
 sg13g2_fill_2 FILLER_42_1623 ();
 sg13g2_decap_8 FILLER_42_1664 ();
 sg13g2_fill_2 FILLER_42_1671 ();
 sg13g2_fill_1 FILLER_42_1673 ();
 sg13g2_decap_8 FILLER_42_1691 ();
 sg13g2_decap_8 FILLER_42_1698 ();
 sg13g2_decap_8 FILLER_42_1705 ();
 sg13g2_decap_8 FILLER_42_1712 ();
 sg13g2_fill_2 FILLER_42_1719 ();
 sg13g2_decap_4 FILLER_42_1724 ();
 sg13g2_fill_1 FILLER_42_1728 ();
 sg13g2_decap_4 FILLER_42_1746 ();
 sg13g2_fill_1 FILLER_42_1750 ();
 sg13g2_fill_1 FILLER_42_1768 ();
 sg13g2_decap_8 FILLER_42_1795 ();
 sg13g2_fill_2 FILLER_42_1802 ();
 sg13g2_decap_8 FILLER_42_1808 ();
 sg13g2_decap_8 FILLER_42_1815 ();
 sg13g2_decap_8 FILLER_42_1822 ();
 sg13g2_decap_8 FILLER_42_1829 ();
 sg13g2_decap_4 FILLER_42_1836 ();
 sg13g2_fill_1 FILLER_42_1840 ();
 sg13g2_fill_2 FILLER_42_1858 ();
 sg13g2_fill_2 FILLER_42_1864 ();
 sg13g2_fill_2 FILLER_42_1871 ();
 sg13g2_decap_8 FILLER_42_1900 ();
 sg13g2_fill_1 FILLER_42_1920 ();
 sg13g2_fill_2 FILLER_42_1934 ();
 sg13g2_fill_1 FILLER_42_1961 ();
 sg13g2_decap_8 FILLER_42_1967 ();
 sg13g2_decap_8 FILLER_42_1974 ();
 sg13g2_decap_4 FILLER_42_1981 ();
 sg13g2_fill_2 FILLER_42_1995 ();
 sg13g2_fill_1 FILLER_42_1997 ();
 sg13g2_decap_4 FILLER_42_2002 ();
 sg13g2_fill_2 FILLER_42_2011 ();
 sg13g2_fill_1 FILLER_42_2013 ();
 sg13g2_fill_2 FILLER_42_2019 ();
 sg13g2_fill_1 FILLER_42_2025 ();
 sg13g2_fill_2 FILLER_42_2052 ();
 sg13g2_fill_1 FILLER_42_2089 ();
 sg13g2_fill_2 FILLER_42_2120 ();
 sg13g2_decap_8 FILLER_42_2127 ();
 sg13g2_fill_2 FILLER_42_2143 ();
 sg13g2_fill_1 FILLER_42_2145 ();
 sg13g2_decap_4 FILLER_42_2189 ();
 sg13g2_fill_2 FILLER_42_2193 ();
 sg13g2_fill_1 FILLER_42_2224 ();
 sg13g2_fill_2 FILLER_42_2269 ();
 sg13g2_fill_2 FILLER_42_2347 ();
 sg13g2_fill_2 FILLER_42_2379 ();
 sg13g2_fill_1 FILLER_42_2381 ();
 sg13g2_decap_8 FILLER_42_2441 ();
 sg13g2_decap_4 FILLER_42_2448 ();
 sg13g2_fill_1 FILLER_42_2456 ();
 sg13g2_fill_1 FILLER_42_2483 ();
 sg13g2_fill_1 FILLER_42_2510 ();
 sg13g2_fill_1 FILLER_42_2537 ();
 sg13g2_fill_1 FILLER_42_2564 ();
 sg13g2_fill_2 FILLER_42_2575 ();
 sg13g2_decap_8 FILLER_42_2581 ();
 sg13g2_decap_8 FILLER_42_2588 ();
 sg13g2_decap_8 FILLER_42_2595 ();
 sg13g2_decap_8 FILLER_42_2602 ();
 sg13g2_decap_8 FILLER_42_2609 ();
 sg13g2_decap_8 FILLER_42_2616 ();
 sg13g2_decap_8 FILLER_42_2623 ();
 sg13g2_decap_8 FILLER_42_2630 ();
 sg13g2_decap_8 FILLER_42_2637 ();
 sg13g2_decap_8 FILLER_42_2644 ();
 sg13g2_decap_8 FILLER_42_2651 ();
 sg13g2_decap_8 FILLER_42_2658 ();
 sg13g2_decap_4 FILLER_42_2665 ();
 sg13g2_fill_1 FILLER_42_2669 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_14 ();
 sg13g2_fill_2 FILLER_43_20 ();
 sg13g2_fill_2 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_29 ();
 sg13g2_fill_1 FILLER_43_34 ();
 sg13g2_fill_2 FILLER_43_39 ();
 sg13g2_fill_1 FILLER_43_41 ();
 sg13g2_fill_1 FILLER_43_77 ();
 sg13g2_fill_1 FILLER_43_130 ();
 sg13g2_fill_1 FILLER_43_139 ();
 sg13g2_fill_2 FILLER_43_196 ();
 sg13g2_fill_1 FILLER_43_198 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_fill_1 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_264 ();
 sg13g2_decap_4 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_290 ();
 sg13g2_fill_1 FILLER_43_305 ();
 sg13g2_fill_2 FILLER_43_319 ();
 sg13g2_decap_8 FILLER_43_326 ();
 sg13g2_fill_2 FILLER_43_344 ();
 sg13g2_fill_1 FILLER_43_358 ();
 sg13g2_fill_2 FILLER_43_392 ();
 sg13g2_decap_4 FILLER_43_399 ();
 sg13g2_fill_1 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_408 ();
 sg13g2_decap_8 FILLER_43_415 ();
 sg13g2_fill_2 FILLER_43_422 ();
 sg13g2_fill_1 FILLER_43_424 ();
 sg13g2_decap_8 FILLER_43_442 ();
 sg13g2_fill_2 FILLER_43_449 ();
 sg13g2_decap_8 FILLER_43_468 ();
 sg13g2_decap_8 FILLER_43_475 ();
 sg13g2_decap_8 FILLER_43_482 ();
 sg13g2_decap_8 FILLER_43_489 ();
 sg13g2_decap_4 FILLER_43_496 ();
 sg13g2_fill_1 FILLER_43_500 ();
 sg13g2_decap_8 FILLER_43_535 ();
 sg13g2_decap_8 FILLER_43_542 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_fill_1 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_fill_2 FILLER_43_617 ();
 sg13g2_fill_1 FILLER_43_629 ();
 sg13g2_fill_2 FILLER_43_647 ();
 sg13g2_fill_1 FILLER_43_649 ();
 sg13g2_decap_4 FILLER_43_704 ();
 sg13g2_fill_1 FILLER_43_708 ();
 sg13g2_decap_4 FILLER_43_714 ();
 sg13g2_fill_1 FILLER_43_718 ();
 sg13g2_fill_2 FILLER_43_755 ();
 sg13g2_fill_1 FILLER_43_757 ();
 sg13g2_fill_2 FILLER_43_801 ();
 sg13g2_decap_4 FILLER_43_813 ();
 sg13g2_fill_2 FILLER_43_817 ();
 sg13g2_fill_2 FILLER_43_846 ();
 sg13g2_fill_1 FILLER_43_856 ();
 sg13g2_decap_8 FILLER_43_913 ();
 sg13g2_fill_1 FILLER_43_920 ();
 sg13g2_fill_2 FILLER_43_947 ();
 sg13g2_fill_2 FILLER_43_959 ();
 sg13g2_fill_1 FILLER_43_961 ();
 sg13g2_fill_2 FILLER_43_966 ();
 sg13g2_fill_1 FILLER_43_968 ();
 sg13g2_fill_2 FILLER_43_990 ();
 sg13g2_fill_1 FILLER_43_992 ();
 sg13g2_fill_1 FILLER_43_1034 ();
 sg13g2_decap_8 FILLER_43_1040 ();
 sg13g2_fill_1 FILLER_43_1047 ();
 sg13g2_decap_8 FILLER_43_1092 ();
 sg13g2_decap_8 FILLER_43_1104 ();
 sg13g2_fill_1 FILLER_43_1141 ();
 sg13g2_fill_1 FILLER_43_1168 ();
 sg13g2_fill_1 FILLER_43_1195 ();
 sg13g2_fill_2 FILLER_43_1217 ();
 sg13g2_fill_1 FILLER_43_1224 ();
 sg13g2_fill_1 FILLER_43_1249 ();
 sg13g2_fill_1 FILLER_43_1268 ();
 sg13g2_decap_8 FILLER_43_1297 ();
 sg13g2_decap_4 FILLER_43_1304 ();
 sg13g2_fill_2 FILLER_43_1324 ();
 sg13g2_fill_2 FILLER_43_1331 ();
 sg13g2_fill_1 FILLER_43_1333 ();
 sg13g2_fill_1 FILLER_43_1341 ();
 sg13g2_decap_4 FILLER_43_1372 ();
 sg13g2_fill_1 FILLER_43_1412 ();
 sg13g2_fill_2 FILLER_43_1443 ();
 sg13g2_decap_8 FILLER_43_1448 ();
 sg13g2_decap_4 FILLER_43_1461 ();
 sg13g2_fill_1 FILLER_43_1465 ();
 sg13g2_fill_2 FILLER_43_1490 ();
 sg13g2_fill_1 FILLER_43_1498 ();
 sg13g2_fill_2 FILLER_43_1509 ();
 sg13g2_fill_2 FILLER_43_1537 ();
 sg13g2_decap_4 FILLER_43_1544 ();
 sg13g2_fill_2 FILLER_43_1548 ();
 sg13g2_fill_1 FILLER_43_1563 ();
 sg13g2_fill_1 FILLER_43_1598 ();
 sg13g2_fill_2 FILLER_43_1602 ();
 sg13g2_fill_1 FILLER_43_1604 ();
 sg13g2_fill_2 FILLER_43_1608 ();
 sg13g2_fill_1 FILLER_43_1610 ();
 sg13g2_decap_4 FILLER_43_1620 ();
 sg13g2_fill_1 FILLER_43_1624 ();
 sg13g2_fill_2 FILLER_43_1630 ();
 sg13g2_fill_1 FILLER_43_1632 ();
 sg13g2_decap_8 FILLER_43_1659 ();
 sg13g2_fill_2 FILLER_43_1666 ();
 sg13g2_fill_1 FILLER_43_1668 ();
 sg13g2_decap_8 FILLER_43_1699 ();
 sg13g2_decap_8 FILLER_43_1706 ();
 sg13g2_decap_8 FILLER_43_1713 ();
 sg13g2_decap_8 FILLER_43_1729 ();
 sg13g2_decap_8 FILLER_43_1736 ();
 sg13g2_decap_8 FILLER_43_1743 ();
 sg13g2_decap_4 FILLER_43_1750 ();
 sg13g2_fill_1 FILLER_43_1754 ();
 sg13g2_fill_1 FILLER_43_1781 ();
 sg13g2_decap_4 FILLER_43_1789 ();
 sg13g2_fill_2 FILLER_43_1793 ();
 sg13g2_fill_2 FILLER_43_1799 ();
 sg13g2_fill_1 FILLER_43_1801 ();
 sg13g2_decap_8 FILLER_43_1812 ();
 sg13g2_decap_8 FILLER_43_1819 ();
 sg13g2_decap_8 FILLER_43_1826 ();
 sg13g2_decap_8 FILLER_43_1833 ();
 sg13g2_decap_8 FILLER_43_1840 ();
 sg13g2_fill_2 FILLER_43_1855 ();
 sg13g2_fill_1 FILLER_43_1857 ();
 sg13g2_fill_1 FILLER_43_1879 ();
 sg13g2_fill_2 FILLER_43_1885 ();
 sg13g2_decap_4 FILLER_43_1893 ();
 sg13g2_fill_1 FILLER_43_1901 ();
 sg13g2_decap_4 FILLER_43_1918 ();
 sg13g2_fill_2 FILLER_43_1959 ();
 sg13g2_decap_8 FILLER_43_1965 ();
 sg13g2_decap_8 FILLER_43_1972 ();
 sg13g2_fill_1 FILLER_43_1979 ();
 sg13g2_fill_2 FILLER_43_2034 ();
 sg13g2_fill_1 FILLER_43_2036 ();
 sg13g2_decap_8 FILLER_43_2050 ();
 sg13g2_decap_4 FILLER_43_2057 ();
 sg13g2_fill_2 FILLER_43_2061 ();
 sg13g2_fill_1 FILLER_43_2076 ();
 sg13g2_fill_1 FILLER_43_2087 ();
 sg13g2_fill_1 FILLER_43_2093 ();
 sg13g2_fill_2 FILLER_43_2098 ();
 sg13g2_decap_8 FILLER_43_2104 ();
 sg13g2_decap_8 FILLER_43_2111 ();
 sg13g2_fill_2 FILLER_43_2118 ();
 sg13g2_fill_1 FILLER_43_2124 ();
 sg13g2_fill_2 FILLER_43_2151 ();
 sg13g2_fill_1 FILLER_43_2183 ();
 sg13g2_fill_2 FILLER_43_2188 ();
 sg13g2_fill_1 FILLER_43_2194 ();
 sg13g2_fill_2 FILLER_43_2212 ();
 sg13g2_fill_1 FILLER_43_2224 ();
 sg13g2_fill_1 FILLER_43_2254 ();
 sg13g2_fill_2 FILLER_43_2271 ();
 sg13g2_fill_1 FILLER_43_2295 ();
 sg13g2_fill_1 FILLER_43_2312 ();
 sg13g2_fill_1 FILLER_43_2359 ();
 sg13g2_fill_2 FILLER_43_2374 ();
 sg13g2_fill_2 FILLER_43_2442 ();
 sg13g2_fill_1 FILLER_43_2444 ();
 sg13g2_fill_2 FILLER_43_2497 ();
 sg13g2_fill_1 FILLER_43_2532 ();
 sg13g2_decap_8 FILLER_43_2603 ();
 sg13g2_decap_8 FILLER_43_2610 ();
 sg13g2_decap_8 FILLER_43_2617 ();
 sg13g2_decap_8 FILLER_43_2624 ();
 sg13g2_decap_8 FILLER_43_2631 ();
 sg13g2_decap_8 FILLER_43_2638 ();
 sg13g2_decap_8 FILLER_43_2645 ();
 sg13g2_decap_8 FILLER_43_2652 ();
 sg13g2_decap_8 FILLER_43_2659 ();
 sg13g2_decap_4 FILLER_43_2666 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_8 FILLER_44_42 ();
 sg13g2_fill_2 FILLER_44_49 ();
 sg13g2_decap_8 FILLER_44_58 ();
 sg13g2_fill_1 FILLER_44_65 ();
 sg13g2_fill_2 FILLER_44_114 ();
 sg13g2_decap_4 FILLER_44_151 ();
 sg13g2_decap_4 FILLER_44_170 ();
 sg13g2_decap_8 FILLER_44_178 ();
 sg13g2_decap_8 FILLER_44_185 ();
 sg13g2_decap_8 FILLER_44_192 ();
 sg13g2_decap_4 FILLER_44_199 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_fill_1 FILLER_44_235 ();
 sg13g2_decap_4 FILLER_44_276 ();
 sg13g2_fill_1 FILLER_44_284 ();
 sg13g2_fill_2 FILLER_44_289 ();
 sg13g2_fill_2 FILLER_44_353 ();
 sg13g2_fill_1 FILLER_44_395 ();
 sg13g2_fill_2 FILLER_44_427 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_1 FILLER_44_438 ();
 sg13g2_fill_2 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_490 ();
 sg13g2_decap_8 FILLER_44_497 ();
 sg13g2_fill_2 FILLER_44_504 ();
 sg13g2_fill_1 FILLER_44_506 ();
 sg13g2_fill_1 FILLER_44_520 ();
 sg13g2_decap_8 FILLER_44_547 ();
 sg13g2_decap_8 FILLER_44_554 ();
 sg13g2_decap_8 FILLER_44_561 ();
 sg13g2_decap_8 FILLER_44_568 ();
 sg13g2_decap_8 FILLER_44_575 ();
 sg13g2_fill_2 FILLER_44_592 ();
 sg13g2_fill_1 FILLER_44_594 ();
 sg13g2_fill_2 FILLER_44_598 ();
 sg13g2_fill_1 FILLER_44_600 ();
 sg13g2_fill_2 FILLER_44_657 ();
 sg13g2_fill_1 FILLER_44_659 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_fill_2 FILLER_44_702 ();
 sg13g2_fill_2 FILLER_44_735 ();
 sg13g2_decap_8 FILLER_44_786 ();
 sg13g2_decap_4 FILLER_44_793 ();
 sg13g2_fill_1 FILLER_44_797 ();
 sg13g2_fill_1 FILLER_44_856 ();
 sg13g2_fill_1 FILLER_44_878 ();
 sg13g2_fill_1 FILLER_44_889 ();
 sg13g2_fill_2 FILLER_44_950 ();
 sg13g2_decap_8 FILLER_44_978 ();
 sg13g2_decap_4 FILLER_44_1006 ();
 sg13g2_decap_8 FILLER_44_1014 ();
 sg13g2_decap_8 FILLER_44_1026 ();
 sg13g2_decap_8 FILLER_44_1033 ();
 sg13g2_decap_4 FILLER_44_1040 ();
 sg13g2_fill_2 FILLER_44_1044 ();
 sg13g2_fill_1 FILLER_44_1051 ();
 sg13g2_fill_2 FILLER_44_1078 ();
 sg13g2_fill_2 FILLER_44_1084 ();
 sg13g2_decap_4 FILLER_44_1112 ();
 sg13g2_fill_2 FILLER_44_1124 ();
 sg13g2_decap_8 FILLER_44_1130 ();
 sg13g2_decap_8 FILLER_44_1137 ();
 sg13g2_decap_4 FILLER_44_1153 ();
 sg13g2_fill_2 FILLER_44_1157 ();
 sg13g2_fill_1 FILLER_44_1163 ();
 sg13g2_fill_1 FILLER_44_1168 ();
 sg13g2_fill_1 FILLER_44_1174 ();
 sg13g2_fill_2 FILLER_44_1179 ();
 sg13g2_fill_2 FILLER_44_1185 ();
 sg13g2_decap_4 FILLER_44_1195 ();
 sg13g2_fill_1 FILLER_44_1199 ();
 sg13g2_fill_1 FILLER_44_1224 ();
 sg13g2_fill_1 FILLER_44_1244 ();
 sg13g2_fill_1 FILLER_44_1255 ();
 sg13g2_decap_8 FILLER_44_1305 ();
 sg13g2_decap_4 FILLER_44_1312 ();
 sg13g2_fill_2 FILLER_44_1316 ();
 sg13g2_decap_4 FILLER_44_1329 ();
 sg13g2_fill_1 FILLER_44_1333 ();
 sg13g2_fill_1 FILLER_44_1348 ();
 sg13g2_decap_8 FILLER_44_1353 ();
 sg13g2_decap_8 FILLER_44_1360 ();
 sg13g2_decap_8 FILLER_44_1367 ();
 sg13g2_decap_8 FILLER_44_1388 ();
 sg13g2_decap_4 FILLER_44_1395 ();
 sg13g2_fill_1 FILLER_44_1399 ();
 sg13g2_decap_4 FILLER_44_1404 ();
 sg13g2_decap_8 FILLER_44_1412 ();
 sg13g2_fill_2 FILLER_44_1428 ();
 sg13g2_fill_1 FILLER_44_1448 ();
 sg13g2_fill_1 FILLER_44_1454 ();
 sg13g2_fill_1 FILLER_44_1469 ();
 sg13g2_fill_2 FILLER_44_1477 ();
 sg13g2_fill_2 FILLER_44_1490 ();
 sg13g2_fill_1 FILLER_44_1504 ();
 sg13g2_fill_1 FILLER_44_1516 ();
 sg13g2_fill_2 FILLER_44_1534 ();
 sg13g2_decap_4 FILLER_44_1549 ();
 sg13g2_fill_2 FILLER_44_1569 ();
 sg13g2_decap_4 FILLER_44_1587 ();
 sg13g2_fill_1 FILLER_44_1605 ();
 sg13g2_fill_2 FILLER_44_1621 ();
 sg13g2_decap_8 FILLER_44_1662 ();
 sg13g2_fill_2 FILLER_44_1669 ();
 sg13g2_decap_4 FILLER_44_1679 ();
 sg13g2_fill_2 FILLER_44_1683 ();
 sg13g2_fill_1 FILLER_44_1711 ();
 sg13g2_fill_2 FILLER_44_1723 ();
 sg13g2_decap_8 FILLER_44_1781 ();
 sg13g2_decap_8 FILLER_44_1824 ();
 sg13g2_decap_8 FILLER_44_1831 ();
 sg13g2_decap_8 FILLER_44_1838 ();
 sg13g2_fill_1 FILLER_44_1850 ();
 sg13g2_fill_1 FILLER_44_1862 ();
 sg13g2_fill_1 FILLER_44_1886 ();
 sg13g2_fill_1 FILLER_44_1891 ();
 sg13g2_fill_1 FILLER_44_1901 ();
 sg13g2_fill_2 FILLER_44_1932 ();
 sg13g2_fill_2 FILLER_44_1942 ();
 sg13g2_fill_1 FILLER_44_1944 ();
 sg13g2_decap_4 FILLER_44_1953 ();
 sg13g2_fill_1 FILLER_44_1957 ();
 sg13g2_decap_8 FILLER_44_1967 ();
 sg13g2_fill_2 FILLER_44_1974 ();
 sg13g2_fill_1 FILLER_44_2011 ();
 sg13g2_fill_2 FILLER_44_2025 ();
 sg13g2_fill_2 FILLER_44_2061 ();
 sg13g2_fill_1 FILLER_44_2063 ();
 sg13g2_fill_2 FILLER_44_2129 ();
 sg13g2_fill_1 FILLER_44_2151 ();
 sg13g2_fill_2 FILLER_44_2208 ();
 sg13g2_fill_1 FILLER_44_2256 ();
 sg13g2_fill_1 FILLER_44_2293 ();
 sg13g2_fill_2 FILLER_44_2386 ();
 sg13g2_decap_4 FILLER_44_2401 ();
 sg13g2_fill_1 FILLER_44_2405 ();
 sg13g2_fill_1 FILLER_44_2432 ();
 sg13g2_fill_1 FILLER_44_2439 ();
 sg13g2_fill_2 FILLER_44_2480 ();
 sg13g2_fill_1 FILLER_44_2591 ();
 sg13g2_decap_8 FILLER_44_2618 ();
 sg13g2_decap_8 FILLER_44_2625 ();
 sg13g2_decap_8 FILLER_44_2632 ();
 sg13g2_decap_8 FILLER_44_2639 ();
 sg13g2_decap_8 FILLER_44_2646 ();
 sg13g2_decap_8 FILLER_44_2653 ();
 sg13g2_decap_8 FILLER_44_2660 ();
 sg13g2_fill_2 FILLER_44_2667 ();
 sg13g2_fill_1 FILLER_44_2669 ();
 sg13g2_fill_1 FILLER_45_38 ();
 sg13g2_fill_1 FILLER_45_59 ();
 sg13g2_fill_2 FILLER_45_64 ();
 sg13g2_fill_2 FILLER_45_107 ();
 sg13g2_fill_2 FILLER_45_114 ();
 sg13g2_decap_4 FILLER_45_133 ();
 sg13g2_fill_2 FILLER_45_151 ();
 sg13g2_decap_4 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_162 ();
 sg13g2_fill_2 FILLER_45_176 ();
 sg13g2_decap_8 FILLER_45_204 ();
 sg13g2_fill_1 FILLER_45_211 ();
 sg13g2_decap_8 FILLER_45_216 ();
 sg13g2_decap_4 FILLER_45_223 ();
 sg13g2_fill_1 FILLER_45_227 ();
 sg13g2_decap_8 FILLER_45_234 ();
 sg13g2_decap_8 FILLER_45_241 ();
 sg13g2_decap_8 FILLER_45_248 ();
 sg13g2_fill_2 FILLER_45_255 ();
 sg13g2_fill_1 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_302 ();
 sg13g2_fill_2 FILLER_45_306 ();
 sg13g2_fill_1 FILLER_45_334 ();
 sg13g2_fill_1 FILLER_45_345 ();
 sg13g2_decap_4 FILLER_45_387 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_fill_2 FILLER_45_409 ();
 sg13g2_fill_2 FILLER_45_419 ();
 sg13g2_fill_1 FILLER_45_421 ();
 sg13g2_decap_4 FILLER_45_455 ();
 sg13g2_fill_1 FILLER_45_459 ();
 sg13g2_fill_2 FILLER_45_486 ();
 sg13g2_fill_1 FILLER_45_488 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_fill_1 FILLER_45_504 ();
 sg13g2_fill_1 FILLER_45_518 ();
 sg13g2_decap_4 FILLER_45_600 ();
 sg13g2_fill_2 FILLER_45_604 ();
 sg13g2_decap_4 FILLER_45_629 ();
 sg13g2_fill_1 FILLER_45_648 ();
 sg13g2_decap_4 FILLER_45_668 ();
 sg13g2_decap_8 FILLER_45_698 ();
 sg13g2_fill_2 FILLER_45_705 ();
 sg13g2_fill_1 FILLER_45_707 ();
 sg13g2_fill_1 FILLER_45_713 ();
 sg13g2_fill_2 FILLER_45_733 ();
 sg13g2_fill_1 FILLER_45_754 ();
 sg13g2_fill_2 FILLER_45_774 ();
 sg13g2_fill_2 FILLER_45_827 ();
 sg13g2_fill_1 FILLER_45_859 ();
 sg13g2_fill_2 FILLER_45_886 ();
 sg13g2_fill_1 FILLER_45_888 ();
 sg13g2_fill_1 FILLER_45_989 ();
 sg13g2_decap_8 FILLER_45_995 ();
 sg13g2_decap_4 FILLER_45_1002 ();
 sg13g2_decap_8 FILLER_45_1011 ();
 sg13g2_decap_4 FILLER_45_1054 ();
 sg13g2_fill_1 FILLER_45_1058 ();
 sg13g2_fill_2 FILLER_45_1064 ();
 sg13g2_fill_1 FILLER_45_1087 ();
 sg13g2_decap_8 FILLER_45_1097 ();
 sg13g2_decap_8 FILLER_45_1104 ();
 sg13g2_fill_1 FILLER_45_1146 ();
 sg13g2_decap_8 FILLER_45_1152 ();
 sg13g2_fill_1 FILLER_45_1167 ();
 sg13g2_fill_2 FILLER_45_1173 ();
 sg13g2_fill_1 FILLER_45_1175 ();
 sg13g2_fill_2 FILLER_45_1185 ();
 sg13g2_fill_1 FILLER_45_1187 ();
 sg13g2_decap_4 FILLER_45_1192 ();
 sg13g2_fill_1 FILLER_45_1196 ();
 sg13g2_fill_1 FILLER_45_1269 ();
 sg13g2_fill_1 FILLER_45_1275 ();
 sg13g2_decap_8 FILLER_45_1290 ();
 sg13g2_decap_8 FILLER_45_1297 ();
 sg13g2_decap_4 FILLER_45_1308 ();
 sg13g2_fill_2 FILLER_45_1312 ();
 sg13g2_fill_2 FILLER_45_1318 ();
 sg13g2_fill_2 FILLER_45_1329 ();
 sg13g2_fill_1 FILLER_45_1331 ();
 sg13g2_decap_8 FILLER_45_1363 ();
 sg13g2_decap_4 FILLER_45_1370 ();
 sg13g2_fill_2 FILLER_45_1374 ();
 sg13g2_fill_2 FILLER_45_1380 ();
 sg13g2_fill_2 FILLER_45_1389 ();
 sg13g2_fill_2 FILLER_45_1417 ();
 sg13g2_fill_1 FILLER_45_1419 ();
 sg13g2_decap_4 FILLER_45_1424 ();
 sg13g2_fill_2 FILLER_45_1428 ();
 sg13g2_fill_1 FILLER_45_1479 ();
 sg13g2_fill_1 FILLER_45_1492 ();
 sg13g2_fill_2 FILLER_45_1501 ();
 sg13g2_fill_2 FILLER_45_1513 ();
 sg13g2_fill_2 FILLER_45_1526 ();
 sg13g2_decap_8 FILLER_45_1541 ();
 sg13g2_decap_4 FILLER_45_1548 ();
 sg13g2_decap_8 FILLER_45_1557 ();
 sg13g2_decap_8 FILLER_45_1564 ();
 sg13g2_fill_1 FILLER_45_1571 ();
 sg13g2_decap_8 FILLER_45_1576 ();
 sg13g2_decap_4 FILLER_45_1583 ();
 sg13g2_decap_4 FILLER_45_1594 ();
 sg13g2_decap_4 FILLER_45_1602 ();
 sg13g2_fill_1 FILLER_45_1606 ();
 sg13g2_decap_8 FILLER_45_1612 ();
 sg13g2_decap_8 FILLER_45_1619 ();
 sg13g2_fill_2 FILLER_45_1626 ();
 sg13g2_fill_1 FILLER_45_1628 ();
 sg13g2_decap_8 FILLER_45_1633 ();
 sg13g2_decap_4 FILLER_45_1640 ();
 sg13g2_fill_1 FILLER_45_1644 ();
 sg13g2_decap_8 FILLER_45_1649 ();
 sg13g2_decap_8 FILLER_45_1656 ();
 sg13g2_decap_8 FILLER_45_1663 ();
 sg13g2_fill_1 FILLER_45_1670 ();
 sg13g2_fill_1 FILLER_45_1678 ();
 sg13g2_decap_8 FILLER_45_1692 ();
 sg13g2_decap_8 FILLER_45_1699 ();
 sg13g2_fill_1 FILLER_45_1706 ();
 sg13g2_fill_1 FILLER_45_1711 ();
 sg13g2_fill_2 FILLER_45_1755 ();
 sg13g2_fill_2 FILLER_45_1761 ();
 sg13g2_decap_4 FILLER_45_1773 ();
 sg13g2_fill_1 FILLER_45_1781 ();
 sg13g2_fill_2 FILLER_45_1787 ();
 sg13g2_decap_8 FILLER_45_1799 ();
 sg13g2_decap_4 FILLER_45_1832 ();
 sg13g2_fill_1 FILLER_45_1836 ();
 sg13g2_decap_8 FILLER_45_1860 ();
 sg13g2_decap_4 FILLER_45_1877 ();
 sg13g2_fill_1 FILLER_45_1887 ();
 sg13g2_fill_1 FILLER_45_1892 ();
 sg13g2_fill_1 FILLER_45_1898 ();
 sg13g2_decap_4 FILLER_45_1908 ();
 sg13g2_fill_1 FILLER_45_1912 ();
 sg13g2_fill_2 FILLER_45_1927 ();
 sg13g2_fill_1 FILLER_45_1939 ();
 sg13g2_decap_8 FILLER_45_1965 ();
 sg13g2_decap_8 FILLER_45_1972 ();
 sg13g2_decap_4 FILLER_45_1979 ();
 sg13g2_fill_2 FILLER_45_1983 ();
 sg13g2_fill_2 FILLER_45_1994 ();
 sg13g2_fill_1 FILLER_45_2000 ();
 sg13g2_fill_2 FILLER_45_2073 ();
 sg13g2_fill_2 FILLER_45_2080 ();
 sg13g2_fill_2 FILLER_45_2097 ();
 sg13g2_fill_1 FILLER_45_2099 ();
 sg13g2_fill_2 FILLER_45_2126 ();
 sg13g2_fill_2 FILLER_45_2140 ();
 sg13g2_fill_1 FILLER_45_2142 ();
 sg13g2_fill_1 FILLER_45_2148 ();
 sg13g2_fill_1 FILLER_45_2248 ();
 sg13g2_fill_1 FILLER_45_2273 ();
 sg13g2_fill_1 FILLER_45_2311 ();
 sg13g2_fill_1 FILLER_45_2356 ();
 sg13g2_decap_4 FILLER_45_2419 ();
 sg13g2_fill_2 FILLER_45_2423 ();
 sg13g2_decap_4 FILLER_45_2435 ();
 sg13g2_fill_1 FILLER_45_2444 ();
 sg13g2_decap_8 FILLER_45_2449 ();
 sg13g2_decap_8 FILLER_45_2456 ();
 sg13g2_fill_1 FILLER_45_2463 ();
 sg13g2_fill_2 FILLER_45_2477 ();
 sg13g2_fill_1 FILLER_45_2479 ();
 sg13g2_decap_8 FILLER_45_2484 ();
 sg13g2_decap_4 FILLER_45_2491 ();
 sg13g2_fill_1 FILLER_45_2495 ();
 sg13g2_fill_1 FILLER_45_2499 ();
 sg13g2_decap_4 FILLER_45_2581 ();
 sg13g2_fill_2 FILLER_45_2585 ();
 sg13g2_decap_8 FILLER_45_2613 ();
 sg13g2_decap_8 FILLER_45_2620 ();
 sg13g2_decap_8 FILLER_45_2627 ();
 sg13g2_decap_8 FILLER_45_2634 ();
 sg13g2_decap_8 FILLER_45_2641 ();
 sg13g2_decap_8 FILLER_45_2648 ();
 sg13g2_decap_8 FILLER_45_2655 ();
 sg13g2_decap_8 FILLER_45_2662 ();
 sg13g2_fill_1 FILLER_45_2669 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_4 ();
 sg13g2_fill_1 FILLER_46_48 ();
 sg13g2_fill_2 FILLER_46_72 ();
 sg13g2_fill_1 FILLER_46_74 ();
 sg13g2_fill_2 FILLER_46_102 ();
 sg13g2_fill_2 FILLER_46_114 ();
 sg13g2_fill_1 FILLER_46_116 ();
 sg13g2_fill_2 FILLER_46_248 ();
 sg13g2_decap_4 FILLER_46_280 ();
 sg13g2_fill_1 FILLER_46_284 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_304 ();
 sg13g2_fill_1 FILLER_46_314 ();
 sg13g2_fill_2 FILLER_46_319 ();
 sg13g2_fill_2 FILLER_46_342 ();
 sg13g2_fill_2 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_380 ();
 sg13g2_fill_1 FILLER_46_394 ();
 sg13g2_fill_2 FILLER_46_410 ();
 sg13g2_fill_1 FILLER_46_412 ();
 sg13g2_fill_2 FILLER_46_453 ();
 sg13g2_fill_1 FILLER_46_486 ();
 sg13g2_fill_1 FILLER_46_539 ();
 sg13g2_fill_2 FILLER_46_570 ();
 sg13g2_fill_2 FILLER_46_576 ();
 sg13g2_fill_1 FILLER_46_598 ();
 sg13g2_decap_4 FILLER_46_622 ();
 sg13g2_fill_1 FILLER_46_626 ();
 sg13g2_decap_4 FILLER_46_631 ();
 sg13g2_decap_4 FILLER_46_641 ();
 sg13g2_fill_1 FILLER_46_690 ();
 sg13g2_decap_8 FILLER_46_695 ();
 sg13g2_decap_8 FILLER_46_702 ();
 sg13g2_decap_8 FILLER_46_709 ();
 sg13g2_decap_8 FILLER_46_716 ();
 sg13g2_decap_4 FILLER_46_723 ();
 sg13g2_fill_2 FILLER_46_727 ();
 sg13g2_decap_4 FILLER_46_742 ();
 sg13g2_decap_8 FILLER_46_750 ();
 sg13g2_decap_8 FILLER_46_757 ();
 sg13g2_fill_2 FILLER_46_780 ();
 sg13g2_fill_1 FILLER_46_862 ();
 sg13g2_decap_8 FILLER_46_897 ();
 sg13g2_decap_8 FILLER_46_933 ();
 sg13g2_decap_8 FILLER_46_940 ();
 sg13g2_fill_2 FILLER_46_947 ();
 sg13g2_fill_1 FILLER_46_949 ();
 sg13g2_fill_2 FILLER_46_980 ();
 sg13g2_fill_2 FILLER_46_999 ();
 sg13g2_decap_4 FILLER_46_1009 ();
 sg13g2_fill_1 FILLER_46_1013 ();
 sg13g2_decap_8 FILLER_46_1050 ();
 sg13g2_fill_2 FILLER_46_1057 ();
 sg13g2_decap_4 FILLER_46_1064 ();
 sg13g2_fill_1 FILLER_46_1093 ();
 sg13g2_fill_2 FILLER_46_1098 ();
 sg13g2_fill_1 FILLER_46_1109 ();
 sg13g2_decap_8 FILLER_46_1145 ();
 sg13g2_decap_8 FILLER_46_1157 ();
 sg13g2_decap_8 FILLER_46_1164 ();
 sg13g2_decap_8 FILLER_46_1171 ();
 sg13g2_fill_1 FILLER_46_1178 ();
 sg13g2_fill_2 FILLER_46_1210 ();
 sg13g2_fill_2 FILLER_46_1242 ();
 sg13g2_fill_2 FILLER_46_1281 ();
 sg13g2_fill_1 FILLER_46_1283 ();
 sg13g2_fill_2 FILLER_46_1288 ();
 sg13g2_fill_2 FILLER_46_1294 ();
 sg13g2_fill_1 FILLER_46_1296 ();
 sg13g2_fill_2 FILLER_46_1348 ();
 sg13g2_fill_2 FILLER_46_1396 ();
 sg13g2_decap_8 FILLER_46_1411 ();
 sg13g2_decap_8 FILLER_46_1418 ();
 sg13g2_decap_8 FILLER_46_1425 ();
 sg13g2_decap_4 FILLER_46_1432 ();
 sg13g2_fill_2 FILLER_46_1436 ();
 sg13g2_fill_2 FILLER_46_1453 ();
 sg13g2_fill_2 FILLER_46_1467 ();
 sg13g2_fill_1 FILLER_46_1498 ();
 sg13g2_fill_2 FILLER_46_1505 ();
 sg13g2_decap_4 FILLER_46_1514 ();
 sg13g2_fill_2 FILLER_46_1518 ();
 sg13g2_fill_2 FILLER_46_1538 ();
 sg13g2_decap_8 FILLER_46_1550 ();
 sg13g2_decap_8 FILLER_46_1557 ();
 sg13g2_fill_2 FILLER_46_1564 ();
 sg13g2_fill_1 FILLER_46_1566 ();
 sg13g2_decap_8 FILLER_46_1573 ();
 sg13g2_decap_8 FILLER_46_1580 ();
 sg13g2_fill_2 FILLER_46_1587 ();
 sg13g2_fill_1 FILLER_46_1589 ();
 sg13g2_decap_8 FILLER_46_1610 ();
 sg13g2_decap_8 FILLER_46_1617 ();
 sg13g2_fill_1 FILLER_46_1624 ();
 sg13g2_decap_8 FILLER_46_1630 ();
 sg13g2_decap_8 FILLER_46_1637 ();
 sg13g2_fill_2 FILLER_46_1644 ();
 sg13g2_fill_1 FILLER_46_1646 ();
 sg13g2_decap_4 FILLER_46_1651 ();
 sg13g2_fill_2 FILLER_46_1655 ();
 sg13g2_decap_4 FILLER_46_1666 ();
 sg13g2_fill_1 FILLER_46_1693 ();
 sg13g2_fill_1 FILLER_46_1705 ();
 sg13g2_fill_2 FILLER_46_1719 ();
 sg13g2_fill_1 FILLER_46_1730 ();
 sg13g2_decap_8 FILLER_46_1757 ();
 sg13g2_fill_1 FILLER_46_1764 ();
 sg13g2_fill_2 FILLER_46_1791 ();
 sg13g2_fill_1 FILLER_46_1793 ();
 sg13g2_fill_1 FILLER_46_1803 ();
 sg13g2_fill_1 FILLER_46_1830 ();
 sg13g2_fill_2 FILLER_46_1836 ();
 sg13g2_fill_1 FILLER_46_1838 ();
 sg13g2_decap_8 FILLER_46_1854 ();
 sg13g2_fill_2 FILLER_46_1904 ();
 sg13g2_fill_1 FILLER_46_1906 ();
 sg13g2_fill_2 FILLER_46_1973 ();
 sg13g2_decap_8 FILLER_46_1983 ();
 sg13g2_decap_4 FILLER_46_1990 ();
 sg13g2_fill_1 FILLER_46_2009 ();
 sg13g2_fill_1 FILLER_46_2028 ();
 sg13g2_fill_2 FILLER_46_2071 ();
 sg13g2_fill_1 FILLER_46_2078 ();
 sg13g2_fill_1 FILLER_46_2096 ();
 sg13g2_fill_2 FILLER_46_2102 ();
 sg13g2_fill_1 FILLER_46_2110 ();
 sg13g2_fill_1 FILLER_46_2128 ();
 sg13g2_fill_1 FILLER_46_2155 ();
 sg13g2_fill_1 FILLER_46_2160 ();
 sg13g2_fill_1 FILLER_46_2186 ();
 sg13g2_fill_2 FILLER_46_2219 ();
 sg13g2_fill_2 FILLER_46_2293 ();
 sg13g2_fill_1 FILLER_46_2397 ();
 sg13g2_fill_2 FILLER_46_2417 ();
 sg13g2_fill_2 FILLER_46_2423 ();
 sg13g2_fill_1 FILLER_46_2425 ();
 sg13g2_decap_8 FILLER_46_2462 ();
 sg13g2_fill_1 FILLER_46_2469 ();
 sg13g2_fill_1 FILLER_46_2526 ();
 sg13g2_fill_1 FILLER_46_2550 ();
 sg13g2_fill_2 FILLER_46_2557 ();
 sg13g2_fill_2 FILLER_46_2565 ();
 sg13g2_fill_2 FILLER_46_2603 ();
 sg13g2_fill_1 FILLER_46_2605 ();
 sg13g2_decap_8 FILLER_46_2610 ();
 sg13g2_decap_8 FILLER_46_2617 ();
 sg13g2_decap_8 FILLER_46_2624 ();
 sg13g2_decap_8 FILLER_46_2631 ();
 sg13g2_decap_8 FILLER_46_2638 ();
 sg13g2_decap_8 FILLER_46_2645 ();
 sg13g2_decap_8 FILLER_46_2652 ();
 sg13g2_decap_8 FILLER_46_2659 ();
 sg13g2_decap_4 FILLER_46_2666 ();
 sg13g2_decap_4 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_113 ();
 sg13g2_fill_2 FILLER_47_119 ();
 sg13g2_fill_1 FILLER_47_142 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_fill_1 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_214 ();
 sg13g2_fill_1 FILLER_47_216 ();
 sg13g2_fill_2 FILLER_47_228 ();
 sg13g2_fill_1 FILLER_47_240 ();
 sg13g2_fill_1 FILLER_47_374 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_fill_2 FILLER_47_441 ();
 sg13g2_fill_1 FILLER_47_443 ();
 sg13g2_fill_2 FILLER_47_448 ();
 sg13g2_decap_4 FILLER_47_455 ();
 sg13g2_fill_2 FILLER_47_459 ();
 sg13g2_decap_4 FILLER_47_465 ();
 sg13g2_fill_2 FILLER_47_499 ();
 sg13g2_fill_2 FILLER_47_506 ();
 sg13g2_fill_1 FILLER_47_508 ();
 sg13g2_fill_2 FILLER_47_514 ();
 sg13g2_fill_2 FILLER_47_550 ();
 sg13g2_fill_2 FILLER_47_591 ();
 sg13g2_fill_1 FILLER_47_609 ();
 sg13g2_fill_2 FILLER_47_614 ();
 sg13g2_fill_1 FILLER_47_626 ();
 sg13g2_decap_8 FILLER_47_631 ();
 sg13g2_fill_2 FILLER_47_638 ();
 sg13g2_fill_2 FILLER_47_654 ();
 sg13g2_fill_1 FILLER_47_656 ();
 sg13g2_fill_2 FILLER_47_683 ();
 sg13g2_fill_2 FILLER_47_700 ();
 sg13g2_decap_4 FILLER_47_726 ();
 sg13g2_decap_8 FILLER_47_738 ();
 sg13g2_decap_4 FILLER_47_745 ();
 sg13g2_fill_2 FILLER_47_753 ();
 sg13g2_fill_1 FILLER_47_773 ();
 sg13g2_fill_1 FILLER_47_806 ();
 sg13g2_fill_1 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_930 ();
 sg13g2_decap_8 FILLER_47_937 ();
 sg13g2_decap_4 FILLER_47_954 ();
 sg13g2_decap_8 FILLER_47_962 ();
 sg13g2_fill_1 FILLER_47_969 ();
 sg13g2_fill_1 FILLER_47_1014 ();
 sg13g2_decap_8 FILLER_47_1020 ();
 sg13g2_fill_2 FILLER_47_1027 ();
 sg13g2_decap_4 FILLER_47_1037 ();
 sg13g2_fill_2 FILLER_47_1041 ();
 sg13g2_fill_2 FILLER_47_1107 ();
 sg13g2_decap_4 FILLER_47_1122 ();
 sg13g2_fill_1 FILLER_47_1138 ();
 sg13g2_fill_2 FILLER_47_1148 ();
 sg13g2_decap_4 FILLER_47_1180 ();
 sg13g2_fill_1 FILLER_47_1184 ();
 sg13g2_decap_4 FILLER_47_1193 ();
 sg13g2_fill_1 FILLER_47_1206 ();
 sg13g2_fill_2 FILLER_47_1215 ();
 sg13g2_fill_2 FILLER_47_1221 ();
 sg13g2_fill_2 FILLER_47_1231 ();
 sg13g2_fill_1 FILLER_47_1268 ();
 sg13g2_decap_4 FILLER_47_1310 ();
 sg13g2_decap_4 FILLER_47_1319 ();
 sg13g2_decap_4 FILLER_47_1327 ();
 sg13g2_fill_2 FILLER_47_1331 ();
 sg13g2_fill_1 FILLER_47_1337 ();
 sg13g2_decap_4 FILLER_47_1426 ();
 sg13g2_fill_2 FILLER_47_1430 ();
 sg13g2_fill_2 FILLER_47_1467 ();
 sg13g2_decap_4 FILLER_47_1525 ();
 sg13g2_fill_1 FILLER_47_1529 ();
 sg13g2_decap_4 FILLER_47_1572 ();
 sg13g2_fill_2 FILLER_47_1576 ();
 sg13g2_decap_4 FILLER_47_1581 ();
 sg13g2_fill_2 FILLER_47_1585 ();
 sg13g2_fill_2 FILLER_47_1596 ();
 sg13g2_decap_4 FILLER_47_1608 ();
 sg13g2_fill_1 FILLER_47_1612 ();
 sg13g2_fill_2 FILLER_47_1620 ();
 sg13g2_fill_1 FILLER_47_1622 ();
 sg13g2_fill_1 FILLER_47_1641 ();
 sg13g2_fill_1 FILLER_47_1652 ();
 sg13g2_fill_1 FILLER_47_1657 ();
 sg13g2_decap_4 FILLER_47_1668 ();
 sg13g2_fill_1 FILLER_47_1688 ();
 sg13g2_fill_2 FILLER_47_1693 ();
 sg13g2_fill_1 FILLER_47_1700 ();
 sg13g2_decap_4 FILLER_47_1706 ();
 sg13g2_decap_4 FILLER_47_1715 ();
 sg13g2_decap_4 FILLER_47_1724 ();
 sg13g2_fill_1 FILLER_47_1741 ();
 sg13g2_decap_4 FILLER_47_1751 ();
 sg13g2_fill_1 FILLER_47_1758 ();
 sg13g2_decap_4 FILLER_47_1765 ();
 sg13g2_fill_1 FILLER_47_1769 ();
 sg13g2_decap_4 FILLER_47_1779 ();
 sg13g2_fill_2 FILLER_47_1783 ();
 sg13g2_fill_2 FILLER_47_1815 ();
 sg13g2_fill_1 FILLER_47_1817 ();
 sg13g2_fill_2 FILLER_47_1834 ();
 sg13g2_fill_1 FILLER_47_1860 ();
 sg13g2_fill_2 FILLER_47_1885 ();
 sg13g2_fill_1 FILLER_47_1887 ();
 sg13g2_fill_2 FILLER_47_1902 ();
 sg13g2_fill_1 FILLER_47_1938 ();
 sg13g2_fill_1 FILLER_47_1944 ();
 sg13g2_fill_2 FILLER_47_1993 ();
 sg13g2_fill_1 FILLER_47_2000 ();
 sg13g2_fill_2 FILLER_47_2027 ();
 sg13g2_decap_4 FILLER_47_2035 ();
 sg13g2_fill_2 FILLER_47_2039 ();
 sg13g2_fill_1 FILLER_47_2110 ();
 sg13g2_fill_1 FILLER_47_2157 ();
 sg13g2_fill_2 FILLER_47_2196 ();
 sg13g2_fill_1 FILLER_47_2351 ();
 sg13g2_fill_1 FILLER_47_2365 ();
 sg13g2_fill_1 FILLER_47_2373 ();
 sg13g2_fill_1 FILLER_47_2393 ();
 sg13g2_fill_1 FILLER_47_2407 ();
 sg13g2_fill_1 FILLER_47_2412 ();
 sg13g2_fill_1 FILLER_47_2439 ();
 sg13g2_fill_2 FILLER_47_2455 ();
 sg13g2_fill_2 FILLER_47_2461 ();
 sg13g2_decap_4 FILLER_47_2473 ();
 sg13g2_fill_2 FILLER_47_2487 ();
 sg13g2_fill_2 FILLER_47_2499 ();
 sg13g2_decap_4 FILLER_47_2569 ();
 sg13g2_fill_2 FILLER_47_2573 ();
 sg13g2_fill_2 FILLER_47_2595 ();
 sg13g2_fill_1 FILLER_47_2597 ();
 sg13g2_decap_8 FILLER_47_2624 ();
 sg13g2_decap_8 FILLER_47_2631 ();
 sg13g2_decap_8 FILLER_47_2638 ();
 sg13g2_decap_8 FILLER_47_2645 ();
 sg13g2_decap_8 FILLER_47_2652 ();
 sg13g2_decap_8 FILLER_47_2659 ();
 sg13g2_decap_4 FILLER_47_2666 ();
 sg13g2_fill_2 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_2 ();
 sg13g2_fill_1 FILLER_48_8 ();
 sg13g2_fill_2 FILLER_48_44 ();
 sg13g2_decap_8 FILLER_48_61 ();
 sg13g2_decap_8 FILLER_48_68 ();
 sg13g2_fill_2 FILLER_48_75 ();
 sg13g2_fill_2 FILLER_48_119 ();
 sg13g2_fill_2 FILLER_48_164 ();
 sg13g2_fill_2 FILLER_48_196 ();
 sg13g2_fill_1 FILLER_48_198 ();
 sg13g2_fill_1 FILLER_48_220 ();
 sg13g2_fill_2 FILLER_48_250 ();
 sg13g2_fill_2 FILLER_48_257 ();
 sg13g2_fill_1 FILLER_48_264 ();
 sg13g2_fill_2 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_357 ();
 sg13g2_fill_1 FILLER_48_362 ();
 sg13g2_decap_8 FILLER_48_367 ();
 sg13g2_fill_1 FILLER_48_374 ();
 sg13g2_fill_2 FILLER_48_447 ();
 sg13g2_fill_1 FILLER_48_449 ();
 sg13g2_decap_8 FILLER_48_457 ();
 sg13g2_fill_2 FILLER_48_464 ();
 sg13g2_fill_1 FILLER_48_466 ();
 sg13g2_decap_8 FILLER_48_475 ();
 sg13g2_decap_8 FILLER_48_482 ();
 sg13g2_decap_8 FILLER_48_489 ();
 sg13g2_decap_4 FILLER_48_496 ();
 sg13g2_fill_2 FILLER_48_504 ();
 sg13g2_fill_1 FILLER_48_506 ();
 sg13g2_fill_1 FILLER_48_511 ();
 sg13g2_fill_1 FILLER_48_538 ();
 sg13g2_fill_2 FILLER_48_545 ();
 sg13g2_fill_1 FILLER_48_563 ();
 sg13g2_fill_2 FILLER_48_569 ();
 sg13g2_fill_2 FILLER_48_576 ();
 sg13g2_fill_1 FILLER_48_617 ();
 sg13g2_fill_2 FILLER_48_631 ();
 sg13g2_decap_8 FILLER_48_643 ();
 sg13g2_decap_8 FILLER_48_650 ();
 sg13g2_fill_1 FILLER_48_657 ();
 sg13g2_fill_1 FILLER_48_672 ();
 sg13g2_fill_2 FILLER_48_697 ();
 sg13g2_fill_2 FILLER_48_732 ();
 sg13g2_fill_2 FILLER_48_772 ();
 sg13g2_fill_1 FILLER_48_781 ();
 sg13g2_fill_1 FILLER_48_853 ();
 sg13g2_fill_2 FILLER_48_924 ();
 sg13g2_fill_1 FILLER_48_926 ();
 sg13g2_fill_1 FILLER_48_931 ();
 sg13g2_fill_1 FILLER_48_968 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_4 FILLER_48_1001 ();
 sg13g2_fill_2 FILLER_48_1009 ();
 sg13g2_fill_1 FILLER_48_1015 ();
 sg13g2_fill_1 FILLER_48_1052 ();
 sg13g2_fill_2 FILLER_48_1079 ();
 sg13g2_fill_1 FILLER_48_1107 ();
 sg13g2_fill_2 FILLER_48_1113 ();
 sg13g2_decap_8 FILLER_48_1146 ();
 sg13g2_decap_8 FILLER_48_1153 ();
 sg13g2_fill_2 FILLER_48_1160 ();
 sg13g2_fill_1 FILLER_48_1162 ();
 sg13g2_decap_4 FILLER_48_1167 ();
 sg13g2_fill_1 FILLER_48_1171 ();
 sg13g2_decap_4 FILLER_48_1176 ();
 sg13g2_fill_1 FILLER_48_1180 ();
 sg13g2_fill_2 FILLER_48_1206 ();
 sg13g2_fill_1 FILLER_48_1225 ();
 sg13g2_fill_2 FILLER_48_1255 ();
 sg13g2_decap_4 FILLER_48_1305 ();
 sg13g2_fill_1 FILLER_48_1309 ();
 sg13g2_decap_8 FILLER_48_1314 ();
 sg13g2_decap_8 FILLER_48_1321 ();
 sg13g2_decap_8 FILLER_48_1328 ();
 sg13g2_fill_2 FILLER_48_1347 ();
 sg13g2_fill_1 FILLER_48_1349 ();
 sg13g2_fill_1 FILLER_48_1374 ();
 sg13g2_decap_8 FILLER_48_1412 ();
 sg13g2_decap_8 FILLER_48_1423 ();
 sg13g2_fill_2 FILLER_48_1430 ();
 sg13g2_fill_1 FILLER_48_1432 ();
 sg13g2_fill_1 FILLER_48_1437 ();
 sg13g2_decap_4 FILLER_48_1447 ();
 sg13g2_fill_2 FILLER_48_1459 ();
 sg13g2_fill_1 FILLER_48_1470 ();
 sg13g2_fill_2 FILLER_48_1492 ();
 sg13g2_fill_1 FILLER_48_1512 ();
 sg13g2_decap_8 FILLER_48_1525 ();
 sg13g2_fill_2 FILLER_48_1532 ();
 sg13g2_fill_2 FILLER_48_1587 ();
 sg13g2_fill_2 FILLER_48_1594 ();
 sg13g2_fill_1 FILLER_48_1596 ();
 sg13g2_fill_2 FILLER_48_1602 ();
 sg13g2_decap_8 FILLER_48_1614 ();
 sg13g2_fill_2 FILLER_48_1621 ();
 sg13g2_fill_1 FILLER_48_1623 ();
 sg13g2_decap_4 FILLER_48_1637 ();
 sg13g2_fill_1 FILLER_48_1641 ();
 sg13g2_fill_1 FILLER_48_1654 ();
 sg13g2_decap_4 FILLER_48_1665 ();
 sg13g2_decap_4 FILLER_48_1687 ();
 sg13g2_fill_2 FILLER_48_1707 ();
 sg13g2_fill_1 FILLER_48_1709 ();
 sg13g2_decap_8 FILLER_48_1715 ();
 sg13g2_fill_1 FILLER_48_1722 ();
 sg13g2_fill_1 FILLER_48_1727 ();
 sg13g2_fill_2 FILLER_48_1759 ();
 sg13g2_fill_1 FILLER_48_1765 ();
 sg13g2_fill_1 FILLER_48_1792 ();
 sg13g2_fill_2 FILLER_48_1802 ();
 sg13g2_fill_1 FILLER_48_1804 ();
 sg13g2_decap_4 FILLER_48_1811 ();
 sg13g2_decap_8 FILLER_48_1823 ();
 sg13g2_decap_8 FILLER_48_1830 ();
 sg13g2_fill_2 FILLER_48_1837 ();
 sg13g2_fill_1 FILLER_48_1863 ();
 sg13g2_fill_1 FILLER_48_1869 ();
 sg13g2_fill_1 FILLER_48_1905 ();
 sg13g2_fill_1 FILLER_48_1931 ();
 sg13g2_fill_1 FILLER_48_1938 ();
 sg13g2_fill_1 FILLER_48_1948 ();
 sg13g2_fill_1 FILLER_48_1966 ();
 sg13g2_fill_1 FILLER_48_1978 ();
 sg13g2_fill_1 FILLER_48_1984 ();
 sg13g2_fill_1 FILLER_48_2011 ();
 sg13g2_fill_2 FILLER_48_2038 ();
 sg13g2_decap_4 FILLER_48_2076 ();
 sg13g2_fill_2 FILLER_48_2080 ();
 sg13g2_decap_4 FILLER_48_2095 ();
 sg13g2_fill_1 FILLER_48_2099 ();
 sg13g2_fill_1 FILLER_48_2118 ();
 sg13g2_fill_1 FILLER_48_2178 ();
 sg13g2_fill_2 FILLER_48_2214 ();
 sg13g2_fill_2 FILLER_48_2297 ();
 sg13g2_fill_1 FILLER_48_2338 ();
 sg13g2_fill_1 FILLER_48_2348 ();
 sg13g2_fill_1 FILLER_48_2371 ();
 sg13g2_fill_1 FILLER_48_2403 ();
 sg13g2_fill_2 FILLER_48_2440 ();
 sg13g2_fill_1 FILLER_48_2442 ();
 sg13g2_fill_2 FILLER_48_2477 ();
 sg13g2_fill_1 FILLER_48_2499 ();
 sg13g2_fill_1 FILLER_48_2556 ();
 sg13g2_fill_2 FILLER_48_2567 ();
 sg13g2_fill_2 FILLER_48_2579 ();
 sg13g2_fill_2 FILLER_48_2607 ();
 sg13g2_fill_1 FILLER_48_2609 ();
 sg13g2_decap_8 FILLER_48_2614 ();
 sg13g2_decap_8 FILLER_48_2621 ();
 sg13g2_decap_8 FILLER_48_2628 ();
 sg13g2_decap_8 FILLER_48_2635 ();
 sg13g2_decap_8 FILLER_48_2642 ();
 sg13g2_decap_8 FILLER_48_2649 ();
 sg13g2_decap_8 FILLER_48_2656 ();
 sg13g2_decap_8 FILLER_48_2663 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_4 ();
 sg13g2_fill_1 FILLER_49_56 ();
 sg13g2_fill_2 FILLER_49_91 ();
 sg13g2_decap_8 FILLER_49_97 ();
 sg13g2_fill_2 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_fill_2 FILLER_49_121 ();
 sg13g2_fill_1 FILLER_49_127 ();
 sg13g2_fill_1 FILLER_49_132 ();
 sg13g2_fill_1 FILLER_49_155 ();
 sg13g2_fill_2 FILLER_49_186 ();
 sg13g2_fill_2 FILLER_49_201 ();
 sg13g2_fill_1 FILLER_49_203 ();
 sg13g2_decap_8 FILLER_49_209 ();
 sg13g2_fill_1 FILLER_49_256 ();
 sg13g2_fill_1 FILLER_49_262 ();
 sg13g2_fill_1 FILLER_49_268 ();
 sg13g2_fill_1 FILLER_49_275 ();
 sg13g2_fill_1 FILLER_49_281 ();
 sg13g2_fill_1 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_293 ();
 sg13g2_fill_1 FILLER_49_300 ();
 sg13g2_fill_2 FILLER_49_310 ();
 sg13g2_fill_1 FILLER_49_319 ();
 sg13g2_fill_2 FILLER_49_328 ();
 sg13g2_fill_1 FILLER_49_336 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_372 ();
 sg13g2_decap_8 FILLER_49_379 ();
 sg13g2_fill_1 FILLER_49_386 ();
 sg13g2_fill_1 FILLER_49_392 ();
 sg13g2_fill_2 FILLER_49_397 ();
 sg13g2_fill_1 FILLER_49_404 ();
 sg13g2_fill_1 FILLER_49_410 ();
 sg13g2_fill_1 FILLER_49_421 ();
 sg13g2_fill_1 FILLER_49_430 ();
 sg13g2_fill_2 FILLER_49_439 ();
 sg13g2_fill_2 FILLER_49_446 ();
 sg13g2_fill_1 FILLER_49_448 ();
 sg13g2_decap_4 FILLER_49_497 ();
 sg13g2_fill_2 FILLER_49_501 ();
 sg13g2_fill_2 FILLER_49_555 ();
 sg13g2_fill_1 FILLER_49_577 ();
 sg13g2_fill_1 FILLER_49_605 ();
 sg13g2_fill_2 FILLER_49_623 ();
 sg13g2_decap_4 FILLER_49_650 ();
 sg13g2_fill_2 FILLER_49_669 ();
 sg13g2_fill_1 FILLER_49_697 ();
 sg13g2_fill_1 FILLER_49_706 ();
 sg13g2_fill_2 FILLER_49_778 ();
 sg13g2_fill_1 FILLER_49_822 ();
 sg13g2_fill_1 FILLER_49_834 ();
 sg13g2_fill_1 FILLER_49_853 ();
 sg13g2_decap_4 FILLER_49_890 ();
 sg13g2_fill_1 FILLER_49_898 ();
 sg13g2_fill_2 FILLER_49_914 ();
 sg13g2_fill_1 FILLER_49_916 ();
 sg13g2_fill_2 FILLER_49_947 ();
 sg13g2_fill_1 FILLER_49_970 ();
 sg13g2_fill_2 FILLER_49_985 ();
 sg13g2_fill_1 FILLER_49_987 ();
 sg13g2_fill_2 FILLER_49_1013 ();
 sg13g2_fill_2 FILLER_49_1030 ();
 sg13g2_fill_1 FILLER_49_1036 ();
 sg13g2_decap_8 FILLER_49_1041 ();
 sg13g2_decap_8 FILLER_49_1048 ();
 sg13g2_fill_2 FILLER_49_1055 ();
 sg13g2_fill_2 FILLER_49_1078 ();
 sg13g2_fill_2 FILLER_49_1085 ();
 sg13g2_decap_4 FILLER_49_1091 ();
 sg13g2_fill_1 FILLER_49_1095 ();
 sg13g2_fill_1 FILLER_49_1127 ();
 sg13g2_fill_2 FILLER_49_1132 ();
 sg13g2_fill_1 FILLER_49_1134 ();
 sg13g2_fill_2 FILLER_49_1176 ();
 sg13g2_fill_2 FILLER_49_1186 ();
 sg13g2_fill_1 FILLER_49_1196 ();
 sg13g2_fill_1 FILLER_49_1221 ();
 sg13g2_fill_1 FILLER_49_1236 ();
 sg13g2_fill_2 FILLER_49_1267 ();
 sg13g2_fill_2 FILLER_49_1278 ();
 sg13g2_fill_1 FILLER_49_1293 ();
 sg13g2_decap_4 FILLER_49_1299 ();
 sg13g2_fill_1 FILLER_49_1303 ();
 sg13g2_decap_8 FILLER_49_1308 ();
 sg13g2_fill_2 FILLER_49_1338 ();
 sg13g2_fill_1 FILLER_49_1370 ();
 sg13g2_fill_2 FILLER_49_1397 ();
 sg13g2_fill_1 FILLER_49_1425 ();
 sg13g2_decap_8 FILLER_49_1462 ();
 sg13g2_fill_1 FILLER_49_1469 ();
 sg13g2_fill_2 FILLER_49_1503 ();
 sg13g2_decap_4 FILLER_49_1522 ();
 sg13g2_fill_2 FILLER_49_1526 ();
 sg13g2_fill_2 FILLER_49_1602 ();
 sg13g2_fill_1 FILLER_49_1604 ();
 sg13g2_decap_8 FILLER_49_1613 ();
 sg13g2_decap_4 FILLER_49_1627 ();
 sg13g2_fill_1 FILLER_49_1631 ();
 sg13g2_fill_1 FILLER_49_1637 ();
 sg13g2_decap_8 FILLER_49_1660 ();
 sg13g2_decap_8 FILLER_49_1667 ();
 sg13g2_fill_1 FILLER_49_1674 ();
 sg13g2_decap_8 FILLER_49_1679 ();
 sg13g2_decap_4 FILLER_49_1686 ();
 sg13g2_fill_1 FILLER_49_1690 ();
 sg13g2_decap_8 FILLER_49_1705 ();
 sg13g2_decap_8 FILLER_49_1712 ();
 sg13g2_decap_8 FILLER_49_1719 ();
 sg13g2_decap_8 FILLER_49_1730 ();
 sg13g2_fill_2 FILLER_49_1737 ();
 sg13g2_decap_4 FILLER_49_1743 ();
 sg13g2_decap_8 FILLER_49_1780 ();
 sg13g2_decap_4 FILLER_49_1787 ();
 sg13g2_fill_2 FILLER_49_1791 ();
 sg13g2_decap_4 FILLER_49_1822 ();
 sg13g2_fill_1 FILLER_49_1826 ();
 sg13g2_decap_8 FILLER_49_1831 ();
 sg13g2_fill_2 FILLER_49_1838 ();
 sg13g2_fill_2 FILLER_49_1878 ();
 sg13g2_fill_2 FILLER_49_1884 ();
 sg13g2_fill_1 FILLER_49_1886 ();
 sg13g2_fill_2 FILLER_49_1892 ();
 sg13g2_fill_1 FILLER_49_1894 ();
 sg13g2_fill_2 FILLER_49_1898 ();
 sg13g2_fill_1 FILLER_49_1900 ();
 sg13g2_decap_8 FILLER_49_1906 ();
 sg13g2_decap_4 FILLER_49_1913 ();
 sg13g2_fill_1 FILLER_49_1938 ();
 sg13g2_fill_1 FILLER_49_1945 ();
 sg13g2_fill_1 FILLER_49_1951 ();
 sg13g2_decap_8 FILLER_49_2032 ();
 sg13g2_fill_1 FILLER_49_2039 ();
 sg13g2_fill_1 FILLER_49_2045 ();
 sg13g2_decap_4 FILLER_49_2050 ();
 sg13g2_fill_2 FILLER_49_2059 ();
 sg13g2_fill_1 FILLER_49_2061 ();
 sg13g2_decap_4 FILLER_49_2070 ();
 sg13g2_decap_4 FILLER_49_2117 ();
 sg13g2_fill_2 FILLER_49_2125 ();
 sg13g2_fill_1 FILLER_49_2127 ();
 sg13g2_fill_2 FILLER_49_2132 ();
 sg13g2_fill_1 FILLER_49_2134 ();
 sg13g2_fill_1 FILLER_49_2152 ();
 sg13g2_fill_1 FILLER_49_2162 ();
 sg13g2_fill_2 FILLER_49_2169 ();
 sg13g2_fill_1 FILLER_49_2187 ();
 sg13g2_fill_2 FILLER_49_2326 ();
 sg13g2_fill_2 FILLER_49_2334 ();
 sg13g2_fill_1 FILLER_49_2354 ();
 sg13g2_fill_1 FILLER_49_2451 ();
 sg13g2_fill_1 FILLER_49_2462 ();
 sg13g2_fill_1 FILLER_49_2473 ();
 sg13g2_decap_4 FILLER_49_2500 ();
 sg13g2_fill_1 FILLER_49_2504 ();
 sg13g2_fill_2 FILLER_49_2533 ();
 sg13g2_fill_1 FILLER_49_2539 ();
 sg13g2_fill_1 FILLER_49_2552 ();
 sg13g2_decap_8 FILLER_49_2604 ();
 sg13g2_decap_8 FILLER_49_2611 ();
 sg13g2_decap_8 FILLER_49_2618 ();
 sg13g2_decap_8 FILLER_49_2625 ();
 sg13g2_decap_8 FILLER_49_2632 ();
 sg13g2_decap_8 FILLER_49_2639 ();
 sg13g2_decap_8 FILLER_49_2646 ();
 sg13g2_decap_8 FILLER_49_2653 ();
 sg13g2_decap_8 FILLER_49_2660 ();
 sg13g2_fill_2 FILLER_49_2667 ();
 sg13g2_fill_1 FILLER_49_2669 ();
 sg13g2_decap_4 FILLER_50_0 ();
 sg13g2_fill_2 FILLER_50_4 ();
 sg13g2_fill_1 FILLER_50_44 ();
 sg13g2_fill_1 FILLER_50_53 ();
 sg13g2_fill_1 FILLER_50_88 ();
 sg13g2_fill_2 FILLER_50_102 ();
 sg13g2_fill_2 FILLER_50_107 ();
 sg13g2_fill_2 FILLER_50_114 ();
 sg13g2_decap_8 FILLER_50_120 ();
 sg13g2_fill_1 FILLER_50_127 ();
 sg13g2_fill_1 FILLER_50_132 ();
 sg13g2_decap_4 FILLER_50_178 ();
 sg13g2_fill_2 FILLER_50_192 ();
 sg13g2_decap_4 FILLER_50_220 ();
 sg13g2_fill_2 FILLER_50_237 ();
 sg13g2_fill_1 FILLER_50_268 ();
 sg13g2_fill_2 FILLER_50_278 ();
 sg13g2_fill_2 FILLER_50_306 ();
 sg13g2_fill_1 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_332 ();
 sg13g2_fill_1 FILLER_50_381 ();
 sg13g2_fill_2 FILLER_50_386 ();
 sg13g2_fill_1 FILLER_50_392 ();
 sg13g2_fill_2 FILLER_50_397 ();
 sg13g2_decap_8 FILLER_50_407 ();
 sg13g2_decap_8 FILLER_50_414 ();
 sg13g2_decap_4 FILLER_50_421 ();
 sg13g2_fill_2 FILLER_50_507 ();
 sg13g2_fill_1 FILLER_50_509 ();
 sg13g2_fill_1 FILLER_50_540 ();
 sg13g2_fill_2 FILLER_50_581 ();
 sg13g2_fill_1 FILLER_50_596 ();
 sg13g2_fill_2 FILLER_50_611 ();
 sg13g2_fill_1 FILLER_50_659 ();
 sg13g2_fill_2 FILLER_50_666 ();
 sg13g2_fill_1 FILLER_50_668 ();
 sg13g2_fill_2 FILLER_50_683 ();
 sg13g2_fill_1 FILLER_50_690 ();
 sg13g2_fill_1 FILLER_50_700 ();
 sg13g2_fill_1 FILLER_50_737 ();
 sg13g2_fill_2 FILLER_50_765 ();
 sg13g2_fill_2 FILLER_50_772 ();
 sg13g2_fill_1 FILLER_50_829 ();
 sg13g2_fill_1 FILLER_50_843 ();
 sg13g2_fill_1 FILLER_50_847 ();
 sg13g2_fill_1 FILLER_50_851 ();
 sg13g2_fill_2 FILLER_50_860 ();
 sg13g2_fill_1 FILLER_50_865 ();
 sg13g2_fill_2 FILLER_50_897 ();
 sg13g2_fill_1 FILLER_50_899 ();
 sg13g2_fill_2 FILLER_50_930 ();
 sg13g2_fill_2 FILLER_50_972 ();
 sg13g2_fill_2 FILLER_50_1021 ();
 sg13g2_fill_1 FILLER_50_1023 ();
 sg13g2_fill_2 FILLER_50_1050 ();
 sg13g2_decap_8 FILLER_50_1056 ();
 sg13g2_fill_2 FILLER_50_1066 ();
 sg13g2_decap_8 FILLER_50_1072 ();
 sg13g2_fill_2 FILLER_50_1079 ();
 sg13g2_fill_1 FILLER_50_1081 ();
 sg13g2_decap_8 FILLER_50_1087 ();
 sg13g2_decap_8 FILLER_50_1094 ();
 sg13g2_fill_2 FILLER_50_1101 ();
 sg13g2_decap_4 FILLER_50_1120 ();
 sg13g2_fill_2 FILLER_50_1160 ();
 sg13g2_fill_1 FILLER_50_1204 ();
 sg13g2_fill_1 FILLER_50_1234 ();
 sg13g2_fill_2 FILLER_50_1240 ();
 sg13g2_fill_2 FILLER_50_1246 ();
 sg13g2_decap_4 FILLER_50_1298 ();
 sg13g2_fill_1 FILLER_50_1307 ();
 sg13g2_fill_1 FILLER_50_1316 ();
 sg13g2_fill_2 FILLER_50_1322 ();
 sg13g2_fill_2 FILLER_50_1346 ();
 sg13g2_fill_1 FILLER_50_1356 ();
 sg13g2_fill_2 FILLER_50_1365 ();
 sg13g2_fill_1 FILLER_50_1381 ();
 sg13g2_fill_1 FILLER_50_1400 ();
 sg13g2_fill_2 FILLER_50_1407 ();
 sg13g2_fill_1 FILLER_50_1409 ();
 sg13g2_decap_4 FILLER_50_1414 ();
 sg13g2_fill_1 FILLER_50_1418 ();
 sg13g2_decap_4 FILLER_50_1450 ();
 sg13g2_fill_1 FILLER_50_1490 ();
 sg13g2_fill_2 FILLER_50_1499 ();
 sg13g2_fill_1 FILLER_50_1509 ();
 sg13g2_decap_4 FILLER_50_1514 ();
 sg13g2_fill_1 FILLER_50_1518 ();
 sg13g2_decap_8 FILLER_50_1523 ();
 sg13g2_fill_2 FILLER_50_1530 ();
 sg13g2_fill_1 FILLER_50_1543 ();
 sg13g2_fill_1 FILLER_50_1553 ();
 sg13g2_fill_2 FILLER_50_1558 ();
 sg13g2_fill_1 FILLER_50_1570 ();
 sg13g2_fill_1 FILLER_50_1581 ();
 sg13g2_fill_2 FILLER_50_1591 ();
 sg13g2_fill_1 FILLER_50_1598 ();
 sg13g2_fill_2 FILLER_50_1604 ();
 sg13g2_fill_2 FILLER_50_1610 ();
 sg13g2_fill_2 FILLER_50_1617 ();
 sg13g2_fill_1 FILLER_50_1619 ();
 sg13g2_decap_8 FILLER_50_1625 ();
 sg13g2_decap_4 FILLER_50_1632 ();
 sg13g2_fill_2 FILLER_50_1636 ();
 sg13g2_fill_1 FILLER_50_1658 ();
 sg13g2_decap_4 FILLER_50_1664 ();
 sg13g2_decap_8 FILLER_50_1673 ();
 sg13g2_decap_8 FILLER_50_1680 ();
 sg13g2_fill_2 FILLER_50_1687 ();
 sg13g2_fill_1 FILLER_50_1689 ();
 sg13g2_decap_8 FILLER_50_1718 ();
 sg13g2_decap_8 FILLER_50_1725 ();
 sg13g2_decap_8 FILLER_50_1732 ();
 sg13g2_fill_2 FILLER_50_1739 ();
 sg13g2_fill_1 FILLER_50_1741 ();
 sg13g2_fill_2 FILLER_50_1747 ();
 sg13g2_fill_2 FILLER_50_1753 ();
 sg13g2_fill_1 FILLER_50_1784 ();
 sg13g2_decap_4 FILLER_50_1818 ();
 sg13g2_fill_1 FILLER_50_1822 ();
 sg13g2_fill_2 FILLER_50_1829 ();
 sg13g2_fill_1 FILLER_50_1831 ();
 sg13g2_fill_1 FILLER_50_1847 ();
 sg13g2_fill_1 FILLER_50_1858 ();
 sg13g2_fill_1 FILLER_50_1864 ();
 sg13g2_decap_4 FILLER_50_1875 ();
 sg13g2_fill_1 FILLER_50_1879 ();
 sg13g2_fill_1 FILLER_50_1884 ();
 sg13g2_fill_1 FILLER_50_1908 ();
 sg13g2_fill_2 FILLER_50_1914 ();
 sg13g2_decap_4 FILLER_50_1921 ();
 sg13g2_fill_1 FILLER_50_1925 ();
 sg13g2_decap_4 FILLER_50_1952 ();
 sg13g2_fill_1 FILLER_50_1956 ();
 sg13g2_fill_2 FILLER_50_1973 ();
 sg13g2_fill_1 FILLER_50_1983 ();
 sg13g2_fill_2 FILLER_50_1989 ();
 sg13g2_fill_2 FILLER_50_1995 ();
 sg13g2_fill_1 FILLER_50_2004 ();
 sg13g2_decap_8 FILLER_50_2042 ();
 sg13g2_decap_4 FILLER_50_2049 ();
 sg13g2_fill_2 FILLER_50_2079 ();
 sg13g2_fill_2 FILLER_50_2094 ();
 sg13g2_decap_8 FILLER_50_2127 ();
 sg13g2_decap_4 FILLER_50_2134 ();
 sg13g2_fill_2 FILLER_50_2138 ();
 sg13g2_fill_1 FILLER_50_2143 ();
 sg13g2_fill_1 FILLER_50_2191 ();
 sg13g2_fill_1 FILLER_50_2221 ();
 sg13g2_fill_2 FILLER_50_2241 ();
 sg13g2_fill_1 FILLER_50_2262 ();
 sg13g2_fill_2 FILLER_50_2268 ();
 sg13g2_fill_1 FILLER_50_2298 ();
 sg13g2_fill_2 FILLER_50_2379 ();
 sg13g2_fill_2 FILLER_50_2388 ();
 sg13g2_fill_2 FILLER_50_2413 ();
 sg13g2_fill_1 FILLER_50_2432 ();
 sg13g2_fill_1 FILLER_50_2459 ();
 sg13g2_fill_1 FILLER_50_2523 ();
 sg13g2_fill_1 FILLER_50_2577 ();
 sg13g2_fill_2 FILLER_50_2591 ();
 sg13g2_decap_8 FILLER_50_2623 ();
 sg13g2_decap_8 FILLER_50_2630 ();
 sg13g2_decap_8 FILLER_50_2637 ();
 sg13g2_decap_8 FILLER_50_2644 ();
 sg13g2_decap_8 FILLER_50_2651 ();
 sg13g2_decap_8 FILLER_50_2658 ();
 sg13g2_decap_4 FILLER_50_2665 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_37 ();
 sg13g2_fill_1 FILLER_51_43 ();
 sg13g2_fill_1 FILLER_51_49 ();
 sg13g2_fill_2 FILLER_51_53 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_fill_1 FILLER_51_69 ();
 sg13g2_fill_1 FILLER_51_83 ();
 sg13g2_fill_1 FILLER_51_94 ();
 sg13g2_fill_1 FILLER_51_103 ();
 sg13g2_fill_2 FILLER_51_135 ();
 sg13g2_decap_4 FILLER_51_150 ();
 sg13g2_fill_2 FILLER_51_163 ();
 sg13g2_fill_1 FILLER_51_165 ();
 sg13g2_fill_2 FILLER_51_203 ();
 sg13g2_decap_4 FILLER_51_214 ();
 sg13g2_fill_2 FILLER_51_218 ();
 sg13g2_fill_1 FILLER_51_235 ();
 sg13g2_fill_2 FILLER_51_254 ();
 sg13g2_fill_2 FILLER_51_275 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_fill_1 FILLER_51_283 ();
 sg13g2_fill_1 FILLER_51_315 ();
 sg13g2_fill_1 FILLER_51_323 ();
 sg13g2_fill_1 FILLER_51_328 ();
 sg13g2_fill_1 FILLER_51_339 ();
 sg13g2_fill_1 FILLER_51_361 ();
 sg13g2_fill_1 FILLER_51_370 ();
 sg13g2_decap_8 FILLER_51_407 ();
 sg13g2_decap_8 FILLER_51_414 ();
 sg13g2_decap_4 FILLER_51_421 ();
 sg13g2_fill_1 FILLER_51_425 ();
 sg13g2_fill_1 FILLER_51_469 ();
 sg13g2_fill_1 FILLER_51_476 ();
 sg13g2_fill_1 FILLER_51_483 ();
 sg13g2_fill_1 FILLER_51_490 ();
 sg13g2_decap_8 FILLER_51_496 ();
 sg13g2_decap_4 FILLER_51_503 ();
 sg13g2_fill_1 FILLER_51_507 ();
 sg13g2_fill_1 FILLER_51_554 ();
 sg13g2_fill_1 FILLER_51_611 ();
 sg13g2_fill_1 FILLER_51_633 ();
 sg13g2_decap_8 FILLER_51_652 ();
 sg13g2_fill_2 FILLER_51_710 ();
 sg13g2_fill_1 FILLER_51_712 ();
 sg13g2_fill_2 FILLER_51_718 ();
 sg13g2_fill_1 FILLER_51_728 ();
 sg13g2_fill_1 FILLER_51_768 ();
 sg13g2_fill_2 FILLER_51_842 ();
 sg13g2_fill_1 FILLER_51_875 ();
 sg13g2_decap_8 FILLER_51_925 ();
 sg13g2_decap_8 FILLER_51_932 ();
 sg13g2_decap_8 FILLER_51_939 ();
 sg13g2_decap_4 FILLER_51_946 ();
 sg13g2_fill_2 FILLER_51_950 ();
 sg13g2_decap_4 FILLER_51_956 ();
 sg13g2_fill_1 FILLER_51_960 ();
 sg13g2_fill_2 FILLER_51_975 ();
 sg13g2_fill_1 FILLER_51_977 ();
 sg13g2_fill_2 FILLER_51_992 ();
 sg13g2_fill_1 FILLER_51_994 ();
 sg13g2_fill_2 FILLER_51_1021 ();
 sg13g2_fill_1 FILLER_51_1023 ();
 sg13g2_decap_4 FILLER_51_1045 ();
 sg13g2_fill_2 FILLER_51_1049 ();
 sg13g2_fill_1 FILLER_51_1056 ();
 sg13g2_fill_1 FILLER_51_1069 ();
 sg13g2_fill_2 FILLER_51_1075 ();
 sg13g2_fill_1 FILLER_51_1077 ();
 sg13g2_fill_2 FILLER_51_1084 ();
 sg13g2_fill_1 FILLER_51_1086 ();
 sg13g2_decap_4 FILLER_51_1113 ();
 sg13g2_fill_1 FILLER_51_1121 ();
 sg13g2_fill_1 FILLER_51_1168 ();
 sg13g2_fill_1 FILLER_51_1202 ();
 sg13g2_fill_2 FILLER_51_1206 ();
 sg13g2_fill_2 FILLER_51_1219 ();
 sg13g2_fill_1 FILLER_51_1256 ();
 sg13g2_fill_1 FILLER_51_1284 ();
 sg13g2_fill_2 FILLER_51_1290 ();
 sg13g2_decap_4 FILLER_51_1313 ();
 sg13g2_fill_1 FILLER_51_1317 ();
 sg13g2_fill_1 FILLER_51_1328 ();
 sg13g2_fill_2 FILLER_51_1352 ();
 sg13g2_fill_2 FILLER_51_1371 ();
 sg13g2_fill_2 FILLER_51_1384 ();
 sg13g2_fill_2 FILLER_51_1411 ();
 sg13g2_decap_8 FILLER_51_1418 ();
 sg13g2_decap_4 FILLER_51_1425 ();
 sg13g2_decap_8 FILLER_51_1433 ();
 sg13g2_fill_2 FILLER_51_1440 ();
 sg13g2_decap_4 FILLER_51_1475 ();
 sg13g2_fill_2 FILLER_51_1479 ();
 sg13g2_fill_2 FILLER_51_1485 ();
 sg13g2_fill_1 FILLER_51_1487 ();
 sg13g2_fill_1 FILLER_51_1495 ();
 sg13g2_decap_8 FILLER_51_1518 ();
 sg13g2_fill_2 FILLER_51_1535 ();
 sg13g2_fill_1 FILLER_51_1548 ();
 sg13g2_fill_1 FILLER_51_1567 ();
 sg13g2_fill_1 FILLER_51_1591 ();
 sg13g2_fill_1 FILLER_51_1609 ();
 sg13g2_fill_2 FILLER_51_1631 ();
 sg13g2_fill_1 FILLER_51_1633 ();
 sg13g2_fill_2 FILLER_51_1644 ();
 sg13g2_fill_2 FILLER_51_1653 ();
 sg13g2_fill_1 FILLER_51_1655 ();
 sg13g2_decap_8 FILLER_51_1662 ();
 sg13g2_fill_1 FILLER_51_1669 ();
 sg13g2_fill_1 FILLER_51_1697 ();
 sg13g2_decap_4 FILLER_51_1713 ();
 sg13g2_fill_2 FILLER_51_1721 ();
 sg13g2_fill_2 FILLER_51_1754 ();
 sg13g2_fill_1 FILLER_51_1756 ();
 sg13g2_fill_2 FILLER_51_1767 ();
 sg13g2_fill_1 FILLER_51_1769 ();
 sg13g2_decap_4 FILLER_51_1774 ();
 sg13g2_fill_2 FILLER_51_1778 ();
 sg13g2_fill_2 FILLER_51_1790 ();
 sg13g2_fill_2 FILLER_51_1800 ();
 sg13g2_fill_2 FILLER_51_1811 ();
 sg13g2_fill_2 FILLER_51_1818 ();
 sg13g2_fill_1 FILLER_51_1820 ();
 sg13g2_fill_1 FILLER_51_1831 ();
 sg13g2_fill_2 FILLER_51_1872 ();
 sg13g2_decap_4 FILLER_51_1879 ();
 sg13g2_fill_2 FILLER_51_1883 ();
 sg13g2_fill_2 FILLER_51_1900 ();
 sg13g2_fill_1 FILLER_51_1902 ();
 sg13g2_fill_2 FILLER_51_1906 ();
 sg13g2_fill_2 FILLER_51_1913 ();
 sg13g2_fill_1 FILLER_51_1915 ();
 sg13g2_fill_1 FILLER_51_1931 ();
 sg13g2_fill_1 FILLER_51_1937 ();
 sg13g2_fill_1 FILLER_51_1943 ();
 sg13g2_fill_1 FILLER_51_1949 ();
 sg13g2_fill_2 FILLER_51_1954 ();
 sg13g2_fill_1 FILLER_51_1956 ();
 sg13g2_fill_2 FILLER_51_1960 ();
 sg13g2_fill_2 FILLER_51_1991 ();
 sg13g2_decap_4 FILLER_51_2039 ();
 sg13g2_fill_1 FILLER_51_2043 ();
 sg13g2_decap_8 FILLER_51_2048 ();
 sg13g2_fill_1 FILLER_51_2055 ();
 sg13g2_fill_1 FILLER_51_2060 ();
 sg13g2_decap_8 FILLER_51_2112 ();
 sg13g2_decap_4 FILLER_51_2119 ();
 sg13g2_fill_2 FILLER_51_2123 ();
 sg13g2_decap_4 FILLER_51_2130 ();
 sg13g2_fill_1 FILLER_51_2142 ();
 sg13g2_fill_1 FILLER_51_2169 ();
 sg13g2_fill_1 FILLER_51_2306 ();
 sg13g2_fill_2 FILLER_51_2323 ();
 sg13g2_fill_1 FILLER_51_2361 ();
 sg13g2_fill_2 FILLER_51_2379 ();
 sg13g2_fill_2 FILLER_51_2411 ();
 sg13g2_fill_1 FILLER_51_2443 ();
 sg13g2_fill_2 FILLER_51_2479 ();
 sg13g2_fill_2 FILLER_51_2491 ();
 sg13g2_fill_2 FILLER_51_2497 ();
 sg13g2_fill_2 FILLER_51_2505 ();
 sg13g2_fill_2 FILLER_51_2513 ();
 sg13g2_fill_1 FILLER_51_2515 ();
 sg13g2_fill_1 FILLER_51_2530 ();
 sg13g2_fill_1 FILLER_51_2546 ();
 sg13g2_fill_2 FILLER_51_2552 ();
 sg13g2_fill_1 FILLER_51_2554 ();
 sg13g2_fill_2 FILLER_51_2566 ();
 sg13g2_decap_8 FILLER_51_2634 ();
 sg13g2_decap_8 FILLER_51_2641 ();
 sg13g2_decap_8 FILLER_51_2648 ();
 sg13g2_decap_8 FILLER_51_2655 ();
 sg13g2_decap_8 FILLER_51_2662 ();
 sg13g2_fill_1 FILLER_51_2669 ();
 sg13g2_decap_4 FILLER_52_0 ();
 sg13g2_decap_4 FILLER_52_44 ();
 sg13g2_fill_2 FILLER_52_48 ();
 sg13g2_decap_8 FILLER_52_53 ();
 sg13g2_fill_2 FILLER_52_60 ();
 sg13g2_fill_1 FILLER_52_62 ();
 sg13g2_decap_4 FILLER_52_68 ();
 sg13g2_decap_4 FILLER_52_140 ();
 sg13g2_fill_2 FILLER_52_144 ();
 sg13g2_fill_1 FILLER_52_150 ();
 sg13g2_decap_4 FILLER_52_187 ();
 sg13g2_fill_1 FILLER_52_191 ();
 sg13g2_decap_4 FILLER_52_198 ();
 sg13g2_fill_1 FILLER_52_202 ();
 sg13g2_fill_1 FILLER_52_209 ();
 sg13g2_decap_8 FILLER_52_214 ();
 sg13g2_fill_2 FILLER_52_221 ();
 sg13g2_fill_1 FILLER_52_223 ();
 sg13g2_decap_4 FILLER_52_238 ();
 sg13g2_fill_1 FILLER_52_242 ();
 sg13g2_decap_4 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_255 ();
 sg13g2_fill_1 FILLER_52_267 ();
 sg13g2_fill_1 FILLER_52_273 ();
 sg13g2_fill_1 FILLER_52_285 ();
 sg13g2_fill_2 FILLER_52_294 ();
 sg13g2_fill_1 FILLER_52_296 ();
 sg13g2_fill_2 FILLER_52_313 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_fill_2 FILLER_52_348 ();
 sg13g2_fill_2 FILLER_52_365 ();
 sg13g2_fill_1 FILLER_52_367 ();
 sg13g2_fill_1 FILLER_52_379 ();
 sg13g2_fill_1 FILLER_52_398 ();
 sg13g2_fill_2 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_449 ();
 sg13g2_fill_1 FILLER_52_482 ();
 sg13g2_decap_8 FILLER_52_491 ();
 sg13g2_decap_8 FILLER_52_498 ();
 sg13g2_fill_1 FILLER_52_522 ();
 sg13g2_fill_1 FILLER_52_532 ();
 sg13g2_fill_2 FILLER_52_582 ();
 sg13g2_fill_2 FILLER_52_601 ();
 sg13g2_fill_2 FILLER_52_612 ();
 sg13g2_decap_8 FILLER_52_626 ();
 sg13g2_decap_4 FILLER_52_633 ();
 sg13g2_fill_2 FILLER_52_666 ();
 sg13g2_fill_1 FILLER_52_673 ();
 sg13g2_fill_1 FILLER_52_716 ();
 sg13g2_fill_2 FILLER_52_803 ();
 sg13g2_fill_1 FILLER_52_836 ();
 sg13g2_fill_1 FILLER_52_858 ();
 sg13g2_decap_8 FILLER_52_926 ();
 sg13g2_decap_8 FILLER_52_933 ();
 sg13g2_decap_8 FILLER_52_940 ();
 sg13g2_fill_2 FILLER_52_947 ();
 sg13g2_decap_8 FILLER_52_955 ();
 sg13g2_decap_4 FILLER_52_962 ();
 sg13g2_fill_1 FILLER_52_966 ();
 sg13g2_decap_4 FILLER_52_997 ();
 sg13g2_fill_2 FILLER_52_1001 ();
 sg13g2_fill_1 FILLER_52_1076 ();
 sg13g2_fill_2 FILLER_52_1087 ();
 sg13g2_fill_1 FILLER_52_1089 ();
 sg13g2_fill_2 FILLER_52_1120 ();
 sg13g2_fill_1 FILLER_52_1208 ();
 sg13g2_fill_1 FILLER_52_1251 ();
 sg13g2_fill_2 FILLER_52_1261 ();
 sg13g2_fill_2 FILLER_52_1293 ();
 sg13g2_fill_2 FILLER_52_1299 ();
 sg13g2_fill_1 FILLER_52_1301 ();
 sg13g2_decap_4 FILLER_52_1311 ();
 sg13g2_fill_1 FILLER_52_1315 ();
 sg13g2_fill_1 FILLER_52_1321 ();
 sg13g2_fill_1 FILLER_52_1336 ();
 sg13g2_fill_1 FILLER_52_1342 ();
 sg13g2_decap_8 FILLER_52_1354 ();
 sg13g2_fill_2 FILLER_52_1361 ();
 sg13g2_fill_2 FILLER_52_1372 ();
 sg13g2_fill_2 FILLER_52_1384 ();
 sg13g2_fill_1 FILLER_52_1404 ();
 sg13g2_fill_2 FILLER_52_1410 ();
 sg13g2_fill_1 FILLER_52_1412 ();
 sg13g2_fill_2 FILLER_52_1428 ();
 sg13g2_fill_1 FILLER_52_1430 ();
 sg13g2_decap_8 FILLER_52_1466 ();
 sg13g2_decap_8 FILLER_52_1473 ();
 sg13g2_fill_1 FILLER_52_1480 ();
 sg13g2_decap_8 FILLER_52_1510 ();
 sg13g2_fill_1 FILLER_52_1554 ();
 sg13g2_fill_1 FILLER_52_1573 ();
 sg13g2_fill_1 FILLER_52_1604 ();
 sg13g2_decap_4 FILLER_52_1619 ();
 sg13g2_fill_2 FILLER_52_1644 ();
 sg13g2_fill_1 FILLER_52_1664 ();
 sg13g2_fill_1 FILLER_52_1670 ();
 sg13g2_fill_1 FILLER_52_1679 ();
 sg13g2_fill_2 FILLER_52_1694 ();
 sg13g2_fill_2 FILLER_52_1700 ();
 sg13g2_fill_1 FILLER_52_1707 ();
 sg13g2_decap_8 FILLER_52_1713 ();
 sg13g2_decap_8 FILLER_52_1720 ();
 sg13g2_decap_4 FILLER_52_1727 ();
 sg13g2_fill_2 FILLER_52_1731 ();
 sg13g2_decap_8 FILLER_52_1737 ();
 sg13g2_fill_2 FILLER_52_1744 ();
 sg13g2_decap_8 FILLER_52_1750 ();
 sg13g2_decap_8 FILLER_52_1757 ();
 sg13g2_decap_4 FILLER_52_1764 ();
 sg13g2_fill_1 FILLER_52_1768 ();
 sg13g2_fill_2 FILLER_52_1783 ();
 sg13g2_fill_1 FILLER_52_1785 ();
 sg13g2_decap_8 FILLER_52_1864 ();
 sg13g2_decap_8 FILLER_52_1892 ();
 sg13g2_fill_2 FILLER_52_1977 ();
 sg13g2_fill_2 FILLER_52_2034 ();
 sg13g2_decap_4 FILLER_52_2078 ();
 sg13g2_fill_1 FILLER_52_2086 ();
 sg13g2_fill_2 FILLER_52_2090 ();
 sg13g2_fill_1 FILLER_52_2092 ();
 sg13g2_decap_4 FILLER_52_2101 ();
 sg13g2_decap_8 FILLER_52_2115 ();
 sg13g2_fill_2 FILLER_52_2122 ();
 sg13g2_fill_1 FILLER_52_2124 ();
 sg13g2_fill_1 FILLER_52_2183 ();
 sg13g2_fill_1 FILLER_52_2233 ();
 sg13g2_fill_1 FILLER_52_2273 ();
 sg13g2_fill_2 FILLER_52_2369 ();
 sg13g2_decap_4 FILLER_52_2410 ();
 sg13g2_decap_4 FILLER_52_2424 ();
 sg13g2_decap_4 FILLER_52_2440 ();
 sg13g2_fill_2 FILLER_52_2444 ();
 sg13g2_fill_1 FILLER_52_2481 ();
 sg13g2_fill_2 FILLER_52_2488 ();
 sg13g2_fill_2 FILLER_52_2496 ();
 sg13g2_fill_2 FILLER_52_2502 ();
 sg13g2_fill_1 FILLER_52_2504 ();
 sg13g2_fill_2 FILLER_52_2537 ();
 sg13g2_fill_1 FILLER_52_2539 ();
 sg13g2_fill_2 FILLER_52_2550 ();
 sg13g2_fill_2 FILLER_52_2584 ();
 sg13g2_fill_1 FILLER_52_2586 ();
 sg13g2_decap_4 FILLER_52_2597 ();
 sg13g2_fill_1 FILLER_52_2601 ();
 sg13g2_decap_8 FILLER_52_2628 ();
 sg13g2_decap_8 FILLER_52_2635 ();
 sg13g2_decap_8 FILLER_52_2642 ();
 sg13g2_decap_8 FILLER_52_2649 ();
 sg13g2_decap_8 FILLER_52_2656 ();
 sg13g2_decap_8 FILLER_52_2663 ();
 sg13g2_fill_2 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_36 ();
 sg13g2_fill_1 FILLER_53_52 ();
 sg13g2_decap_8 FILLER_53_57 ();
 sg13g2_decap_4 FILLER_53_64 ();
 sg13g2_fill_1 FILLER_53_68 ();
 sg13g2_fill_1 FILLER_53_126 ();
 sg13g2_fill_1 FILLER_53_132 ();
 sg13g2_fill_2 FILLER_53_144 ();
 sg13g2_fill_1 FILLER_53_146 ();
 sg13g2_decap_4 FILLER_53_177 ();
 sg13g2_decap_8 FILLER_53_185 ();
 sg13g2_fill_2 FILLER_53_205 ();
 sg13g2_fill_2 FILLER_53_215 ();
 sg13g2_fill_1 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_255 ();
 sg13g2_fill_2 FILLER_53_259 ();
 sg13g2_fill_1 FILLER_53_265 ();
 sg13g2_fill_1 FILLER_53_343 ();
 sg13g2_fill_2 FILLER_53_370 ();
 sg13g2_decap_8 FILLER_53_440 ();
 sg13g2_fill_2 FILLER_53_447 ();
 sg13g2_fill_1 FILLER_53_449 ();
 sg13g2_decap_8 FILLER_53_467 ();
 sg13g2_decap_4 FILLER_53_474 ();
 sg13g2_decap_4 FILLER_53_486 ();
 sg13g2_decap_8 FILLER_53_496 ();
 sg13g2_decap_4 FILLER_53_511 ();
 sg13g2_fill_1 FILLER_53_515 ();
 sg13g2_fill_1 FILLER_53_522 ();
 sg13g2_fill_1 FILLER_53_531 ();
 sg13g2_fill_2 FILLER_53_559 ();
 sg13g2_decap_4 FILLER_53_602 ();
 sg13g2_fill_1 FILLER_53_606 ();
 sg13g2_fill_2 FILLER_53_611 ();
 sg13g2_fill_1 FILLER_53_613 ();
 sg13g2_fill_2 FILLER_53_623 ();
 sg13g2_fill_1 FILLER_53_625 ();
 sg13g2_decap_8 FILLER_53_631 ();
 sg13g2_fill_1 FILLER_53_638 ();
 sg13g2_fill_2 FILLER_53_646 ();
 sg13g2_fill_1 FILLER_53_700 ();
 sg13g2_fill_2 FILLER_53_707 ();
 sg13g2_fill_1 FILLER_53_823 ();
 sg13g2_fill_2 FILLER_53_835 ();
 sg13g2_decap_8 FILLER_53_890 ();
 sg13g2_fill_2 FILLER_53_897 ();
 sg13g2_fill_1 FILLER_53_899 ();
 sg13g2_decap_4 FILLER_53_930 ();
 sg13g2_fill_1 FILLER_53_934 ();
 sg13g2_decap_8 FILLER_53_964 ();
 sg13g2_decap_8 FILLER_53_971 ();
 sg13g2_decap_8 FILLER_53_978 ();
 sg13g2_decap_8 FILLER_53_989 ();
 sg13g2_decap_8 FILLER_53_996 ();
 sg13g2_fill_2 FILLER_53_1008 ();
 sg13g2_fill_1 FILLER_53_1010 ();
 sg13g2_fill_2 FILLER_53_1147 ();
 sg13g2_fill_2 FILLER_53_1153 ();
 sg13g2_fill_2 FILLER_53_1162 ();
 sg13g2_fill_2 FILLER_53_1185 ();
 sg13g2_fill_2 FILLER_53_1220 ();
 sg13g2_fill_1 FILLER_53_1226 ();
 sg13g2_fill_1 FILLER_53_1232 ();
 sg13g2_fill_2 FILLER_53_1243 ();
 sg13g2_fill_2 FILLER_53_1249 ();
 sg13g2_decap_8 FILLER_53_1257 ();
 sg13g2_decap_4 FILLER_53_1269 ();
 sg13g2_decap_4 FILLER_53_1322 ();
 sg13g2_fill_1 FILLER_53_1345 ();
 sg13g2_decap_4 FILLER_53_1357 ();
 sg13g2_fill_1 FILLER_53_1361 ();
 sg13g2_decap_8 FILLER_53_1366 ();
 sg13g2_decap_4 FILLER_53_1373 ();
 sg13g2_fill_2 FILLER_53_1382 ();
 sg13g2_decap_4 FILLER_53_1388 ();
 sg13g2_fill_2 FILLER_53_1392 ();
 sg13g2_decap_8 FILLER_53_1400 ();
 sg13g2_fill_2 FILLER_53_1413 ();
 sg13g2_fill_2 FILLER_53_1420 ();
 sg13g2_fill_2 FILLER_53_1426 ();
 sg13g2_fill_1 FILLER_53_1428 ();
 sg13g2_decap_8 FILLER_53_1458 ();
 sg13g2_decap_8 FILLER_53_1465 ();
 sg13g2_decap_4 FILLER_53_1472 ();
 sg13g2_fill_2 FILLER_53_1502 ();
 sg13g2_fill_1 FILLER_53_1504 ();
 sg13g2_decap_4 FILLER_53_1526 ();
 sg13g2_fill_1 FILLER_53_1530 ();
 sg13g2_fill_2 FILLER_53_1549 ();
 sg13g2_fill_2 FILLER_53_1556 ();
 sg13g2_fill_1 FILLER_53_1567 ();
 sg13g2_fill_1 FILLER_53_1590 ();
 sg13g2_fill_1 FILLER_53_1604 ();
 sg13g2_fill_1 FILLER_53_1613 ();
 sg13g2_fill_2 FILLER_53_1641 ();
 sg13g2_decap_8 FILLER_53_1651 ();
 sg13g2_fill_1 FILLER_53_1665 ();
 sg13g2_fill_2 FILLER_53_1676 ();
 sg13g2_fill_1 FILLER_53_1678 ();
 sg13g2_fill_1 FILLER_53_1684 ();
 sg13g2_fill_1 FILLER_53_1697 ();
 sg13g2_fill_1 FILLER_53_1705 ();
 sg13g2_decap_4 FILLER_53_1711 ();
 sg13g2_decap_8 FILLER_53_1719 ();
 sg13g2_fill_2 FILLER_53_1726 ();
 sg13g2_fill_1 FILLER_53_1728 ();
 sg13g2_fill_1 FILLER_53_1734 ();
 sg13g2_fill_2 FILLER_53_1774 ();
 sg13g2_fill_2 FILLER_53_1802 ();
 sg13g2_fill_1 FILLER_53_1830 ();
 sg13g2_fill_2 FILLER_53_1844 ();
 sg13g2_fill_1 FILLER_53_1854 ();
 sg13g2_fill_1 FILLER_53_1869 ();
 sg13g2_fill_1 FILLER_53_1874 ();
 sg13g2_decap_4 FILLER_53_1885 ();
 sg13g2_fill_1 FILLER_53_1889 ();
 sg13g2_decap_8 FILLER_53_1900 ();
 sg13g2_decap_4 FILLER_53_1907 ();
 sg13g2_fill_2 FILLER_53_1911 ();
 sg13g2_fill_1 FILLER_53_1917 ();
 sg13g2_fill_2 FILLER_53_1987 ();
 sg13g2_fill_1 FILLER_53_1994 ();
 sg13g2_fill_1 FILLER_53_2004 ();
 sg13g2_fill_1 FILLER_53_2010 ();
 sg13g2_fill_1 FILLER_53_2015 ();
 sg13g2_fill_2 FILLER_53_2076 ();
 sg13g2_fill_1 FILLER_53_2078 ();
 sg13g2_decap_8 FILLER_53_2144 ();
 sg13g2_decap_8 FILLER_53_2151 ();
 sg13g2_fill_2 FILLER_53_2162 ();
 sg13g2_fill_1 FILLER_53_2164 ();
 sg13g2_fill_1 FILLER_53_2207 ();
 sg13g2_fill_2 FILLER_53_2372 ();
 sg13g2_fill_2 FILLER_53_2410 ();
 sg13g2_fill_1 FILLER_53_2412 ();
 sg13g2_fill_1 FILLER_53_2439 ();
 sg13g2_fill_2 FILLER_53_2447 ();
 sg13g2_decap_8 FILLER_53_2469 ();
 sg13g2_fill_2 FILLER_53_2476 ();
 sg13g2_decap_8 FILLER_53_2481 ();
 sg13g2_decap_8 FILLER_53_2488 ();
 sg13g2_decap_4 FILLER_53_2495 ();
 sg13g2_fill_2 FILLER_53_2499 ();
 sg13g2_fill_2 FILLER_53_2505 ();
 sg13g2_fill_1 FILLER_53_2517 ();
 sg13g2_decap_8 FILLER_53_2616 ();
 sg13g2_decap_8 FILLER_53_2623 ();
 sg13g2_decap_8 FILLER_53_2630 ();
 sg13g2_decap_8 FILLER_53_2637 ();
 sg13g2_decap_8 FILLER_53_2644 ();
 sg13g2_decap_8 FILLER_53_2651 ();
 sg13g2_decap_8 FILLER_53_2658 ();
 sg13g2_decap_4 FILLER_53_2665 ();
 sg13g2_fill_1 FILLER_53_2669 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_fill_2 FILLER_54_25 ();
 sg13g2_fill_1 FILLER_54_27 ();
 sg13g2_fill_1 FILLER_54_33 ();
 sg13g2_decap_8 FILLER_54_62 ();
 sg13g2_fill_1 FILLER_54_69 ();
 sg13g2_fill_2 FILLER_54_78 ();
 sg13g2_fill_1 FILLER_54_111 ();
 sg13g2_decap_4 FILLER_54_174 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_1 FILLER_54_185 ();
 sg13g2_decap_4 FILLER_54_191 ();
 sg13g2_fill_2 FILLER_54_195 ();
 sg13g2_fill_2 FILLER_54_209 ();
 sg13g2_fill_1 FILLER_54_272 ();
 sg13g2_fill_1 FILLER_54_278 ();
 sg13g2_fill_2 FILLER_54_283 ();
 sg13g2_fill_1 FILLER_54_313 ();
 sg13g2_fill_2 FILLER_54_325 ();
 sg13g2_fill_1 FILLER_54_348 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_fill_2 FILLER_54_399 ();
 sg13g2_fill_1 FILLER_54_401 ();
 sg13g2_decap_4 FILLER_54_431 ();
 sg13g2_fill_2 FILLER_54_465 ();
 sg13g2_fill_1 FILLER_54_467 ();
 sg13g2_decap_4 FILLER_54_477 ();
 sg13g2_fill_1 FILLER_54_481 ();
 sg13g2_decap_4 FILLER_54_518 ();
 sg13g2_fill_1 FILLER_54_522 ();
 sg13g2_fill_2 FILLER_54_531 ();
 sg13g2_fill_2 FILLER_54_547 ();
 sg13g2_decap_8 FILLER_54_592 ();
 sg13g2_fill_1 FILLER_54_599 ();
 sg13g2_decap_4 FILLER_54_604 ();
 sg13g2_decap_4 FILLER_54_634 ();
 sg13g2_fill_2 FILLER_54_638 ();
 sg13g2_fill_1 FILLER_54_666 ();
 sg13g2_fill_1 FILLER_54_708 ();
 sg13g2_fill_1 FILLER_54_745 ();
 sg13g2_fill_2 FILLER_54_758 ();
 sg13g2_fill_2 FILLER_54_775 ();
 sg13g2_fill_2 FILLER_54_793 ();
 sg13g2_fill_1 FILLER_54_809 ();
 sg13g2_fill_1 FILLER_54_839 ();
 sg13g2_fill_2 FILLER_54_886 ();
 sg13g2_fill_1 FILLER_54_888 ();
 sg13g2_fill_2 FILLER_54_899 ();
 sg13g2_fill_2 FILLER_54_905 ();
 sg13g2_fill_1 FILLER_54_907 ();
 sg13g2_fill_2 FILLER_54_918 ();
 sg13g2_fill_2 FILLER_54_926 ();
 sg13g2_fill_1 FILLER_54_942 ();
 sg13g2_decap_8 FILLER_54_969 ();
 sg13g2_decap_8 FILLER_54_976 ();
 sg13g2_decap_8 FILLER_54_983 ();
 sg13g2_decap_4 FILLER_54_990 ();
 sg13g2_fill_1 FILLER_54_994 ();
 sg13g2_decap_8 FILLER_54_999 ();
 sg13g2_decap_4 FILLER_54_1006 ();
 sg13g2_fill_1 FILLER_54_1010 ();
 sg13g2_decap_8 FILLER_54_1064 ();
 sg13g2_decap_8 FILLER_54_1086 ();
 sg13g2_fill_1 FILLER_54_1093 ();
 sg13g2_decap_4 FILLER_54_1102 ();
 sg13g2_fill_1 FILLER_54_1106 ();
 sg13g2_fill_2 FILLER_54_1117 ();
 sg13g2_fill_1 FILLER_54_1123 ();
 sg13g2_fill_2 FILLER_54_1153 ();
 sg13g2_fill_2 FILLER_54_1160 ();
 sg13g2_fill_1 FILLER_54_1232 ();
 sg13g2_decap_8 FILLER_54_1248 ();
 sg13g2_decap_8 FILLER_54_1255 ();
 sg13g2_decap_8 FILLER_54_1262 ();
 sg13g2_fill_2 FILLER_54_1269 ();
 sg13g2_fill_2 FILLER_54_1281 ();
 sg13g2_fill_1 FILLER_54_1283 ();
 sg13g2_fill_1 FILLER_54_1300 ();
 sg13g2_decap_8 FILLER_54_1314 ();
 sg13g2_fill_2 FILLER_54_1336 ();
 sg13g2_fill_1 FILLER_54_1338 ();
 sg13g2_decap_8 FILLER_54_1355 ();
 sg13g2_fill_1 FILLER_54_1362 ();
 sg13g2_fill_2 FILLER_54_1373 ();
 sg13g2_fill_1 FILLER_54_1383 ();
 sg13g2_fill_2 FILLER_54_1405 ();
 sg13g2_decap_4 FILLER_54_1421 ();
 sg13g2_fill_1 FILLER_54_1425 ();
 sg13g2_decap_8 FILLER_54_1459 ();
 sg13g2_decap_8 FILLER_54_1466 ();
 sg13g2_decap_8 FILLER_54_1473 ();
 sg13g2_fill_1 FILLER_54_1480 ();
 sg13g2_fill_1 FILLER_54_1504 ();
 sg13g2_decap_4 FILLER_54_1509 ();
 sg13g2_fill_2 FILLER_54_1513 ();
 sg13g2_fill_1 FILLER_54_1533 ();
 sg13g2_decap_8 FILLER_54_1553 ();
 sg13g2_fill_2 FILLER_54_1560 ();
 sg13g2_decap_8 FILLER_54_1571 ();
 sg13g2_decap_4 FILLER_54_1578 ();
 sg13g2_fill_1 FILLER_54_1582 ();
 sg13g2_fill_1 FILLER_54_1600 ();
 sg13g2_decap_8 FILLER_54_1606 ();
 sg13g2_fill_1 FILLER_54_1613 ();
 sg13g2_decap_4 FILLER_54_1618 ();
 sg13g2_fill_1 FILLER_54_1622 ();
 sg13g2_fill_2 FILLER_54_1627 ();
 sg13g2_fill_1 FILLER_54_1629 ();
 sg13g2_fill_2 FILLER_54_1657 ();
 sg13g2_fill_2 FILLER_54_1664 ();
 sg13g2_fill_1 FILLER_54_1666 ();
 sg13g2_fill_1 FILLER_54_1680 ();
 sg13g2_fill_1 FILLER_54_1692 ();
 sg13g2_fill_1 FILLER_54_1698 ();
 sg13g2_fill_1 FILLER_54_1712 ();
 sg13g2_decap_8 FILLER_54_1730 ();
 sg13g2_fill_2 FILLER_54_1737 ();
 sg13g2_fill_1 FILLER_54_1739 ();
 sg13g2_decap_8 FILLER_54_1744 ();
 sg13g2_decap_4 FILLER_54_1751 ();
 sg13g2_fill_2 FILLER_54_1755 ();
 sg13g2_fill_1 FILLER_54_1761 ();
 sg13g2_fill_1 FILLER_54_1778 ();
 sg13g2_fill_2 FILLER_54_1789 ();
 sg13g2_fill_1 FILLER_54_1791 ();
 sg13g2_decap_8 FILLER_54_1826 ();
 sg13g2_decap_8 FILLER_54_1833 ();
 sg13g2_decap_4 FILLER_54_1840 ();
 sg13g2_fill_1 FILLER_54_1844 ();
 sg13g2_decap_4 FILLER_54_1848 ();
 sg13g2_fill_1 FILLER_54_1852 ();
 sg13g2_fill_1 FILLER_54_1858 ();
 sg13g2_fill_1 FILLER_54_1892 ();
 sg13g2_decap_4 FILLER_54_1897 ();
 sg13g2_fill_2 FILLER_54_1901 ();
 sg13g2_fill_2 FILLER_54_1916 ();
 sg13g2_fill_1 FILLER_54_1931 ();
 sg13g2_fill_1 FILLER_54_1948 ();
 sg13g2_fill_1 FILLER_54_1968 ();
 sg13g2_fill_1 FILLER_54_1979 ();
 sg13g2_fill_1 FILLER_54_2001 ();
 sg13g2_fill_1 FILLER_54_2016 ();
 sg13g2_fill_1 FILLER_54_2034 ();
 sg13g2_fill_2 FILLER_54_2066 ();
 sg13g2_fill_1 FILLER_54_2068 ();
 sg13g2_decap_4 FILLER_54_2095 ();
 sg13g2_fill_1 FILLER_54_2099 ();
 sg13g2_fill_2 FILLER_54_2105 ();
 sg13g2_fill_1 FILLER_54_2112 ();
 sg13g2_decap_8 FILLER_54_2154 ();
 sg13g2_decap_4 FILLER_54_2161 ();
 sg13g2_fill_2 FILLER_54_2165 ();
 sg13g2_fill_2 FILLER_54_2170 ();
 sg13g2_fill_2 FILLER_54_2185 ();
 sg13g2_fill_1 FILLER_54_2191 ();
 sg13g2_fill_1 FILLER_54_2223 ();
 sg13g2_fill_1 FILLER_54_2247 ();
 sg13g2_fill_2 FILLER_54_2258 ();
 sg13g2_fill_2 FILLER_54_2264 ();
 sg13g2_fill_1 FILLER_54_2281 ();
 sg13g2_fill_1 FILLER_54_2296 ();
 sg13g2_fill_2 FILLER_54_2353 ();
 sg13g2_fill_1 FILLER_54_2365 ();
 sg13g2_fill_1 FILLER_54_2372 ();
 sg13g2_fill_1 FILLER_54_2383 ();
 sg13g2_fill_1 FILLER_54_2390 ();
 sg13g2_fill_2 FILLER_54_2397 ();
 sg13g2_fill_1 FILLER_54_2440 ();
 sg13g2_decap_8 FILLER_54_2467 ();
 sg13g2_decap_8 FILLER_54_2474 ();
 sg13g2_fill_2 FILLER_54_2481 ();
 sg13g2_fill_1 FILLER_54_2497 ();
 sg13g2_fill_2 FILLER_54_2509 ();
 sg13g2_fill_1 FILLER_54_2535 ();
 sg13g2_fill_1 FILLER_54_2550 ();
 sg13g2_fill_1 FILLER_54_2555 ();
 sg13g2_fill_2 FILLER_54_2595 ();
 sg13g2_fill_1 FILLER_54_2597 ();
 sg13g2_fill_1 FILLER_54_2624 ();
 sg13g2_decap_8 FILLER_54_2629 ();
 sg13g2_decap_8 FILLER_54_2636 ();
 sg13g2_decap_8 FILLER_54_2643 ();
 sg13g2_decap_8 FILLER_54_2650 ();
 sg13g2_decap_8 FILLER_54_2657 ();
 sg13g2_decap_4 FILLER_54_2664 ();
 sg13g2_fill_2 FILLER_54_2668 ();
 sg13g2_fill_2 FILLER_55_3 ();
 sg13g2_fill_1 FILLER_55_13 ();
 sg13g2_decap_4 FILLER_55_18 ();
 sg13g2_fill_2 FILLER_55_30 ();
 sg13g2_fill_1 FILLER_55_56 ();
 sg13g2_fill_2 FILLER_55_67 ();
 sg13g2_fill_2 FILLER_55_87 ();
 sg13g2_decap_8 FILLER_55_97 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_decap_8 FILLER_55_111 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_decap_4 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_162 ();
 sg13g2_fill_2 FILLER_55_203 ();
 sg13g2_fill_1 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_211 ();
 sg13g2_fill_1 FILLER_55_213 ();
 sg13g2_fill_1 FILLER_55_218 ();
 sg13g2_fill_2 FILLER_55_250 ();
 sg13g2_fill_1 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_312 ();
 sg13g2_fill_1 FILLER_55_349 ();
 sg13g2_fill_2 FILLER_55_355 ();
 sg13g2_fill_2 FILLER_55_384 ();
 sg13g2_decap_4 FILLER_55_395 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_decap_4 FILLER_55_409 ();
 sg13g2_fill_2 FILLER_55_413 ();
 sg13g2_decap_4 FILLER_55_421 ();
 sg13g2_fill_1 FILLER_55_425 ();
 sg13g2_fill_1 FILLER_55_432 ();
 sg13g2_fill_1 FILLER_55_463 ();
 sg13g2_fill_1 FILLER_55_470 ();
 sg13g2_fill_2 FILLER_55_479 ();
 sg13g2_fill_1 FILLER_55_481 ();
 sg13g2_fill_2 FILLER_55_488 ();
 sg13g2_fill_2 FILLER_55_498 ();
 sg13g2_fill_2 FILLER_55_504 ();
 sg13g2_fill_2 FILLER_55_512 ();
 sg13g2_decap_4 FILLER_55_522 ();
 sg13g2_fill_2 FILLER_55_561 ();
 sg13g2_fill_1 FILLER_55_563 ();
 sg13g2_fill_2 FILLER_55_577 ();
 sg13g2_fill_1 FILLER_55_579 ();
 sg13g2_fill_1 FILLER_55_590 ();
 sg13g2_fill_2 FILLER_55_621 ();
 sg13g2_decap_8 FILLER_55_627 ();
 sg13g2_decap_8 FILLER_55_634 ();
 sg13g2_decap_4 FILLER_55_641 ();
 sg13g2_fill_1 FILLER_55_645 ();
 sg13g2_decap_4 FILLER_55_655 ();
 sg13g2_fill_1 FILLER_55_659 ();
 sg13g2_fill_1 FILLER_55_665 ();
 sg13g2_decap_4 FILLER_55_670 ();
 sg13g2_fill_2 FILLER_55_674 ();
 sg13g2_fill_2 FILLER_55_701 ();
 sg13g2_fill_2 FILLER_55_709 ();
 sg13g2_fill_2 FILLER_55_753 ();
 sg13g2_fill_1 FILLER_55_829 ();
 sg13g2_fill_1 FILLER_55_842 ();
 sg13g2_fill_1 FILLER_55_853 ();
 sg13g2_fill_2 FILLER_55_933 ();
 sg13g2_fill_1 FILLER_55_952 ();
 sg13g2_decap_8 FILLER_55_1011 ();
 sg13g2_decap_8 FILLER_55_1018 ();
 sg13g2_decap_8 FILLER_55_1025 ();
 sg13g2_decap_8 FILLER_55_1032 ();
 sg13g2_decap_8 FILLER_55_1039 ();
 sg13g2_decap_8 FILLER_55_1046 ();
 sg13g2_fill_2 FILLER_55_1053 ();
 sg13g2_decap_8 FILLER_55_1077 ();
 sg13g2_fill_2 FILLER_55_1084 ();
 sg13g2_decap_8 FILLER_55_1096 ();
 sg13g2_fill_2 FILLER_55_1103 ();
 sg13g2_fill_1 FILLER_55_1126 ();
 sg13g2_fill_1 FILLER_55_1132 ();
 sg13g2_fill_1 FILLER_55_1159 ();
 sg13g2_fill_1 FILLER_55_1169 ();
 sg13g2_fill_2 FILLER_55_1178 ();
 sg13g2_fill_2 FILLER_55_1198 ();
 sg13g2_fill_1 FILLER_55_1242 ();
 sg13g2_decap_4 FILLER_55_1247 ();
 sg13g2_fill_2 FILLER_55_1255 ();
 sg13g2_fill_2 FILLER_55_1287 ();
 sg13g2_fill_1 FILLER_55_1289 ();
 sg13g2_fill_1 FILLER_55_1316 ();
 sg13g2_decap_8 FILLER_55_1325 ();
 sg13g2_fill_2 FILLER_55_1344 ();
 sg13g2_fill_1 FILLER_55_1346 ();
 sg13g2_fill_1 FILLER_55_1364 ();
 sg13g2_fill_2 FILLER_55_1375 ();
 sg13g2_fill_1 FILLER_55_1377 ();
 sg13g2_decap_4 FILLER_55_1413 ();
 sg13g2_decap_8 FILLER_55_1427 ();
 sg13g2_fill_2 FILLER_55_1434 ();
 sg13g2_decap_4 FILLER_55_1446 ();
 sg13g2_fill_1 FILLER_55_1455 ();
 sg13g2_fill_1 FILLER_55_1461 ();
 sg13g2_fill_2 FILLER_55_1467 ();
 sg13g2_fill_2 FILLER_55_1473 ();
 sg13g2_fill_1 FILLER_55_1478 ();
 sg13g2_fill_1 FILLER_55_1492 ();
 sg13g2_fill_1 FILLER_55_1498 ();
 sg13g2_decap_4 FILLER_55_1567 ();
 sg13g2_fill_1 FILLER_55_1571 ();
 sg13g2_decap_4 FILLER_55_1584 ();
 sg13g2_fill_2 FILLER_55_1588 ();
 sg13g2_decap_8 FILLER_55_1614 ();
 sg13g2_decap_4 FILLER_55_1621 ();
 sg13g2_fill_2 FILLER_55_1625 ();
 sg13g2_decap_8 FILLER_55_1655 ();
 sg13g2_decap_8 FILLER_55_1662 ();
 sg13g2_decap_8 FILLER_55_1669 ();
 sg13g2_fill_2 FILLER_55_1676 ();
 sg13g2_decap_8 FILLER_55_1698 ();
 sg13g2_fill_2 FILLER_55_1705 ();
 sg13g2_decap_8 FILLER_55_1711 ();
 sg13g2_decap_4 FILLER_55_1718 ();
 sg13g2_fill_2 FILLER_55_1722 ();
 sg13g2_decap_4 FILLER_55_1728 ();
 sg13g2_fill_1 FILLER_55_1732 ();
 sg13g2_fill_2 FILLER_55_1763 ();
 sg13g2_fill_1 FILLER_55_1765 ();
 sg13g2_fill_2 FILLER_55_1774 ();
 sg13g2_fill_1 FILLER_55_1776 ();
 sg13g2_decap_8 FILLER_55_1821 ();
 sg13g2_decap_4 FILLER_55_1828 ();
 sg13g2_fill_1 FILLER_55_1832 ();
 sg13g2_decap_4 FILLER_55_1837 ();
 sg13g2_fill_1 FILLER_55_1841 ();
 sg13g2_fill_1 FILLER_55_1852 ();
 sg13g2_decap_4 FILLER_55_1861 ();
 sg13g2_fill_1 FILLER_55_1880 ();
 sg13g2_fill_1 FILLER_55_1899 ();
 sg13g2_fill_2 FILLER_55_1913 ();
 sg13g2_fill_1 FILLER_55_1915 ();
 sg13g2_decap_4 FILLER_55_1930 ();
 sg13g2_fill_1 FILLER_55_1948 ();
 sg13g2_fill_1 FILLER_55_1952 ();
 sg13g2_fill_2 FILLER_55_1957 ();
 sg13g2_fill_1 FILLER_55_2006 ();
 sg13g2_fill_2 FILLER_55_2021 ();
 sg13g2_fill_1 FILLER_55_2035 ();
 sg13g2_fill_1 FILLER_55_2045 ();
 sg13g2_fill_1 FILLER_55_2101 ();
 sg13g2_fill_2 FILLER_55_2128 ();
 sg13g2_fill_2 FILLER_55_2135 ();
 sg13g2_fill_1 FILLER_55_2137 ();
 sg13g2_fill_1 FILLER_55_2232 ();
 sg13g2_fill_1 FILLER_55_2240 ();
 sg13g2_fill_2 FILLER_55_2323 ();
 sg13g2_fill_1 FILLER_55_2345 ();
 sg13g2_fill_1 FILLER_55_2352 ();
 sg13g2_fill_1 FILLER_55_2379 ();
 sg13g2_fill_1 FILLER_55_2406 ();
 sg13g2_fill_2 FILLER_55_2413 ();
 sg13g2_fill_1 FILLER_55_2415 ();
 sg13g2_fill_2 FILLER_55_2420 ();
 sg13g2_fill_1 FILLER_55_2422 ();
 sg13g2_decap_8 FILLER_55_2427 ();
 sg13g2_decap_8 FILLER_55_2434 ();
 sg13g2_fill_2 FILLER_55_2441 ();
 sg13g2_fill_2 FILLER_55_2448 ();
 sg13g2_fill_1 FILLER_55_2450 ();
 sg13g2_decap_8 FILLER_55_2461 ();
 sg13g2_fill_2 FILLER_55_2468 ();
 sg13g2_decap_4 FILLER_55_2522 ();
 sg13g2_fill_2 FILLER_55_2552 ();
 sg13g2_fill_1 FILLER_55_2569 ();
 sg13g2_fill_1 FILLER_55_2576 ();
 sg13g2_fill_1 FILLER_55_2593 ();
 sg13g2_fill_1 FILLER_55_2598 ();
 sg13g2_decap_8 FILLER_55_2625 ();
 sg13g2_decap_8 FILLER_55_2632 ();
 sg13g2_decap_8 FILLER_55_2639 ();
 sg13g2_decap_8 FILLER_55_2646 ();
 sg13g2_decap_8 FILLER_55_2653 ();
 sg13g2_decap_8 FILLER_55_2660 ();
 sg13g2_fill_2 FILLER_55_2667 ();
 sg13g2_fill_1 FILLER_55_2669 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_64 ();
 sg13g2_fill_2 FILLER_56_73 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_fill_1 FILLER_56_89 ();
 sg13g2_fill_1 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_112 ();
 sg13g2_decap_8 FILLER_56_119 ();
 sg13g2_decap_4 FILLER_56_126 ();
 sg13g2_fill_2 FILLER_56_135 ();
 sg13g2_decap_4 FILLER_56_145 ();
 sg13g2_fill_2 FILLER_56_179 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_decap_4 FILLER_56_192 ();
 sg13g2_fill_2 FILLER_56_215 ();
 sg13g2_fill_2 FILLER_56_239 ();
 sg13g2_fill_1 FILLER_56_241 ();
 sg13g2_fill_2 FILLER_56_246 ();
 sg13g2_fill_1 FILLER_56_252 ();
 sg13g2_fill_2 FILLER_56_257 ();
 sg13g2_fill_1 FILLER_56_310 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_decap_8 FILLER_56_374 ();
 sg13g2_fill_1 FILLER_56_381 ();
 sg13g2_decap_8 FILLER_56_412 ();
 sg13g2_decap_8 FILLER_56_419 ();
 sg13g2_fill_2 FILLER_56_426 ();
 sg13g2_fill_1 FILLER_56_518 ();
 sg13g2_fill_1 FILLER_56_527 ();
 sg13g2_fill_1 FILLER_56_536 ();
 sg13g2_decap_8 FILLER_56_543 ();
 sg13g2_decap_4 FILLER_56_550 ();
 sg13g2_fill_2 FILLER_56_567 ();
 sg13g2_fill_1 FILLER_56_569 ();
 sg13g2_fill_2 FILLER_56_578 ();
 sg13g2_fill_1 FILLER_56_580 ();
 sg13g2_fill_2 FILLER_56_591 ();
 sg13g2_decap_4 FILLER_56_619 ();
 sg13g2_decap_8 FILLER_56_633 ();
 sg13g2_decap_4 FILLER_56_640 ();
 sg13g2_fill_1 FILLER_56_644 ();
 sg13g2_fill_2 FILLER_56_668 ();
 sg13g2_fill_1 FILLER_56_670 ();
 sg13g2_fill_2 FILLER_56_703 ();
 sg13g2_fill_1 FILLER_56_788 ();
 sg13g2_fill_1 FILLER_56_825 ();
 sg13g2_fill_2 FILLER_56_831 ();
 sg13g2_fill_2 FILLER_56_842 ();
 sg13g2_fill_1 FILLER_56_848 ();
 sg13g2_fill_2 FILLER_56_904 ();
 sg13g2_fill_1 FILLER_56_906 ();
 sg13g2_decap_8 FILLER_56_912 ();
 sg13g2_fill_2 FILLER_56_947 ();
 sg13g2_fill_2 FILLER_56_957 ();
 sg13g2_fill_2 FILLER_56_1012 ();
 sg13g2_fill_1 FILLER_56_1054 ();
 sg13g2_fill_2 FILLER_56_1199 ();
 sg13g2_fill_2 FILLER_56_1258 ();
 sg13g2_fill_1 FILLER_56_1260 ();
 sg13g2_fill_2 FILLER_56_1287 ();
 sg13g2_fill_1 FILLER_56_1293 ();
 sg13g2_fill_2 FILLER_56_1298 ();
 sg13g2_fill_2 FILLER_56_1304 ();
 sg13g2_fill_1 FILLER_56_1317 ();
 sg13g2_fill_1 FILLER_56_1353 ();
 sg13g2_fill_2 FILLER_56_1377 ();
 sg13g2_fill_1 FILLER_56_1379 ();
 sg13g2_decap_4 FILLER_56_1412 ();
 sg13g2_decap_8 FILLER_56_1426 ();
 sg13g2_decap_8 FILLER_56_1433 ();
 sg13g2_fill_2 FILLER_56_1440 ();
 sg13g2_fill_1 FILLER_56_1528 ();
 sg13g2_fill_1 FILLER_56_1534 ();
 sg13g2_decap_8 FILLER_56_1547 ();
 sg13g2_decap_8 FILLER_56_1554 ();
 sg13g2_fill_2 FILLER_56_1561 ();
 sg13g2_decap_4 FILLER_56_1567 ();
 sg13g2_decap_4 FILLER_56_1581 ();
 sg13g2_fill_1 FILLER_56_1590 ();
 sg13g2_fill_1 FILLER_56_1609 ();
 sg13g2_fill_2 FILLER_56_1624 ();
 sg13g2_decap_4 FILLER_56_1631 ();
 sg13g2_decap_8 FILLER_56_1644 ();
 sg13g2_fill_2 FILLER_56_1651 ();
 sg13g2_fill_1 FILLER_56_1653 ();
 sg13g2_decap_4 FILLER_56_1667 ();
 sg13g2_fill_1 FILLER_56_1671 ();
 sg13g2_fill_2 FILLER_56_1682 ();
 sg13g2_fill_1 FILLER_56_1684 ();
 sg13g2_fill_2 FILLER_56_1711 ();
 sg13g2_fill_1 FILLER_56_1713 ();
 sg13g2_decap_8 FILLER_56_1723 ();
 sg13g2_fill_2 FILLER_56_1730 ();
 sg13g2_fill_1 FILLER_56_1732 ();
 sg13g2_decap_4 FILLER_56_1738 ();
 sg13g2_decap_8 FILLER_56_1756 ();
 sg13g2_decap_8 FILLER_56_1763 ();
 sg13g2_decap_8 FILLER_56_1770 ();
 sg13g2_fill_1 FILLER_56_1789 ();
 sg13g2_fill_1 FILLER_56_1799 ();
 sg13g2_decap_8 FILLER_56_1809 ();
 sg13g2_fill_1 FILLER_56_1816 ();
 sg13g2_fill_2 FILLER_56_1821 ();
 sg13g2_fill_1 FILLER_56_1853 ();
 sg13g2_fill_2 FILLER_56_1887 ();
 sg13g2_fill_2 FILLER_56_1902 ();
 sg13g2_fill_1 FILLER_56_1909 ();
 sg13g2_fill_1 FILLER_56_1918 ();
 sg13g2_fill_2 FILLER_56_1928 ();
 sg13g2_fill_2 FILLER_56_1935 ();
 sg13g2_fill_2 FILLER_56_1944 ();
 sg13g2_fill_1 FILLER_56_1959 ();
 sg13g2_fill_1 FILLER_56_1990 ();
 sg13g2_fill_1 FILLER_56_1999 ();
 sg13g2_fill_1 FILLER_56_2018 ();
 sg13g2_fill_2 FILLER_56_2052 ();
 sg13g2_fill_1 FILLER_56_2054 ();
 sg13g2_decap_4 FILLER_56_2098 ();
 sg13g2_fill_2 FILLER_56_2102 ();
 sg13g2_decap_4 FILLER_56_2112 ();
 sg13g2_fill_1 FILLER_56_2116 ();
 sg13g2_decap_4 FILLER_56_2121 ();
 sg13g2_fill_1 FILLER_56_2125 ();
 sg13g2_fill_2 FILLER_56_2152 ();
 sg13g2_fill_1 FILLER_56_2154 ();
 sg13g2_decap_4 FILLER_56_2162 ();
 sg13g2_fill_1 FILLER_56_2166 ();
 sg13g2_fill_2 FILLER_56_2179 ();
 sg13g2_fill_1 FILLER_56_2200 ();
 sg13g2_fill_1 FILLER_56_2206 ();
 sg13g2_fill_1 FILLER_56_2223 ();
 sg13g2_fill_1 FILLER_56_2230 ();
 sg13g2_fill_1 FILLER_56_2242 ();
 sg13g2_fill_2 FILLER_56_2295 ();
 sg13g2_fill_2 FILLER_56_2355 ();
 sg13g2_fill_1 FILLER_56_2357 ();
 sg13g2_fill_2 FILLER_56_2378 ();
 sg13g2_fill_1 FILLER_56_2380 ();
 sg13g2_decap_8 FILLER_56_2411 ();
 sg13g2_decap_8 FILLER_56_2418 ();
 sg13g2_fill_2 FILLER_56_2425 ();
 sg13g2_fill_2 FILLER_56_2443 ();
 sg13g2_fill_1 FILLER_56_2445 ();
 sg13g2_decap_4 FILLER_56_2456 ();
 sg13g2_fill_1 FILLER_56_2460 ();
 sg13g2_decap_4 FILLER_56_2471 ();
 sg13g2_fill_1 FILLER_56_2475 ();
 sg13g2_decap_4 FILLER_56_2480 ();
 sg13g2_decap_4 FILLER_56_2501 ();
 sg13g2_fill_2 FILLER_56_2509 ();
 sg13g2_decap_8 FILLER_56_2517 ();
 sg13g2_decap_8 FILLER_56_2524 ();
 sg13g2_decap_8 FILLER_56_2531 ();
 sg13g2_decap_8 FILLER_56_2538 ();
 sg13g2_decap_8 FILLER_56_2545 ();
 sg13g2_decap_8 FILLER_56_2575 ();
 sg13g2_decap_4 FILLER_56_2582 ();
 sg13g2_fill_2 FILLER_56_2596 ();
 sg13g2_fill_1 FILLER_56_2598 ();
 sg13g2_decap_8 FILLER_56_2629 ();
 sg13g2_decap_8 FILLER_56_2636 ();
 sg13g2_decap_8 FILLER_56_2643 ();
 sg13g2_decap_8 FILLER_56_2650 ();
 sg13g2_decap_8 FILLER_56_2657 ();
 sg13g2_decap_4 FILLER_56_2664 ();
 sg13g2_fill_2 FILLER_56_2668 ();
 sg13g2_fill_1 FILLER_57_0 ();
 sg13g2_fill_1 FILLER_57_90 ();
 sg13g2_fill_1 FILLER_57_122 ();
 sg13g2_decap_8 FILLER_57_128 ();
 sg13g2_decap_8 FILLER_57_135 ();
 sg13g2_decap_8 FILLER_57_142 ();
 sg13g2_decap_8 FILLER_57_149 ();
 sg13g2_decap_4 FILLER_57_156 ();
 sg13g2_decap_8 FILLER_57_164 ();
 sg13g2_decap_8 FILLER_57_171 ();
 sg13g2_fill_2 FILLER_57_178 ();
 sg13g2_fill_1 FILLER_57_180 ();
 sg13g2_decap_4 FILLER_57_207 ();
 sg13g2_decap_4 FILLER_57_219 ();
 sg13g2_fill_2 FILLER_57_223 ();
 sg13g2_decap_8 FILLER_57_234 ();
 sg13g2_fill_2 FILLER_57_241 ();
 sg13g2_decap_4 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_262 ();
 sg13g2_fill_1 FILLER_57_267 ();
 sg13g2_fill_1 FILLER_57_272 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_fill_1 FILLER_57_309 ();
 sg13g2_fill_1 FILLER_57_327 ();
 sg13g2_decap_4 FILLER_57_398 ();
 sg13g2_fill_1 FILLER_57_402 ();
 sg13g2_decap_4 FILLER_57_447 ();
 sg13g2_fill_2 FILLER_57_457 ();
 sg13g2_decap_4 FILLER_57_467 ();
 sg13g2_fill_1 FILLER_57_471 ();
 sg13g2_decap_4 FILLER_57_476 ();
 sg13g2_fill_2 FILLER_57_480 ();
 sg13g2_decap_8 FILLER_57_487 ();
 sg13g2_decap_4 FILLER_57_494 ();
 sg13g2_fill_1 FILLER_57_498 ();
 sg13g2_fill_2 FILLER_57_503 ();
 sg13g2_fill_2 FILLER_57_513 ();
 sg13g2_decap_8 FILLER_57_521 ();
 sg13g2_decap_8 FILLER_57_528 ();
 sg13g2_fill_2 FILLER_57_535 ();
 sg13g2_fill_1 FILLER_57_537 ();
 sg13g2_decap_4 FILLER_57_551 ();
 sg13g2_fill_1 FILLER_57_555 ();
 sg13g2_fill_2 FILLER_57_566 ();
 sg13g2_fill_2 FILLER_57_594 ();
 sg13g2_fill_1 FILLER_57_596 ();
 sg13g2_fill_1 FILLER_57_601 ();
 sg13g2_decap_8 FILLER_57_606 ();
 sg13g2_decap_4 FILLER_57_613 ();
 sg13g2_fill_1 FILLER_57_617 ();
 sg13g2_fill_2 FILLER_57_644 ();
 sg13g2_fill_1 FILLER_57_676 ();
 sg13g2_fill_2 FILLER_57_697 ();
 sg13g2_fill_2 FILLER_57_733 ();
 sg13g2_fill_1 FILLER_57_746 ();
 sg13g2_fill_1 FILLER_57_789 ();
 sg13g2_fill_1 FILLER_57_825 ();
 sg13g2_fill_1 FILLER_57_856 ();
 sg13g2_fill_2 FILLER_57_861 ();
 sg13g2_fill_1 FILLER_57_873 ();
 sg13g2_fill_1 FILLER_57_878 ();
 sg13g2_fill_2 FILLER_57_905 ();
 sg13g2_fill_2 FILLER_57_911 ();
 sg13g2_decap_4 FILLER_57_918 ();
 sg13g2_decap_4 FILLER_57_962 ();
 sg13g2_fill_1 FILLER_57_996 ();
 sg13g2_fill_1 FILLER_57_1001 ();
 sg13g2_fill_1 FILLER_57_1011 ();
 sg13g2_fill_1 FILLER_57_1038 ();
 sg13g2_fill_1 FILLER_57_1049 ();
 sg13g2_fill_1 FILLER_57_1071 ();
 sg13g2_decap_8 FILLER_57_1076 ();
 sg13g2_decap_8 FILLER_57_1083 ();
 sg13g2_fill_2 FILLER_57_1090 ();
 sg13g2_fill_1 FILLER_57_1092 ();
 sg13g2_fill_2 FILLER_57_1149 ();
 sg13g2_fill_2 FILLER_57_1176 ();
 sg13g2_fill_1 FILLER_57_1190 ();
 sg13g2_decap_8 FILLER_57_1240 ();
 sg13g2_fill_2 FILLER_57_1247 ();
 sg13g2_fill_1 FILLER_57_1253 ();
 sg13g2_fill_1 FILLER_57_1302 ();
 sg13g2_decap_8 FILLER_57_1311 ();
 sg13g2_decap_4 FILLER_57_1318 ();
 sg13g2_fill_1 FILLER_57_1327 ();
 sg13g2_fill_1 FILLER_57_1340 ();
 sg13g2_fill_2 FILLER_57_1357 ();
 sg13g2_fill_1 FILLER_57_1363 ();
 sg13g2_fill_1 FILLER_57_1368 ();
 sg13g2_fill_1 FILLER_57_1374 ();
 sg13g2_decap_4 FILLER_57_1379 ();
 sg13g2_decap_4 FILLER_57_1387 ();
 sg13g2_fill_1 FILLER_57_1395 ();
 sg13g2_fill_2 FILLER_57_1402 ();
 sg13g2_fill_1 FILLER_57_1409 ();
 sg13g2_fill_2 FILLER_57_1436 ();
 sg13g2_fill_1 FILLER_57_1438 ();
 sg13g2_decap_8 FILLER_57_1457 ();
 sg13g2_decap_8 FILLER_57_1464 ();
 sg13g2_fill_2 FILLER_57_1471 ();
 sg13g2_decap_4 FILLER_57_1482 ();
 sg13g2_fill_1 FILLER_57_1486 ();
 sg13g2_fill_1 FILLER_57_1522 ();
 sg13g2_fill_2 FILLER_57_1563 ();
 sg13g2_decap_8 FILLER_57_1570 ();
 sg13g2_decap_8 FILLER_57_1577 ();
 sg13g2_fill_1 FILLER_57_1584 ();
 sg13g2_decap_4 FILLER_57_1599 ();
 sg13g2_fill_1 FILLER_57_1603 ();
 sg13g2_decap_4 FILLER_57_1608 ();
 sg13g2_fill_2 FILLER_57_1622 ();
 sg13g2_fill_1 FILLER_57_1624 ();
 sg13g2_decap_8 FILLER_57_1628 ();
 sg13g2_decap_4 FILLER_57_1641 ();
 sg13g2_decap_4 FILLER_57_1649 ();
 sg13g2_decap_8 FILLER_57_1657 ();
 sg13g2_decap_8 FILLER_57_1664 ();
 sg13g2_decap_8 FILLER_57_1671 ();
 sg13g2_decap_8 FILLER_57_1678 ();
 sg13g2_fill_1 FILLER_57_1703 ();
 sg13g2_decap_8 FILLER_57_1718 ();
 sg13g2_decap_4 FILLER_57_1725 ();
 sg13g2_fill_2 FILLER_57_1729 ();
 sg13g2_fill_1 FILLER_57_1744 ();
 sg13g2_fill_2 FILLER_57_1771 ();
 sg13g2_decap_8 FILLER_57_1778 ();
 sg13g2_decap_8 FILLER_57_1785 ();
 sg13g2_decap_8 FILLER_57_1792 ();
 sg13g2_decap_8 FILLER_57_1799 ();
 sg13g2_decap_8 FILLER_57_1806 ();
 sg13g2_fill_1 FILLER_57_1813 ();
 sg13g2_decap_8 FILLER_57_1819 ();
 sg13g2_decap_8 FILLER_57_1826 ();
 sg13g2_decap_4 FILLER_57_1833 ();
 sg13g2_fill_2 FILLER_57_1837 ();
 sg13g2_fill_1 FILLER_57_1844 ();
 sg13g2_fill_1 FILLER_57_1856 ();
 sg13g2_fill_1 FILLER_57_1863 ();
 sg13g2_fill_1 FILLER_57_1875 ();
 sg13g2_decap_4 FILLER_57_1907 ();
 sg13g2_fill_1 FILLER_57_1911 ();
 sg13g2_decap_4 FILLER_57_1921 ();
 sg13g2_fill_2 FILLER_57_1925 ();
 sg13g2_fill_2 FILLER_57_1931 ();
 sg13g2_fill_1 FILLER_57_1954 ();
 sg13g2_fill_1 FILLER_57_1960 ();
 sg13g2_fill_1 FILLER_57_1994 ();
 sg13g2_fill_2 FILLER_57_2092 ();
 sg13g2_fill_2 FILLER_57_2099 ();
 sg13g2_decap_4 FILLER_57_2106 ();
 sg13g2_decap_4 FILLER_57_2115 ();
 sg13g2_decap_4 FILLER_57_2128 ();
 sg13g2_fill_2 FILLER_57_2132 ();
 sg13g2_fill_2 FILLER_57_2138 ();
 sg13g2_fill_1 FILLER_57_2140 ();
 sg13g2_fill_1 FILLER_57_2150 ();
 sg13g2_fill_1 FILLER_57_2157 ();
 sg13g2_fill_1 FILLER_57_2191 ();
 sg13g2_fill_2 FILLER_57_2221 ();
 sg13g2_fill_2 FILLER_57_2228 ();
 sg13g2_fill_1 FILLER_57_2239 ();
 sg13g2_fill_1 FILLER_57_2245 ();
 sg13g2_fill_2 FILLER_57_2251 ();
 sg13g2_fill_2 FILLER_57_2283 ();
 sg13g2_fill_1 FILLER_57_2290 ();
 sg13g2_fill_1 FILLER_57_2334 ();
 sg13g2_decap_8 FILLER_57_2355 ();
 sg13g2_fill_2 FILLER_57_2362 ();
 sg13g2_fill_2 FILLER_57_2369 ();
 sg13g2_decap_4 FILLER_57_2388 ();
 sg13g2_fill_1 FILLER_57_2392 ();
 sg13g2_decap_8 FILLER_57_2397 ();
 sg13g2_fill_1 FILLER_57_2404 ();
 sg13g2_fill_2 FILLER_57_2471 ();
 sg13g2_fill_1 FILLER_57_2473 ();
 sg13g2_decap_4 FILLER_57_2500 ();
 sg13g2_fill_1 FILLER_57_2504 ();
 sg13g2_decap_4 FILLER_57_2510 ();
 sg13g2_fill_1 FILLER_57_2523 ();
 sg13g2_fill_1 FILLER_57_2559 ();
 sg13g2_decap_8 FILLER_57_2565 ();
 sg13g2_decap_8 FILLER_57_2582 ();
 sg13g2_decap_8 FILLER_57_2599 ();
 sg13g2_fill_2 FILLER_57_2606 ();
 sg13g2_fill_1 FILLER_57_2608 ();
 sg13g2_decap_8 FILLER_57_2613 ();
 sg13g2_decap_8 FILLER_57_2620 ();
 sg13g2_decap_8 FILLER_57_2627 ();
 sg13g2_decap_8 FILLER_57_2634 ();
 sg13g2_decap_8 FILLER_57_2641 ();
 sg13g2_decap_8 FILLER_57_2648 ();
 sg13g2_decap_8 FILLER_57_2655 ();
 sg13g2_decap_8 FILLER_57_2662 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_fill_1 FILLER_58_76 ();
 sg13g2_fill_2 FILLER_58_100 ();
 sg13g2_fill_2 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_144 ();
 sg13g2_fill_2 FILLER_58_150 ();
 sg13g2_fill_2 FILLER_58_157 ();
 sg13g2_fill_2 FILLER_58_163 ();
 sg13g2_decap_4 FILLER_58_169 ();
 sg13g2_decap_8 FILLER_58_177 ();
 sg13g2_decap_4 FILLER_58_184 ();
 sg13g2_decap_8 FILLER_58_218 ();
 sg13g2_decap_8 FILLER_58_225 ();
 sg13g2_decap_4 FILLER_58_232 ();
 sg13g2_fill_1 FILLER_58_236 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_249 ();
 sg13g2_fill_1 FILLER_58_255 ();
 sg13g2_fill_1 FILLER_58_261 ();
 sg13g2_fill_1 FILLER_58_280 ();
 sg13g2_fill_2 FILLER_58_285 ();
 sg13g2_fill_2 FILLER_58_298 ();
 sg13g2_fill_1 FILLER_58_300 ();
 sg13g2_fill_2 FILLER_58_344 ();
 sg13g2_fill_2 FILLER_58_356 ();
 sg13g2_decap_8 FILLER_58_388 ();
 sg13g2_decap_8 FILLER_58_395 ();
 sg13g2_fill_1 FILLER_58_402 ();
 sg13g2_fill_1 FILLER_58_411 ();
 sg13g2_fill_1 FILLER_58_450 ();
 sg13g2_fill_2 FILLER_58_463 ();
 sg13g2_decap_8 FILLER_58_500 ();
 sg13g2_decap_8 FILLER_58_507 ();
 sg13g2_fill_1 FILLER_58_514 ();
 sg13g2_decap_8 FILLER_58_519 ();
 sg13g2_decap_4 FILLER_58_526 ();
 sg13g2_fill_2 FILLER_58_530 ();
 sg13g2_fill_1 FILLER_58_536 ();
 sg13g2_fill_2 FILLER_58_607 ();
 sg13g2_fill_1 FILLER_58_609 ();
 sg13g2_decap_8 FILLER_58_614 ();
 sg13g2_decap_4 FILLER_58_621 ();
 sg13g2_fill_2 FILLER_58_788 ();
 sg13g2_fill_1 FILLER_58_847 ();
 sg13g2_fill_2 FILLER_58_890 ();
 sg13g2_fill_2 FILLER_58_960 ();
 sg13g2_decap_8 FILLER_58_1005 ();
 sg13g2_fill_2 FILLER_58_1012 ();
 sg13g2_decap_4 FILLER_58_1024 ();
 sg13g2_fill_2 FILLER_58_1028 ();
 sg13g2_fill_2 FILLER_58_1081 ();
 sg13g2_fill_1 FILLER_58_1083 ();
 sg13g2_decap_8 FILLER_58_1136 ();
 sg13g2_decap_4 FILLER_58_1143 ();
 sg13g2_fill_2 FILLER_58_1147 ();
 sg13g2_fill_1 FILLER_58_1185 ();
 sg13g2_fill_1 FILLER_58_1206 ();
 sg13g2_fill_2 FILLER_58_1210 ();
 sg13g2_fill_2 FILLER_58_1232 ();
 sg13g2_fill_1 FILLER_58_1234 ();
 sg13g2_fill_2 FILLER_58_1240 ();
 sg13g2_fill_2 FILLER_58_1253 ();
 sg13g2_fill_1 FILLER_58_1259 ();
 sg13g2_decap_4 FILLER_58_1274 ();
 sg13g2_fill_1 FILLER_58_1278 ();
 sg13g2_decap_4 FILLER_58_1284 ();
 sg13g2_fill_1 FILLER_58_1304 ();
 sg13g2_fill_2 FILLER_58_1313 ();
 sg13g2_fill_1 FILLER_58_1315 ();
 sg13g2_decap_4 FILLER_58_1321 ();
 sg13g2_fill_2 FILLER_58_1333 ();
 sg13g2_fill_2 FILLER_58_1343 ();
 sg13g2_decap_4 FILLER_58_1359 ();
 sg13g2_fill_1 FILLER_58_1363 ();
 sg13g2_decap_4 FILLER_58_1368 ();
 sg13g2_fill_1 FILLER_58_1372 ();
 sg13g2_fill_2 FILLER_58_1382 ();
 sg13g2_fill_1 FILLER_58_1403 ();
 sg13g2_decap_4 FILLER_58_1434 ();
 sg13g2_fill_2 FILLER_58_1438 ();
 sg13g2_fill_2 FILLER_58_1444 ();
 sg13g2_decap_8 FILLER_58_1451 ();
 sg13g2_decap_8 FILLER_58_1458 ();
 sg13g2_fill_2 FILLER_58_1465 ();
 sg13g2_fill_1 FILLER_58_1467 ();
 sg13g2_decap_8 FILLER_58_1477 ();
 sg13g2_fill_1 FILLER_58_1484 ();
 sg13g2_decap_4 FILLER_58_1511 ();
 sg13g2_fill_1 FILLER_58_1515 ();
 sg13g2_fill_1 FILLER_58_1524 ();
 sg13g2_fill_1 FILLER_58_1560 ();
 sg13g2_fill_1 FILLER_58_1565 ();
 sg13g2_fill_2 FILLER_58_1570 ();
 sg13g2_decap_8 FILLER_58_1584 ();
 sg13g2_fill_1 FILLER_58_1591 ();
 sg13g2_decap_4 FILLER_58_1596 ();
 sg13g2_fill_2 FILLER_58_1600 ();
 sg13g2_decap_4 FILLER_58_1607 ();
 sg13g2_decap_8 FILLER_58_1615 ();
 sg13g2_fill_1 FILLER_58_1622 ();
 sg13g2_decap_8 FILLER_58_1636 ();
 sg13g2_decap_8 FILLER_58_1643 ();
 sg13g2_decap_8 FILLER_58_1650 ();
 sg13g2_fill_2 FILLER_58_1657 ();
 sg13g2_fill_1 FILLER_58_1659 ();
 sg13g2_decap_4 FILLER_58_1666 ();
 sg13g2_fill_1 FILLER_58_1700 ();
 sg13g2_fill_2 FILLER_58_1721 ();
 sg13g2_decap_8 FILLER_58_1739 ();
 sg13g2_fill_2 FILLER_58_1746 ();
 sg13g2_fill_1 FILLER_58_1748 ();
 sg13g2_decap_4 FILLER_58_1771 ();
 sg13g2_fill_1 FILLER_58_1784 ();
 sg13g2_decap_8 FILLER_58_1794 ();
 sg13g2_decap_8 FILLER_58_1801 ();
 sg13g2_fill_2 FILLER_58_1808 ();
 sg13g2_fill_1 FILLER_58_1810 ();
 sg13g2_decap_4 FILLER_58_1851 ();
 sg13g2_fill_1 FILLER_58_1859 ();
 sg13g2_fill_1 FILLER_58_1882 ();
 sg13g2_decap_4 FILLER_58_1909 ();
 sg13g2_fill_1 FILLER_58_1913 ();
 sg13g2_decap_4 FILLER_58_1920 ();
 sg13g2_fill_2 FILLER_58_1924 ();
 sg13g2_fill_2 FILLER_58_1945 ();
 sg13g2_fill_2 FILLER_58_2030 ();
 sg13g2_fill_1 FILLER_58_2032 ();
 sg13g2_fill_2 FILLER_58_2047 ();
 sg13g2_fill_2 FILLER_58_2079 ();
 sg13g2_fill_1 FILLER_58_2086 ();
 sg13g2_fill_2 FILLER_58_2092 ();
 sg13g2_fill_1 FILLER_58_2098 ();
 sg13g2_fill_2 FILLER_58_2142 ();
 sg13g2_fill_1 FILLER_58_2144 ();
 sg13g2_fill_2 FILLER_58_2151 ();
 sg13g2_fill_2 FILLER_58_2169 ();
 sg13g2_fill_1 FILLER_58_2182 ();
 sg13g2_fill_2 FILLER_58_2198 ();
 sg13g2_fill_1 FILLER_58_2204 ();
 sg13g2_fill_1 FILLER_58_2209 ();
 sg13g2_fill_2 FILLER_58_2249 ();
 sg13g2_fill_1 FILLER_58_2261 ();
 sg13g2_fill_1 FILLER_58_2271 ();
 sg13g2_fill_2 FILLER_58_2277 ();
 sg13g2_fill_2 FILLER_58_2313 ();
 sg13g2_fill_1 FILLER_58_2327 ();
 sg13g2_fill_2 FILLER_58_2338 ();
 sg13g2_fill_1 FILLER_58_2345 ();
 sg13g2_fill_2 FILLER_58_2351 ();
 sg13g2_fill_2 FILLER_58_2362 ();
 sg13g2_decap_4 FILLER_58_2373 ();
 sg13g2_fill_1 FILLER_58_2404 ();
 sg13g2_fill_1 FILLER_58_2431 ();
 sg13g2_fill_2 FILLER_58_2452 ();
 sg13g2_decap_4 FILLER_58_2460 ();
 sg13g2_decap_8 FILLER_58_2496 ();
 sg13g2_fill_2 FILLER_58_2503 ();
 sg13g2_fill_1 FILLER_58_2505 ();
 sg13g2_decap_8 FILLER_58_2610 ();
 sg13g2_decap_8 FILLER_58_2617 ();
 sg13g2_decap_8 FILLER_58_2624 ();
 sg13g2_decap_8 FILLER_58_2631 ();
 sg13g2_decap_8 FILLER_58_2638 ();
 sg13g2_decap_8 FILLER_58_2645 ();
 sg13g2_decap_8 FILLER_58_2652 ();
 sg13g2_decap_8 FILLER_58_2659 ();
 sg13g2_decap_4 FILLER_58_2666 ();
 sg13g2_fill_1 FILLER_59_24 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_83 ();
 sg13g2_decap_4 FILLER_59_120 ();
 sg13g2_fill_2 FILLER_59_150 ();
 sg13g2_fill_1 FILLER_59_183 ();
 sg13g2_fill_2 FILLER_59_219 ();
 sg13g2_fill_2 FILLER_59_251 ();
 sg13g2_decap_8 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_285 ();
 sg13g2_decap_4 FILLER_59_292 ();
 sg13g2_fill_2 FILLER_59_296 ();
 sg13g2_fill_2 FILLER_59_306 ();
 sg13g2_fill_1 FILLER_59_308 ();
 sg13g2_fill_1 FILLER_59_315 ();
 sg13g2_fill_1 FILLER_59_323 ();
 sg13g2_decap_4 FILLER_59_328 ();
 sg13g2_fill_1 FILLER_59_332 ();
 sg13g2_fill_2 FILLER_59_338 ();
 sg13g2_fill_1 FILLER_59_348 ();
 sg13g2_fill_2 FILLER_59_354 ();
 sg13g2_decap_4 FILLER_59_361 ();
 sg13g2_fill_1 FILLER_59_369 ();
 sg13g2_decap_8 FILLER_59_374 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_4 FILLER_59_388 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_2 FILLER_59_397 ();
 sg13g2_fill_2 FILLER_59_416 ();
 sg13g2_fill_1 FILLER_59_418 ();
 sg13g2_fill_2 FILLER_59_437 ();
 sg13g2_fill_1 FILLER_59_439 ();
 sg13g2_fill_2 FILLER_59_445 ();
 sg13g2_fill_1 FILLER_59_447 ();
 sg13g2_fill_1 FILLER_59_478 ();
 sg13g2_fill_2 FILLER_59_523 ();
 sg13g2_fill_2 FILLER_59_578 ();
 sg13g2_fill_2 FILLER_59_642 ();
 sg13g2_fill_1 FILLER_59_644 ();
 sg13g2_fill_2 FILLER_59_690 ();
 sg13g2_fill_2 FILLER_59_739 ();
 sg13g2_fill_1 FILLER_59_824 ();
 sg13g2_fill_1 FILLER_59_835 ();
 sg13g2_fill_2 FILLER_59_859 ();
 sg13g2_fill_2 FILLER_59_902 ();
 sg13g2_fill_2 FILLER_59_913 ();
 sg13g2_fill_2 FILLER_59_936 ();
 sg13g2_decap_8 FILLER_59_950 ();
 sg13g2_decap_8 FILLER_59_957 ();
 sg13g2_fill_1 FILLER_59_964 ();
 sg13g2_decap_4 FILLER_59_976 ();
 sg13g2_decap_4 FILLER_59_984 ();
 sg13g2_fill_2 FILLER_59_988 ();
 sg13g2_decap_8 FILLER_59_1007 ();
 sg13g2_fill_1 FILLER_59_1014 ();
 sg13g2_fill_2 FILLER_59_1068 ();
 sg13g2_fill_1 FILLER_59_1106 ();
 sg13g2_decap_4 FILLER_59_1111 ();
 sg13g2_fill_2 FILLER_59_1125 ();
 sg13g2_fill_1 FILLER_59_1127 ();
 sg13g2_decap_8 FILLER_59_1132 ();
 sg13g2_decap_8 FILLER_59_1139 ();
 sg13g2_decap_8 FILLER_59_1146 ();
 sg13g2_fill_2 FILLER_59_1153 ();
 sg13g2_fill_2 FILLER_59_1225 ();
 sg13g2_fill_1 FILLER_59_1237 ();
 sg13g2_fill_1 FILLER_59_1252 ();
 sg13g2_fill_1 FILLER_59_1261 ();
 sg13g2_fill_2 FILLER_59_1276 ();
 sg13g2_decap_4 FILLER_59_1282 ();
 sg13g2_decap_4 FILLER_59_1291 ();
 sg13g2_fill_1 FILLER_59_1295 ();
 sg13g2_decap_8 FILLER_59_1313 ();
 sg13g2_decap_4 FILLER_59_1324 ();
 sg13g2_fill_2 FILLER_59_1328 ();
 sg13g2_fill_1 FILLER_59_1340 ();
 sg13g2_fill_1 FILLER_59_1387 ();
 sg13g2_fill_2 FILLER_59_1409 ();
 sg13g2_fill_2 FILLER_59_1416 ();
 sg13g2_fill_1 FILLER_59_1418 ();
 sg13g2_decap_4 FILLER_59_1445 ();
 sg13g2_fill_1 FILLER_59_1449 ();
 sg13g2_fill_2 FILLER_59_1454 ();
 sg13g2_decap_4 FILLER_59_1468 ();
 sg13g2_decap_8 FILLER_59_1476 ();
 sg13g2_decap_8 FILLER_59_1483 ();
 sg13g2_decap_8 FILLER_59_1495 ();
 sg13g2_decap_4 FILLER_59_1502 ();
 sg13g2_fill_1 FILLER_59_1506 ();
 sg13g2_decap_4 FILLER_59_1510 ();
 sg13g2_fill_2 FILLER_59_1518 ();
 sg13g2_fill_2 FILLER_59_1528 ();
 sg13g2_fill_1 FILLER_59_1539 ();
 sg13g2_decap_8 FILLER_59_1546 ();
 sg13g2_decap_8 FILLER_59_1553 ();
 sg13g2_decap_8 FILLER_59_1560 ();
 sg13g2_decap_8 FILLER_59_1567 ();
 sg13g2_decap_8 FILLER_59_1579 ();
 sg13g2_fill_2 FILLER_59_1586 ();
 sg13g2_fill_1 FILLER_59_1618 ();
 sg13g2_fill_2 FILLER_59_1624 ();
 sg13g2_fill_2 FILLER_59_1632 ();
 sg13g2_fill_2 FILLER_59_1644 ();
 sg13g2_fill_1 FILLER_59_1646 ();
 sg13g2_fill_1 FILLER_59_1656 ();
 sg13g2_fill_2 FILLER_59_1666 ();
 sg13g2_fill_2 FILLER_59_1673 ();
 sg13g2_fill_1 FILLER_59_1675 ();
 sg13g2_fill_1 FILLER_59_1681 ();
 sg13g2_fill_1 FILLER_59_1691 ();
 sg13g2_fill_1 FILLER_59_1759 ();
 sg13g2_fill_1 FILLER_59_1769 ();
 sg13g2_fill_2 FILLER_59_1774 ();
 sg13g2_fill_1 FILLER_59_1781 ();
 sg13g2_decap_4 FILLER_59_1795 ();
 sg13g2_fill_2 FILLER_59_1799 ();
 sg13g2_fill_2 FILLER_59_1805 ();
 sg13g2_decap_8 FILLER_59_1812 ();
 sg13g2_fill_1 FILLER_59_1819 ();
 sg13g2_decap_4 FILLER_59_1829 ();
 sg13g2_fill_2 FILLER_59_1833 ();
 sg13g2_decap_4 FILLER_59_1843 ();
 sg13g2_fill_2 FILLER_59_1847 ();
 sg13g2_decap_8 FILLER_59_1859 ();
 sg13g2_fill_2 FILLER_59_1866 ();
 sg13g2_decap_4 FILLER_59_1878 ();
 sg13g2_fill_2 FILLER_59_1882 ();
 sg13g2_fill_2 FILLER_59_1888 ();
 sg13g2_decap_8 FILLER_59_1894 ();
 sg13g2_decap_4 FILLER_59_1901 ();
 sg13g2_fill_2 FILLER_59_1905 ();
 sg13g2_decap_8 FILLER_59_1995 ();
 sg13g2_decap_4 FILLER_59_2002 ();
 sg13g2_fill_2 FILLER_59_2006 ();
 sg13g2_fill_1 FILLER_59_2044 ();
 sg13g2_fill_1 FILLER_59_2050 ();
 sg13g2_fill_1 FILLER_59_2056 ();
 sg13g2_fill_1 FILLER_59_2061 ();
 sg13g2_fill_1 FILLER_59_2066 ();
 sg13g2_decap_8 FILLER_59_2072 ();
 sg13g2_decap_8 FILLER_59_2079 ();
 sg13g2_fill_2 FILLER_59_2086 ();
 sg13g2_fill_1 FILLER_59_2088 ();
 sg13g2_decap_8 FILLER_59_2135 ();
 sg13g2_decap_8 FILLER_59_2142 ();
 sg13g2_fill_1 FILLER_59_2149 ();
 sg13g2_fill_2 FILLER_59_2162 ();
 sg13g2_fill_1 FILLER_59_2171 ();
 sg13g2_fill_1 FILLER_59_2177 ();
 sg13g2_fill_1 FILLER_59_2183 ();
 sg13g2_fill_1 FILLER_59_2270 ();
 sg13g2_fill_1 FILLER_59_2279 ();
 sg13g2_fill_1 FILLER_59_2315 ();
 sg13g2_fill_1 FILLER_59_2320 ();
 sg13g2_fill_2 FILLER_59_2383 ();
 sg13g2_fill_2 FILLER_59_2390 ();
 sg13g2_decap_8 FILLER_59_2400 ();
 sg13g2_fill_1 FILLER_59_2413 ();
 sg13g2_fill_1 FILLER_59_2418 ();
 sg13g2_fill_1 FILLER_59_2423 ();
 sg13g2_fill_1 FILLER_59_2434 ();
 sg13g2_fill_1 FILLER_59_2448 ();
 sg13g2_fill_2 FILLER_59_2475 ();
 sg13g2_fill_1 FILLER_59_2477 ();
 sg13g2_fill_2 FILLER_59_2495 ();
 sg13g2_fill_1 FILLER_59_2497 ();
 sg13g2_decap_4 FILLER_59_2516 ();
 sg13g2_fill_1 FILLER_59_2535 ();
 sg13g2_fill_1 FILLER_59_2541 ();
 sg13g2_fill_2 FILLER_59_2551 ();
 sg13g2_fill_1 FILLER_59_2558 ();
 sg13g2_fill_1 FILLER_59_2563 ();
 sg13g2_fill_2 FILLER_59_2577 ();
 sg13g2_fill_1 FILLER_59_2579 ();
 sg13g2_decap_8 FILLER_59_2606 ();
 sg13g2_decap_8 FILLER_59_2613 ();
 sg13g2_decap_8 FILLER_59_2620 ();
 sg13g2_decap_8 FILLER_59_2627 ();
 sg13g2_decap_8 FILLER_59_2634 ();
 sg13g2_decap_8 FILLER_59_2641 ();
 sg13g2_decap_8 FILLER_59_2648 ();
 sg13g2_decap_8 FILLER_59_2655 ();
 sg13g2_decap_8 FILLER_59_2662 ();
 sg13g2_fill_1 FILLER_59_2669 ();
 sg13g2_fill_1 FILLER_60_13 ();
 sg13g2_fill_2 FILLER_60_73 ();
 sg13g2_fill_2 FILLER_60_89 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_2 FILLER_60_112 ();
 sg13g2_fill_2 FILLER_60_119 ();
 sg13g2_fill_2 FILLER_60_157 ();
 sg13g2_decap_8 FILLER_60_216 ();
 sg13g2_decap_4 FILLER_60_223 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_decap_4 FILLER_60_299 ();
 sg13g2_fill_2 FILLER_60_303 ();
 sg13g2_decap_4 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_366 ();
 sg13g2_decap_8 FILLER_60_372 ();
 sg13g2_decap_4 FILLER_60_379 ();
 sg13g2_fill_1 FILLER_60_388 ();
 sg13g2_fill_1 FILLER_60_402 ();
 sg13g2_fill_1 FILLER_60_458 ();
 sg13g2_fill_1 FILLER_60_495 ();
 sg13g2_fill_2 FILLER_60_501 ();
 sg13g2_fill_1 FILLER_60_525 ();
 sg13g2_fill_2 FILLER_60_532 ();
 sg13g2_fill_1 FILLER_60_539 ();
 sg13g2_fill_2 FILLER_60_566 ();
 sg13g2_decap_8 FILLER_60_576 ();
 sg13g2_decap_4 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_587 ();
 sg13g2_decap_4 FILLER_60_594 ();
 sg13g2_fill_2 FILLER_60_634 ();
 sg13g2_fill_1 FILLER_60_636 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_decap_8 FILLER_60_708 ();
 sg13g2_decap_8 FILLER_60_720 ();
 sg13g2_fill_1 FILLER_60_753 ();
 sg13g2_fill_1 FILLER_60_758 ();
 sg13g2_fill_1 FILLER_60_814 ();
 sg13g2_decap_4 FILLER_60_866 ();
 sg13g2_fill_1 FILLER_60_876 ();
 sg13g2_fill_2 FILLER_60_885 ();
 sg13g2_fill_1 FILLER_60_887 ();
 sg13g2_fill_1 FILLER_60_900 ();
 sg13g2_decap_8 FILLER_60_983 ();
 sg13g2_decap_8 FILLER_60_990 ();
 sg13g2_fill_2 FILLER_60_997 ();
 sg13g2_decap_8 FILLER_60_1009 ();
 sg13g2_decap_8 FILLER_60_1016 ();
 sg13g2_fill_2 FILLER_60_1023 ();
 sg13g2_fill_1 FILLER_60_1025 ();
 sg13g2_decap_8 FILLER_60_1030 ();
 sg13g2_decap_4 FILLER_60_1037 ();
 sg13g2_fill_2 FILLER_60_1077 ();
 sg13g2_fill_1 FILLER_60_1079 ();
 sg13g2_decap_8 FILLER_60_1101 ();
 sg13g2_decap_4 FILLER_60_1108 ();
 sg13g2_fill_1 FILLER_60_1112 ();
 sg13g2_fill_2 FILLER_60_1121 ();
 sg13g2_decap_8 FILLER_60_1144 ();
 sg13g2_fill_1 FILLER_60_1151 ();
 sg13g2_fill_1 FILLER_60_1185 ();
 sg13g2_fill_1 FILLER_60_1194 ();
 sg13g2_decap_4 FILLER_60_1199 ();
 sg13g2_fill_1 FILLER_60_1203 ();
 sg13g2_decap_4 FILLER_60_1217 ();
 sg13g2_fill_1 FILLER_60_1243 ();
 sg13g2_fill_1 FILLER_60_1249 ();
 sg13g2_fill_1 FILLER_60_1260 ();
 sg13g2_fill_1 FILLER_60_1266 ();
 sg13g2_decap_8 FILLER_60_1298 ();
 sg13g2_fill_1 FILLER_60_1305 ();
 sg13g2_decap_4 FILLER_60_1335 ();
 sg13g2_decap_8 FILLER_60_1342 ();
 sg13g2_decap_4 FILLER_60_1349 ();
 sg13g2_fill_1 FILLER_60_1362 ();
 sg13g2_decap_8 FILLER_60_1367 ();
 sg13g2_fill_1 FILLER_60_1374 ();
 sg13g2_fill_1 FILLER_60_1383 ();
 sg13g2_fill_1 FILLER_60_1388 ();
 sg13g2_fill_1 FILLER_60_1405 ();
 sg13g2_fill_1 FILLER_60_1415 ();
 sg13g2_decap_4 FILLER_60_1421 ();
 sg13g2_fill_1 FILLER_60_1425 ();
 sg13g2_fill_2 FILLER_60_1443 ();
 sg13g2_fill_1 FILLER_60_1445 ();
 sg13g2_fill_2 FILLER_60_1464 ();
 sg13g2_decap_8 FILLER_60_1476 ();
 sg13g2_fill_1 FILLER_60_1483 ();
 sg13g2_decap_4 FILLER_60_1493 ();
 sg13g2_fill_2 FILLER_60_1501 ();
 sg13g2_decap_8 FILLER_60_1507 ();
 sg13g2_decap_8 FILLER_60_1514 ();
 sg13g2_decap_8 FILLER_60_1521 ();
 sg13g2_decap_8 FILLER_60_1528 ();
 sg13g2_decap_8 FILLER_60_1535 ();
 sg13g2_decap_8 FILLER_60_1542 ();
 sg13g2_decap_8 FILLER_60_1549 ();
 sg13g2_decap_8 FILLER_60_1556 ();
 sg13g2_fill_2 FILLER_60_1563 ();
 sg13g2_fill_1 FILLER_60_1565 ();
 sg13g2_fill_2 FILLER_60_1578 ();
 sg13g2_fill_1 FILLER_60_1580 ();
 sg13g2_decap_8 FILLER_60_1585 ();
 sg13g2_fill_2 FILLER_60_1592 ();
 sg13g2_decap_8 FILLER_60_1598 ();
 sg13g2_decap_4 FILLER_60_1605 ();
 sg13g2_fill_1 FILLER_60_1609 ();
 sg13g2_fill_1 FILLER_60_1623 ();
 sg13g2_fill_2 FILLER_60_1640 ();
 sg13g2_fill_1 FILLER_60_1642 ();
 sg13g2_fill_1 FILLER_60_1658 ();
 sg13g2_fill_1 FILLER_60_1672 ();
 sg13g2_fill_2 FILLER_60_1678 ();
 sg13g2_decap_4 FILLER_60_1708 ();
 sg13g2_fill_2 FILLER_60_1717 ();
 sg13g2_fill_1 FILLER_60_1719 ();
 sg13g2_fill_1 FILLER_60_1749 ();
 sg13g2_fill_2 FILLER_60_1768 ();
 sg13g2_fill_1 FILLER_60_1770 ();
 sg13g2_fill_1 FILLER_60_1780 ();
 sg13g2_fill_1 FILLER_60_1790 ();
 sg13g2_fill_2 FILLER_60_1795 ();
 sg13g2_fill_2 FILLER_60_1811 ();
 sg13g2_decap_8 FILLER_60_1817 ();
 sg13g2_decap_8 FILLER_60_1824 ();
 sg13g2_decap_8 FILLER_60_1831 ();
 sg13g2_decap_8 FILLER_60_1838 ();
 sg13g2_fill_2 FILLER_60_1845 ();
 sg13g2_decap_8 FILLER_60_1903 ();
 sg13g2_decap_4 FILLER_60_1910 ();
 sg13g2_decap_4 FILLER_60_1920 ();
 sg13g2_fill_1 FILLER_60_1924 ();
 sg13g2_fill_1 FILLER_60_1950 ();
 sg13g2_decap_8 FILLER_60_1992 ();
 sg13g2_decap_4 FILLER_60_1999 ();
 sg13g2_decap_4 FILLER_60_2012 ();
 sg13g2_fill_1 FILLER_60_2029 ();
 sg13g2_decap_8 FILLER_60_2056 ();
 sg13g2_decap_8 FILLER_60_2063 ();
 sg13g2_fill_2 FILLER_60_2070 ();
 sg13g2_fill_1 FILLER_60_2100 ();
 sg13g2_fill_1 FILLER_60_2127 ();
 sg13g2_decap_4 FILLER_60_2132 ();
 sg13g2_fill_1 FILLER_60_2136 ();
 sg13g2_decap_8 FILLER_60_2141 ();
 sg13g2_decap_8 FILLER_60_2148 ();
 sg13g2_decap_4 FILLER_60_2155 ();
 sg13g2_fill_1 FILLER_60_2159 ();
 sg13g2_fill_2 FILLER_60_2182 ();
 sg13g2_fill_2 FILLER_60_2230 ();
 sg13g2_fill_1 FILLER_60_2236 ();
 sg13g2_fill_2 FILLER_60_2301 ();
 sg13g2_fill_2 FILLER_60_2310 ();
 sg13g2_decap_8 FILLER_60_2395 ();
 sg13g2_decap_8 FILLER_60_2402 ();
 sg13g2_decap_4 FILLER_60_2422 ();
 sg13g2_fill_1 FILLER_60_2426 ();
 sg13g2_fill_2 FILLER_60_2433 ();
 sg13g2_fill_2 FILLER_60_2440 ();
 sg13g2_decap_4 FILLER_60_2463 ();
 sg13g2_fill_1 FILLER_60_2535 ();
 sg13g2_decap_8 FILLER_60_2615 ();
 sg13g2_decap_8 FILLER_60_2622 ();
 sg13g2_decap_8 FILLER_60_2629 ();
 sg13g2_decap_8 FILLER_60_2636 ();
 sg13g2_decap_8 FILLER_60_2643 ();
 sg13g2_decap_8 FILLER_60_2650 ();
 sg13g2_decap_8 FILLER_60_2657 ();
 sg13g2_decap_4 FILLER_60_2664 ();
 sg13g2_fill_2 FILLER_60_2668 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_27 ();
 sg13g2_fill_1 FILLER_61_38 ();
 sg13g2_fill_1 FILLER_61_80 ();
 sg13g2_fill_2 FILLER_61_107 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_fill_2 FILLER_61_140 ();
 sg13g2_fill_1 FILLER_61_152 ();
 sg13g2_fill_1 FILLER_61_158 ();
 sg13g2_fill_1 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_175 ();
 sg13g2_fill_2 FILLER_61_187 ();
 sg13g2_fill_1 FILLER_61_308 ();
 sg13g2_fill_1 FILLER_61_321 ();
 sg13g2_fill_2 FILLER_61_348 ();
 sg13g2_fill_1 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_61_356 ();
 sg13g2_fill_1 FILLER_61_420 ();
 sg13g2_fill_1 FILLER_61_427 ();
 sg13g2_fill_1 FILLER_61_456 ();
 sg13g2_fill_2 FILLER_61_475 ();
 sg13g2_fill_1 FILLER_61_482 ();
 sg13g2_fill_1 FILLER_61_514 ();
 sg13g2_fill_2 FILLER_61_521 ();
 sg13g2_fill_1 FILLER_61_536 ();
 sg13g2_fill_1 FILLER_61_542 ();
 sg13g2_fill_2 FILLER_61_548 ();
 sg13g2_fill_2 FILLER_61_554 ();
 sg13g2_fill_2 FILLER_61_586 ();
 sg13g2_fill_1 FILLER_61_588 ();
 sg13g2_decap_4 FILLER_61_594 ();
 sg13g2_fill_2 FILLER_61_598 ();
 sg13g2_fill_1 FILLER_61_639 ();
 sg13g2_fill_1 FILLER_61_648 ();
 sg13g2_fill_1 FILLER_61_659 ();
 sg13g2_fill_1 FILLER_61_686 ();
 sg13g2_fill_1 FILLER_61_718 ();
 sg13g2_fill_2 FILLER_61_755 ();
 sg13g2_decap_4 FILLER_61_763 ();
 sg13g2_fill_2 FILLER_61_767 ();
 sg13g2_decap_4 FILLER_61_794 ();
 sg13g2_fill_2 FILLER_61_809 ();
 sg13g2_decap_4 FILLER_61_870 ();
 sg13g2_fill_1 FILLER_61_874 ();
 sg13g2_fill_2 FILLER_61_880 ();
 sg13g2_fill_2 FILLER_61_901 ();
 sg13g2_fill_1 FILLER_61_903 ();
 sg13g2_fill_2 FILLER_61_923 ();
 sg13g2_fill_1 FILLER_61_982 ();
 sg13g2_fill_1 FILLER_61_1031 ();
 sg13g2_fill_1 FILLER_61_1036 ();
 sg13g2_fill_2 FILLER_61_1047 ();
 sg13g2_fill_1 FILLER_61_1053 ();
 sg13g2_fill_2 FILLER_61_1093 ();
 sg13g2_fill_2 FILLER_61_1131 ();
 sg13g2_fill_1 FILLER_61_1133 ();
 sg13g2_decap_8 FILLER_61_1170 ();
 sg13g2_decap_4 FILLER_61_1177 ();
 sg13g2_fill_1 FILLER_61_1181 ();
 sg13g2_decap_4 FILLER_61_1188 ();
 sg13g2_fill_2 FILLER_61_1192 ();
 sg13g2_fill_1 FILLER_61_1241 ();
 sg13g2_fill_2 FILLER_61_1268 ();
 sg13g2_fill_1 FILLER_61_1270 ();
 sg13g2_fill_2 FILLER_61_1274 ();
 sg13g2_decap_8 FILLER_61_1280 ();
 sg13g2_decap_8 FILLER_61_1287 ();
 sg13g2_decap_4 FILLER_61_1294 ();
 sg13g2_fill_1 FILLER_61_1305 ();
 sg13g2_fill_1 FILLER_61_1343 ();
 sg13g2_decap_8 FILLER_61_1348 ();
 sg13g2_decap_8 FILLER_61_1355 ();
 sg13g2_decap_8 FILLER_61_1362 ();
 sg13g2_decap_8 FILLER_61_1369 ();
 sg13g2_decap_4 FILLER_61_1376 ();
 sg13g2_fill_2 FILLER_61_1380 ();
 sg13g2_decap_4 FILLER_61_1386 ();
 sg13g2_fill_2 FILLER_61_1390 ();
 sg13g2_decap_4 FILLER_61_1396 ();
 sg13g2_fill_2 FILLER_61_1400 ();
 sg13g2_fill_2 FILLER_61_1411 ();
 sg13g2_fill_1 FILLER_61_1418 ();
 sg13g2_fill_1 FILLER_61_1423 ();
 sg13g2_decap_8 FILLER_61_1432 ();
 sg13g2_fill_2 FILLER_61_1443 ();
 sg13g2_fill_1 FILLER_61_1471 ();
 sg13g2_fill_1 FILLER_61_1485 ();
 sg13g2_fill_2 FILLER_61_1490 ();
 sg13g2_fill_2 FILLER_61_1497 ();
 sg13g2_decap_8 FILLER_61_1503 ();
 sg13g2_decap_8 FILLER_61_1510 ();
 sg13g2_decap_4 FILLER_61_1517 ();
 sg13g2_fill_2 FILLER_61_1525 ();
 sg13g2_fill_1 FILLER_61_1527 ();
 sg13g2_fill_1 FILLER_61_1552 ();
 sg13g2_decap_4 FILLER_61_1590 ();
 sg13g2_decap_8 FILLER_61_1602 ();
 sg13g2_fill_2 FILLER_61_1609 ();
 sg13g2_decap_8 FILLER_61_1615 ();
 sg13g2_fill_1 FILLER_61_1635 ();
 sg13g2_fill_2 FILLER_61_1649 ();
 sg13g2_fill_1 FILLER_61_1659 ();
 sg13g2_fill_1 FILLER_61_1699 ();
 sg13g2_fill_2 FILLER_61_1705 ();
 sg13g2_fill_2 FILLER_61_1712 ();
 sg13g2_decap_8 FILLER_61_1732 ();
 sg13g2_fill_1 FILLER_61_1739 ();
 sg13g2_decap_4 FILLER_61_1754 ();
 sg13g2_fill_2 FILLER_61_1762 ();
 sg13g2_fill_2 FILLER_61_1769 ();
 sg13g2_decap_4 FILLER_61_1776 ();
 sg13g2_fill_1 FILLER_61_1825 ();
 sg13g2_decap_8 FILLER_61_1830 ();
 sg13g2_fill_2 FILLER_61_1837 ();
 sg13g2_decap_8 FILLER_61_1872 ();
 sg13g2_fill_2 FILLER_61_1879 ();
 sg13g2_decap_8 FILLER_61_1894 ();
 sg13g2_decap_8 FILLER_61_1901 ();
 sg13g2_fill_2 FILLER_61_1908 ();
 sg13g2_fill_1 FILLER_61_1910 ();
 sg13g2_fill_1 FILLER_61_1935 ();
 sg13g2_fill_1 FILLER_61_1948 ();
 sg13g2_fill_2 FILLER_61_1962 ();
 sg13g2_fill_1 FILLER_61_1972 ();
 sg13g2_fill_1 FILLER_61_1981 ();
 sg13g2_fill_1 FILLER_61_1986 ();
 sg13g2_fill_1 FILLER_61_1992 ();
 sg13g2_fill_1 FILLER_61_1997 ();
 sg13g2_fill_1 FILLER_61_2076 ();
 sg13g2_fill_1 FILLER_61_2103 ();
 sg13g2_fill_2 FILLER_61_2121 ();
 sg13g2_fill_2 FILLER_61_2165 ();
 sg13g2_fill_1 FILLER_61_2167 ();
 sg13g2_fill_2 FILLER_61_2173 ();
 sg13g2_fill_1 FILLER_61_2186 ();
 sg13g2_fill_2 FILLER_61_2192 ();
 sg13g2_fill_2 FILLER_61_2198 ();
 sg13g2_fill_1 FILLER_61_2205 ();
 sg13g2_fill_1 FILLER_61_2210 ();
 sg13g2_fill_1 FILLER_61_2226 ();
 sg13g2_fill_1 FILLER_61_2235 ();
 sg13g2_fill_1 FILLER_61_2248 ();
 sg13g2_fill_1 FILLER_61_2267 ();
 sg13g2_fill_2 FILLER_61_2309 ();
 sg13g2_fill_1 FILLER_61_2321 ();
 sg13g2_fill_1 FILLER_61_2328 ();
 sg13g2_fill_2 FILLER_61_2341 ();
 sg13g2_fill_2 FILLER_61_2353 ();
 sg13g2_fill_2 FILLER_61_2373 ();
 sg13g2_fill_2 FILLER_61_2394 ();
 sg13g2_decap_4 FILLER_61_2409 ();
 sg13g2_fill_2 FILLER_61_2413 ();
 sg13g2_fill_2 FILLER_61_2470 ();
 sg13g2_fill_1 FILLER_61_2472 ();
 sg13g2_decap_8 FILLER_61_2533 ();
 sg13g2_decap_8 FILLER_61_2550 ();
 sg13g2_decap_8 FILLER_61_2557 ();
 sg13g2_decap_4 FILLER_61_2564 ();
 sg13g2_fill_2 FILLER_61_2568 ();
 sg13g2_fill_2 FILLER_61_2584 ();
 sg13g2_decap_8 FILLER_61_2612 ();
 sg13g2_decap_8 FILLER_61_2619 ();
 sg13g2_decap_8 FILLER_61_2626 ();
 sg13g2_decap_8 FILLER_61_2633 ();
 sg13g2_decap_8 FILLER_61_2640 ();
 sg13g2_decap_8 FILLER_61_2647 ();
 sg13g2_decap_8 FILLER_61_2654 ();
 sg13g2_decap_8 FILLER_61_2661 ();
 sg13g2_fill_2 FILLER_61_2668 ();
 sg13g2_fill_2 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_74 ();
 sg13g2_fill_2 FILLER_62_86 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_fill_1 FILLER_62_102 ();
 sg13g2_fill_1 FILLER_62_136 ();
 sg13g2_decap_8 FILLER_62_141 ();
 sg13g2_decap_4 FILLER_62_148 ();
 sg13g2_fill_2 FILLER_62_152 ();
 sg13g2_decap_8 FILLER_62_159 ();
 sg13g2_fill_1 FILLER_62_171 ();
 sg13g2_fill_1 FILLER_62_183 ();
 sg13g2_fill_2 FILLER_62_245 ();
 sg13g2_fill_1 FILLER_62_267 ();
 sg13g2_fill_1 FILLER_62_277 ();
 sg13g2_fill_2 FILLER_62_287 ();
 sg13g2_fill_2 FILLER_62_318 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_fill_2 FILLER_62_421 ();
 sg13g2_fill_2 FILLER_62_431 ();
 sg13g2_fill_1 FILLER_62_433 ();
 sg13g2_fill_1 FILLER_62_449 ();
 sg13g2_fill_1 FILLER_62_455 ();
 sg13g2_fill_1 FILLER_62_468 ();
 sg13g2_fill_1 FILLER_62_498 ();
 sg13g2_fill_1 FILLER_62_503 ();
 sg13g2_fill_2 FILLER_62_512 ();
 sg13g2_fill_1 FILLER_62_514 ();
 sg13g2_decap_4 FILLER_62_536 ();
 sg13g2_fill_2 FILLER_62_554 ();
 sg13g2_decap_4 FILLER_62_561 ();
 sg13g2_decap_4 FILLER_62_569 ();
 sg13g2_fill_1 FILLER_62_599 ();
 sg13g2_fill_2 FILLER_62_630 ();
 sg13g2_decap_8 FILLER_62_636 ();
 sg13g2_fill_1 FILLER_62_643 ();
 sg13g2_decap_4 FILLER_62_652 ();
 sg13g2_decap_8 FILLER_62_660 ();
 sg13g2_decap_8 FILLER_62_671 ();
 sg13g2_decap_8 FILLER_62_678 ();
 sg13g2_fill_2 FILLER_62_685 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_758 ();
 sg13g2_decap_4 FILLER_62_765 ();
 sg13g2_fill_2 FILLER_62_775 ();
 sg13g2_fill_2 FILLER_62_782 ();
 sg13g2_fill_1 FILLER_62_789 ();
 sg13g2_fill_2 FILLER_62_858 ();
 sg13g2_decap_4 FILLER_62_865 ();
 sg13g2_fill_2 FILLER_62_876 ();
 sg13g2_fill_1 FILLER_62_913 ();
 sg13g2_decap_8 FILLER_62_931 ();
 sg13g2_fill_2 FILLER_62_938 ();
 sg13g2_fill_1 FILLER_62_940 ();
 sg13g2_decap_4 FILLER_62_950 ();
 sg13g2_decap_4 FILLER_62_959 ();
 sg13g2_fill_2 FILLER_62_967 ();
 sg13g2_fill_1 FILLER_62_973 ();
 sg13g2_fill_2 FILLER_62_978 ();
 sg13g2_fill_1 FILLER_62_988 ();
 sg13g2_fill_2 FILLER_62_1032 ();
 sg13g2_fill_1 FILLER_62_1043 ();
 sg13g2_fill_2 FILLER_62_1061 ();
 sg13g2_fill_1 FILLER_62_1063 ();
 sg13g2_fill_2 FILLER_62_1068 ();
 sg13g2_fill_2 FILLER_62_1096 ();
 sg13g2_fill_1 FILLER_62_1098 ();
 sg13g2_fill_1 FILLER_62_1135 ();
 sg13g2_fill_1 FILLER_62_1176 ();
 sg13g2_fill_1 FILLER_62_1182 ();
 sg13g2_fill_2 FILLER_62_1222 ();
 sg13g2_fill_1 FILLER_62_1224 ();
 sg13g2_decap_8 FILLER_62_1229 ();
 sg13g2_decap_8 FILLER_62_1236 ();
 sg13g2_fill_1 FILLER_62_1243 ();
 sg13g2_fill_1 FILLER_62_1248 ();
 sg13g2_decap_8 FILLER_62_1253 ();
 sg13g2_fill_1 FILLER_62_1260 ();
 sg13g2_decap_4 FILLER_62_1266 ();
 sg13g2_fill_1 FILLER_62_1270 ();
 sg13g2_fill_1 FILLER_62_1277 ();
 sg13g2_decap_8 FILLER_62_1282 ();
 sg13g2_fill_1 FILLER_62_1289 ();
 sg13g2_fill_1 FILLER_62_1300 ();
 sg13g2_fill_1 FILLER_62_1310 ();
 sg13g2_decap_8 FILLER_62_1329 ();
 sg13g2_decap_4 FILLER_62_1336 ();
 sg13g2_fill_1 FILLER_62_1340 ();
 sg13g2_decap_4 FILLER_62_1366 ();
 sg13g2_fill_1 FILLER_62_1370 ();
 sg13g2_fill_2 FILLER_62_1392 ();
 sg13g2_fill_1 FILLER_62_1394 ();
 sg13g2_fill_2 FILLER_62_1407 ();
 sg13g2_fill_2 FILLER_62_1414 ();
 sg13g2_fill_1 FILLER_62_1416 ();
 sg13g2_fill_1 FILLER_62_1426 ();
 sg13g2_decap_4 FILLER_62_1440 ();
 sg13g2_fill_2 FILLER_62_1444 ();
 sg13g2_fill_1 FILLER_62_1462 ();
 sg13g2_fill_1 FILLER_62_1468 ();
 sg13g2_fill_2 FILLER_62_1473 ();
 sg13g2_fill_1 FILLER_62_1505 ();
 sg13g2_fill_1 FILLER_62_1511 ();
 sg13g2_fill_1 FILLER_62_1520 ();
 sg13g2_fill_2 FILLER_62_1525 ();
 sg13g2_fill_1 FILLER_62_1527 ();
 sg13g2_fill_1 FILLER_62_1532 ();
 sg13g2_fill_2 FILLER_62_1585 ();
 sg13g2_decap_8 FILLER_62_1591 ();
 sg13g2_decap_4 FILLER_62_1598 ();
 sg13g2_fill_1 FILLER_62_1602 ();
 sg13g2_decap_8 FILLER_62_1607 ();
 sg13g2_fill_1 FILLER_62_1614 ();
 sg13g2_fill_1 FILLER_62_1629 ();
 sg13g2_decap_8 FILLER_62_1638 ();
 sg13g2_fill_2 FILLER_62_1658 ();
 sg13g2_fill_1 FILLER_62_1660 ();
 sg13g2_fill_2 FILLER_62_1665 ();
 sg13g2_fill_2 FILLER_62_1678 ();
 sg13g2_fill_2 FILLER_62_1694 ();
 sg13g2_fill_1 FILLER_62_1696 ();
 sg13g2_decap_4 FILLER_62_1728 ();
 sg13g2_fill_1 FILLER_62_1732 ();
 sg13g2_fill_2 FILLER_62_1743 ();
 sg13g2_fill_1 FILLER_62_1745 ();
 sg13g2_fill_1 FILLER_62_1751 ();
 sg13g2_fill_1 FILLER_62_1779 ();
 sg13g2_fill_2 FILLER_62_1784 ();
 sg13g2_fill_1 FILLER_62_1786 ();
 sg13g2_fill_1 FILLER_62_1805 ();
 sg13g2_decap_4 FILLER_62_1832 ();
 sg13g2_fill_1 FILLER_62_1836 ();
 sg13g2_decap_4 FILLER_62_1842 ();
 sg13g2_fill_2 FILLER_62_1846 ();
 sg13g2_decap_8 FILLER_62_1865 ();
 sg13g2_decap_8 FILLER_62_1872 ();
 sg13g2_fill_2 FILLER_62_1879 ();
 sg13g2_fill_2 FILLER_62_1902 ();
 sg13g2_fill_2 FILLER_62_1914 ();
 sg13g2_fill_2 FILLER_62_1936 ();
 sg13g2_fill_2 FILLER_62_1946 ();
 sg13g2_fill_1 FILLER_62_1962 ();
 sg13g2_fill_1 FILLER_62_1976 ();
 sg13g2_fill_1 FILLER_62_2003 ();
 sg13g2_fill_2 FILLER_62_2030 ();
 sg13g2_fill_2 FILLER_62_2036 ();
 sg13g2_fill_2 FILLER_62_2043 ();
 sg13g2_fill_1 FILLER_62_2045 ();
 sg13g2_decap_4 FILLER_62_2059 ();
 sg13g2_fill_2 FILLER_62_2105 ();
 sg13g2_fill_2 FILLER_62_2115 ();
 sg13g2_decap_8 FILLER_62_2122 ();
 sg13g2_decap_4 FILLER_62_2159 ();
 sg13g2_fill_2 FILLER_62_2163 ();
 sg13g2_fill_1 FILLER_62_2170 ();
 sg13g2_decap_4 FILLER_62_2180 ();
 sg13g2_fill_1 FILLER_62_2184 ();
 sg13g2_fill_1 FILLER_62_2207 ();
 sg13g2_fill_1 FILLER_62_2212 ();
 sg13g2_fill_1 FILLER_62_2217 ();
 sg13g2_fill_2 FILLER_62_2249 ();
 sg13g2_fill_1 FILLER_62_2292 ();
 sg13g2_decap_8 FILLER_62_2334 ();
 sg13g2_decap_8 FILLER_62_2341 ();
 sg13g2_decap_4 FILLER_62_2348 ();
 sg13g2_fill_2 FILLER_62_2352 ();
 sg13g2_decap_8 FILLER_62_2364 ();
 sg13g2_decap_4 FILLER_62_2371 ();
 sg13g2_fill_1 FILLER_62_2375 ();
 sg13g2_fill_2 FILLER_62_2393 ();
 sg13g2_fill_2 FILLER_62_2453 ();
 sg13g2_fill_2 FILLER_62_2461 ();
 sg13g2_fill_1 FILLER_62_2489 ();
 sg13g2_decap_4 FILLER_62_2499 ();
 sg13g2_fill_1 FILLER_62_2503 ();
 sg13g2_fill_1 FILLER_62_2513 ();
 sg13g2_fill_2 FILLER_62_2542 ();
 sg13g2_fill_1 FILLER_62_2606 ();
 sg13g2_decap_8 FILLER_62_2614 ();
 sg13g2_decap_8 FILLER_62_2621 ();
 sg13g2_decap_8 FILLER_62_2628 ();
 sg13g2_decap_8 FILLER_62_2635 ();
 sg13g2_decap_8 FILLER_62_2642 ();
 sg13g2_decap_8 FILLER_62_2649 ();
 sg13g2_decap_8 FILLER_62_2656 ();
 sg13g2_decap_8 FILLER_62_2663 ();
 sg13g2_fill_1 FILLER_63_0 ();
 sg13g2_fill_1 FILLER_63_27 ();
 sg13g2_fill_1 FILLER_63_38 ();
 sg13g2_fill_1 FILLER_63_43 ();
 sg13g2_fill_2 FILLER_63_78 ();
 sg13g2_decap_8 FILLER_63_83 ();
 sg13g2_decap_8 FILLER_63_90 ();
 sg13g2_decap_8 FILLER_63_97 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_150 ();
 sg13g2_fill_1 FILLER_63_192 ();
 sg13g2_fill_2 FILLER_63_244 ();
 sg13g2_fill_2 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_decap_8 FILLER_63_320 ();
 sg13g2_fill_2 FILLER_63_327 ();
 sg13g2_decap_8 FILLER_63_333 ();
 sg13g2_fill_2 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_4 FILLER_63_385 ();
 sg13g2_decap_4 FILLER_63_398 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_4 FILLER_63_478 ();
 sg13g2_fill_1 FILLER_63_482 ();
 sg13g2_decap_4 FILLER_63_492 ();
 sg13g2_fill_1 FILLER_63_496 ();
 sg13g2_decap_4 FILLER_63_501 ();
 sg13g2_fill_1 FILLER_63_505 ();
 sg13g2_fill_1 FILLER_63_510 ();
 sg13g2_fill_2 FILLER_63_551 ();
 sg13g2_fill_1 FILLER_63_583 ();
 sg13g2_fill_1 FILLER_63_588 ();
 sg13g2_decap_8 FILLER_63_593 ();
 sg13g2_decap_4 FILLER_63_600 ();
 sg13g2_fill_2 FILLER_63_604 ();
 sg13g2_decap_8 FILLER_63_620 ();
 sg13g2_decap_8 FILLER_63_627 ();
 sg13g2_fill_1 FILLER_63_634 ();
 sg13g2_decap_4 FILLER_63_639 ();
 sg13g2_fill_2 FILLER_63_643 ();
 sg13g2_fill_2 FILLER_63_650 ();
 sg13g2_decap_8 FILLER_63_673 ();
 sg13g2_fill_1 FILLER_63_684 ();
 sg13g2_decap_8 FILLER_63_793 ();
 sg13g2_decap_8 FILLER_63_800 ();
 sg13g2_fill_2 FILLER_63_807 ();
 sg13g2_fill_1 FILLER_63_809 ();
 sg13g2_decap_8 FILLER_63_814 ();
 sg13g2_decap_4 FILLER_63_821 ();
 sg13g2_fill_2 FILLER_63_825 ();
 sg13g2_decap_8 FILLER_63_852 ();
 sg13g2_decap_4 FILLER_63_859 ();
 sg13g2_fill_1 FILLER_63_863 ();
 sg13g2_fill_2 FILLER_63_894 ();
 sg13g2_fill_1 FILLER_63_896 ();
 sg13g2_fill_1 FILLER_63_915 ();
 sg13g2_fill_1 FILLER_63_945 ();
 sg13g2_fill_1 FILLER_63_950 ();
 sg13g2_fill_2 FILLER_63_959 ();
 sg13g2_fill_2 FILLER_63_971 ();
 sg13g2_fill_2 FILLER_63_978 ();
 sg13g2_decap_4 FILLER_63_996 ();
 sg13g2_fill_2 FILLER_63_1000 ();
 sg13g2_decap_4 FILLER_63_1039 ();
 sg13g2_fill_1 FILLER_63_1043 ();
 sg13g2_decap_4 FILLER_63_1047 ();
 sg13g2_fill_1 FILLER_63_1051 ();
 sg13g2_fill_2 FILLER_63_1056 ();
 sg13g2_fill_1 FILLER_63_1077 ();
 sg13g2_decap_8 FILLER_63_1104 ();
 sg13g2_fill_2 FILLER_63_1111 ();
 sg13g2_fill_2 FILLER_63_1117 ();
 sg13g2_fill_1 FILLER_63_1119 ();
 sg13g2_decap_8 FILLER_63_1124 ();
 sg13g2_fill_2 FILLER_63_1131 ();
 sg13g2_decap_8 FILLER_63_1138 ();
 sg13g2_decap_8 FILLER_63_1145 ();
 sg13g2_fill_1 FILLER_63_1152 ();
 sg13g2_decap_8 FILLER_63_1157 ();
 sg13g2_decap_8 FILLER_63_1164 ();
 sg13g2_fill_1 FILLER_63_1171 ();
 sg13g2_decap_8 FILLER_63_1176 ();
 sg13g2_decap_8 FILLER_63_1183 ();
 sg13g2_decap_4 FILLER_63_1194 ();
 sg13g2_decap_8 FILLER_63_1201 ();
 sg13g2_decap_4 FILLER_63_1233 ();
 sg13g2_fill_1 FILLER_63_1237 ();
 sg13g2_fill_1 FILLER_63_1271 ();
 sg13g2_fill_1 FILLER_63_1302 ();
 sg13g2_fill_2 FILLER_63_1329 ();
 sg13g2_fill_2 FILLER_63_1338 ();
 sg13g2_fill_1 FILLER_63_1340 ();
 sg13g2_fill_1 FILLER_63_1353 ();
 sg13g2_fill_1 FILLER_63_1359 ();
 sg13g2_fill_1 FILLER_63_1365 ();
 sg13g2_fill_1 FILLER_63_1374 ();
 sg13g2_fill_2 FILLER_63_1388 ();
 sg13g2_fill_2 FILLER_63_1408 ();
 sg13g2_fill_1 FILLER_63_1410 ();
 sg13g2_fill_2 FILLER_63_1415 ();
 sg13g2_decap_4 FILLER_63_1422 ();
 sg13g2_fill_2 FILLER_63_1432 ();
 sg13g2_fill_1 FILLER_63_1434 ();
 sg13g2_fill_1 FILLER_63_1448 ();
 sg13g2_fill_2 FILLER_63_1484 ();
 sg13g2_fill_1 FILLER_63_1545 ();
 sg13g2_fill_2 FILLER_63_1560 ();
 sg13g2_fill_2 FILLER_63_1585 ();
 sg13g2_decap_8 FILLER_63_1592 ();
 sg13g2_decap_8 FILLER_63_1599 ();
 sg13g2_decap_4 FILLER_63_1606 ();
 sg13g2_fill_2 FILLER_63_1610 ();
 sg13g2_decap_4 FILLER_63_1616 ();
 sg13g2_decap_4 FILLER_63_1624 ();
 sg13g2_fill_1 FILLER_63_1628 ();
 sg13g2_fill_1 FILLER_63_1641 ();
 sg13g2_fill_2 FILLER_63_1665 ();
 sg13g2_fill_1 FILLER_63_1698 ();
 sg13g2_fill_2 FILLER_63_1704 ();
 sg13g2_fill_2 FILLER_63_1738 ();
 sg13g2_fill_2 FILLER_63_1750 ();
 sg13g2_decap_4 FILLER_63_1757 ();
 sg13g2_fill_2 FILLER_63_1761 ();
 sg13g2_fill_2 FILLER_63_1776 ();
 sg13g2_fill_1 FILLER_63_1783 ();
 sg13g2_fill_2 FILLER_63_1795 ();
 sg13g2_fill_1 FILLER_63_1802 ();
 sg13g2_decap_8 FILLER_63_1846 ();
 sg13g2_fill_1 FILLER_63_1853 ();
 sg13g2_fill_1 FILLER_63_1885 ();
 sg13g2_decap_4 FILLER_63_1912 ();
 sg13g2_fill_1 FILLER_63_1916 ();
 sg13g2_fill_1 FILLER_63_1931 ();
 sg13g2_decap_8 FILLER_63_1942 ();
 sg13g2_decap_4 FILLER_63_1949 ();
 sg13g2_fill_2 FILLER_63_1953 ();
 sg13g2_fill_1 FILLER_63_2030 ();
 sg13g2_fill_2 FILLER_63_2037 ();
 sg13g2_fill_2 FILLER_63_2065 ();
 sg13g2_fill_2 FILLER_63_2072 ();
 sg13g2_fill_1 FILLER_63_2083 ();
 sg13g2_fill_1 FILLER_63_2088 ();
 sg13g2_fill_1 FILLER_63_2093 ();
 sg13g2_fill_1 FILLER_63_2099 ();
 sg13g2_fill_1 FILLER_63_2105 ();
 sg13g2_fill_1 FILLER_63_2116 ();
 sg13g2_decap_4 FILLER_63_2165 ();
 sg13g2_decap_4 FILLER_63_2179 ();
 sg13g2_fill_1 FILLER_63_2183 ();
 sg13g2_fill_2 FILLER_63_2197 ();
 sg13g2_fill_1 FILLER_63_2199 ();
 sg13g2_fill_1 FILLER_63_2270 ();
 sg13g2_fill_1 FILLER_63_2309 ();
 sg13g2_fill_2 FILLER_63_2317 ();
 sg13g2_fill_1 FILLER_63_2326 ();
 sg13g2_fill_2 FILLER_63_2342 ();
 sg13g2_decap_4 FILLER_63_2349 ();
 sg13g2_decap_4 FILLER_63_2358 ();
 sg13g2_decap_4 FILLER_63_2388 ();
 sg13g2_fill_1 FILLER_63_2434 ();
 sg13g2_fill_1 FILLER_63_2441 ();
 sg13g2_decap_8 FILLER_63_2475 ();
 sg13g2_fill_1 FILLER_63_2482 ();
 sg13g2_decap_4 FILLER_63_2493 ();
 sg13g2_fill_1 FILLER_63_2497 ();
 sg13g2_fill_1 FILLER_63_2507 ();
 sg13g2_fill_1 FILLER_63_2595 ();
 sg13g2_fill_1 FILLER_63_2600 ();
 sg13g2_decap_8 FILLER_63_2627 ();
 sg13g2_decap_8 FILLER_63_2634 ();
 sg13g2_decap_8 FILLER_63_2641 ();
 sg13g2_decap_8 FILLER_63_2648 ();
 sg13g2_decap_8 FILLER_63_2655 ();
 sg13g2_decap_8 FILLER_63_2662 ();
 sg13g2_fill_1 FILLER_63_2669 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_decap_4 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_77 ();
 sg13g2_decap_4 FILLER_64_82 ();
 sg13g2_fill_2 FILLER_64_90 ();
 sg13g2_fill_2 FILLER_64_118 ();
 sg13g2_fill_2 FILLER_64_131 ();
 sg13g2_fill_1 FILLER_64_164 ();
 sg13g2_fill_2 FILLER_64_174 ();
 sg13g2_fill_1 FILLER_64_176 ();
 sg13g2_decap_8 FILLER_64_181 ();
 sg13g2_decap_8 FILLER_64_188 ();
 sg13g2_decap_8 FILLER_64_195 ();
 sg13g2_decap_8 FILLER_64_202 ();
 sg13g2_decap_4 FILLER_64_231 ();
 sg13g2_fill_2 FILLER_64_235 ();
 sg13g2_fill_1 FILLER_64_265 ();
 sg13g2_fill_1 FILLER_64_271 ();
 sg13g2_fill_2 FILLER_64_277 ();
 sg13g2_decap_4 FILLER_64_301 ();
 sg13g2_fill_2 FILLER_64_305 ();
 sg13g2_decap_4 FILLER_64_310 ();
 sg13g2_fill_1 FILLER_64_314 ();
 sg13g2_decap_8 FILLER_64_320 ();
 sg13g2_decap_4 FILLER_64_327 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_decap_8 FILLER_64_342 ();
 sg13g2_decap_4 FILLER_64_349 ();
 sg13g2_fill_2 FILLER_64_358 ();
 sg13g2_fill_1 FILLER_64_360 ();
 sg13g2_decap_4 FILLER_64_378 ();
 sg13g2_fill_2 FILLER_64_386 ();
 sg13g2_decap_8 FILLER_64_397 ();
 sg13g2_decap_8 FILLER_64_413 ();
 sg13g2_decap_8 FILLER_64_420 ();
 sg13g2_decap_8 FILLER_64_427 ();
 sg13g2_fill_1 FILLER_64_434 ();
 sg13g2_decap_4 FILLER_64_439 ();
 sg13g2_decap_8 FILLER_64_446 ();
 sg13g2_decap_4 FILLER_64_453 ();
 sg13g2_decap_4 FILLER_64_465 ();
 sg13g2_fill_1 FILLER_64_469 ();
 sg13g2_fill_2 FILLER_64_496 ();
 sg13g2_fill_1 FILLER_64_498 ();
 sg13g2_decap_8 FILLER_64_504 ();
 sg13g2_fill_2 FILLER_64_511 ();
 sg13g2_fill_1 FILLER_64_521 ();
 sg13g2_fill_1 FILLER_64_526 ();
 sg13g2_fill_1 FILLER_64_532 ();
 sg13g2_fill_2 FILLER_64_538 ();
 sg13g2_fill_1 FILLER_64_540 ();
 sg13g2_fill_1 FILLER_64_547 ();
 sg13g2_decap_4 FILLER_64_553 ();
 sg13g2_decap_8 FILLER_64_561 ();
 sg13g2_decap_8 FILLER_64_568 ();
 sg13g2_decap_8 FILLER_64_575 ();
 sg13g2_decap_8 FILLER_64_582 ();
 sg13g2_decap_8 FILLER_64_589 ();
 sg13g2_decap_8 FILLER_64_596 ();
 sg13g2_decap_8 FILLER_64_603 ();
 sg13g2_fill_2 FILLER_64_610 ();
 sg13g2_fill_2 FILLER_64_648 ();
 sg13g2_fill_1 FILLER_64_694 ();
 sg13g2_decap_8 FILLER_64_703 ();
 sg13g2_fill_1 FILLER_64_710 ();
 sg13g2_decap_8 FILLER_64_719 ();
 sg13g2_decap_8 FILLER_64_726 ();
 sg13g2_fill_2 FILLER_64_733 ();
 sg13g2_fill_2 FILLER_64_760 ();
 sg13g2_fill_1 FILLER_64_766 ();
 sg13g2_fill_1 FILLER_64_787 ();
 sg13g2_fill_1 FILLER_64_798 ();
 sg13g2_fill_1 FILLER_64_825 ();
 sg13g2_fill_1 FILLER_64_832 ();
 sg13g2_fill_1 FILLER_64_838 ();
 sg13g2_fill_2 FILLER_64_854 ();
 sg13g2_decap_8 FILLER_64_859 ();
 sg13g2_decap_8 FILLER_64_866 ();
 sg13g2_decap_4 FILLER_64_888 ();
 sg13g2_fill_2 FILLER_64_918 ();
 sg13g2_fill_1 FILLER_64_959 ();
 sg13g2_fill_1 FILLER_64_986 ();
 sg13g2_fill_1 FILLER_64_1018 ();
 sg13g2_fill_2 FILLER_64_1026 ();
 sg13g2_fill_1 FILLER_64_1038 ();
 sg13g2_decap_8 FILLER_64_1044 ();
 sg13g2_decap_8 FILLER_64_1051 ();
 sg13g2_decap_4 FILLER_64_1058 ();
 sg13g2_fill_1 FILLER_64_1065 ();
 sg13g2_decap_8 FILLER_64_1097 ();
 sg13g2_fill_1 FILLER_64_1104 ();
 sg13g2_decap_8 FILLER_64_1141 ();
 sg13g2_decap_4 FILLER_64_1152 ();
 sg13g2_fill_1 FILLER_64_1156 ();
 sg13g2_decap_4 FILLER_64_1162 ();
 sg13g2_decap_8 FILLER_64_1176 ();
 sg13g2_fill_2 FILLER_64_1183 ();
 sg13g2_fill_1 FILLER_64_1185 ();
 sg13g2_fill_2 FILLER_64_1196 ();
 sg13g2_fill_2 FILLER_64_1223 ();
 sg13g2_fill_2 FILLER_64_1233 ();
 sg13g2_fill_2 FILLER_64_1254 ();
 sg13g2_decap_4 FILLER_64_1260 ();
 sg13g2_fill_2 FILLER_64_1264 ();
 sg13g2_fill_1 FILLER_64_1293 ();
 sg13g2_fill_1 FILLER_64_1299 ();
 sg13g2_fill_2 FILLER_64_1328 ();
 sg13g2_fill_1 FILLER_64_1343 ();
 sg13g2_fill_1 FILLER_64_1357 ();
 sg13g2_fill_1 FILLER_64_1363 ();
 sg13g2_fill_1 FILLER_64_1382 ();
 sg13g2_fill_1 FILLER_64_1388 ();
 sg13g2_fill_1 FILLER_64_1393 ();
 sg13g2_fill_1 FILLER_64_1400 ();
 sg13g2_fill_2 FILLER_64_1406 ();
 sg13g2_fill_2 FILLER_64_1426 ();
 sg13g2_fill_1 FILLER_64_1428 ();
 sg13g2_decap_4 FILLER_64_1434 ();
 sg13g2_fill_1 FILLER_64_1438 ();
 sg13g2_fill_2 FILLER_64_1497 ();
 sg13g2_decap_4 FILLER_64_1552 ();
 sg13g2_fill_1 FILLER_64_1556 ();
 sg13g2_decap_4 FILLER_64_1561 ();
 sg13g2_decap_8 FILLER_64_1586 ();
 sg13g2_decap_8 FILLER_64_1593 ();
 sg13g2_decap_8 FILLER_64_1600 ();
 sg13g2_decap_8 FILLER_64_1607 ();
 sg13g2_decap_4 FILLER_64_1614 ();
 sg13g2_fill_2 FILLER_64_1628 ();
 sg13g2_fill_2 FILLER_64_1638 ();
 sg13g2_fill_1 FILLER_64_1645 ();
 sg13g2_decap_4 FILLER_64_1665 ();
 sg13g2_fill_2 FILLER_64_1690 ();
 sg13g2_fill_1 FILLER_64_1731 ();
 sg13g2_fill_1 FILLER_64_1736 ();
 sg13g2_fill_1 FILLER_64_1743 ();
 sg13g2_decap_4 FILLER_64_1757 ();
 sg13g2_fill_1 FILLER_64_1792 ();
 sg13g2_fill_1 FILLER_64_1797 ();
 sg13g2_fill_1 FILLER_64_1807 ();
 sg13g2_fill_2 FILLER_64_1854 ();
 sg13g2_fill_1 FILLER_64_1856 ();
 sg13g2_decap_4 FILLER_64_1868 ();
 sg13g2_decap_8 FILLER_64_1876 ();
 sg13g2_decap_8 FILLER_64_1883 ();
 sg13g2_decap_4 FILLER_64_1890 ();
 sg13g2_fill_1 FILLER_64_1894 ();
 sg13g2_decap_8 FILLER_64_1899 ();
 sg13g2_decap_4 FILLER_64_1937 ();
 sg13g2_fill_1 FILLER_64_2015 ();
 sg13g2_decap_4 FILLER_64_2042 ();
 sg13g2_fill_2 FILLER_64_2050 ();
 sg13g2_fill_1 FILLER_64_2052 ();
 sg13g2_fill_2 FILLER_64_2057 ();
 sg13g2_fill_1 FILLER_64_2059 ();
 sg13g2_decap_4 FILLER_64_2065 ();
 sg13g2_fill_1 FILLER_64_2069 ();
 sg13g2_decap_8 FILLER_64_2084 ();
 sg13g2_fill_2 FILLER_64_2091 ();
 sg13g2_decap_4 FILLER_64_2097 ();
 sg13g2_fill_1 FILLER_64_2105 ();
 sg13g2_fill_2 FILLER_64_2115 ();
 sg13g2_fill_1 FILLER_64_2117 ();
 sg13g2_fill_2 FILLER_64_2138 ();
 sg13g2_decap_8 FILLER_64_2164 ();
 sg13g2_decap_8 FILLER_64_2171 ();
 sg13g2_fill_1 FILLER_64_2235 ();
 sg13g2_fill_1 FILLER_64_2241 ();
 sg13g2_fill_1 FILLER_64_2262 ();
 sg13g2_decap_8 FILLER_64_2275 ();
 sg13g2_fill_1 FILLER_64_2282 ();
 sg13g2_fill_1 FILLER_64_2294 ();
 sg13g2_fill_1 FILLER_64_2303 ();
 sg13g2_fill_2 FILLER_64_2335 ();
 sg13g2_decap_8 FILLER_64_2359 ();
 sg13g2_fill_2 FILLER_64_2366 ();
 sg13g2_decap_8 FILLER_64_2372 ();
 sg13g2_decap_4 FILLER_64_2379 ();
 sg13g2_fill_2 FILLER_64_2399 ();
 sg13g2_fill_1 FILLER_64_2401 ();
 sg13g2_decap_4 FILLER_64_2406 ();
 sg13g2_fill_2 FILLER_64_2410 ();
 sg13g2_fill_2 FILLER_64_2422 ();
 sg13g2_fill_1 FILLER_64_2457 ();
 sg13g2_fill_2 FILLER_64_2516 ();
 sg13g2_decap_8 FILLER_64_2631 ();
 sg13g2_decap_8 FILLER_64_2638 ();
 sg13g2_decap_8 FILLER_64_2645 ();
 sg13g2_decap_8 FILLER_64_2652 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_4 FILLER_64_2666 ();
 sg13g2_decap_4 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_4 ();
 sg13g2_decap_8 FILLER_65_13 ();
 sg13g2_fill_2 FILLER_65_20 ();
 sg13g2_fill_1 FILLER_65_22 ();
 sg13g2_decap_8 FILLER_65_31 ();
 sg13g2_decap_4 FILLER_65_38 ();
 sg13g2_fill_1 FILLER_65_42 ();
 sg13g2_fill_1 FILLER_65_52 ();
 sg13g2_fill_1 FILLER_65_59 ();
 sg13g2_fill_2 FILLER_65_83 ();
 sg13g2_fill_2 FILLER_65_90 ();
 sg13g2_fill_1 FILLER_65_92 ();
 sg13g2_fill_1 FILLER_65_114 ();
 sg13g2_decap_4 FILLER_65_120 ();
 sg13g2_fill_2 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_194 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_fill_2 FILLER_65_211 ();
 sg13g2_fill_1 FILLER_65_213 ();
 sg13g2_fill_2 FILLER_65_226 ();
 sg13g2_fill_1 FILLER_65_228 ();
 sg13g2_fill_2 FILLER_65_241 ();
 sg13g2_fill_2 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_304 ();
 sg13g2_decap_8 FILLER_65_341 ();
 sg13g2_decap_8 FILLER_65_348 ();
 sg13g2_decap_4 FILLER_65_355 ();
 sg13g2_fill_2 FILLER_65_359 ();
 sg13g2_fill_2 FILLER_65_443 ();
 sg13g2_fill_2 FILLER_65_459 ();
 sg13g2_decap_8 FILLER_65_465 ();
 sg13g2_fill_2 FILLER_65_472 ();
 sg13g2_fill_1 FILLER_65_474 ();
 sg13g2_fill_2 FILLER_65_482 ();
 sg13g2_decap_8 FILLER_65_496 ();
 sg13g2_fill_2 FILLER_65_503 ();
 sg13g2_fill_1 FILLER_65_516 ();
 sg13g2_decap_4 FILLER_65_521 ();
 sg13g2_fill_2 FILLER_65_534 ();
 sg13g2_fill_1 FILLER_65_536 ();
 sg13g2_fill_1 FILLER_65_542 ();
 sg13g2_fill_1 FILLER_65_547 ();
 sg13g2_fill_2 FILLER_65_556 ();
 sg13g2_decap_8 FILLER_65_588 ();
 sg13g2_decap_4 FILLER_65_595 ();
 sg13g2_fill_2 FILLER_65_599 ();
 sg13g2_fill_2 FILLER_65_610 ();
 sg13g2_fill_1 FILLER_65_638 ();
 sg13g2_fill_1 FILLER_65_643 ();
 sg13g2_fill_1 FILLER_65_655 ();
 sg13g2_fill_2 FILLER_65_663 ();
 sg13g2_fill_2 FILLER_65_744 ();
 sg13g2_fill_2 FILLER_65_751 ();
 sg13g2_decap_8 FILLER_65_757 ();
 sg13g2_decap_4 FILLER_65_764 ();
 sg13g2_decap_8 FILLER_65_772 ();
 sg13g2_fill_1 FILLER_65_779 ();
 sg13g2_fill_2 FILLER_65_802 ();
 sg13g2_fill_1 FILLER_65_804 ();
 sg13g2_decap_4 FILLER_65_838 ();
 sg13g2_decap_8 FILLER_65_874 ();
 sg13g2_decap_4 FILLER_65_881 ();
 sg13g2_fill_1 FILLER_65_885 ();
 sg13g2_fill_1 FILLER_65_922 ();
 sg13g2_fill_2 FILLER_65_928 ();
 sg13g2_fill_1 FILLER_65_953 ();
 sg13g2_decap_8 FILLER_65_1020 ();
 sg13g2_fill_1 FILLER_65_1027 ();
 sg13g2_fill_1 FILLER_65_1033 ();
 sg13g2_fill_2 FILLER_65_1039 ();
 sg13g2_fill_1 FILLER_65_1041 ();
 sg13g2_fill_1 FILLER_65_1051 ();
 sg13g2_fill_1 FILLER_65_1064 ();
 sg13g2_fill_1 FILLER_65_1077 ();
 sg13g2_decap_8 FILLER_65_1088 ();
 sg13g2_decap_4 FILLER_65_1105 ();
 sg13g2_fill_1 FILLER_65_1119 ();
 sg13g2_fill_2 FILLER_65_1150 ();
 sg13g2_decap_8 FILLER_65_1169 ();
 sg13g2_decap_8 FILLER_65_1176 ();
 sg13g2_fill_1 FILLER_65_1183 ();
 sg13g2_fill_1 FILLER_65_1214 ();
 sg13g2_fill_1 FILLER_65_1220 ();
 sg13g2_fill_2 FILLER_65_1231 ();
 sg13g2_fill_1 FILLER_65_1233 ();
 sg13g2_decap_4 FILLER_65_1245 ();
 sg13g2_fill_2 FILLER_65_1249 ();
 sg13g2_decap_4 FILLER_65_1259 ();
 sg13g2_fill_2 FILLER_65_1267 ();
 sg13g2_fill_2 FILLER_65_1275 ();
 sg13g2_fill_2 FILLER_65_1283 ();
 sg13g2_fill_1 FILLER_65_1292 ();
 sg13g2_fill_2 FILLER_65_1340 ();
 sg13g2_decap_4 FILLER_65_1346 ();
 sg13g2_decap_8 FILLER_65_1373 ();
 sg13g2_decap_8 FILLER_65_1380 ();
 sg13g2_decap_8 FILLER_65_1398 ();
 sg13g2_fill_2 FILLER_65_1405 ();
 sg13g2_decap_4 FILLER_65_1428 ();
 sg13g2_decap_8 FILLER_65_1437 ();
 sg13g2_decap_8 FILLER_65_1448 ();
 sg13g2_fill_1 FILLER_65_1455 ();
 sg13g2_decap_4 FILLER_65_1461 ();
 sg13g2_fill_2 FILLER_65_1469 ();
 sg13g2_fill_1 FILLER_65_1471 ();
 sg13g2_decap_8 FILLER_65_1497 ();
 sg13g2_decap_4 FILLER_65_1504 ();
 sg13g2_decap_8 FILLER_65_1559 ();
 sg13g2_decap_8 FILLER_65_1566 ();
 sg13g2_decap_8 FILLER_65_1573 ();
 sg13g2_decap_8 FILLER_65_1580 ();
 sg13g2_decap_8 FILLER_65_1587 ();
 sg13g2_decap_8 FILLER_65_1594 ();
 sg13g2_decap_8 FILLER_65_1601 ();
 sg13g2_decap_8 FILLER_65_1608 ();
 sg13g2_fill_2 FILLER_65_1615 ();
 sg13g2_decap_8 FILLER_65_1622 ();
 sg13g2_decap_4 FILLER_65_1676 ();
 sg13g2_fill_2 FILLER_65_1726 ();
 sg13g2_decap_8 FILLER_65_1744 ();
 sg13g2_fill_2 FILLER_65_1756 ();
 sg13g2_decap_4 FILLER_65_1777 ();
 sg13g2_fill_1 FILLER_65_1781 ();
 sg13g2_fill_2 FILLER_65_1796 ();
 sg13g2_fill_1 FILLER_65_1826 ();
 sg13g2_fill_2 FILLER_65_1853 ();
 sg13g2_fill_2 FILLER_65_1859 ();
 sg13g2_decap_8 FILLER_65_1891 ();
 sg13g2_decap_8 FILLER_65_1898 ();
 sg13g2_fill_2 FILLER_65_1905 ();
 sg13g2_fill_1 FILLER_65_1947 ();
 sg13g2_decap_4 FILLER_65_1953 ();
 sg13g2_decap_4 FILLER_65_1966 ();
 sg13g2_decap_8 FILLER_65_1994 ();
 sg13g2_decap_8 FILLER_65_2001 ();
 sg13g2_fill_1 FILLER_65_2008 ();
 sg13g2_fill_1 FILLER_65_2019 ();
 sg13g2_fill_1 FILLER_65_2029 ();
 sg13g2_fill_1 FILLER_65_2034 ();
 sg13g2_fill_2 FILLER_65_2039 ();
 sg13g2_fill_2 FILLER_65_2046 ();
 sg13g2_fill_1 FILLER_65_2048 ();
 sg13g2_decap_4 FILLER_65_2053 ();
 sg13g2_fill_1 FILLER_65_2057 ();
 sg13g2_fill_2 FILLER_65_2075 ();
 sg13g2_fill_1 FILLER_65_2077 ();
 sg13g2_fill_1 FILLER_65_2083 ();
 sg13g2_fill_1 FILLER_65_2088 ();
 sg13g2_fill_1 FILLER_65_2093 ();
 sg13g2_fill_2 FILLER_65_2137 ();
 sg13g2_fill_1 FILLER_65_2139 ();
 sg13g2_decap_4 FILLER_65_2166 ();
 sg13g2_fill_2 FILLER_65_2170 ();
 sg13g2_fill_1 FILLER_65_2181 ();
 sg13g2_decap_4 FILLER_65_2224 ();
 sg13g2_fill_1 FILLER_65_2236 ();
 sg13g2_fill_1 FILLER_65_2247 ();
 sg13g2_fill_1 FILLER_65_2252 ();
 sg13g2_fill_1 FILLER_65_2263 ();
 sg13g2_fill_1 FILLER_65_2268 ();
 sg13g2_decap_4 FILLER_65_2277 ();
 sg13g2_fill_1 FILLER_65_2281 ();
 sg13g2_decap_4 FILLER_65_2309 ();
 sg13g2_fill_2 FILLER_65_2313 ();
 sg13g2_decap_4 FILLER_65_2319 ();
 sg13g2_decap_4 FILLER_65_2337 ();
 sg13g2_fill_2 FILLER_65_2341 ();
 sg13g2_fill_2 FILLER_65_2373 ();
 sg13g2_fill_2 FILLER_65_2401 ();
 sg13g2_fill_1 FILLER_65_2403 ();
 sg13g2_fill_1 FILLER_65_2430 ();
 sg13g2_fill_2 FILLER_65_2483 ();
 sg13g2_fill_1 FILLER_65_2514 ();
 sg13g2_decap_8 FILLER_65_2534 ();
 sg13g2_decap_4 FILLER_65_2541 ();
 sg13g2_fill_1 FILLER_65_2545 ();
 sg13g2_fill_2 FILLER_65_2555 ();
 sg13g2_decap_8 FILLER_65_2620 ();
 sg13g2_decap_8 FILLER_65_2627 ();
 sg13g2_decap_8 FILLER_65_2634 ();
 sg13g2_decap_8 FILLER_65_2641 ();
 sg13g2_decap_8 FILLER_65_2648 ();
 sg13g2_decap_8 FILLER_65_2655 ();
 sg13g2_decap_8 FILLER_65_2662 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_fill_2 FILLER_66_21 ();
 sg13g2_fill_1 FILLER_66_23 ();
 sg13g2_fill_2 FILLER_66_38 ();
 sg13g2_decap_8 FILLER_66_44 ();
 sg13g2_fill_1 FILLER_66_89 ();
 sg13g2_fill_1 FILLER_66_121 ();
 sg13g2_fill_2 FILLER_66_127 ();
 sg13g2_fill_1 FILLER_66_129 ();
 sg13g2_fill_1 FILLER_66_156 ();
 sg13g2_fill_1 FILLER_66_167 ();
 sg13g2_decap_4 FILLER_66_194 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_decap_4 FILLER_66_204 ();
 sg13g2_decap_4 FILLER_66_218 ();
 sg13g2_fill_1 FILLER_66_222 ();
 sg13g2_fill_2 FILLER_66_229 ();
 sg13g2_fill_1 FILLER_66_236 ();
 sg13g2_fill_2 FILLER_66_242 ();
 sg13g2_fill_1 FILLER_66_252 ();
 sg13g2_fill_1 FILLER_66_258 ();
 sg13g2_fill_2 FILLER_66_299 ();
 sg13g2_decap_8 FILLER_66_306 ();
 sg13g2_fill_2 FILLER_66_313 ();
 sg13g2_fill_1 FILLER_66_315 ();
 sg13g2_decap_4 FILLER_66_320 ();
 sg13g2_fill_2 FILLER_66_324 ();
 sg13g2_fill_1 FILLER_66_330 ();
 sg13g2_fill_2 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_359 ();
 sg13g2_decap_8 FILLER_66_363 ();
 sg13g2_decap_4 FILLER_66_370 ();
 sg13g2_fill_2 FILLER_66_461 ();
 sg13g2_fill_1 FILLER_66_479 ();
 sg13g2_fill_2 FILLER_66_499 ();
 sg13g2_fill_2 FILLER_66_518 ();
 sg13g2_fill_1 FILLER_66_535 ();
 sg13g2_fill_1 FILLER_66_562 ();
 sg13g2_fill_2 FILLER_66_567 ();
 sg13g2_fill_1 FILLER_66_569 ();
 sg13g2_fill_2 FILLER_66_574 ();
 sg13g2_decap_4 FILLER_66_581 ();
 sg13g2_fill_2 FILLER_66_585 ();
 sg13g2_fill_2 FILLER_66_591 ();
 sg13g2_fill_2 FILLER_66_619 ();
 sg13g2_fill_2 FILLER_66_708 ();
 sg13g2_fill_1 FILLER_66_713 ();
 sg13g2_decap_8 FILLER_66_725 ();
 sg13g2_fill_2 FILLER_66_732 ();
 sg13g2_fill_1 FILLER_66_734 ();
 sg13g2_fill_2 FILLER_66_740 ();
 sg13g2_fill_2 FILLER_66_752 ();
 sg13g2_fill_1 FILLER_66_754 ();
 sg13g2_decap_4 FILLER_66_765 ();
 sg13g2_fill_2 FILLER_66_769 ();
 sg13g2_fill_2 FILLER_66_776 ();
 sg13g2_fill_1 FILLER_66_778 ();
 sg13g2_fill_2 FILLER_66_819 ();
 sg13g2_fill_1 FILLER_66_866 ();
 sg13g2_fill_2 FILLER_66_872 ();
 sg13g2_decap_4 FILLER_66_878 ();
 sg13g2_fill_1 FILLER_66_882 ();
 sg13g2_decap_4 FILLER_66_888 ();
 sg13g2_fill_1 FILLER_66_892 ();
 sg13g2_fill_1 FILLER_66_904 ();
 sg13g2_fill_1 FILLER_66_914 ();
 sg13g2_fill_2 FILLER_66_954 ();
 sg13g2_fill_2 FILLER_66_961 ();
 sg13g2_fill_1 FILLER_66_966 ();
 sg13g2_decap_8 FILLER_66_1010 ();
 sg13g2_decap_8 FILLER_66_1017 ();
 sg13g2_fill_2 FILLER_66_1060 ();
 sg13g2_fill_1 FILLER_66_1081 ();
 sg13g2_decap_8 FILLER_66_1121 ();
 sg13g2_decap_4 FILLER_66_1128 ();
 sg13g2_fill_1 FILLER_66_1132 ();
 sg13g2_decap_8 FILLER_66_1136 ();
 sg13g2_decap_8 FILLER_66_1143 ();
 sg13g2_decap_4 FILLER_66_1150 ();
 sg13g2_fill_1 FILLER_66_1154 ();
 sg13g2_fill_1 FILLER_66_1173 ();
 sg13g2_fill_1 FILLER_66_1217 ();
 sg13g2_fill_1 FILLER_66_1228 ();
 sg13g2_fill_2 FILLER_66_1253 ();
 sg13g2_fill_1 FILLER_66_1267 ();
 sg13g2_fill_1 FILLER_66_1276 ();
 sg13g2_decap_4 FILLER_66_1312 ();
 sg13g2_decap_4 FILLER_66_1324 ();
 sg13g2_decap_8 FILLER_66_1332 ();
 sg13g2_decap_4 FILLER_66_1339 ();
 sg13g2_decap_4 FILLER_66_1351 ();
 sg13g2_fill_2 FILLER_66_1368 ();
 sg13g2_fill_1 FILLER_66_1370 ();
 sg13g2_decap_8 FILLER_66_1383 ();
 sg13g2_decap_8 FILLER_66_1390 ();
 sg13g2_decap_8 FILLER_66_1397 ();
 sg13g2_fill_1 FILLER_66_1404 ();
 sg13g2_fill_2 FILLER_66_1410 ();
 sg13g2_fill_1 FILLER_66_1420 ();
 sg13g2_decap_8 FILLER_66_1437 ();
 sg13g2_decap_4 FILLER_66_1444 ();
 sg13g2_fill_2 FILLER_66_1448 ();
 sg13g2_decap_8 FILLER_66_1455 ();
 sg13g2_decap_8 FILLER_66_1479 ();
 sg13g2_fill_1 FILLER_66_1486 ();
 sg13g2_fill_1 FILLER_66_1491 ();
 sg13g2_fill_1 FILLER_66_1501 ();
 sg13g2_decap_4 FILLER_66_1521 ();
 sg13g2_fill_2 FILLER_66_1525 ();
 sg13g2_fill_1 FILLER_66_1551 ();
 sg13g2_fill_2 FILLER_66_1574 ();
 sg13g2_decap_8 FILLER_66_1584 ();
 sg13g2_decap_8 FILLER_66_1591 ();
 sg13g2_decap_8 FILLER_66_1598 ();
 sg13g2_decap_8 FILLER_66_1605 ();
 sg13g2_decap_4 FILLER_66_1612 ();
 sg13g2_fill_1 FILLER_66_1632 ();
 sg13g2_fill_2 FILLER_66_1638 ();
 sg13g2_fill_1 FILLER_66_1645 ();
 sg13g2_fill_2 FILLER_66_1651 ();
 sg13g2_fill_2 FILLER_66_1679 ();
 sg13g2_decap_4 FILLER_66_1690 ();
 sg13g2_fill_1 FILLER_66_1702 ();
 sg13g2_decap_4 FILLER_66_1709 ();
 sg13g2_fill_1 FILLER_66_1713 ();
 sg13g2_fill_2 FILLER_66_1719 ();
 sg13g2_fill_1 FILLER_66_1770 ();
 sg13g2_fill_1 FILLER_66_1777 ();
 sg13g2_fill_1 FILLER_66_1795 ();
 sg13g2_fill_2 FILLER_66_1854 ();
 sg13g2_fill_1 FILLER_66_1856 ();
 sg13g2_fill_1 FILLER_66_1890 ();
 sg13g2_fill_1 FILLER_66_1975 ();
 sg13g2_fill_2 FILLER_66_1982 ();
 sg13g2_decap_8 FILLER_66_1988 ();
 sg13g2_fill_2 FILLER_66_1995 ();
 sg13g2_fill_1 FILLER_66_1997 ();
 sg13g2_fill_1 FILLER_66_2035 ();
 sg13g2_fill_2 FILLER_66_2041 ();
 sg13g2_fill_2 FILLER_66_2069 ();
 sg13g2_fill_2 FILLER_66_2075 ();
 sg13g2_fill_1 FILLER_66_2077 ();
 sg13g2_fill_2 FILLER_66_2104 ();
 sg13g2_fill_2 FILLER_66_2116 ();
 sg13g2_fill_1 FILLER_66_2118 ();
 sg13g2_fill_2 FILLER_66_2123 ();
 sg13g2_fill_1 FILLER_66_2129 ();
 sg13g2_fill_1 FILLER_66_2135 ();
 sg13g2_fill_2 FILLER_66_2175 ();
 sg13g2_fill_1 FILLER_66_2177 ();
 sg13g2_decap_8 FILLER_66_2244 ();
 sg13g2_decap_8 FILLER_66_2251 ();
 sg13g2_decap_4 FILLER_66_2258 ();
 sg13g2_fill_2 FILLER_66_2262 ();
 sg13g2_decap_8 FILLER_66_2301 ();
 sg13g2_decap_4 FILLER_66_2308 ();
 sg13g2_fill_1 FILLER_66_2312 ();
 sg13g2_decap_8 FILLER_66_2352 ();
 sg13g2_fill_2 FILLER_66_2359 ();
 sg13g2_fill_1 FILLER_66_2361 ();
 sg13g2_decap_8 FILLER_66_2366 ();
 sg13g2_decap_8 FILLER_66_2373 ();
 sg13g2_fill_1 FILLER_66_2380 ();
 sg13g2_fill_1 FILLER_66_2490 ();
 sg13g2_fill_2 FILLER_66_2501 ();
 sg13g2_fill_2 FILLER_66_2507 ();
 sg13g2_decap_4 FILLER_66_2523 ();
 sg13g2_decap_8 FILLER_66_2533 ();
 sg13g2_decap_4 FILLER_66_2540 ();
 sg13g2_fill_2 FILLER_66_2544 ();
 sg13g2_fill_1 FILLER_66_2584 ();
 sg13g2_fill_2 FILLER_66_2589 ();
 sg13g2_decap_8 FILLER_66_2621 ();
 sg13g2_decap_8 FILLER_66_2628 ();
 sg13g2_decap_8 FILLER_66_2635 ();
 sg13g2_decap_8 FILLER_66_2642 ();
 sg13g2_decap_8 FILLER_66_2649 ();
 sg13g2_decap_8 FILLER_66_2656 ();
 sg13g2_decap_8 FILLER_66_2663 ();
 sg13g2_fill_2 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_33 ();
 sg13g2_fill_1 FILLER_67_42 ();
 sg13g2_fill_2 FILLER_67_73 ();
 sg13g2_fill_1 FILLER_67_75 ();
 sg13g2_fill_1 FILLER_67_86 ();
 sg13g2_decap_8 FILLER_67_128 ();
 sg13g2_decap_8 FILLER_67_139 ();
 sg13g2_decap_4 FILLER_67_146 ();
 sg13g2_fill_1 FILLER_67_154 ();
 sg13g2_fill_1 FILLER_67_160 ();
 sg13g2_fill_1 FILLER_67_175 ();
 sg13g2_fill_1 FILLER_67_181 ();
 sg13g2_decap_4 FILLER_67_186 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_fill_2 FILLER_67_214 ();
 sg13g2_fill_1 FILLER_67_221 ();
 sg13g2_fill_2 FILLER_67_227 ();
 sg13g2_fill_1 FILLER_67_255 ();
 sg13g2_fill_1 FILLER_67_265 ();
 sg13g2_fill_2 FILLER_67_271 ();
 sg13g2_fill_2 FILLER_67_278 ();
 sg13g2_fill_1 FILLER_67_288 ();
 sg13g2_decap_8 FILLER_67_293 ();
 sg13g2_fill_2 FILLER_67_310 ();
 sg13g2_fill_1 FILLER_67_312 ();
 sg13g2_fill_2 FILLER_67_322 ();
 sg13g2_fill_2 FILLER_67_333 ();
 sg13g2_fill_2 FILLER_67_342 ();
 sg13g2_fill_1 FILLER_67_344 ();
 sg13g2_decap_4 FILLER_67_353 ();
 sg13g2_fill_2 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_398 ();
 sg13g2_fill_2 FILLER_67_452 ();
 sg13g2_fill_1 FILLER_67_465 ();
 sg13g2_fill_2 FILLER_67_471 ();
 sg13g2_fill_2 FILLER_67_478 ();
 sg13g2_fill_2 FILLER_67_535 ();
 sg13g2_fill_2 FILLER_67_551 ();
 sg13g2_fill_1 FILLER_67_579 ();
 sg13g2_fill_1 FILLER_67_601 ();
 sg13g2_fill_1 FILLER_67_626 ();
 sg13g2_fill_2 FILLER_67_650 ();
 sg13g2_fill_2 FILLER_67_668 ();
 sg13g2_fill_1 FILLER_67_678 ();
 sg13g2_fill_1 FILLER_67_692 ();
 sg13g2_fill_2 FILLER_67_698 ();
 sg13g2_fill_1 FILLER_67_717 ();
 sg13g2_fill_2 FILLER_67_744 ();
 sg13g2_fill_1 FILLER_67_746 ();
 sg13g2_fill_2 FILLER_67_777 ();
 sg13g2_fill_1 FILLER_67_779 ();
 sg13g2_decap_4 FILLER_67_784 ();
 sg13g2_fill_1 FILLER_67_788 ();
 sg13g2_decap_4 FILLER_67_799 ();
 sg13g2_fill_1 FILLER_67_803 ();
 sg13g2_decap_4 FILLER_67_814 ();
 sg13g2_fill_1 FILLER_67_818 ();
 sg13g2_fill_2 FILLER_67_823 ();
 sg13g2_fill_1 FILLER_67_825 ();
 sg13g2_decap_8 FILLER_67_831 ();
 sg13g2_fill_2 FILLER_67_838 ();
 sg13g2_fill_1 FILLER_67_840 ();
 sg13g2_decap_4 FILLER_67_849 ();
 sg13g2_fill_1 FILLER_67_853 ();
 sg13g2_fill_1 FILLER_67_867 ();
 sg13g2_fill_2 FILLER_67_872 ();
 sg13g2_decap_4 FILLER_67_883 ();
 sg13g2_fill_1 FILLER_67_887 ();
 sg13g2_fill_1 FILLER_67_893 ();
 sg13g2_decap_4 FILLER_67_897 ();
 sg13g2_fill_2 FILLER_67_901 ();
 sg13g2_fill_1 FILLER_67_912 ();
 sg13g2_fill_2 FILLER_67_971 ();
 sg13g2_decap_8 FILLER_67_1012 ();
 sg13g2_fill_2 FILLER_67_1019 ();
 sg13g2_fill_1 FILLER_67_1021 ();
 sg13g2_fill_1 FILLER_67_1089 ();
 sg13g2_fill_2 FILLER_67_1096 ();
 sg13g2_fill_1 FILLER_67_1154 ();
 sg13g2_decap_8 FILLER_67_1168 ();
 sg13g2_fill_1 FILLER_67_1175 ();
 sg13g2_fill_1 FILLER_67_1189 ();
 sg13g2_fill_1 FILLER_67_1224 ();
 sg13g2_fill_2 FILLER_67_1247 ();
 sg13g2_fill_2 FILLER_67_1253 ();
 sg13g2_fill_2 FILLER_67_1260 ();
 sg13g2_decap_8 FILLER_67_1266 ();
 sg13g2_fill_2 FILLER_67_1273 ();
 sg13g2_fill_1 FILLER_67_1275 ();
 sg13g2_decap_4 FILLER_67_1284 ();
 sg13g2_decap_8 FILLER_67_1305 ();
 sg13g2_decap_8 FILLER_67_1312 ();
 sg13g2_decap_8 FILLER_67_1319 ();
 sg13g2_decap_4 FILLER_67_1326 ();
 sg13g2_fill_2 FILLER_67_1369 ();
 sg13g2_decap_4 FILLER_67_1385 ();
 sg13g2_decap_8 FILLER_67_1399 ();
 sg13g2_decap_8 FILLER_67_1406 ();
 sg13g2_decap_8 FILLER_67_1417 ();
 sg13g2_decap_8 FILLER_67_1424 ();
 sg13g2_decap_8 FILLER_67_1431 ();
 sg13g2_fill_1 FILLER_67_1438 ();
 sg13g2_fill_1 FILLER_67_1458 ();
 sg13g2_fill_2 FILLER_67_1464 ();
 sg13g2_decap_8 FILLER_67_1471 ();
 sg13g2_decap_8 FILLER_67_1478 ();
 sg13g2_fill_2 FILLER_67_1498 ();
 sg13g2_fill_2 FILLER_67_1505 ();
 sg13g2_fill_1 FILLER_67_1507 ();
 sg13g2_fill_2 FILLER_67_1512 ();
 sg13g2_fill_1 FILLER_67_1514 ();
 sg13g2_fill_1 FILLER_67_1519 ();
 sg13g2_fill_1 FILLER_67_1525 ();
 sg13g2_fill_1 FILLER_67_1537 ();
 sg13g2_fill_2 FILLER_67_1554 ();
 sg13g2_fill_1 FILLER_67_1556 ();
 sg13g2_fill_1 FILLER_67_1567 ();
 sg13g2_fill_1 FILLER_67_1573 ();
 sg13g2_fill_2 FILLER_67_1579 ();
 sg13g2_fill_2 FILLER_67_1592 ();
 sg13g2_decap_4 FILLER_67_1608 ();
 sg13g2_decap_4 FILLER_67_1640 ();
 sg13g2_fill_1 FILLER_67_1644 ();
 sg13g2_fill_2 FILLER_67_1649 ();
 sg13g2_fill_2 FILLER_67_1660 ();
 sg13g2_decap_8 FILLER_67_1683 ();
 sg13g2_decap_8 FILLER_67_1690 ();
 sg13g2_decap_8 FILLER_67_1697 ();
 sg13g2_decap_4 FILLER_67_1709 ();
 sg13g2_fill_1 FILLER_67_1713 ();
 sg13g2_fill_1 FILLER_67_1734 ();
 sg13g2_fill_1 FILLER_67_1740 ();
 sg13g2_fill_2 FILLER_67_1745 ();
 sg13g2_fill_1 FILLER_67_1752 ();
 sg13g2_fill_2 FILLER_67_1762 ();
 sg13g2_decap_4 FILLER_67_1782 ();
 sg13g2_fill_1 FILLER_67_1796 ();
 sg13g2_fill_1 FILLER_67_1802 ();
 sg13g2_fill_1 FILLER_67_1850 ();
 sg13g2_decap_4 FILLER_67_1856 ();
 sg13g2_fill_2 FILLER_67_1860 ();
 sg13g2_decap_4 FILLER_67_1869 ();
 sg13g2_fill_2 FILLER_67_1877 ();
 sg13g2_fill_1 FILLER_67_1879 ();
 sg13g2_decap_8 FILLER_67_1885 ();
 sg13g2_decap_8 FILLER_67_1892 ();
 sg13g2_fill_1 FILLER_67_1899 ();
 sg13g2_decap_8 FILLER_67_1935 ();
 sg13g2_decap_8 FILLER_67_1942 ();
 sg13g2_decap_4 FILLER_67_1949 ();
 sg13g2_fill_1 FILLER_67_1988 ();
 sg13g2_fill_2 FILLER_67_1994 ();
 sg13g2_fill_1 FILLER_67_1996 ();
 sg13g2_fill_1 FILLER_67_2105 ();
 sg13g2_fill_1 FILLER_67_2139 ();
 sg13g2_fill_2 FILLER_67_2181 ();
 sg13g2_fill_1 FILLER_67_2183 ();
 sg13g2_fill_1 FILLER_67_2195 ();
 sg13g2_fill_2 FILLER_67_2226 ();
 sg13g2_fill_2 FILLER_67_2266 ();
 sg13g2_fill_1 FILLER_67_2304 ();
 sg13g2_fill_1 FILLER_67_2309 ();
 sg13g2_decap_8 FILLER_67_2314 ();
 sg13g2_decap_4 FILLER_67_2321 ();
 sg13g2_fill_1 FILLER_67_2325 ();
 sg13g2_decap_8 FILLER_67_2330 ();
 sg13g2_fill_1 FILLER_67_2363 ();
 sg13g2_decap_8 FILLER_67_2369 ();
 sg13g2_decap_8 FILLER_67_2376 ();
 sg13g2_fill_2 FILLER_67_2383 ();
 sg13g2_fill_1 FILLER_67_2395 ();
 sg13g2_fill_2 FILLER_67_2422 ();
 sg13g2_fill_1 FILLER_67_2424 ();
 sg13g2_fill_1 FILLER_67_2443 ();
 sg13g2_fill_2 FILLER_67_2450 ();
 sg13g2_decap_8 FILLER_67_2463 ();
 sg13g2_decap_8 FILLER_67_2470 ();
 sg13g2_fill_1 FILLER_67_2477 ();
 sg13g2_fill_1 FILLER_67_2484 ();
 sg13g2_fill_1 FILLER_67_2490 ();
 sg13g2_decap_4 FILLER_67_2530 ();
 sg13g2_fill_2 FILLER_67_2534 ();
 sg13g2_fill_1 FILLER_67_2576 ();
 sg13g2_decap_8 FILLER_67_2626 ();
 sg13g2_decap_8 FILLER_67_2633 ();
 sg13g2_decap_8 FILLER_67_2640 ();
 sg13g2_decap_8 FILLER_67_2647 ();
 sg13g2_decap_8 FILLER_67_2654 ();
 sg13g2_decap_8 FILLER_67_2661 ();
 sg13g2_fill_2 FILLER_67_2668 ();
 sg13g2_fill_1 FILLER_68_0 ();
 sg13g2_fill_1 FILLER_68_27 ();
 sg13g2_fill_1 FILLER_68_54 ();
 sg13g2_fill_2 FILLER_68_81 ();
 sg13g2_fill_1 FILLER_68_93 ();
 sg13g2_fill_1 FILLER_68_125 ();
 sg13g2_decap_8 FILLER_68_134 ();
 sg13g2_decap_4 FILLER_68_141 ();
 sg13g2_fill_2 FILLER_68_151 ();
 sg13g2_fill_1 FILLER_68_153 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_4 FILLER_68_166 ();
 sg13g2_fill_1 FILLER_68_170 ();
 sg13g2_decap_4 FILLER_68_175 ();
 sg13g2_fill_1 FILLER_68_211 ();
 sg13g2_fill_1 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_272 ();
 sg13g2_fill_2 FILLER_68_289 ();
 sg13g2_fill_2 FILLER_68_312 ();
 sg13g2_fill_2 FILLER_68_319 ();
 sg13g2_fill_1 FILLER_68_321 ();
 sg13g2_fill_2 FILLER_68_336 ();
 sg13g2_fill_1 FILLER_68_338 ();
 sg13g2_decap_4 FILLER_68_361 ();
 sg13g2_fill_2 FILLER_68_365 ();
 sg13g2_decap_8 FILLER_68_383 ();
 sg13g2_decap_4 FILLER_68_390 ();
 sg13g2_fill_2 FILLER_68_405 ();
 sg13g2_fill_1 FILLER_68_467 ();
 sg13g2_fill_1 FILLER_68_472 ();
 sg13g2_fill_1 FILLER_68_490 ();
 sg13g2_fill_1 FILLER_68_504 ();
 sg13g2_decap_8 FILLER_68_564 ();
 sg13g2_decap_4 FILLER_68_571 ();
 sg13g2_fill_2 FILLER_68_575 ();
 sg13g2_fill_2 FILLER_68_635 ();
 sg13g2_fill_2 FILLER_68_657 ();
 sg13g2_fill_2 FILLER_68_684 ();
 sg13g2_fill_2 FILLER_68_690 ();
 sg13g2_fill_1 FILLER_68_699 ();
 sg13g2_fill_1 FILLER_68_706 ();
 sg13g2_fill_2 FILLER_68_756 ();
 sg13g2_decap_8 FILLER_68_805 ();
 sg13g2_decap_4 FILLER_68_812 ();
 sg13g2_fill_1 FILLER_68_816 ();
 sg13g2_fill_1 FILLER_68_840 ();
 sg13g2_decap_4 FILLER_68_855 ();
 sg13g2_fill_1 FILLER_68_859 ();
 sg13g2_fill_1 FILLER_68_865 ();
 sg13g2_fill_1 FILLER_68_871 ();
 sg13g2_fill_1 FILLER_68_903 ();
 sg13g2_fill_1 FILLER_68_942 ();
 sg13g2_decap_8 FILLER_68_1023 ();
 sg13g2_fill_2 FILLER_68_1030 ();
 sg13g2_decap_4 FILLER_68_1050 ();
 sg13g2_fill_1 FILLER_68_1054 ();
 sg13g2_fill_2 FILLER_68_1176 ();
 sg13g2_fill_1 FILLER_68_1203 ();
 sg13g2_fill_2 FILLER_68_1212 ();
 sg13g2_fill_2 FILLER_68_1233 ();
 sg13g2_fill_2 FILLER_68_1255 ();
 sg13g2_fill_1 FILLER_68_1257 ();
 sg13g2_fill_2 FILLER_68_1262 ();
 sg13g2_fill_2 FILLER_68_1272 ();
 sg13g2_fill_1 FILLER_68_1274 ();
 sg13g2_decap_8 FILLER_68_1280 ();
 sg13g2_decap_8 FILLER_68_1287 ();
 sg13g2_decap_8 FILLER_68_1294 ();
 sg13g2_fill_2 FILLER_68_1301 ();
 sg13g2_fill_1 FILLER_68_1303 ();
 sg13g2_decap_8 FILLER_68_1308 ();
 sg13g2_fill_2 FILLER_68_1315 ();
 sg13g2_fill_1 FILLER_68_1317 ();
 sg13g2_fill_2 FILLER_68_1339 ();
 sg13g2_decap_4 FILLER_68_1346 ();
 sg13g2_decap_8 FILLER_68_1366 ();
 sg13g2_fill_2 FILLER_68_1373 ();
 sg13g2_decap_8 FILLER_68_1379 ();
 sg13g2_fill_2 FILLER_68_1386 ();
 sg13g2_fill_1 FILLER_68_1388 ();
 sg13g2_decap_8 FILLER_68_1393 ();
 sg13g2_decap_8 FILLER_68_1400 ();
 sg13g2_decap_4 FILLER_68_1407 ();
 sg13g2_fill_2 FILLER_68_1411 ();
 sg13g2_decap_8 FILLER_68_1422 ();
 sg13g2_fill_2 FILLER_68_1429 ();
 sg13g2_fill_1 FILLER_68_1431 ();
 sg13g2_decap_4 FILLER_68_1455 ();
 sg13g2_fill_2 FILLER_68_1463 ();
 sg13g2_fill_2 FILLER_68_1473 ();
 sg13g2_fill_1 FILLER_68_1475 ();
 sg13g2_fill_2 FILLER_68_1481 ();
 sg13g2_fill_2 FILLER_68_1493 ();
 sg13g2_fill_2 FILLER_68_1508 ();
 sg13g2_fill_1 FILLER_68_1510 ();
 sg13g2_fill_2 FILLER_68_1519 ();
 sg13g2_fill_1 FILLER_68_1546 ();
 sg13g2_fill_2 FILLER_68_1590 ();
 sg13g2_fill_2 FILLER_68_1598 ();
 sg13g2_fill_1 FILLER_68_1608 ();
 sg13g2_fill_1 FILLER_68_1625 ();
 sg13g2_fill_1 FILLER_68_1634 ();
 sg13g2_decap_4 FILLER_68_1654 ();
 sg13g2_decap_8 FILLER_68_1663 ();
 sg13g2_fill_1 FILLER_68_1670 ();
 sg13g2_decap_8 FILLER_68_1689 ();
 sg13g2_decap_8 FILLER_68_1699 ();
 sg13g2_fill_1 FILLER_68_1706 ();
 sg13g2_fill_2 FILLER_68_1716 ();
 sg13g2_fill_1 FILLER_68_1747 ();
 sg13g2_fill_1 FILLER_68_1760 ();
 sg13g2_fill_1 FILLER_68_1772 ();
 sg13g2_fill_1 FILLER_68_1799 ();
 sg13g2_fill_1 FILLER_68_1847 ();
 sg13g2_fill_2 FILLER_68_1855 ();
 sg13g2_decap_8 FILLER_68_1890 ();
 sg13g2_decap_8 FILLER_68_1897 ();
 sg13g2_fill_2 FILLER_68_1918 ();
 sg13g2_decap_8 FILLER_68_1925 ();
 sg13g2_decap_4 FILLER_68_1942 ();
 sg13g2_fill_1 FILLER_68_1946 ();
 sg13g2_decap_8 FILLER_68_1993 ();
 sg13g2_decap_4 FILLER_68_2000 ();
 sg13g2_fill_1 FILLER_68_2004 ();
 sg13g2_fill_2 FILLER_68_2009 ();
 sg13g2_fill_2 FILLER_68_2015 ();
 sg13g2_fill_1 FILLER_68_2017 ();
 sg13g2_fill_2 FILLER_68_2100 ();
 sg13g2_decap_4 FILLER_68_2108 ();
 sg13g2_fill_1 FILLER_68_2112 ();
 sg13g2_decap_8 FILLER_68_2122 ();
 sg13g2_fill_2 FILLER_68_2134 ();
 sg13g2_fill_1 FILLER_68_2136 ();
 sg13g2_fill_1 FILLER_68_2145 ();
 sg13g2_fill_1 FILLER_68_2199 ();
 sg13g2_fill_1 FILLER_68_2216 ();
 sg13g2_fill_2 FILLER_68_2235 ();
 sg13g2_decap_8 FILLER_68_2317 ();
 sg13g2_decap_8 FILLER_68_2324 ();
 sg13g2_decap_4 FILLER_68_2331 ();
 sg13g2_fill_1 FILLER_68_2335 ();
 sg13g2_fill_2 FILLER_68_2340 ();
 sg13g2_fill_1 FILLER_68_2342 ();
 sg13g2_decap_8 FILLER_68_2369 ();
 sg13g2_fill_1 FILLER_68_2376 ();
 sg13g2_decap_4 FILLER_68_2403 ();
 sg13g2_fill_2 FILLER_68_2407 ();
 sg13g2_fill_1 FILLER_68_2492 ();
 sg13g2_fill_1 FILLER_68_2500 ();
 sg13g2_fill_1 FILLER_68_2507 ();
 sg13g2_fill_2 FILLER_68_2525 ();
 sg13g2_fill_1 FILLER_68_2527 ();
 sg13g2_fill_2 FILLER_68_2570 ();
 sg13g2_fill_2 FILLER_68_2614 ();
 sg13g2_decap_8 FILLER_68_2642 ();
 sg13g2_decap_8 FILLER_68_2649 ();
 sg13g2_decap_8 FILLER_68_2656 ();
 sg13g2_decap_8 FILLER_68_2663 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_fill_1 FILLER_69_11 ();
 sg13g2_fill_1 FILLER_69_16 ();
 sg13g2_fill_1 FILLER_69_27 ();
 sg13g2_fill_1 FILLER_69_42 ();
 sg13g2_fill_2 FILLER_69_47 ();
 sg13g2_fill_1 FILLER_69_49 ();
 sg13g2_fill_2 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_72 ();
 sg13g2_fill_2 FILLER_69_96 ();
 sg13g2_fill_1 FILLER_69_98 ();
 sg13g2_fill_2 FILLER_69_103 ();
 sg13g2_fill_2 FILLER_69_113 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_decap_8 FILLER_69_124 ();
 sg13g2_fill_2 FILLER_69_131 ();
 sg13g2_decap_8 FILLER_69_173 ();
 sg13g2_decap_8 FILLER_69_180 ();
 sg13g2_decap_8 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_212 ();
 sg13g2_fill_1 FILLER_69_238 ();
 sg13g2_fill_1 FILLER_69_247 ();
 sg13g2_fill_2 FILLER_69_254 ();
 sg13g2_fill_2 FILLER_69_261 ();
 sg13g2_fill_2 FILLER_69_280 ();
 sg13g2_fill_1 FILLER_69_282 ();
 sg13g2_decap_4 FILLER_69_315 ();
 sg13g2_fill_2 FILLER_69_319 ();
 sg13g2_decap_4 FILLER_69_326 ();
 sg13g2_fill_1 FILLER_69_330 ();
 sg13g2_fill_2 FILLER_69_337 ();
 sg13g2_fill_1 FILLER_69_339 ();
 sg13g2_fill_2 FILLER_69_434 ();
 sg13g2_fill_1 FILLER_69_436 ();
 sg13g2_decap_8 FILLER_69_563 ();
 sg13g2_fill_2 FILLER_69_570 ();
 sg13g2_fill_1 FILLER_69_572 ();
 sg13g2_decap_4 FILLER_69_577 ();
 sg13g2_fill_1 FILLER_69_581 ();
 sg13g2_fill_2 FILLER_69_608 ();
 sg13g2_fill_2 FILLER_69_625 ();
 sg13g2_fill_1 FILLER_69_660 ();
 sg13g2_fill_1 FILLER_69_700 ();
 sg13g2_decap_8 FILLER_69_708 ();
 sg13g2_decap_4 FILLER_69_719 ();
 sg13g2_fill_2 FILLER_69_723 ();
 sg13g2_decap_4 FILLER_69_735 ();
 sg13g2_fill_2 FILLER_69_739 ();
 sg13g2_fill_2 FILLER_69_754 ();
 sg13g2_fill_2 FILLER_69_766 ();
 sg13g2_fill_2 FILLER_69_776 ();
 sg13g2_decap_4 FILLER_69_788 ();
 sg13g2_fill_2 FILLER_69_797 ();
 sg13g2_decap_4 FILLER_69_807 ();
 sg13g2_decap_4 FILLER_69_841 ();
 sg13g2_decap_4 FILLER_69_868 ();
 sg13g2_decap_4 FILLER_69_898 ();
 sg13g2_fill_2 FILLER_69_902 ();
 sg13g2_fill_1 FILLER_69_913 ();
 sg13g2_fill_1 FILLER_69_928 ();
 sg13g2_fill_1 FILLER_69_937 ();
 sg13g2_fill_2 FILLER_69_989 ();
 sg13g2_decap_8 FILLER_69_1033 ();
 sg13g2_decap_8 FILLER_69_1040 ();
 sg13g2_fill_2 FILLER_69_1047 ();
 sg13g2_fill_2 FILLER_69_1057 ();
 sg13g2_decap_4 FILLER_69_1095 ();
 sg13g2_decap_8 FILLER_69_1149 ();
 sg13g2_fill_1 FILLER_69_1156 ();
 sg13g2_decap_8 FILLER_69_1161 ();
 sg13g2_decap_4 FILLER_69_1168 ();
 sg13g2_fill_2 FILLER_69_1191 ();
 sg13g2_fill_1 FILLER_69_1233 ();
 sg13g2_fill_2 FILLER_69_1248 ();
 sg13g2_fill_1 FILLER_69_1255 ();
 sg13g2_fill_2 FILLER_69_1260 ();
 sg13g2_fill_1 FILLER_69_1262 ();
 sg13g2_fill_2 FILLER_69_1267 ();
 sg13g2_fill_1 FILLER_69_1269 ();
 sg13g2_decap_4 FILLER_69_1275 ();
 sg13g2_fill_2 FILLER_69_1284 ();
 sg13g2_fill_1 FILLER_69_1286 ();
 sg13g2_decap_8 FILLER_69_1295 ();
 sg13g2_decap_8 FILLER_69_1306 ();
 sg13g2_fill_1 FILLER_69_1317 ();
 sg13g2_fill_1 FILLER_69_1323 ();
 sg13g2_fill_1 FILLER_69_1330 ();
 sg13g2_fill_1 FILLER_69_1336 ();
 sg13g2_fill_1 FILLER_69_1342 ();
 sg13g2_fill_1 FILLER_69_1348 ();
 sg13g2_decap_4 FILLER_69_1368 ();
 sg13g2_fill_1 FILLER_69_1372 ();
 sg13g2_fill_2 FILLER_69_1404 ();
 sg13g2_fill_2 FILLER_69_1411 ();
 sg13g2_fill_1 FILLER_69_1413 ();
 sg13g2_fill_1 FILLER_69_1418 ();
 sg13g2_fill_1 FILLER_69_1423 ();
 sg13g2_fill_1 FILLER_69_1434 ();
 sg13g2_fill_1 FILLER_69_1439 ();
 sg13g2_fill_1 FILLER_69_1445 ();
 sg13g2_fill_1 FILLER_69_1452 ();
 sg13g2_decap_8 FILLER_69_1458 ();
 sg13g2_fill_1 FILLER_69_1493 ();
 sg13g2_fill_2 FILLER_69_1509 ();
 sg13g2_fill_1 FILLER_69_1524 ();
 sg13g2_fill_2 FILLER_69_1533 ();
 sg13g2_fill_1 FILLER_69_1535 ();
 sg13g2_decap_4 FILLER_69_1540 ();
 sg13g2_decap_4 FILLER_69_1551 ();
 sg13g2_fill_1 FILLER_69_1559 ();
 sg13g2_fill_1 FILLER_69_1566 ();
 sg13g2_decap_8 FILLER_69_1583 ();
 sg13g2_fill_1 FILLER_69_1595 ();
 sg13g2_fill_2 FILLER_69_1608 ();
 sg13g2_fill_2 FILLER_69_1615 ();
 sg13g2_fill_1 FILLER_69_1629 ();
 sg13g2_fill_1 FILLER_69_1659 ();
 sg13g2_fill_1 FILLER_69_1669 ();
 sg13g2_decap_8 FILLER_69_1682 ();
 sg13g2_decap_4 FILLER_69_1695 ();
 sg13g2_fill_2 FILLER_69_1699 ();
 sg13g2_fill_1 FILLER_69_1708 ();
 sg13g2_fill_2 FILLER_69_1719 ();
 sg13g2_decap_8 FILLER_69_1725 ();
 sg13g2_decap_8 FILLER_69_1732 ();
 sg13g2_fill_2 FILLER_69_1749 ();
 sg13g2_fill_1 FILLER_69_1757 ();
 sg13g2_fill_1 FILLER_69_1779 ();
 sg13g2_fill_1 FILLER_69_1813 ();
 sg13g2_fill_1 FILLER_69_1833 ();
 sg13g2_decap_8 FILLER_69_1847 ();
 sg13g2_decap_4 FILLER_69_1854 ();
 sg13g2_fill_1 FILLER_69_1858 ();
 sg13g2_fill_2 FILLER_69_1889 ();
 sg13g2_decap_4 FILLER_69_1895 ();
 sg13g2_decap_8 FILLER_69_1929 ();
 sg13g2_fill_1 FILLER_69_1951 ();
 sg13g2_decap_8 FILLER_69_1958 ();
 sg13g2_fill_2 FILLER_69_1965 ();
 sg13g2_decap_8 FILLER_69_1971 ();
 sg13g2_fill_2 FILLER_69_2027 ();
 sg13g2_decap_4 FILLER_69_2055 ();
 sg13g2_decap_4 FILLER_69_2083 ();
 sg13g2_fill_1 FILLER_69_2087 ();
 sg13g2_fill_2 FILLER_69_2092 ();
 sg13g2_fill_1 FILLER_69_2094 ();
 sg13g2_fill_1 FILLER_69_2111 ();
 sg13g2_fill_2 FILLER_69_2135 ();
 sg13g2_fill_1 FILLER_69_2142 ();
 sg13g2_fill_1 FILLER_69_2153 ();
 sg13g2_fill_2 FILLER_69_2161 ();
 sg13g2_fill_2 FILLER_69_2175 ();
 sg13g2_fill_1 FILLER_69_2227 ();
 sg13g2_fill_2 FILLER_69_2254 ();
 sg13g2_decap_4 FILLER_69_2266 ();
 sg13g2_fill_1 FILLER_69_2270 ();
 sg13g2_decap_8 FILLER_69_2307 ();
 sg13g2_decap_4 FILLER_69_2314 ();
 sg13g2_fill_2 FILLER_69_2354 ();
 sg13g2_fill_1 FILLER_69_2356 ();
 sg13g2_decap_8 FILLER_69_2393 ();
 sg13g2_fill_2 FILLER_69_2400 ();
 sg13g2_fill_1 FILLER_69_2402 ();
 sg13g2_fill_2 FILLER_69_2413 ();
 sg13g2_fill_1 FILLER_69_2415 ();
 sg13g2_fill_1 FILLER_69_2446 ();
 sg13g2_fill_1 FILLER_69_2487 ();
 sg13g2_fill_2 FILLER_69_2522 ();
 sg13g2_fill_2 FILLER_69_2530 ();
 sg13g2_fill_1 FILLER_69_2546 ();
 sg13g2_decap_8 FILLER_69_2627 ();
 sg13g2_decap_8 FILLER_69_2634 ();
 sg13g2_decap_8 FILLER_69_2641 ();
 sg13g2_decap_8 FILLER_69_2648 ();
 sg13g2_decap_8 FILLER_69_2655 ();
 sg13g2_decap_8 FILLER_69_2662 ();
 sg13g2_fill_1 FILLER_69_2669 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_4 FILLER_70_7 ();
 sg13g2_fill_2 FILLER_70_11 ();
 sg13g2_decap_8 FILLER_70_17 ();
 sg13g2_decap_8 FILLER_70_24 ();
 sg13g2_fill_1 FILLER_70_31 ();
 sg13g2_fill_1 FILLER_70_72 ();
 sg13g2_fill_1 FILLER_70_104 ();
 sg13g2_decap_8 FILLER_70_113 ();
 sg13g2_fill_2 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_fill_2 FILLER_70_128 ();
 sg13g2_fill_1 FILLER_70_130 ();
 sg13g2_fill_2 FILLER_70_176 ();
 sg13g2_fill_1 FILLER_70_178 ();
 sg13g2_fill_2 FILLER_70_184 ();
 sg13g2_fill_2 FILLER_70_215 ();
 sg13g2_fill_1 FILLER_70_217 ();
 sg13g2_fill_2 FILLER_70_256 ();
 sg13g2_fill_1 FILLER_70_268 ();
 sg13g2_fill_1 FILLER_70_283 ();
 sg13g2_fill_2 FILLER_70_290 ();
 sg13g2_fill_2 FILLER_70_297 ();
 sg13g2_fill_2 FILLER_70_304 ();
 sg13g2_decap_8 FILLER_70_312 ();
 sg13g2_fill_2 FILLER_70_319 ();
 sg13g2_decap_4 FILLER_70_341 ();
 sg13g2_fill_1 FILLER_70_345 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_fill_1 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_362 ();
 sg13g2_decap_8 FILLER_70_369 ();
 sg13g2_fill_1 FILLER_70_376 ();
 sg13g2_decap_8 FILLER_70_381 ();
 sg13g2_decap_4 FILLER_70_388 ();
 sg13g2_fill_1 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_fill_2 FILLER_70_404 ();
 sg13g2_fill_2 FILLER_70_410 ();
 sg13g2_fill_1 FILLER_70_412 ();
 sg13g2_fill_2 FILLER_70_439 ();
 sg13g2_decap_8 FILLER_70_454 ();
 sg13g2_decap_4 FILLER_70_461 ();
 sg13g2_fill_1 FILLER_70_465 ();
 sg13g2_decap_4 FILLER_70_470 ();
 sg13g2_decap_8 FILLER_70_478 ();
 sg13g2_decap_8 FILLER_70_485 ();
 sg13g2_decap_4 FILLER_70_492 ();
 sg13g2_fill_2 FILLER_70_496 ();
 sg13g2_fill_1 FILLER_70_502 ();
 sg13g2_decap_4 FILLER_70_510 ();
 sg13g2_fill_2 FILLER_70_514 ();
 sg13g2_fill_2 FILLER_70_529 ();
 sg13g2_fill_1 FILLER_70_531 ();
 sg13g2_decap_8 FILLER_70_558 ();
 sg13g2_decap_8 FILLER_70_565 ();
 sg13g2_decap_8 FILLER_70_572 ();
 sg13g2_decap_8 FILLER_70_579 ();
 sg13g2_decap_4 FILLER_70_586 ();
 sg13g2_decap_4 FILLER_70_598 ();
 sg13g2_fill_2 FILLER_70_641 ();
 sg13g2_fill_2 FILLER_70_652 ();
 sg13g2_fill_1 FILLER_70_669 ();
 sg13g2_decap_8 FILLER_70_683 ();
 sg13g2_fill_2 FILLER_70_690 ();
 sg13g2_decap_8 FILLER_70_726 ();
 sg13g2_fill_2 FILLER_70_733 ();
 sg13g2_fill_1 FILLER_70_735 ();
 sg13g2_decap_8 FILLER_70_764 ();
 sg13g2_decap_8 FILLER_70_771 ();
 sg13g2_fill_2 FILLER_70_778 ();
 sg13g2_fill_1 FILLER_70_780 ();
 sg13g2_fill_2 FILLER_70_833 ();
 sg13g2_fill_1 FILLER_70_835 ();
 sg13g2_fill_1 FILLER_70_846 ();
 sg13g2_fill_2 FILLER_70_882 ();
 sg13g2_fill_1 FILLER_70_888 ();
 sg13g2_fill_2 FILLER_70_903 ();
 sg13g2_fill_1 FILLER_70_905 ();
 sg13g2_fill_1 FILLER_70_912 ();
 sg13g2_decap_4 FILLER_70_919 ();
 sg13g2_fill_1 FILLER_70_941 ();
 sg13g2_fill_1 FILLER_70_951 ();
 sg13g2_fill_2 FILLER_70_984 ();
 sg13g2_decap_4 FILLER_70_1022 ();
 sg13g2_fill_2 FILLER_70_1026 ();
 sg13g2_fill_2 FILLER_70_1036 ();
 sg13g2_fill_1 FILLER_70_1038 ();
 sg13g2_fill_2 FILLER_70_1093 ();
 sg13g2_fill_2 FILLER_70_1113 ();
 sg13g2_decap_8 FILLER_70_1119 ();
 sg13g2_fill_1 FILLER_70_1126 ();
 sg13g2_decap_4 FILLER_70_1131 ();
 sg13g2_decap_8 FILLER_70_1139 ();
 sg13g2_fill_1 FILLER_70_1146 ();
 sg13g2_decap_4 FILLER_70_1173 ();
 sg13g2_fill_2 FILLER_70_1177 ();
 sg13g2_fill_1 FILLER_70_1209 ();
 sg13g2_decap_4 FILLER_70_1227 ();
 sg13g2_decap_4 FILLER_70_1235 ();
 sg13g2_fill_1 FILLER_70_1239 ();
 sg13g2_fill_2 FILLER_70_1252 ();
 sg13g2_fill_1 FILLER_70_1254 ();
 sg13g2_fill_1 FILLER_70_1267 ();
 sg13g2_decap_4 FILLER_70_1272 ();
 sg13g2_fill_1 FILLER_70_1281 ();
 sg13g2_decap_4 FILLER_70_1304 ();
 sg13g2_fill_1 FILLER_70_1308 ();
 sg13g2_fill_1 FILLER_70_1317 ();
 sg13g2_decap_4 FILLER_70_1323 ();
 sg13g2_fill_2 FILLER_70_1327 ();
 sg13g2_fill_1 FILLER_70_1344 ();
 sg13g2_fill_1 FILLER_70_1360 ();
 sg13g2_decap_8 FILLER_70_1367 ();
 sg13g2_fill_1 FILLER_70_1374 ();
 sg13g2_decap_8 FILLER_70_1379 ();
 sg13g2_fill_2 FILLER_70_1386 ();
 sg13g2_fill_1 FILLER_70_1397 ();
 sg13g2_fill_2 FILLER_70_1415 ();
 sg13g2_fill_2 FILLER_70_1446 ();
 sg13g2_decap_8 FILLER_70_1453 ();
 sg13g2_fill_2 FILLER_70_1460 ();
 sg13g2_fill_1 FILLER_70_1462 ();
 sg13g2_fill_1 FILLER_70_1477 ();
 sg13g2_fill_2 FILLER_70_1515 ();
 sg13g2_fill_2 FILLER_70_1538 ();
 sg13g2_fill_1 FILLER_70_1540 ();
 sg13g2_decap_8 FILLER_70_1548 ();
 sg13g2_decap_8 FILLER_70_1555 ();
 sg13g2_decap_8 FILLER_70_1562 ();
 sg13g2_decap_8 FILLER_70_1569 ();
 sg13g2_decap_8 FILLER_70_1576 ();
 sg13g2_decap_8 FILLER_70_1583 ();
 sg13g2_fill_2 FILLER_70_1590 ();
 sg13g2_fill_1 FILLER_70_1592 ();
 sg13g2_fill_1 FILLER_70_1620 ();
 sg13g2_decap_4 FILLER_70_1629 ();
 sg13g2_fill_2 FILLER_70_1633 ();
 sg13g2_fill_1 FILLER_70_1651 ();
 sg13g2_fill_2 FILLER_70_1657 ();
 sg13g2_fill_1 FILLER_70_1659 ();
 sg13g2_fill_2 FILLER_70_1668 ();
 sg13g2_fill_2 FILLER_70_1678 ();
 sg13g2_fill_1 FILLER_70_1680 ();
 sg13g2_decap_4 FILLER_70_1693 ();
 sg13g2_fill_1 FILLER_70_1697 ();
 sg13g2_fill_1 FILLER_70_1702 ();
 sg13g2_decap_4 FILLER_70_1708 ();
 sg13g2_fill_1 FILLER_70_1712 ();
 sg13g2_fill_1 FILLER_70_1728 ();
 sg13g2_fill_1 FILLER_70_1734 ();
 sg13g2_fill_2 FILLER_70_1745 ();
 sg13g2_fill_1 FILLER_70_1747 ();
 sg13g2_fill_2 FILLER_70_1773 ();
 sg13g2_decap_4 FILLER_70_1784 ();
 sg13g2_decap_4 FILLER_70_1803 ();
 sg13g2_decap_4 FILLER_70_1812 ();
 sg13g2_fill_1 FILLER_70_1821 ();
 sg13g2_fill_1 FILLER_70_1843 ();
 sg13g2_decap_8 FILLER_70_1848 ();
 sg13g2_decap_8 FILLER_70_1855 ();
 sg13g2_decap_8 FILLER_70_1862 ();
 sg13g2_decap_8 FILLER_70_1873 ();
 sg13g2_decap_4 FILLER_70_1880 ();
 sg13g2_fill_1 FILLER_70_1884 ();
 sg13g2_fill_1 FILLER_70_1889 ();
 sg13g2_fill_2 FILLER_70_1932 ();
 sg13g2_fill_1 FILLER_70_1960 ();
 sg13g2_fill_2 FILLER_70_1965 ();
 sg13g2_decap_4 FILLER_70_1977 ();
 sg13g2_fill_2 FILLER_70_2017 ();
 sg13g2_fill_1 FILLER_70_2054 ();
 sg13g2_fill_1 FILLER_70_2074 ();
 sg13g2_fill_2 FILLER_70_2109 ();
 sg13g2_fill_1 FILLER_70_2111 ();
 sg13g2_fill_2 FILLER_70_2179 ();
 sg13g2_fill_2 FILLER_70_2249 ();
 sg13g2_fill_2 FILLER_70_2277 ();
 sg13g2_fill_1 FILLER_70_2285 ();
 sg13g2_decap_8 FILLER_70_2321 ();
 sg13g2_decap_8 FILLER_70_2328 ();
 sg13g2_fill_1 FILLER_70_2335 ();
 sg13g2_fill_1 FILLER_70_2352 ();
 sg13g2_decap_4 FILLER_70_2367 ();
 sg13g2_fill_2 FILLER_70_2371 ();
 sg13g2_fill_1 FILLER_70_2384 ();
 sg13g2_decap_8 FILLER_70_2440 ();
 sg13g2_decap_8 FILLER_70_2447 ();
 sg13g2_decap_4 FILLER_70_2454 ();
 sg13g2_fill_2 FILLER_70_2479 ();
 sg13g2_fill_1 FILLER_70_2481 ();
 sg13g2_fill_1 FILLER_70_2585 ();
 sg13g2_decap_8 FILLER_70_2604 ();
 sg13g2_decap_8 FILLER_70_2611 ();
 sg13g2_decap_8 FILLER_70_2618 ();
 sg13g2_decap_8 FILLER_70_2625 ();
 sg13g2_decap_8 FILLER_70_2632 ();
 sg13g2_decap_8 FILLER_70_2639 ();
 sg13g2_decap_8 FILLER_70_2646 ();
 sg13g2_decap_8 FILLER_70_2653 ();
 sg13g2_decap_8 FILLER_70_2660 ();
 sg13g2_fill_2 FILLER_70_2667 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_fill_2 FILLER_71_7 ();
 sg13g2_fill_1 FILLER_71_35 ();
 sg13g2_fill_2 FILLER_71_41 ();
 sg13g2_decap_8 FILLER_71_53 ();
 sg13g2_fill_1 FILLER_71_60 ();
 sg13g2_decap_4 FILLER_71_66 ();
 sg13g2_fill_1 FILLER_71_70 ();
 sg13g2_decap_4 FILLER_71_114 ();
 sg13g2_fill_2 FILLER_71_122 ();
 sg13g2_fill_1 FILLER_71_124 ();
 sg13g2_fill_1 FILLER_71_160 ();
 sg13g2_fill_2 FILLER_71_171 ();
 sg13g2_fill_1 FILLER_71_199 ();
 sg13g2_fill_2 FILLER_71_209 ();
 sg13g2_fill_2 FILLER_71_255 ();
 sg13g2_fill_1 FILLER_71_257 ();
 sg13g2_fill_2 FILLER_71_271 ();
 sg13g2_decap_8 FILLER_71_278 ();
 sg13g2_decap_8 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_306 ();
 sg13g2_fill_1 FILLER_71_313 ();
 sg13g2_decap_4 FILLER_71_323 ();
 sg13g2_fill_2 FILLER_71_331 ();
 sg13g2_fill_1 FILLER_71_333 ();
 sg13g2_decap_8 FILLER_71_369 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_1 FILLER_71_378 ();
 sg13g2_decap_4 FILLER_71_388 ();
 sg13g2_fill_1 FILLER_71_396 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_71_409 ();
 sg13g2_decap_4 FILLER_71_416 ();
 sg13g2_fill_1 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_425 ();
 sg13g2_fill_1 FILLER_71_427 ();
 sg13g2_decap_4 FILLER_71_442 ();
 sg13g2_decap_8 FILLER_71_463 ();
 sg13g2_decap_8 FILLER_71_470 ();
 sg13g2_decap_8 FILLER_71_477 ();
 sg13g2_decap_8 FILLER_71_484 ();
 sg13g2_fill_2 FILLER_71_499 ();
 sg13g2_fill_1 FILLER_71_501 ();
 sg13g2_decap_8 FILLER_71_512 ();
 sg13g2_decap_8 FILLER_71_519 ();
 sg13g2_fill_2 FILLER_71_526 ();
 sg13g2_fill_1 FILLER_71_528 ();
 sg13g2_fill_2 FILLER_71_533 ();
 sg13g2_fill_1 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_558 ();
 sg13g2_decap_4 FILLER_71_565 ();
 sg13g2_decap_8 FILLER_71_572 ();
 sg13g2_fill_2 FILLER_71_579 ();
 sg13g2_fill_2 FILLER_71_598 ();
 sg13g2_fill_1 FILLER_71_615 ();
 sg13g2_fill_2 FILLER_71_660 ();
 sg13g2_fill_2 FILLER_71_666 ();
 sg13g2_fill_1 FILLER_71_668 ();
 sg13g2_decap_8 FILLER_71_695 ();
 sg13g2_decap_8 FILLER_71_702 ();
 sg13g2_fill_1 FILLER_71_779 ();
 sg13g2_decap_8 FILLER_71_806 ();
 sg13g2_fill_2 FILLER_71_813 ();
 sg13g2_fill_2 FILLER_71_819 ();
 sg13g2_fill_1 FILLER_71_821 ();
 sg13g2_fill_2 FILLER_71_832 ();
 sg13g2_fill_2 FILLER_71_839 ();
 sg13g2_fill_1 FILLER_71_841 ();
 sg13g2_fill_1 FILLER_71_852 ();
 sg13g2_decap_4 FILLER_71_879 ();
 sg13g2_fill_2 FILLER_71_883 ();
 sg13g2_decap_8 FILLER_71_911 ();
 sg13g2_decap_8 FILLER_71_918 ();
 sg13g2_fill_2 FILLER_71_925 ();
 sg13g2_fill_1 FILLER_71_927 ();
 sg13g2_decap_4 FILLER_71_934 ();
 sg13g2_fill_1 FILLER_71_938 ();
 sg13g2_decap_8 FILLER_71_987 ();
 sg13g2_decap_4 FILLER_71_994 ();
 sg13g2_fill_2 FILLER_71_998 ();
 sg13g2_decap_8 FILLER_71_1008 ();
 sg13g2_fill_1 FILLER_71_1015 ();
 sg13g2_decap_4 FILLER_71_1055 ();
 sg13g2_fill_1 FILLER_71_1059 ();
 sg13g2_fill_1 FILLER_71_1088 ();
 sg13g2_decap_8 FILLER_71_1106 ();
 sg13g2_decap_8 FILLER_71_1113 ();
 sg13g2_fill_1 FILLER_71_1137 ();
 sg13g2_fill_1 FILLER_71_1174 ();
 sg13g2_fill_1 FILLER_71_1179 ();
 sg13g2_fill_1 FILLER_71_1225 ();
 sg13g2_fill_2 FILLER_71_1248 ();
 sg13g2_fill_1 FILLER_71_1250 ();
 sg13g2_decap_4 FILLER_71_1296 ();
 sg13g2_fill_1 FILLER_71_1310 ();
 sg13g2_fill_2 FILLER_71_1329 ();
 sg13g2_decap_8 FILLER_71_1361 ();
 sg13g2_decap_8 FILLER_71_1368 ();
 sg13g2_fill_1 FILLER_71_1401 ();
 sg13g2_fill_1 FILLER_71_1406 ();
 sg13g2_decap_4 FILLER_71_1416 ();
 sg13g2_fill_2 FILLER_71_1434 ();
 sg13g2_fill_1 FILLER_71_1441 ();
 sg13g2_fill_1 FILLER_71_1452 ();
 sg13g2_fill_2 FILLER_71_1458 ();
 sg13g2_fill_1 FILLER_71_1460 ();
 sg13g2_fill_1 FILLER_71_1488 ();
 sg13g2_fill_1 FILLER_71_1494 ();
 sg13g2_fill_1 FILLER_71_1499 ();
 sg13g2_fill_2 FILLER_71_1503 ();
 sg13g2_fill_1 FILLER_71_1509 ();
 sg13g2_fill_2 FILLER_71_1514 ();
 sg13g2_fill_1 FILLER_71_1516 ();
 sg13g2_fill_2 FILLER_71_1530 ();
 sg13g2_decap_8 FILLER_71_1543 ();
 sg13g2_decap_8 FILLER_71_1554 ();
 sg13g2_fill_1 FILLER_71_1561 ();
 sg13g2_fill_1 FILLER_71_1566 ();
 sg13g2_fill_2 FILLER_71_1572 ();
 sg13g2_fill_1 FILLER_71_1574 ();
 sg13g2_decap_8 FILLER_71_1579 ();
 sg13g2_decap_4 FILLER_71_1586 ();
 sg13g2_fill_2 FILLER_71_1590 ();
 sg13g2_fill_1 FILLER_71_1616 ();
 sg13g2_fill_1 FILLER_71_1632 ();
 sg13g2_fill_2 FILLER_71_1643 ();
 sg13g2_fill_1 FILLER_71_1645 ();
 sg13g2_fill_1 FILLER_71_1657 ();
 sg13g2_decap_8 FILLER_71_1664 ();
 sg13g2_decap_8 FILLER_71_1686 ();
 sg13g2_fill_2 FILLER_71_1693 ();
 sg13g2_fill_1 FILLER_71_1695 ();
 sg13g2_fill_2 FILLER_71_1709 ();
 sg13g2_fill_1 FILLER_71_1711 ();
 sg13g2_decap_8 FILLER_71_1729 ();
 sg13g2_decap_4 FILLER_71_1736 ();
 sg13g2_fill_1 FILLER_71_1740 ();
 sg13g2_fill_1 FILLER_71_1745 ();
 sg13g2_fill_2 FILLER_71_1751 ();
 sg13g2_decap_4 FILLER_71_1769 ();
 sg13g2_fill_2 FILLER_71_1773 ();
 sg13g2_fill_2 FILLER_71_1780 ();
 sg13g2_fill_1 FILLER_71_1782 ();
 sg13g2_decap_8 FILLER_71_1845 ();
 sg13g2_decap_8 FILLER_71_1852 ();
 sg13g2_decap_8 FILLER_71_1859 ();
 sg13g2_decap_8 FILLER_71_1866 ();
 sg13g2_decap_8 FILLER_71_1873 ();
 sg13g2_decap_8 FILLER_71_1880 ();
 sg13g2_fill_1 FILLER_71_1887 ();
 sg13g2_fill_1 FILLER_71_1940 ();
 sg13g2_fill_2 FILLER_71_1967 ();
 sg13g2_fill_1 FILLER_71_1995 ();
 sg13g2_fill_2 FILLER_71_2041 ();
 sg13g2_fill_1 FILLER_71_2050 ();
 sg13g2_fill_1 FILLER_71_2069 ();
 sg13g2_fill_1 FILLER_71_2078 ();
 sg13g2_decap_4 FILLER_71_2087 ();
 sg13g2_fill_1 FILLER_71_2091 ();
 sg13g2_fill_1 FILLER_71_2097 ();
 sg13g2_fill_2 FILLER_71_2145 ();
 sg13g2_fill_1 FILLER_71_2212 ();
 sg13g2_fill_1 FILLER_71_2235 ();
 sg13g2_fill_2 FILLER_71_2240 ();
 sg13g2_decap_8 FILLER_71_2252 ();
 sg13g2_fill_1 FILLER_71_2259 ();
 sg13g2_decap_4 FILLER_71_2264 ();
 sg13g2_fill_2 FILLER_71_2279 ();
 sg13g2_fill_1 FILLER_71_2281 ();
 sg13g2_decap_4 FILLER_71_2292 ();
 sg13g2_fill_2 FILLER_71_2296 ();
 sg13g2_decap_8 FILLER_71_2302 ();
 sg13g2_fill_2 FILLER_71_2309 ();
 sg13g2_fill_1 FILLER_71_2311 ();
 sg13g2_fill_1 FILLER_71_2316 ();
 sg13g2_decap_8 FILLER_71_2333 ();
 sg13g2_decap_4 FILLER_71_2340 ();
 sg13g2_fill_2 FILLER_71_2344 ();
 sg13g2_fill_1 FILLER_71_2358 ();
 sg13g2_decap_8 FILLER_71_2385 ();
 sg13g2_fill_1 FILLER_71_2392 ();
 sg13g2_fill_2 FILLER_71_2407 ();
 sg13g2_fill_1 FILLER_71_2409 ();
 sg13g2_fill_1 FILLER_71_2436 ();
 sg13g2_fill_2 FILLER_71_2450 ();
 sg13g2_fill_2 FILLER_71_2462 ();
 sg13g2_decap_8 FILLER_71_2470 ();
 sg13g2_decap_4 FILLER_71_2477 ();
 sg13g2_fill_1 FILLER_71_2515 ();
 sg13g2_fill_1 FILLER_71_2547 ();
 sg13g2_fill_1 FILLER_71_2552 ();
 sg13g2_fill_2 FILLER_71_2568 ();
 sg13g2_fill_1 FILLER_71_2570 ();
 sg13g2_decap_8 FILLER_71_2587 ();
 sg13g2_fill_1 FILLER_71_2594 ();
 sg13g2_decap_8 FILLER_71_2621 ();
 sg13g2_decap_8 FILLER_71_2628 ();
 sg13g2_decap_8 FILLER_71_2635 ();
 sg13g2_decap_8 FILLER_71_2642 ();
 sg13g2_decap_8 FILLER_71_2649 ();
 sg13g2_decap_8 FILLER_71_2656 ();
 sg13g2_decap_8 FILLER_71_2663 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_85 ();
 sg13g2_fill_1 FILLER_72_87 ();
 sg13g2_fill_2 FILLER_72_93 ();
 sg13g2_fill_2 FILLER_72_117 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_fill_1 FILLER_72_161 ();
 sg13g2_fill_2 FILLER_72_192 ();
 sg13g2_fill_1 FILLER_72_194 ();
 sg13g2_fill_2 FILLER_72_203 ();
 sg13g2_decap_4 FILLER_72_214 ();
 sg13g2_fill_1 FILLER_72_218 ();
 sg13g2_decap_4 FILLER_72_224 ();
 sg13g2_fill_2 FILLER_72_228 ();
 sg13g2_decap_4 FILLER_72_255 ();
 sg13g2_fill_2 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_265 ();
 sg13g2_decap_4 FILLER_72_302 ();
 sg13g2_fill_2 FILLER_72_356 ();
 sg13g2_fill_1 FILLER_72_358 ();
 sg13g2_fill_2 FILLER_72_364 ();
 sg13g2_fill_1 FILLER_72_379 ();
 sg13g2_decap_4 FILLER_72_410 ();
 sg13g2_decap_8 FILLER_72_418 ();
 sg13g2_decap_4 FILLER_72_425 ();
 sg13g2_decap_4 FILLER_72_433 ();
 sg13g2_fill_1 FILLER_72_437 ();
 sg13g2_decap_8 FILLER_72_486 ();
 sg13g2_decap_8 FILLER_72_493 ();
 sg13g2_fill_1 FILLER_72_500 ();
 sg13g2_decap_4 FILLER_72_542 ();
 sg13g2_fill_2 FILLER_72_546 ();
 sg13g2_decap_8 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_570 ();
 sg13g2_fill_2 FILLER_72_581 ();
 sg13g2_fill_1 FILLER_72_583 ();
 sg13g2_fill_2 FILLER_72_589 ();
 sg13g2_fill_1 FILLER_72_625 ();
 sg13g2_fill_1 FILLER_72_640 ();
 sg13g2_fill_2 FILLER_72_654 ();
 sg13g2_fill_1 FILLER_72_662 ();
 sg13g2_decap_4 FILLER_72_705 ();
 sg13g2_decap_4 FILLER_72_775 ();
 sg13g2_decap_8 FILLER_72_810 ();
 sg13g2_fill_2 FILLER_72_817 ();
 sg13g2_fill_2 FILLER_72_872 ();
 sg13g2_fill_1 FILLER_72_874 ();
 sg13g2_fill_2 FILLER_72_889 ();
 sg13g2_fill_2 FILLER_72_953 ();
 sg13g2_fill_1 FILLER_72_985 ();
 sg13g2_decap_4 FILLER_72_1022 ();
 sg13g2_fill_1 FILLER_72_1026 ();
 sg13g2_decap_4 FILLER_72_1031 ();
 sg13g2_decap_8 FILLER_72_1064 ();
 sg13g2_decap_8 FILLER_72_1071 ();
 sg13g2_fill_2 FILLER_72_1137 ();
 sg13g2_fill_1 FILLER_72_1139 ();
 sg13g2_decap_4 FILLER_72_1150 ();
 sg13g2_fill_1 FILLER_72_1154 ();
 sg13g2_decap_4 FILLER_72_1159 ();
 sg13g2_decap_8 FILLER_72_1167 ();
 sg13g2_decap_8 FILLER_72_1174 ();
 sg13g2_decap_4 FILLER_72_1181 ();
 sg13g2_decap_4 FILLER_72_1189 ();
 sg13g2_decap_8 FILLER_72_1227 ();
 sg13g2_decap_4 FILLER_72_1234 ();
 sg13g2_fill_2 FILLER_72_1238 ();
 sg13g2_decap_4 FILLER_72_1257 ();
 sg13g2_fill_2 FILLER_72_1266 ();
 sg13g2_fill_1 FILLER_72_1268 ();
 sg13g2_fill_1 FILLER_72_1291 ();
 sg13g2_fill_1 FILLER_72_1297 ();
 sg13g2_fill_2 FILLER_72_1324 ();
 sg13g2_fill_2 FILLER_72_1347 ();
 sg13g2_fill_1 FILLER_72_1349 ();
 sg13g2_decap_8 FILLER_72_1355 ();
 sg13g2_decap_8 FILLER_72_1362 ();
 sg13g2_decap_4 FILLER_72_1369 ();
 sg13g2_fill_1 FILLER_72_1386 ();
 sg13g2_fill_1 FILLER_72_1392 ();
 sg13g2_fill_1 FILLER_72_1400 ();
 sg13g2_fill_1 FILLER_72_1405 ();
 sg13g2_fill_2 FILLER_72_1442 ();
 sg13g2_fill_1 FILLER_72_1448 ();
 sg13g2_decap_8 FILLER_72_1453 ();
 sg13g2_decap_8 FILLER_72_1460 ();
 sg13g2_fill_2 FILLER_72_1467 ();
 sg13g2_fill_2 FILLER_72_1491 ();
 sg13g2_fill_1 FILLER_72_1510 ();
 sg13g2_fill_1 FILLER_72_1515 ();
 sg13g2_fill_1 FILLER_72_1525 ();
 sg13g2_fill_2 FILLER_72_1539 ();
 sg13g2_fill_2 FILLER_72_1571 ();
 sg13g2_decap_8 FILLER_72_1578 ();
 sg13g2_decap_4 FILLER_72_1585 ();
 sg13g2_fill_1 FILLER_72_1589 ();
 sg13g2_decap_4 FILLER_72_1594 ();
 sg13g2_fill_2 FILLER_72_1618 ();
 sg13g2_decap_8 FILLER_72_1625 ();
 sg13g2_decap_4 FILLER_72_1632 ();
 sg13g2_decap_8 FILLER_72_1640 ();
 sg13g2_fill_2 FILLER_72_1647 ();
 sg13g2_fill_1 FILLER_72_1649 ();
 sg13g2_decap_8 FILLER_72_1654 ();
 sg13g2_fill_1 FILLER_72_1661 ();
 sg13g2_decap_4 FILLER_72_1666 ();
 sg13g2_fill_2 FILLER_72_1670 ();
 sg13g2_fill_2 FILLER_72_1686 ();
 sg13g2_decap_8 FILLER_72_1695 ();
 sg13g2_fill_2 FILLER_72_1717 ();
 sg13g2_decap_8 FILLER_72_1723 ();
 sg13g2_decap_8 FILLER_72_1730 ();
 sg13g2_fill_1 FILLER_72_1737 ();
 sg13g2_fill_1 FILLER_72_1743 ();
 sg13g2_decap_4 FILLER_72_1749 ();
 sg13g2_fill_1 FILLER_72_1753 ();
 sg13g2_fill_1 FILLER_72_1759 ();
 sg13g2_fill_2 FILLER_72_1773 ();
 sg13g2_fill_1 FILLER_72_1775 ();
 sg13g2_fill_2 FILLER_72_1799 ();
 sg13g2_fill_1 FILLER_72_1801 ();
 sg13g2_fill_1 FILLER_72_1807 ();
 sg13g2_fill_1 FILLER_72_1839 ();
 sg13g2_decap_8 FILLER_72_1850 ();
 sg13g2_decap_8 FILLER_72_1857 ();
 sg13g2_decap_8 FILLER_72_1864 ();
 sg13g2_decap_8 FILLER_72_1871 ();
 sg13g2_decap_8 FILLER_72_1878 ();
 sg13g2_decap_8 FILLER_72_1885 ();
 sg13g2_decap_4 FILLER_72_1892 ();
 sg13g2_fill_1 FILLER_72_1896 ();
 sg13g2_fill_1 FILLER_72_1907 ();
 sg13g2_decap_4 FILLER_72_1912 ();
 sg13g2_fill_2 FILLER_72_1926 ();
 sg13g2_fill_1 FILLER_72_1928 ();
 sg13g2_fill_2 FILLER_72_1955 ();
 sg13g2_fill_1 FILLER_72_1977 ();
 sg13g2_fill_1 FILLER_72_1992 ();
 sg13g2_fill_2 FILLER_72_2022 ();
 sg13g2_fill_1 FILLER_72_2024 ();
 sg13g2_fill_1 FILLER_72_2029 ();
 sg13g2_fill_1 FILLER_72_2060 ();
 sg13g2_fill_2 FILLER_72_2071 ();
 sg13g2_fill_1 FILLER_72_2097 ();
 sg13g2_fill_2 FILLER_72_2120 ();
 sg13g2_decap_8 FILLER_72_2126 ();
 sg13g2_fill_1 FILLER_72_2133 ();
 sg13g2_fill_2 FILLER_72_2160 ();
 sg13g2_fill_1 FILLER_72_2162 ();
 sg13g2_decap_8 FILLER_72_2167 ();
 sg13g2_fill_1 FILLER_72_2182 ();
 sg13g2_fill_2 FILLER_72_2258 ();
 sg13g2_decap_8 FILLER_72_2265 ();
 sg13g2_decap_4 FILLER_72_2272 ();
 sg13g2_fill_1 FILLER_72_2276 ();
 sg13g2_decap_8 FILLER_72_2287 ();
 sg13g2_decap_4 FILLER_72_2298 ();
 sg13g2_fill_1 FILLER_72_2302 ();
 sg13g2_decap_4 FILLER_72_2338 ();
 sg13g2_decap_8 FILLER_72_2357 ();
 sg13g2_fill_2 FILLER_72_2364 ();
 sg13g2_fill_1 FILLER_72_2376 ();
 sg13g2_decap_4 FILLER_72_2389 ();
 sg13g2_fill_1 FILLER_72_2393 ();
 sg13g2_decap_4 FILLER_72_2404 ();
 sg13g2_fill_1 FILLER_72_2408 ();
 sg13g2_fill_2 FILLER_72_2475 ();
 sg13g2_decap_4 FILLER_72_2487 ();
 sg13g2_fill_1 FILLER_72_2491 ();
 sg13g2_decap_8 FILLER_72_2512 ();
 sg13g2_fill_1 FILLER_72_2519 ();
 sg13g2_fill_2 FILLER_72_2530 ();
 sg13g2_fill_2 FILLER_72_2554 ();
 sg13g2_fill_2 FILLER_72_2569 ();
 sg13g2_decap_8 FILLER_72_2581 ();
 sg13g2_decap_8 FILLER_72_2614 ();
 sg13g2_decap_8 FILLER_72_2621 ();
 sg13g2_decap_8 FILLER_72_2628 ();
 sg13g2_decap_8 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2642 ();
 sg13g2_decap_8 FILLER_72_2649 ();
 sg13g2_decap_8 FILLER_72_2656 ();
 sg13g2_decap_8 FILLER_72_2663 ();
 sg13g2_fill_1 FILLER_73_0 ();
 sg13g2_fill_1 FILLER_73_5 ();
 sg13g2_fill_1 FILLER_73_32 ();
 sg13g2_fill_1 FILLER_73_51 ();
 sg13g2_decap_4 FILLER_73_57 ();
 sg13g2_decap_8 FILLER_73_65 ();
 sg13g2_decap_4 FILLER_73_72 ();
 sg13g2_fill_2 FILLER_73_110 ();
 sg13g2_decap_8 FILLER_73_117 ();
 sg13g2_decap_8 FILLER_73_124 ();
 sg13g2_fill_1 FILLER_73_131 ();
 sg13g2_decap_8 FILLER_73_136 ();
 sg13g2_decap_8 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_150 ();
 sg13g2_decap_4 FILLER_73_156 ();
 sg13g2_fill_2 FILLER_73_183 ();
 sg13g2_decap_4 FILLER_73_189 ();
 sg13g2_fill_2 FILLER_73_236 ();
 sg13g2_fill_1 FILLER_73_238 ();
 sg13g2_fill_1 FILLER_73_288 ();
 sg13g2_fill_2 FILLER_73_294 ();
 sg13g2_fill_1 FILLER_73_296 ();
 sg13g2_fill_2 FILLER_73_314 ();
 sg13g2_fill_2 FILLER_73_337 ();
 sg13g2_decap_8 FILLER_73_374 ();
 sg13g2_decap_8 FILLER_73_425 ();
 sg13g2_fill_2 FILLER_73_432 ();
 sg13g2_fill_1 FILLER_73_439 ();
 sg13g2_fill_1 FILLER_73_444 ();
 sg13g2_fill_1 FILLER_73_449 ();
 sg13g2_fill_1 FILLER_73_454 ();
 sg13g2_fill_1 FILLER_73_459 ();
 sg13g2_fill_2 FILLER_73_506 ();
 sg13g2_fill_2 FILLER_73_542 ();
 sg13g2_fill_1 FILLER_73_544 ();
 sg13g2_decap_4 FILLER_73_550 ();
 sg13g2_fill_2 FILLER_73_554 ();
 sg13g2_decap_4 FILLER_73_568 ();
 sg13g2_fill_2 FILLER_73_607 ();
 sg13g2_fill_2 FILLER_73_616 ();
 sg13g2_fill_2 FILLER_73_657 ();
 sg13g2_fill_1 FILLER_73_685 ();
 sg13g2_fill_2 FILLER_73_690 ();
 sg13g2_fill_1 FILLER_73_692 ();
 sg13g2_decap_8 FILLER_73_697 ();
 sg13g2_fill_1 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_709 ();
 sg13g2_fill_2 FILLER_73_736 ();
 sg13g2_decap_8 FILLER_73_776 ();
 sg13g2_decap_8 FILLER_73_783 ();
 sg13g2_fill_1 FILLER_73_790 ();
 sg13g2_decap_4 FILLER_73_801 ();
 sg13g2_decap_8 FILLER_73_815 ();
 sg13g2_fill_2 FILLER_73_822 ();
 sg13g2_fill_1 FILLER_73_824 ();
 sg13g2_fill_1 FILLER_73_835 ();
 sg13g2_fill_2 FILLER_73_953 ();
 sg13g2_fill_2 FILLER_73_961 ();
 sg13g2_decap_4 FILLER_73_976 ();
 sg13g2_fill_2 FILLER_73_980 ();
 sg13g2_fill_2 FILLER_73_1038 ();
 sg13g2_fill_1 FILLER_73_1106 ();
 sg13g2_fill_1 FILLER_73_1133 ();
 sg13g2_fill_2 FILLER_73_1160 ();
 sg13g2_decap_8 FILLER_73_1166 ();
 sg13g2_decap_8 FILLER_73_1173 ();
 sg13g2_decap_8 FILLER_73_1180 ();
 sg13g2_decap_8 FILLER_73_1187 ();
 sg13g2_decap_8 FILLER_73_1194 ();
 sg13g2_fill_1 FILLER_73_1201 ();
 sg13g2_decap_8 FILLER_73_1225 ();
 sg13g2_decap_8 FILLER_73_1232 ();
 sg13g2_fill_2 FILLER_73_1239 ();
 sg13g2_fill_1 FILLER_73_1241 ();
 sg13g2_decap_4 FILLER_73_1246 ();
 sg13g2_fill_1 FILLER_73_1250 ();
 sg13g2_decap_8 FILLER_73_1257 ();
 sg13g2_fill_2 FILLER_73_1273 ();
 sg13g2_fill_1 FILLER_73_1275 ();
 sg13g2_fill_2 FILLER_73_1281 ();
 sg13g2_fill_2 FILLER_73_1288 ();
 sg13g2_fill_1 FILLER_73_1290 ();
 sg13g2_decap_8 FILLER_73_1295 ();
 sg13g2_fill_2 FILLER_73_1302 ();
 sg13g2_decap_8 FILLER_73_1313 ();
 sg13g2_fill_2 FILLER_73_1320 ();
 sg13g2_fill_1 FILLER_73_1322 ();
 sg13g2_decap_4 FILLER_73_1326 ();
 sg13g2_fill_1 FILLER_73_1336 ();
 sg13g2_decap_8 FILLER_73_1349 ();
 sg13g2_decap_4 FILLER_73_1356 ();
 sg13g2_decap_8 FILLER_73_1368 ();
 sg13g2_fill_1 FILLER_73_1375 ();
 sg13g2_fill_2 FILLER_73_1397 ();
 sg13g2_fill_1 FILLER_73_1399 ();
 sg13g2_fill_2 FILLER_73_1404 ();
 sg13g2_fill_1 FILLER_73_1406 ();
 sg13g2_fill_2 FILLER_73_1426 ();
 sg13g2_decap_8 FILLER_73_1465 ();
 sg13g2_decap_4 FILLER_73_1472 ();
 sg13g2_fill_2 FILLER_73_1476 ();
 sg13g2_decap_4 FILLER_73_1485 ();
 sg13g2_fill_1 FILLER_73_1492 ();
 sg13g2_fill_2 FILLER_73_1503 ();
 sg13g2_fill_1 FILLER_73_1505 ();
 sg13g2_fill_1 FILLER_73_1519 ();
 sg13g2_decap_8 FILLER_73_1565 ();
 sg13g2_decap_4 FILLER_73_1572 ();
 sg13g2_fill_1 FILLER_73_1576 ();
 sg13g2_fill_1 FILLER_73_1582 ();
 sg13g2_fill_2 FILLER_73_1587 ();
 sg13g2_fill_1 FILLER_73_1598 ();
 sg13g2_fill_2 FILLER_73_1607 ();
 sg13g2_fill_2 FILLER_73_1619 ();
 sg13g2_fill_1 FILLER_73_1633 ();
 sg13g2_decap_8 FILLER_73_1640 ();
 sg13g2_fill_1 FILLER_73_1647 ();
 sg13g2_decap_4 FILLER_73_1653 ();
 sg13g2_fill_2 FILLER_73_1657 ();
 sg13g2_decap_8 FILLER_73_1678 ();
 sg13g2_fill_1 FILLER_73_1685 ();
 sg13g2_decap_8 FILLER_73_1691 ();
 sg13g2_decap_8 FILLER_73_1698 ();
 sg13g2_fill_2 FILLER_73_1705 ();
 sg13g2_fill_2 FILLER_73_1717 ();
 sg13g2_decap_8 FILLER_73_1734 ();
 sg13g2_decap_4 FILLER_73_1741 ();
 sg13g2_decap_4 FILLER_73_1765 ();
 sg13g2_fill_2 FILLER_73_1769 ();
 sg13g2_fill_2 FILLER_73_1794 ();
 sg13g2_fill_1 FILLER_73_1802 ();
 sg13g2_fill_1 FILLER_73_1809 ();
 sg13g2_decap_8 FILLER_73_1856 ();
 sg13g2_decap_8 FILLER_73_1863 ();
 sg13g2_fill_1 FILLER_73_1870 ();
 sg13g2_fill_1 FILLER_73_1929 ();
 sg13g2_fill_2 FILLER_73_1940 ();
 sg13g2_decap_8 FILLER_73_1956 ();
 sg13g2_fill_2 FILLER_73_1963 ();
 sg13g2_decap_8 FILLER_73_1991 ();
 sg13g2_decap_8 FILLER_73_1998 ();
 sg13g2_fill_2 FILLER_73_2005 ();
 sg13g2_fill_1 FILLER_73_2017 ();
 sg13g2_fill_2 FILLER_73_2087 ();
 sg13g2_fill_1 FILLER_73_2089 ();
 sg13g2_fill_1 FILLER_73_2120 ();
 sg13g2_decap_4 FILLER_73_2127 ();
 sg13g2_fill_1 FILLER_73_2136 ();
 sg13g2_fill_2 FILLER_73_2141 ();
 sg13g2_decap_8 FILLER_73_2147 ();
 sg13g2_decap_4 FILLER_73_2169 ();
 sg13g2_fill_2 FILLER_73_2186 ();
 sg13g2_decap_8 FILLER_73_2242 ();
 sg13g2_fill_2 FILLER_73_2392 ();
 sg13g2_fill_1 FILLER_73_2394 ();
 sg13g2_decap_8 FILLER_73_2421 ();
 sg13g2_fill_2 FILLER_73_2428 ();
 sg13g2_fill_1 FILLER_73_2430 ();
 sg13g2_decap_8 FILLER_73_2435 ();
 sg13g2_decap_8 FILLER_73_2442 ();
 sg13g2_decap_4 FILLER_73_2449 ();
 sg13g2_fill_1 FILLER_73_2457 ();
 sg13g2_fill_2 FILLER_73_2468 ();
 sg13g2_fill_1 FILLER_73_2539 ();
 sg13g2_decap_4 FILLER_73_2576 ();
 sg13g2_fill_1 FILLER_73_2580 ();
 sg13g2_decap_8 FILLER_73_2617 ();
 sg13g2_decap_8 FILLER_73_2624 ();
 sg13g2_decap_8 FILLER_73_2631 ();
 sg13g2_decap_8 FILLER_73_2638 ();
 sg13g2_decap_8 FILLER_73_2645 ();
 sg13g2_decap_8 FILLER_73_2652 ();
 sg13g2_decap_8 FILLER_73_2659 ();
 sg13g2_decap_4 FILLER_73_2666 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_38 ();
 sg13g2_fill_1 FILLER_74_42 ();
 sg13g2_fill_2 FILLER_74_48 ();
 sg13g2_fill_1 FILLER_74_76 ();
 sg13g2_fill_1 FILLER_74_81 ();
 sg13g2_fill_2 FILLER_74_103 ();
 sg13g2_fill_2 FILLER_74_110 ();
 sg13g2_fill_1 FILLER_74_112 ();
 sg13g2_fill_1 FILLER_74_118 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_decap_4 FILLER_74_180 ();
 sg13g2_fill_1 FILLER_74_184 ();
 sg13g2_fill_1 FILLER_74_200 ();
 sg13g2_fill_1 FILLER_74_209 ();
 sg13g2_fill_1 FILLER_74_214 ();
 sg13g2_fill_2 FILLER_74_241 ();
 sg13g2_fill_1 FILLER_74_248 ();
 sg13g2_fill_2 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_303 ();
 sg13g2_decap_8 FILLER_74_310 ();
 sg13g2_decap_4 FILLER_74_317 ();
 sg13g2_fill_1 FILLER_74_321 ();
 sg13g2_fill_1 FILLER_74_327 ();
 sg13g2_decap_4 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_371 ();
 sg13g2_decap_8 FILLER_74_376 ();
 sg13g2_fill_2 FILLER_74_418 ();
 sg13g2_fill_1 FILLER_74_420 ();
 sg13g2_decap_8 FILLER_74_426 ();
 sg13g2_fill_2 FILLER_74_433 ();
 sg13g2_fill_1 FILLER_74_435 ();
 sg13g2_fill_1 FILLER_74_462 ();
 sg13g2_decap_8 FILLER_74_502 ();
 sg13g2_decap_4 FILLER_74_509 ();
 sg13g2_fill_1 FILLER_74_513 ();
 sg13g2_fill_2 FILLER_74_523 ();
 sg13g2_fill_1 FILLER_74_525 ();
 sg13g2_fill_2 FILLER_74_531 ();
 sg13g2_decap_8 FILLER_74_546 ();
 sg13g2_decap_4 FILLER_74_553 ();
 sg13g2_fill_1 FILLER_74_557 ();
 sg13g2_fill_1 FILLER_74_591 ();
 sg13g2_fill_2 FILLER_74_600 ();
 sg13g2_fill_1 FILLER_74_621 ();
 sg13g2_fill_1 FILLER_74_642 ();
 sg13g2_fill_2 FILLER_74_652 ();
 sg13g2_fill_1 FILLER_74_659 ();
 sg13g2_fill_1 FILLER_74_664 ();
 sg13g2_fill_1 FILLER_74_675 ();
 sg13g2_fill_2 FILLER_74_684 ();
 sg13g2_decap_4 FILLER_74_712 ();
 sg13g2_fill_2 FILLER_74_742 ();
 sg13g2_fill_2 FILLER_74_770 ();
 sg13g2_fill_1 FILLER_74_772 ();
 sg13g2_fill_2 FILLER_74_799 ();
 sg13g2_fill_1 FILLER_74_801 ();
 sg13g2_fill_2 FILLER_74_828 ();
 sg13g2_fill_2 FILLER_74_882 ();
 sg13g2_fill_1 FILLER_74_938 ();
 sg13g2_fill_2 FILLER_74_943 ();
 sg13g2_decap_8 FILLER_74_969 ();
 sg13g2_fill_1 FILLER_74_976 ();
 sg13g2_decap_4 FILLER_74_999 ();
 sg13g2_fill_2 FILLER_74_1009 ();
 sg13g2_fill_1 FILLER_74_1011 ();
 sg13g2_decap_8 FILLER_74_1026 ();
 sg13g2_decap_4 FILLER_74_1033 ();
 sg13g2_decap_4 FILLER_74_1067 ();
 sg13g2_fill_1 FILLER_74_1071 ();
 sg13g2_fill_2 FILLER_74_1088 ();
 sg13g2_fill_1 FILLER_74_1090 ();
 sg13g2_decap_4 FILLER_74_1095 ();
 sg13g2_fill_1 FILLER_74_1099 ();
 sg13g2_fill_1 FILLER_74_1140 ();
 sg13g2_fill_1 FILLER_74_1151 ();
 sg13g2_decap_8 FILLER_74_1181 ();
 sg13g2_decap_8 FILLER_74_1188 ();
 sg13g2_fill_1 FILLER_74_1195 ();
 sg13g2_fill_1 FILLER_74_1226 ();
 sg13g2_fill_2 FILLER_74_1236 ();
 sg13g2_fill_1 FILLER_74_1238 ();
 sg13g2_decap_8 FILLER_74_1243 ();
 sg13g2_fill_2 FILLER_74_1259 ();
 sg13g2_fill_1 FILLER_74_1276 ();
 sg13g2_fill_2 FILLER_74_1287 ();
 sg13g2_fill_1 FILLER_74_1289 ();
 sg13g2_decap_8 FILLER_74_1295 ();
 sg13g2_decap_8 FILLER_74_1302 ();
 sg13g2_decap_8 FILLER_74_1309 ();
 sg13g2_decap_8 FILLER_74_1316 ();
 sg13g2_fill_2 FILLER_74_1323 ();
 sg13g2_fill_1 FILLER_74_1325 ();
 sg13g2_fill_2 FILLER_74_1337 ();
 sg13g2_decap_4 FILLER_74_1344 ();
 sg13g2_fill_1 FILLER_74_1348 ();
 sg13g2_decap_4 FILLER_74_1354 ();
 sg13g2_decap_8 FILLER_74_1362 ();
 sg13g2_fill_2 FILLER_74_1369 ();
 sg13g2_fill_1 FILLER_74_1371 ();
 sg13g2_fill_1 FILLER_74_1409 ();
 sg13g2_fill_2 FILLER_74_1414 ();
 sg13g2_fill_1 FILLER_74_1416 ();
 sg13g2_fill_1 FILLER_74_1421 ();
 sg13g2_fill_1 FILLER_74_1427 ();
 sg13g2_fill_1 FILLER_74_1432 ();
 sg13g2_fill_1 FILLER_74_1442 ();
 sg13g2_decap_8 FILLER_74_1449 ();
 sg13g2_fill_2 FILLER_74_1460 ();
 sg13g2_fill_2 FILLER_74_1471 ();
 sg13g2_fill_1 FILLER_74_1473 ();
 sg13g2_fill_2 FILLER_74_1524 ();
 sg13g2_decap_4 FILLER_74_1530 ();
 sg13g2_decap_4 FILLER_74_1537 ();
 sg13g2_fill_1 FILLER_74_1545 ();
 sg13g2_decap_8 FILLER_74_1552 ();
 sg13g2_fill_1 FILLER_74_1559 ();
 sg13g2_decap_8 FILLER_74_1584 ();
 sg13g2_fill_1 FILLER_74_1591 ();
 sg13g2_fill_1 FILLER_74_1601 ();
 sg13g2_fill_2 FILLER_74_1623 ();
 sg13g2_fill_1 FILLER_74_1625 ();
 sg13g2_fill_2 FILLER_74_1636 ();
 sg13g2_fill_1 FILLER_74_1643 ();
 sg13g2_decap_4 FILLER_74_1651 ();
 sg13g2_fill_2 FILLER_74_1655 ();
 sg13g2_fill_1 FILLER_74_1666 ();
 sg13g2_fill_2 FILLER_74_1672 ();
 sg13g2_fill_1 FILLER_74_1678 ();
 sg13g2_fill_2 FILLER_74_1687 ();
 sg13g2_decap_8 FILLER_74_1695 ();
 sg13g2_fill_2 FILLER_74_1702 ();
 sg13g2_decap_4 FILLER_74_1709 ();
 sg13g2_fill_2 FILLER_74_1717 ();
 sg13g2_fill_1 FILLER_74_1719 ();
 sg13g2_fill_2 FILLER_74_1723 ();
 sg13g2_fill_1 FILLER_74_1725 ();
 sg13g2_fill_2 FILLER_74_1759 ();
 sg13g2_fill_1 FILLER_74_1761 ();
 sg13g2_fill_1 FILLER_74_1766 ();
 sg13g2_fill_1 FILLER_74_1776 ();
 sg13g2_fill_1 FILLER_74_1792 ();
 sg13g2_fill_2 FILLER_74_1816 ();
 sg13g2_decap_8 FILLER_74_1856 ();
 sg13g2_decap_8 FILLER_74_1863 ();
 sg13g2_decap_8 FILLER_74_1870 ();
 sg13g2_fill_2 FILLER_74_1877 ();
 sg13g2_decap_8 FILLER_74_1893 ();
 sg13g2_decap_4 FILLER_74_1900 ();
 sg13g2_fill_1 FILLER_74_1904 ();
 sg13g2_fill_1 FILLER_74_1909 ();
 sg13g2_fill_1 FILLER_74_1920 ();
 sg13g2_decap_4 FILLER_74_1953 ();
 sg13g2_decap_8 FILLER_74_1961 ();
 sg13g2_decap_8 FILLER_74_1978 ();
 sg13g2_fill_1 FILLER_74_1985 ();
 sg13g2_decap_8 FILLER_74_1996 ();
 sg13g2_fill_2 FILLER_74_2003 ();
 sg13g2_fill_2 FILLER_74_2009 ();
 sg13g2_fill_1 FILLER_74_2011 ();
 sg13g2_fill_2 FILLER_74_2038 ();
 sg13g2_fill_1 FILLER_74_2040 ();
 sg13g2_fill_2 FILLER_74_2080 ();
 sg13g2_fill_2 FILLER_74_2092 ();
 sg13g2_fill_1 FILLER_74_2094 ();
 sg13g2_fill_2 FILLER_74_2126 ();
 sg13g2_fill_2 FILLER_74_2132 ();
 sg13g2_fill_1 FILLER_74_2134 ();
 sg13g2_decap_8 FILLER_74_2175 ();
 sg13g2_decap_4 FILLER_74_2182 ();
 sg13g2_fill_1 FILLER_74_2203 ();
 sg13g2_fill_2 FILLER_74_2239 ();
 sg13g2_fill_1 FILLER_74_2266 ();
 sg13g2_fill_2 FILLER_74_2289 ();
 sg13g2_decap_8 FILLER_74_2295 ();
 sg13g2_fill_2 FILLER_74_2302 ();
 sg13g2_decap_4 FILLER_74_2323 ();
 sg13g2_fill_2 FILLER_74_2332 ();
 sg13g2_fill_1 FILLER_74_2366 ();
 sg13g2_fill_2 FILLER_74_2420 ();
 sg13g2_decap_8 FILLER_74_2432 ();
 sg13g2_decap_4 FILLER_74_2439 ();
 sg13g2_decap_4 FILLER_74_2455 ();
 sg13g2_fill_2 FILLER_74_2459 ();
 sg13g2_decap_4 FILLER_74_2491 ();
 sg13g2_fill_2 FILLER_74_2495 ();
 sg13g2_fill_1 FILLER_74_2523 ();
 sg13g2_fill_1 FILLER_74_2534 ();
 sg13g2_fill_2 FILLER_74_2539 ();
 sg13g2_decap_4 FILLER_74_2545 ();
 sg13g2_fill_2 FILLER_74_2549 ();
 sg13g2_decap_4 FILLER_74_2561 ();
 sg13g2_decap_4 FILLER_74_2571 ();
 sg13g2_fill_2 FILLER_74_2575 ();
 sg13g2_fill_2 FILLER_74_2591 ();
 sg13g2_fill_1 FILLER_74_2593 ();
 sg13g2_decap_8 FILLER_74_2606 ();
 sg13g2_decap_8 FILLER_74_2613 ();
 sg13g2_decap_8 FILLER_74_2620 ();
 sg13g2_decap_8 FILLER_74_2627 ();
 sg13g2_decap_8 FILLER_74_2634 ();
 sg13g2_decap_8 FILLER_74_2641 ();
 sg13g2_decap_8 FILLER_74_2648 ();
 sg13g2_decap_8 FILLER_74_2655 ();
 sg13g2_decap_8 FILLER_74_2662 ();
 sg13g2_fill_1 FILLER_74_2669 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_4 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_15 ();
 sg13g2_fill_2 FILLER_75_22 ();
 sg13g2_fill_1 FILLER_75_24 ();
 sg13g2_decap_8 FILLER_75_30 ();
 sg13g2_decap_8 FILLER_75_37 ();
 sg13g2_decap_8 FILLER_75_44 ();
 sg13g2_fill_2 FILLER_75_82 ();
 sg13g2_fill_1 FILLER_75_89 ();
 sg13g2_decap_4 FILLER_75_121 ();
 sg13g2_fill_1 FILLER_75_125 ();
 sg13g2_fill_2 FILLER_75_151 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_180 ();
 sg13g2_fill_2 FILLER_75_187 ();
 sg13g2_fill_1 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_230 ();
 sg13g2_decap_8 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_244 ();
 sg13g2_decap_8 FILLER_75_251 ();
 sg13g2_decap_8 FILLER_75_258 ();
 sg13g2_decap_4 FILLER_75_265 ();
 sg13g2_fill_2 FILLER_75_269 ();
 sg13g2_fill_1 FILLER_75_279 ();
 sg13g2_fill_2 FILLER_75_295 ();
 sg13g2_decap_8 FILLER_75_318 ();
 sg13g2_fill_2 FILLER_75_325 ();
 sg13g2_fill_1 FILLER_75_327 ();
 sg13g2_decap_8 FILLER_75_362 ();
 sg13g2_decap_4 FILLER_75_369 ();
 sg13g2_fill_1 FILLER_75_378 ();
 sg13g2_decap_4 FILLER_75_383 ();
 sg13g2_fill_1 FILLER_75_387 ();
 sg13g2_fill_2 FILLER_75_394 ();
 sg13g2_decap_8 FILLER_75_456 ();
 sg13g2_fill_2 FILLER_75_463 ();
 sg13g2_fill_2 FILLER_75_491 ();
 sg13g2_fill_1 FILLER_75_493 ();
 sg13g2_fill_2 FILLER_75_502 ();
 sg13g2_fill_1 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_510 ();
 sg13g2_fill_2 FILLER_75_517 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_decap_4 FILLER_75_530 ();
 sg13g2_fill_2 FILLER_75_534 ();
 sg13g2_fill_2 FILLER_75_546 ();
 sg13g2_fill_1 FILLER_75_548 ();
 sg13g2_fill_1 FILLER_75_566 ();
 sg13g2_fill_2 FILLER_75_601 ();
 sg13g2_fill_2 FILLER_75_613 ();
 sg13g2_fill_1 FILLER_75_622 ();
 sg13g2_fill_2 FILLER_75_663 ();
 sg13g2_decap_8 FILLER_75_701 ();
 sg13g2_decap_8 FILLER_75_708 ();
 sg13g2_fill_2 FILLER_75_715 ();
 sg13g2_fill_1 FILLER_75_717 ();
 sg13g2_fill_1 FILLER_75_722 ();
 sg13g2_fill_2 FILLER_75_762 ();
 sg13g2_fill_1 FILLER_75_764 ();
 sg13g2_decap_8 FILLER_75_795 ();
 sg13g2_fill_1 FILLER_75_802 ();
 sg13g2_fill_1 FILLER_75_835 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_fill_2 FILLER_75_847 ();
 sg13g2_fill_1 FILLER_75_857 ();
 sg13g2_decap_4 FILLER_75_906 ();
 sg13g2_decap_8 FILLER_75_914 ();
 sg13g2_decap_8 FILLER_75_921 ();
 sg13g2_fill_2 FILLER_75_928 ();
 sg13g2_decap_8 FILLER_75_935 ();
 sg13g2_decap_8 FILLER_75_942 ();
 sg13g2_decap_4 FILLER_75_949 ();
 sg13g2_fill_1 FILLER_75_963 ();
 sg13g2_decap_8 FILLER_75_974 ();
 sg13g2_fill_2 FILLER_75_981 ();
 sg13g2_fill_1 FILLER_75_983 ();
 sg13g2_decap_4 FILLER_75_1000 ();
 sg13g2_fill_2 FILLER_75_1004 ();
 sg13g2_decap_8 FILLER_75_1038 ();
 sg13g2_fill_2 FILLER_75_1045 ();
 sg13g2_fill_1 FILLER_75_1070 ();
 sg13g2_decap_8 FILLER_75_1097 ();
 sg13g2_decap_8 FILLER_75_1104 ();
 sg13g2_decap_4 FILLER_75_1111 ();
 sg13g2_fill_1 FILLER_75_1115 ();
 sg13g2_decap_4 FILLER_75_1136 ();
 sg13g2_fill_1 FILLER_75_1140 ();
 sg13g2_decap_8 FILLER_75_1145 ();
 sg13g2_decap_8 FILLER_75_1159 ();
 sg13g2_decap_8 FILLER_75_1166 ();
 sg13g2_decap_8 FILLER_75_1173 ();
 sg13g2_decap_8 FILLER_75_1180 ();
 sg13g2_decap_4 FILLER_75_1187 ();
 sg13g2_fill_1 FILLER_75_1191 ();
 sg13g2_fill_2 FILLER_75_1200 ();
 sg13g2_fill_1 FILLER_75_1202 ();
 sg13g2_fill_1 FILLER_75_1212 ();
 sg13g2_fill_1 FILLER_75_1223 ();
 sg13g2_fill_2 FILLER_75_1234 ();
 sg13g2_decap_4 FILLER_75_1240 ();
 sg13g2_fill_1 FILLER_75_1244 ();
 sg13g2_fill_1 FILLER_75_1286 ();
 sg13g2_decap_4 FILLER_75_1292 ();
 sg13g2_fill_1 FILLER_75_1296 ();
 sg13g2_decap_8 FILLER_75_1301 ();
 sg13g2_decap_4 FILLER_75_1308 ();
 sg13g2_fill_2 FILLER_75_1316 ();
 sg13g2_fill_2 FILLER_75_1321 ();
 sg13g2_fill_1 FILLER_75_1323 ();
 sg13g2_decap_4 FILLER_75_1339 ();
 sg13g2_fill_1 FILLER_75_1343 ();
 sg13g2_fill_2 FILLER_75_1348 ();
 sg13g2_fill_1 FILLER_75_1350 ();
 sg13g2_decap_4 FILLER_75_1355 ();
 sg13g2_fill_2 FILLER_75_1367 ();
 sg13g2_fill_2 FILLER_75_1386 ();
 sg13g2_decap_4 FILLER_75_1398 ();
 sg13g2_fill_2 FILLER_75_1406 ();
 sg13g2_decap_8 FILLER_75_1414 ();
 sg13g2_decap_4 FILLER_75_1421 ();
 sg13g2_fill_2 FILLER_75_1455 ();
 sg13g2_fill_2 FILLER_75_1460 ();
 sg13g2_fill_2 FILLER_75_1470 ();
 sg13g2_fill_1 FILLER_75_1516 ();
 sg13g2_fill_2 FILLER_75_1531 ();
 sg13g2_fill_1 FILLER_75_1533 ();
 sg13g2_decap_4 FILLER_75_1572 ();
 sg13g2_decap_8 FILLER_75_1582 ();
 sg13g2_decap_8 FILLER_75_1589 ();
 sg13g2_decap_4 FILLER_75_1596 ();
 sg13g2_fill_1 FILLER_75_1619 ();
 sg13g2_decap_8 FILLER_75_1624 ();
 sg13g2_fill_2 FILLER_75_1631 ();
 sg13g2_fill_2 FILLER_75_1638 ();
 sg13g2_fill_2 FILLER_75_1658 ();
 sg13g2_fill_1 FILLER_75_1660 ();
 sg13g2_fill_2 FILLER_75_1697 ();
 sg13g2_fill_1 FILLER_75_1699 ();
 sg13g2_decap_8 FILLER_75_1706 ();
 sg13g2_fill_1 FILLER_75_1713 ();
 sg13g2_fill_1 FILLER_75_1718 ();
 sg13g2_fill_2 FILLER_75_1725 ();
 sg13g2_decap_8 FILLER_75_1731 ();
 sg13g2_decap_4 FILLER_75_1738 ();
 sg13g2_fill_2 FILLER_75_1742 ();
 sg13g2_fill_2 FILLER_75_1759 ();
 sg13g2_decap_4 FILLER_75_1766 ();
 sg13g2_fill_2 FILLER_75_1784 ();
 sg13g2_decap_8 FILLER_75_1851 ();
 sg13g2_decap_8 FILLER_75_1858 ();
 sg13g2_decap_8 FILLER_75_1865 ();
 sg13g2_decap_8 FILLER_75_1872 ();
 sg13g2_decap_4 FILLER_75_1879 ();
 sg13g2_fill_2 FILLER_75_1883 ();
 sg13g2_fill_1 FILLER_75_1889 ();
 sg13g2_fill_2 FILLER_75_1959 ();
 sg13g2_fill_1 FILLER_75_1961 ();
 sg13g2_fill_2 FILLER_75_1967 ();
 sg13g2_fill_2 FILLER_75_1979 ();
 sg13g2_fill_1 FILLER_75_1981 ();
 sg13g2_decap_8 FILLER_75_1986 ();
 sg13g2_decap_8 FILLER_75_1993 ();
 sg13g2_decap_8 FILLER_75_2010 ();
 sg13g2_decap_8 FILLER_75_2017 ();
 sg13g2_fill_2 FILLER_75_2024 ();
 sg13g2_fill_1 FILLER_75_2026 ();
 sg13g2_fill_1 FILLER_75_2037 ();
 sg13g2_decap_4 FILLER_75_2042 ();
 sg13g2_decap_4 FILLER_75_2049 ();
 sg13g2_fill_2 FILLER_75_2062 ();
 sg13g2_fill_1 FILLER_75_2064 ();
 sg13g2_fill_2 FILLER_75_2069 ();
 sg13g2_fill_2 FILLER_75_2089 ();
 sg13g2_fill_1 FILLER_75_2095 ();
 sg13g2_fill_1 FILLER_75_2101 ();
 sg13g2_decap_8 FILLER_75_2120 ();
 sg13g2_fill_1 FILLER_75_2127 ();
 sg13g2_fill_1 FILLER_75_2141 ();
 sg13g2_fill_1 FILLER_75_2160 ();
 sg13g2_decap_4 FILLER_75_2171 ();
 sg13g2_decap_8 FILLER_75_2180 ();
 sg13g2_fill_2 FILLER_75_2187 ();
 sg13g2_fill_1 FILLER_75_2189 ();
 sg13g2_fill_1 FILLER_75_2195 ();
 sg13g2_fill_2 FILLER_75_2212 ();
 sg13g2_fill_1 FILLER_75_2214 ();
 sg13g2_fill_2 FILLER_75_2225 ();
 sg13g2_fill_2 FILLER_75_2263 ();
 sg13g2_decap_4 FILLER_75_2314 ();
 sg13g2_fill_2 FILLER_75_2318 ();
 sg13g2_fill_2 FILLER_75_2356 ();
 sg13g2_decap_4 FILLER_75_2368 ();
 sg13g2_fill_2 FILLER_75_2404 ();
 sg13g2_decap_4 FILLER_75_2410 ();
 sg13g2_fill_2 FILLER_75_2414 ();
 sg13g2_decap_8 FILLER_75_2442 ();
 sg13g2_decap_8 FILLER_75_2449 ();
 sg13g2_fill_2 FILLER_75_2468 ();
 sg13g2_decap_8 FILLER_75_2490 ();
 sg13g2_decap_4 FILLER_75_2511 ();
 sg13g2_fill_2 FILLER_75_2519 ();
 sg13g2_fill_1 FILLER_75_2521 ();
 sg13g2_decap_4 FILLER_75_2528 ();
 sg13g2_decap_8 FILLER_75_2546 ();
 sg13g2_decap_8 FILLER_75_2553 ();
 sg13g2_decap_4 FILLER_75_2560 ();
 sg13g2_fill_2 FILLER_75_2600 ();
 sg13g2_decap_8 FILLER_75_2606 ();
 sg13g2_decap_8 FILLER_75_2613 ();
 sg13g2_decap_8 FILLER_75_2620 ();
 sg13g2_decap_8 FILLER_75_2627 ();
 sg13g2_decap_8 FILLER_75_2634 ();
 sg13g2_decap_8 FILLER_75_2641 ();
 sg13g2_decap_8 FILLER_75_2648 ();
 sg13g2_decap_8 FILLER_75_2655 ();
 sg13g2_decap_8 FILLER_75_2662 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_fill_1 FILLER_76_7 ();
 sg13g2_fill_1 FILLER_76_83 ();
 sg13g2_fill_1 FILLER_76_89 ();
 sg13g2_fill_2 FILLER_76_95 ();
 sg13g2_fill_2 FILLER_76_101 ();
 sg13g2_decap_4 FILLER_76_115 ();
 sg13g2_fill_2 FILLER_76_150 ();
 sg13g2_fill_2 FILLER_76_167 ();
 sg13g2_fill_1 FILLER_76_175 ();
 sg13g2_decap_4 FILLER_76_229 ();
 sg13g2_fill_1 FILLER_76_233 ();
 sg13g2_decap_8 FILLER_76_253 ();
 sg13g2_decap_4 FILLER_76_260 ();
 sg13g2_fill_1 FILLER_76_264 ();
 sg13g2_fill_2 FILLER_76_285 ();
 sg13g2_fill_1 FILLER_76_287 ();
 sg13g2_fill_1 FILLER_76_296 ();
 sg13g2_decap_8 FILLER_76_318 ();
 sg13g2_decap_8 FILLER_76_325 ();
 sg13g2_decap_8 FILLER_76_332 ();
 sg13g2_decap_8 FILLER_76_343 ();
 sg13g2_decap_8 FILLER_76_350 ();
 sg13g2_decap_4 FILLER_76_357 ();
 sg13g2_fill_1 FILLER_76_402 ();
 sg13g2_fill_1 FILLER_76_407 ();
 sg13g2_decap_4 FILLER_76_413 ();
 sg13g2_fill_2 FILLER_76_417 ();
 sg13g2_fill_1 FILLER_76_423 ();
 sg13g2_fill_2 FILLER_76_428 ();
 sg13g2_fill_1 FILLER_76_434 ();
 sg13g2_fill_2 FILLER_76_439 ();
 sg13g2_fill_2 FILLER_76_445 ();
 sg13g2_fill_2 FILLER_76_451 ();
 sg13g2_fill_2 FILLER_76_462 ();
 sg13g2_fill_1 FILLER_76_468 ();
 sg13g2_fill_1 FILLER_76_473 ();
 sg13g2_fill_1 FILLER_76_480 ();
 sg13g2_fill_1 FILLER_76_499 ();
 sg13g2_decap_8 FILLER_76_508 ();
 sg13g2_decap_4 FILLER_76_515 ();
 sg13g2_fill_1 FILLER_76_523 ();
 sg13g2_decap_8 FILLER_76_534 ();
 sg13g2_decap_4 FILLER_76_541 ();
 sg13g2_fill_2 FILLER_76_545 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_fill_1 FILLER_76_564 ();
 sg13g2_fill_2 FILLER_76_581 ();
 sg13g2_fill_1 FILLER_76_589 ();
 sg13g2_fill_1 FILLER_76_600 ();
 sg13g2_fill_1 FILLER_76_606 ();
 sg13g2_fill_1 FILLER_76_612 ();
 sg13g2_fill_1 FILLER_76_628 ();
 sg13g2_fill_1 FILLER_76_659 ();
 sg13g2_fill_1 FILLER_76_688 ();
 sg13g2_decap_8 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_702 ();
 sg13g2_decap_8 FILLER_76_709 ();
 sg13g2_decap_8 FILLER_76_716 ();
 sg13g2_decap_4 FILLER_76_723 ();
 sg13g2_fill_1 FILLER_76_727 ();
 sg13g2_fill_2 FILLER_76_732 ();
 sg13g2_fill_1 FILLER_76_734 ();
 sg13g2_fill_2 FILLER_76_745 ();
 sg13g2_fill_2 FILLER_76_788 ();
 sg13g2_fill_2 FILLER_76_804 ();
 sg13g2_fill_1 FILLER_76_806 ();
 sg13g2_fill_2 FILLER_76_815 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_fill_2 FILLER_76_834 ();
 sg13g2_fill_1 FILLER_76_836 ();
 sg13g2_fill_2 FILLER_76_853 ();
 sg13g2_fill_1 FILLER_76_871 ();
 sg13g2_decap_8 FILLER_76_876 ();
 sg13g2_decap_8 FILLER_76_883 ();
 sg13g2_fill_1 FILLER_76_890 ();
 sg13g2_decap_8 FILLER_76_907 ();
 sg13g2_fill_1 FILLER_76_924 ();
 sg13g2_fill_1 FILLER_76_931 ();
 sg13g2_fill_1 FILLER_76_938 ();
 sg13g2_fill_1 FILLER_76_945 ();
 sg13g2_fill_2 FILLER_76_972 ();
 sg13g2_decap_4 FILLER_76_1000 ();
 sg13g2_decap_4 FILLER_76_1014 ();
 sg13g2_decap_8 FILLER_76_1022 ();
 sg13g2_decap_4 FILLER_76_1029 ();
 sg13g2_fill_2 FILLER_76_1033 ();
 sg13g2_fill_2 FILLER_76_1039 ();
 sg13g2_fill_1 FILLER_76_1041 ();
 sg13g2_decap_4 FILLER_76_1054 ();
 sg13g2_fill_1 FILLER_76_1058 ();
 sg13g2_decap_8 FILLER_76_1065 ();
 sg13g2_decap_4 FILLER_76_1072 ();
 sg13g2_fill_2 FILLER_76_1076 ();
 sg13g2_decap_8 FILLER_76_1088 ();
 sg13g2_decap_8 FILLER_76_1095 ();
 sg13g2_decap_8 FILLER_76_1102 ();
 sg13g2_fill_2 FILLER_76_1127 ();
 sg13g2_fill_1 FILLER_76_1129 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_fill_2 FILLER_76_1180 ();
 sg13g2_fill_1 FILLER_76_1182 ();
 sg13g2_fill_1 FILLER_76_1194 ();
 sg13g2_fill_2 FILLER_76_1211 ();
 sg13g2_fill_1 FILLER_76_1213 ();
 sg13g2_fill_2 FILLER_76_1247 ();
 sg13g2_fill_1 FILLER_76_1266 ();
 sg13g2_decap_4 FILLER_76_1302 ();
 sg13g2_fill_1 FILLER_76_1351 ();
 sg13g2_fill_2 FILLER_76_1360 ();
 sg13g2_fill_1 FILLER_76_1362 ();
 sg13g2_fill_1 FILLER_76_1396 ();
 sg13g2_decap_4 FILLER_76_1411 ();
 sg13g2_fill_1 FILLER_76_1415 ();
 sg13g2_fill_2 FILLER_76_1502 ();
 sg13g2_fill_2 FILLER_76_1513 ();
 sg13g2_fill_1 FILLER_76_1528 ();
 sg13g2_fill_1 FILLER_76_1535 ();
 sg13g2_fill_1 FILLER_76_1572 ();
 sg13g2_fill_1 FILLER_76_1585 ();
 sg13g2_fill_2 FILLER_76_1589 ();
 sg13g2_fill_1 FILLER_76_1599 ();
 sg13g2_fill_2 FILLER_76_1631 ();
 sg13g2_fill_1 FILLER_76_1662 ();
 sg13g2_fill_2 FILLER_76_1673 ();
 sg13g2_fill_1 FILLER_76_1675 ();
 sg13g2_fill_1 FILLER_76_1691 ();
 sg13g2_decap_4 FILLER_76_1698 ();
 sg13g2_fill_2 FILLER_76_1717 ();
 sg13g2_fill_1 FILLER_76_1719 ();
 sg13g2_fill_1 FILLER_76_1725 ();
 sg13g2_fill_2 FILLER_76_1741 ();
 sg13g2_fill_1 FILLER_76_1743 ();
 sg13g2_decap_8 FILLER_76_1773 ();
 sg13g2_decap_4 FILLER_76_1784 ();
 sg13g2_fill_1 FILLER_76_1851 ();
 sg13g2_fill_1 FILLER_76_1902 ();
 sg13g2_fill_1 FILLER_76_1907 ();
 sg13g2_fill_1 FILLER_76_1914 ();
 sg13g2_fill_1 FILLER_76_1921 ();
 sg13g2_fill_1 FILLER_76_1948 ();
 sg13g2_fill_1 FILLER_76_1975 ();
 sg13g2_decap_4 FILLER_76_2002 ();
 sg13g2_fill_2 FILLER_76_2006 ();
 sg13g2_decap_4 FILLER_76_2022 ();
 sg13g2_decap_4 FILLER_76_2036 ();
 sg13g2_decap_8 FILLER_76_2050 ();
 sg13g2_decap_4 FILLER_76_2057 ();
 sg13g2_fill_2 FILLER_76_2066 ();
 sg13g2_fill_1 FILLER_76_2068 ();
 sg13g2_fill_1 FILLER_76_2131 ();
 sg13g2_fill_1 FILLER_76_2136 ();
 sg13g2_fill_1 FILLER_76_2142 ();
 sg13g2_decap_8 FILLER_76_2169 ();
 sg13g2_decap_8 FILLER_76_2176 ();
 sg13g2_decap_8 FILLER_76_2183 ();
 sg13g2_decap_8 FILLER_76_2190 ();
 sg13g2_fill_1 FILLER_76_2217 ();
 sg13g2_decap_4 FILLER_76_2223 ();
 sg13g2_decap_4 FILLER_76_2247 ();
 sg13g2_fill_1 FILLER_76_2251 ();
 sg13g2_fill_2 FILLER_76_2292 ();
 sg13g2_fill_1 FILLER_76_2294 ();
 sg13g2_decap_4 FILLER_76_2299 ();
 sg13g2_fill_2 FILLER_76_2303 ();
 sg13g2_decap_4 FILLER_76_2310 ();
 sg13g2_fill_2 FILLER_76_2314 ();
 sg13g2_fill_1 FILLER_76_2326 ();
 sg13g2_fill_1 FILLER_76_2333 ();
 sg13g2_fill_2 FILLER_76_2338 ();
 sg13g2_fill_1 FILLER_76_2346 ();
 sg13g2_fill_2 FILLER_76_2357 ();
 sg13g2_decap_8 FILLER_76_2369 ();
 sg13g2_fill_1 FILLER_76_2386 ();
 sg13g2_decap_4 FILLER_76_2397 ();
 sg13g2_fill_2 FILLER_76_2401 ();
 sg13g2_decap_8 FILLER_76_2467 ();
 sg13g2_fill_2 FILLER_76_2503 ();
 sg13g2_fill_1 FILLER_76_2505 ();
 sg13g2_decap_4 FILLER_76_2516 ();
 sg13g2_decap_8 FILLER_76_2530 ();
 sg13g2_fill_2 FILLER_76_2563 ();
 sg13g2_fill_1 FILLER_76_2565 ();
 sg13g2_decap_8 FILLER_76_2582 ();
 sg13g2_fill_2 FILLER_76_2589 ();
 sg13g2_decap_8 FILLER_76_2617 ();
 sg13g2_decap_8 FILLER_76_2624 ();
 sg13g2_decap_8 FILLER_76_2631 ();
 sg13g2_decap_8 FILLER_76_2638 ();
 sg13g2_decap_8 FILLER_76_2645 ();
 sg13g2_decap_8 FILLER_76_2652 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_21 ();
 sg13g2_fill_1 FILLER_77_27 ();
 sg13g2_fill_2 FILLER_77_48 ();
 sg13g2_fill_1 FILLER_77_50 ();
 sg13g2_fill_1 FILLER_77_74 ();
 sg13g2_decap_8 FILLER_77_99 ();
 sg13g2_fill_1 FILLER_77_116 ();
 sg13g2_fill_1 FILLER_77_122 ();
 sg13g2_fill_1 FILLER_77_133 ();
 sg13g2_fill_1 FILLER_77_203 ();
 sg13g2_fill_1 FILLER_77_223 ();
 sg13g2_fill_2 FILLER_77_227 ();
 sg13g2_fill_2 FILLER_77_269 ();
 sg13g2_fill_2 FILLER_77_274 ();
 sg13g2_fill_1 FILLER_77_276 ();
 sg13g2_fill_1 FILLER_77_282 ();
 sg13g2_fill_1 FILLER_77_291 ();
 sg13g2_decap_4 FILLER_77_297 ();
 sg13g2_fill_2 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_324 ();
 sg13g2_decap_8 FILLER_77_331 ();
 sg13g2_decap_8 FILLER_77_338 ();
 sg13g2_decap_8 FILLER_77_345 ();
 sg13g2_decap_8 FILLER_77_352 ();
 sg13g2_fill_2 FILLER_77_359 ();
 sg13g2_fill_1 FILLER_77_369 ();
 sg13g2_fill_2 FILLER_77_395 ();
 sg13g2_decap_4 FILLER_77_437 ();
 sg13g2_fill_2 FILLER_77_441 ();
 sg13g2_fill_1 FILLER_77_474 ();
 sg13g2_decap_4 FILLER_77_519 ();
 sg13g2_fill_2 FILLER_77_523 ();
 sg13g2_decap_8 FILLER_77_555 ();
 sg13g2_fill_1 FILLER_77_609 ();
 sg13g2_fill_1 FILLER_77_632 ();
 sg13g2_fill_1 FILLER_77_637 ();
 sg13g2_fill_1 FILLER_77_643 ();
 sg13g2_fill_2 FILLER_77_649 ();
 sg13g2_fill_2 FILLER_77_683 ();
 sg13g2_fill_2 FILLER_77_693 ();
 sg13g2_fill_1 FILLER_77_700 ();
 sg13g2_fill_1 FILLER_77_706 ();
 sg13g2_decap_8 FILLER_77_711 ();
 sg13g2_decap_8 FILLER_77_718 ();
 sg13g2_decap_8 FILLER_77_725 ();
 sg13g2_decap_4 FILLER_77_732 ();
 sg13g2_fill_2 FILLER_77_740 ();
 sg13g2_fill_2 FILLER_77_752 ();
 sg13g2_fill_1 FILLER_77_754 ();
 sg13g2_fill_2 FILLER_77_765 ();
 sg13g2_fill_1 FILLER_77_767 ();
 sg13g2_decap_4 FILLER_77_778 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_858 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_decap_4 FILLER_77_908 ();
 sg13g2_fill_2 FILLER_77_912 ();
 sg13g2_fill_1 FILLER_77_957 ();
 sg13g2_fill_1 FILLER_77_977 ();
 sg13g2_fill_2 FILLER_77_1004 ();
 sg13g2_fill_2 FILLER_77_1016 ();
 sg13g2_fill_1 FILLER_77_1018 ();
 sg13g2_decap_4 FILLER_77_1055 ();
 sg13g2_fill_1 FILLER_77_1059 ();
 sg13g2_decap_4 FILLER_77_1096 ();
 sg13g2_fill_2 FILLER_77_1100 ();
 sg13g2_fill_2 FILLER_77_1122 ();
 sg13g2_decap_4 FILLER_77_1175 ();
 sg13g2_fill_2 FILLER_77_1223 ();
 sg13g2_fill_2 FILLER_77_1230 ();
 sg13g2_fill_2 FILLER_77_1261 ();
 sg13g2_fill_1 FILLER_77_1305 ();
 sg13g2_fill_2 FILLER_77_1311 ();
 sg13g2_fill_1 FILLER_77_1313 ();
 sg13g2_fill_1 FILLER_77_1323 ();
 sg13g2_fill_1 FILLER_77_1363 ();
 sg13g2_decap_4 FILLER_77_1391 ();
 sg13g2_fill_1 FILLER_77_1407 ();
 sg13g2_fill_1 FILLER_77_1475 ();
 sg13g2_fill_1 FILLER_77_1489 ();
 sg13g2_decap_4 FILLER_77_1544 ();
 sg13g2_fill_2 FILLER_77_1548 ();
 sg13g2_decap_4 FILLER_77_1554 ();
 sg13g2_fill_2 FILLER_77_1558 ();
 sg13g2_fill_2 FILLER_77_1566 ();
 sg13g2_fill_1 FILLER_77_1568 ();
 sg13g2_decap_4 FILLER_77_1575 ();
 sg13g2_fill_2 FILLER_77_1579 ();
 sg13g2_fill_1 FILLER_77_1585 ();
 sg13g2_fill_1 FILLER_77_1608 ();
 sg13g2_fill_2 FILLER_77_1630 ();
 sg13g2_fill_1 FILLER_77_1661 ();
 sg13g2_fill_1 FILLER_77_1709 ();
 sg13g2_fill_1 FILLER_77_1732 ();
 sg13g2_fill_1 FILLER_77_1738 ();
 sg13g2_fill_1 FILLER_77_1747 ();
 sg13g2_decap_4 FILLER_77_1772 ();
 sg13g2_fill_2 FILLER_77_1817 ();
 sg13g2_fill_2 FILLER_77_1824 ();
 sg13g2_fill_1 FILLER_77_1830 ();
 sg13g2_fill_2 FILLER_77_1841 ();
 sg13g2_decap_8 FILLER_77_1847 ();
 sg13g2_decap_8 FILLER_77_1854 ();
 sg13g2_fill_1 FILLER_77_1891 ();
 sg13g2_fill_2 FILLER_77_1928 ();
 sg13g2_fill_1 FILLER_77_1930 ();
 sg13g2_fill_1 FILLER_77_1957 ();
 sg13g2_fill_2 FILLER_77_1968 ();
 sg13g2_fill_2 FILLER_77_1976 ();
 sg13g2_fill_2 FILLER_77_2004 ();
 sg13g2_fill_1 FILLER_77_2006 ();
 sg13g2_fill_2 FILLER_77_2033 ();
 sg13g2_fill_1 FILLER_77_2035 ();
 sg13g2_fill_2 FILLER_77_2046 ();
 sg13g2_decap_8 FILLER_77_2074 ();
 sg13g2_fill_1 FILLER_77_2081 ();
 sg13g2_fill_1 FILLER_77_2086 ();
 sg13g2_fill_2 FILLER_77_2140 ();
 sg13g2_decap_8 FILLER_77_2168 ();
 sg13g2_fill_1 FILLER_77_2175 ();
 sg13g2_fill_2 FILLER_77_2202 ();
 sg13g2_fill_1 FILLER_77_2218 ();
 sg13g2_fill_1 FILLER_77_2245 ();
 sg13g2_fill_1 FILLER_77_2256 ();
 sg13g2_fill_1 FILLER_77_2267 ();
 sg13g2_fill_1 FILLER_77_2278 ();
 sg13g2_decap_4 FILLER_77_2289 ();
 sg13g2_decap_8 FILLER_77_2297 ();
 sg13g2_fill_2 FILLER_77_2304 ();
 sg13g2_decap_4 FILLER_77_2342 ();
 sg13g2_fill_1 FILLER_77_2346 ();
 sg13g2_decap_8 FILLER_77_2377 ();
 sg13g2_decap_8 FILLER_77_2384 ();
 sg13g2_decap_8 FILLER_77_2401 ();
 sg13g2_decap_4 FILLER_77_2408 ();
 sg13g2_fill_1 FILLER_77_2412 ();
 sg13g2_fill_2 FILLER_77_2439 ();
 sg13g2_fill_1 FILLER_77_2445 ();
 sg13g2_decap_8 FILLER_77_2472 ();
 sg13g2_decap_4 FILLER_77_2479 ();
 sg13g2_decap_4 FILLER_77_2549 ();
 sg13g2_fill_1 FILLER_77_2553 ();
 sg13g2_decap_4 FILLER_77_2577 ();
 sg13g2_fill_1 FILLER_77_2581 ();
 sg13g2_decap_8 FILLER_77_2608 ();
 sg13g2_decap_8 FILLER_77_2615 ();
 sg13g2_decap_8 FILLER_77_2622 ();
 sg13g2_decap_8 FILLER_77_2629 ();
 sg13g2_decap_8 FILLER_77_2636 ();
 sg13g2_decap_8 FILLER_77_2643 ();
 sg13g2_decap_8 FILLER_77_2650 ();
 sg13g2_decap_8 FILLER_77_2657 ();
 sg13g2_decap_4 FILLER_77_2664 ();
 sg13g2_fill_2 FILLER_77_2668 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_decap_4 FILLER_78_38 ();
 sg13g2_fill_2 FILLER_78_55 ();
 sg13g2_fill_1 FILLER_78_57 ();
 sg13g2_fill_2 FILLER_78_146 ();
 sg13g2_fill_1 FILLER_78_152 ();
 sg13g2_fill_2 FILLER_78_235 ();
 sg13g2_fill_1 FILLER_78_242 ();
 sg13g2_fill_1 FILLER_78_269 ();
 sg13g2_fill_1 FILLER_78_275 ();
 sg13g2_fill_1 FILLER_78_302 ();
 sg13g2_fill_1 FILLER_78_334 ();
 sg13g2_decap_8 FILLER_78_348 ();
 sg13g2_decap_8 FILLER_78_355 ();
 sg13g2_fill_1 FILLER_78_362 ();
 sg13g2_fill_2 FILLER_78_480 ();
 sg13g2_fill_1 FILLER_78_482 ();
 sg13g2_decap_8 FILLER_78_489 ();
 sg13g2_fill_1 FILLER_78_496 ();
 sg13g2_fill_1 FILLER_78_528 ();
 sg13g2_decap_8 FILLER_78_555 ();
 sg13g2_fill_1 FILLER_78_620 ();
 sg13g2_fill_2 FILLER_78_647 ();
 sg13g2_fill_2 FILLER_78_675 ();
 sg13g2_fill_1 FILLER_78_683 ();
 sg13g2_fill_2 FILLER_78_694 ();
 sg13g2_fill_1 FILLER_78_696 ();
 sg13g2_decap_4 FILLER_78_723 ();
 sg13g2_fill_2 FILLER_78_727 ();
 sg13g2_fill_2 FILLER_78_755 ();
 sg13g2_fill_1 FILLER_78_757 ();
 sg13g2_decap_4 FILLER_78_784 ();
 sg13g2_fill_2 FILLER_78_788 ();
 sg13g2_fill_1 FILLER_78_882 ();
 sg13g2_fill_1 FILLER_78_909 ();
 sg13g2_fill_2 FILLER_78_972 ();
 sg13g2_decap_4 FILLER_78_1014 ();
 sg13g2_fill_1 FILLER_78_1018 ();
 sg13g2_fill_1 FILLER_78_1075 ();
 sg13g2_fill_1 FILLER_78_1086 ();
 sg13g2_fill_2 FILLER_78_1113 ();
 sg13g2_fill_1 FILLER_78_1141 ();
 sg13g2_fill_2 FILLER_78_1152 ();
 sg13g2_decap_4 FILLER_78_1180 ();
 sg13g2_fill_1 FILLER_78_1184 ();
 sg13g2_fill_2 FILLER_78_1211 ();
 sg13g2_fill_1 FILLER_78_1213 ();
 sg13g2_fill_2 FILLER_78_1242 ();
 sg13g2_fill_2 FILLER_78_1278 ();
 sg13g2_fill_1 FILLER_78_1288 ();
 sg13g2_fill_1 FILLER_78_1294 ();
 sg13g2_fill_1 FILLER_78_1300 ();
 sg13g2_fill_1 FILLER_78_1306 ();
 sg13g2_fill_2 FILLER_78_1312 ();
 sg13g2_fill_1 FILLER_78_1319 ();
 sg13g2_fill_1 FILLER_78_1333 ();
 sg13g2_fill_1 FILLER_78_1339 ();
 sg13g2_fill_1 FILLER_78_1345 ();
 sg13g2_fill_1 FILLER_78_1361 ();
 sg13g2_fill_1 FILLER_78_1371 ();
 sg13g2_fill_1 FILLER_78_1376 ();
 sg13g2_fill_2 FILLER_78_1396 ();
 sg13g2_fill_2 FILLER_78_1403 ();
 sg13g2_decap_4 FILLER_78_1423 ();
 sg13g2_fill_1 FILLER_78_1427 ();
 sg13g2_fill_1 FILLER_78_1438 ();
 sg13g2_fill_1 FILLER_78_1444 ();
 sg13g2_fill_2 FILLER_78_1475 ();
 sg13g2_fill_1 FILLER_78_1477 ();
 sg13g2_fill_1 FILLER_78_1518 ();
 sg13g2_fill_2 FILLER_78_1529 ();
 sg13g2_fill_2 FILLER_78_1557 ();
 sg13g2_decap_8 FILLER_78_1563 ();
 sg13g2_decap_8 FILLER_78_1570 ();
 sg13g2_fill_2 FILLER_78_1577 ();
 sg13g2_decap_4 FILLER_78_1597 ();
 sg13g2_fill_2 FILLER_78_1606 ();
 sg13g2_fill_2 FILLER_78_1670 ();
 sg13g2_fill_1 FILLER_78_1680 ();
 sg13g2_fill_1 FILLER_78_1700 ();
 sg13g2_fill_1 FILLER_78_1706 ();
 sg13g2_fill_2 FILLER_78_1739 ();
 sg13g2_fill_1 FILLER_78_1746 ();
 sg13g2_fill_1 FILLER_78_1751 ();
 sg13g2_fill_2 FILLER_78_1802 ();
 sg13g2_fill_1 FILLER_78_1804 ();
 sg13g2_fill_1 FILLER_78_1818 ();
 sg13g2_decap_8 FILLER_78_1841 ();
 sg13g2_fill_1 FILLER_78_1848 ();
 sg13g2_decap_4 FILLER_78_1854 ();
 sg13g2_fill_1 FILLER_78_1910 ();
 sg13g2_fill_1 FILLER_78_1964 ();
 sg13g2_fill_1 FILLER_78_1991 ();
 sg13g2_fill_1 FILLER_78_2006 ();
 sg13g2_fill_1 FILLER_78_2056 ();
 sg13g2_fill_2 FILLER_78_2083 ();
 sg13g2_fill_2 FILLER_78_2095 ();
 sg13g2_decap_8 FILLER_78_2161 ();
 sg13g2_decap_8 FILLER_78_2168 ();
 sg13g2_decap_4 FILLER_78_2241 ();
 sg13g2_fill_2 FILLER_78_2245 ();
 sg13g2_fill_1 FILLER_78_2277 ();
 sg13g2_decap_4 FILLER_78_2282 ();
 sg13g2_fill_1 FILLER_78_2352 ();
 sg13g2_decap_8 FILLER_78_2383 ();
 sg13g2_fill_1 FILLER_78_2420 ();
 sg13g2_decap_8 FILLER_78_2425 ();
 sg13g2_fill_2 FILLER_78_2432 ();
 sg13g2_fill_1 FILLER_78_2434 ();
 sg13g2_decap_8 FILLER_78_2465 ();
 sg13g2_fill_1 FILLER_78_2472 ();
 sg13g2_fill_1 FILLER_78_2511 ();
 sg13g2_decap_4 FILLER_78_2538 ();
 sg13g2_decap_4 FILLER_78_2552 ();
 sg13g2_decap_8 FILLER_78_2582 ();
 sg13g2_fill_1 FILLER_78_2589 ();
 sg13g2_decap_8 FILLER_78_2594 ();
 sg13g2_decap_8 FILLER_78_2601 ();
 sg13g2_decap_8 FILLER_78_2608 ();
 sg13g2_decap_8 FILLER_78_2615 ();
 sg13g2_decap_8 FILLER_78_2622 ();
 sg13g2_decap_8 FILLER_78_2629 ();
 sg13g2_decap_8 FILLER_78_2636 ();
 sg13g2_decap_8 FILLER_78_2643 ();
 sg13g2_decap_8 FILLER_78_2650 ();
 sg13g2_decap_8 FILLER_78_2657 ();
 sg13g2_decap_4 FILLER_78_2664 ();
 sg13g2_fill_2 FILLER_78_2668 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_fill_1 FILLER_79_15 ();
 sg13g2_fill_1 FILLER_79_20 ();
 sg13g2_fill_1 FILLER_79_108 ();
 sg13g2_fill_2 FILLER_79_175 ();
 sg13g2_fill_1 FILLER_79_191 ();
 sg13g2_fill_1 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_79_203 ();
 sg13g2_fill_1 FILLER_79_211 ();
 sg13g2_fill_1 FILLER_79_253 ();
 sg13g2_fill_1 FILLER_79_268 ();
 sg13g2_fill_1 FILLER_79_277 ();
 sg13g2_fill_2 FILLER_79_287 ();
 sg13g2_fill_1 FILLER_79_289 ();
 sg13g2_decap_8 FILLER_79_325 ();
 sg13g2_decap_8 FILLER_79_332 ();
 sg13g2_fill_1 FILLER_79_339 ();
 sg13g2_decap_8 FILLER_79_353 ();
 sg13g2_decap_4 FILLER_79_360 ();
 sg13g2_fill_1 FILLER_79_364 ();
 sg13g2_fill_2 FILLER_79_399 ();
 sg13g2_decap_4 FILLER_79_431 ();
 sg13g2_fill_2 FILLER_79_439 ();
 sg13g2_fill_1 FILLER_79_441 ();
 sg13g2_fill_2 FILLER_79_446 ();
 sg13g2_fill_1 FILLER_79_448 ();
 sg13g2_fill_2 FILLER_79_453 ();
 sg13g2_fill_1 FILLER_79_455 ();
 sg13g2_decap_4 FILLER_79_504 ();
 sg13g2_fill_1 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_513 ();
 sg13g2_fill_1 FILLER_79_520 ();
 sg13g2_fill_1 FILLER_79_525 ();
 sg13g2_decap_4 FILLER_79_565 ();
 sg13g2_fill_1 FILLER_79_569 ();
 sg13g2_fill_1 FILLER_79_574 ();
 sg13g2_decap_4 FILLER_79_607 ();
 sg13g2_fill_2 FILLER_79_637 ();
 sg13g2_fill_2 FILLER_79_675 ();
 sg13g2_fill_1 FILLER_79_687 ();
 sg13g2_fill_2 FILLER_79_695 ();
 sg13g2_fill_1 FILLER_79_701 ();
 sg13g2_fill_2 FILLER_79_728 ();
 sg13g2_fill_1 FILLER_79_756 ();
 sg13g2_fill_2 FILLER_79_797 ();
 sg13g2_fill_1 FILLER_79_799 ();
 sg13g2_decap_8 FILLER_79_832 ();
 sg13g2_fill_1 FILLER_79_839 ();
 sg13g2_decap_8 FILLER_79_876 ();
 sg13g2_fill_2 FILLER_79_942 ();
 sg13g2_fill_1 FILLER_79_980 ();
 sg13g2_fill_2 FILLER_79_985 ();
 sg13g2_fill_2 FILLER_79_1075 ();
 sg13g2_fill_2 FILLER_79_1091 ();
 sg13g2_decap_8 FILLER_79_1097 ();
 sg13g2_fill_1 FILLER_79_1104 ();
 sg13g2_decap_4 FILLER_79_1131 ();
 sg13g2_fill_1 FILLER_79_1135 ();
 sg13g2_fill_1 FILLER_79_1162 ();
 sg13g2_decap_8 FILLER_79_1180 ();
 sg13g2_decap_4 FILLER_79_1187 ();
 sg13g2_decap_4 FILLER_79_1195 ();
 sg13g2_fill_1 FILLER_79_1199 ();
 sg13g2_fill_2 FILLER_79_1204 ();
 sg13g2_fill_1 FILLER_79_1206 ();
 sg13g2_fill_2 FILLER_79_1216 ();
 sg13g2_fill_2 FILLER_79_1222 ();
 sg13g2_fill_1 FILLER_79_1224 ();
 sg13g2_decap_4 FILLER_79_1230 ();
 sg13g2_fill_2 FILLER_79_1234 ();
 sg13g2_fill_2 FILLER_79_1252 ();
 sg13g2_fill_1 FILLER_79_1254 ();
 sg13g2_fill_1 FILLER_79_1259 ();
 sg13g2_fill_1 FILLER_79_1295 ();
 sg13g2_fill_1 FILLER_79_1309 ();
 sg13g2_fill_1 FILLER_79_1314 ();
 sg13g2_fill_1 FILLER_79_1319 ();
 sg13g2_fill_2 FILLER_79_1324 ();
 sg13g2_fill_2 FILLER_79_1336 ();
 sg13g2_fill_2 FILLER_79_1342 ();
 sg13g2_fill_1 FILLER_79_1344 ();
 sg13g2_fill_2 FILLER_79_1350 ();
 sg13g2_fill_1 FILLER_79_1352 ();
 sg13g2_fill_2 FILLER_79_1358 ();
 sg13g2_decap_8 FILLER_79_1390 ();
 sg13g2_fill_1 FILLER_79_1397 ();
 sg13g2_fill_1 FILLER_79_1424 ();
 sg13g2_fill_2 FILLER_79_1434 ();
 sg13g2_fill_1 FILLER_79_1440 ();
 sg13g2_fill_1 FILLER_79_1446 ();
 sg13g2_fill_1 FILLER_79_1452 ();
 sg13g2_fill_1 FILLER_79_1458 ();
 sg13g2_decap_8 FILLER_79_1464 ();
 sg13g2_decap_4 FILLER_79_1476 ();
 sg13g2_decap_4 FILLER_79_1492 ();
 sg13g2_decap_8 FILLER_79_1505 ();
 sg13g2_decap_8 FILLER_79_1512 ();
 sg13g2_decap_8 FILLER_79_1558 ();
 sg13g2_decap_8 FILLER_79_1565 ();
 sg13g2_decap_8 FILLER_79_1572 ();
 sg13g2_decap_8 FILLER_79_1579 ();
 sg13g2_decap_8 FILLER_79_1586 ();
 sg13g2_fill_2 FILLER_79_1593 ();
 sg13g2_fill_2 FILLER_79_1617 ();
 sg13g2_fill_1 FILLER_79_1628 ();
 sg13g2_decap_8 FILLER_79_1647 ();
 sg13g2_fill_2 FILLER_79_1695 ();
 sg13g2_decap_4 FILLER_79_1705 ();
 sg13g2_fill_1 FILLER_79_1717 ();
 sg13g2_fill_1 FILLER_79_1743 ();
 sg13g2_fill_2 FILLER_79_1772 ();
 sg13g2_fill_1 FILLER_79_1787 ();
 sg13g2_fill_1 FILLER_79_1798 ();
 sg13g2_decap_4 FILLER_79_1808 ();
 sg13g2_fill_2 FILLER_79_1812 ();
 sg13g2_fill_1 FILLER_79_1818 ();
 sg13g2_fill_1 FILLER_79_1824 ();
 sg13g2_fill_2 FILLER_79_1829 ();
 sg13g2_decap_8 FILLER_79_1857 ();
 sg13g2_decap_4 FILLER_79_1864 ();
 sg13g2_fill_1 FILLER_79_1868 ();
 sg13g2_decap_4 FILLER_79_1897 ();
 sg13g2_fill_1 FILLER_79_1901 ();
 sg13g2_decap_8 FILLER_79_1912 ();
 sg13g2_decap_4 FILLER_79_1945 ();
 sg13g2_fill_1 FILLER_79_1949 ();
 sg13g2_decap_4 FILLER_79_1986 ();
 sg13g2_decap_8 FILLER_79_2000 ();
 sg13g2_fill_1 FILLER_79_2007 ();
 sg13g2_decap_4 FILLER_79_2012 ();
 sg13g2_fill_2 FILLER_79_2056 ();
 sg13g2_decap_4 FILLER_79_2084 ();
 sg13g2_fill_1 FILLER_79_2088 ();
 sg13g2_fill_2 FILLER_79_2115 ();
 sg13g2_decap_8 FILLER_79_2151 ();
 sg13g2_decap_8 FILLER_79_2158 ();
 sg13g2_decap_4 FILLER_79_2165 ();
 sg13g2_decap_4 FILLER_79_2177 ();
 sg13g2_fill_1 FILLER_79_2181 ();
 sg13g2_fill_1 FILLER_79_2186 ();
 sg13g2_decap_4 FILLER_79_2191 ();
 sg13g2_decap_8 FILLER_79_2205 ();
 sg13g2_fill_2 FILLER_79_2212 ();
 sg13g2_decap_4 FILLER_79_2218 ();
 sg13g2_fill_1 FILLER_79_2222 ();
 sg13g2_decap_8 FILLER_79_2233 ();
 sg13g2_fill_2 FILLER_79_2240 ();
 sg13g2_decap_8 FILLER_79_2268 ();
 sg13g2_fill_2 FILLER_79_2275 ();
 sg13g2_decap_8 FILLER_79_2303 ();
 sg13g2_fill_1 FILLER_79_2350 ();
 sg13g2_decap_8 FILLER_79_2361 ();
 sg13g2_decap_8 FILLER_79_2407 ();
 sg13g2_decap_4 FILLER_79_2414 ();
 sg13g2_decap_4 FILLER_79_2432 ();
 sg13g2_fill_2 FILLER_79_2456 ();
 sg13g2_fill_1 FILLER_79_2458 ();
 sg13g2_fill_2 FILLER_79_2495 ();
 sg13g2_fill_2 FILLER_79_2501 ();
 sg13g2_fill_2 FILLER_79_2513 ();
 sg13g2_fill_1 FILLER_79_2515 ();
 sg13g2_decap_4 FILLER_79_2546 ();
 sg13g2_fill_2 FILLER_79_2550 ();
 sg13g2_decap_8 FILLER_79_2582 ();
 sg13g2_decap_8 FILLER_79_2589 ();
 sg13g2_decap_8 FILLER_79_2596 ();
 sg13g2_decap_8 FILLER_79_2603 ();
 sg13g2_decap_8 FILLER_79_2610 ();
 sg13g2_decap_8 FILLER_79_2617 ();
 sg13g2_decap_8 FILLER_79_2624 ();
 sg13g2_decap_8 FILLER_79_2631 ();
 sg13g2_decap_8 FILLER_79_2638 ();
 sg13g2_decap_8 FILLER_79_2645 ();
 sg13g2_decap_8 FILLER_79_2652 ();
 sg13g2_decap_8 FILLER_79_2659 ();
 sg13g2_decap_4 FILLER_79_2666 ();
 sg13g2_fill_2 FILLER_80_0 ();
 sg13g2_fill_2 FILLER_80_28 ();
 sg13g2_fill_1 FILLER_80_30 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_4 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_57 ();
 sg13g2_decap_8 FILLER_80_64 ();
 sg13g2_decap_4 FILLER_80_71 ();
 sg13g2_fill_1 FILLER_80_137 ();
 sg13g2_fill_1 FILLER_80_176 ();
 sg13g2_fill_2 FILLER_80_200 ();
 sg13g2_fill_1 FILLER_80_212 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_fill_2 FILLER_80_262 ();
 sg13g2_fill_1 FILLER_80_286 ();
 sg13g2_decap_8 FILLER_80_291 ();
 sg13g2_decap_4 FILLER_80_298 ();
 sg13g2_fill_1 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_307 ();
 sg13g2_decap_8 FILLER_80_314 ();
 sg13g2_decap_4 FILLER_80_321 ();
 sg13g2_fill_1 FILLER_80_325 ();
 sg13g2_decap_4 FILLER_80_331 ();
 sg13g2_fill_1 FILLER_80_335 ();
 sg13g2_fill_2 FILLER_80_355 ();
 sg13g2_fill_1 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_fill_1 FILLER_80_424 ();
 sg13g2_decap_8 FILLER_80_435 ();
 sg13g2_decap_8 FILLER_80_442 ();
 sg13g2_decap_8 FILLER_80_449 ();
 sg13g2_fill_2 FILLER_80_456 ();
 sg13g2_fill_1 FILLER_80_458 ();
 sg13g2_decap_8 FILLER_80_471 ();
 sg13g2_decap_8 FILLER_80_478 ();
 sg13g2_decap_4 FILLER_80_485 ();
 sg13g2_fill_2 FILLER_80_489 ();
 sg13g2_decap_8 FILLER_80_517 ();
 sg13g2_decap_8 FILLER_80_524 ();
 sg13g2_decap_4 FILLER_80_531 ();
 sg13g2_decap_8 FILLER_80_539 ();
 sg13g2_fill_2 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_552 ();
 sg13g2_decap_8 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_4 FILLER_80_573 ();
 sg13g2_decap_4 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_fill_2 FILLER_80_616 ();
 sg13g2_fill_1 FILLER_80_618 ();
 sg13g2_decap_4 FILLER_80_623 ();
 sg13g2_fill_1 FILLER_80_627 ();
 sg13g2_decap_8 FILLER_80_632 ();
 sg13g2_decap_8 FILLER_80_639 ();
 sg13g2_fill_2 FILLER_80_646 ();
 sg13g2_fill_1 FILLER_80_648 ();
 sg13g2_fill_2 FILLER_80_653 ();
 sg13g2_fill_1 FILLER_80_655 ();
 sg13g2_decap_4 FILLER_80_660 ();
 sg13g2_fill_2 FILLER_80_664 ();
 sg13g2_decap_4 FILLER_80_718 ();
 sg13g2_fill_1 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_740 ();
 sg13g2_decap_8 FILLER_80_747 ();
 sg13g2_decap_8 FILLER_80_754 ();
 sg13g2_decap_8 FILLER_80_761 ();
 sg13g2_decap_8 FILLER_80_772 ();
 sg13g2_decap_8 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_786 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_800 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_fill_2 FILLER_80_857 ();
 sg13g2_fill_1 FILLER_80_863 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_fill_2 FILLER_80_889 ();
 sg13g2_fill_1 FILLER_80_891 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_914 ();
 sg13g2_decap_4 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_929 ();
 sg13g2_decap_8 FILLER_80_936 ();
 sg13g2_decap_8 FILLER_80_943 ();
 sg13g2_fill_2 FILLER_80_950 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_fill_2 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_976 ();
 sg13g2_fill_2 FILLER_80_983 ();
 sg13g2_fill_1 FILLER_80_985 ();
 sg13g2_decap_4 FILLER_80_991 ();
 sg13g2_decap_4 FILLER_80_999 ();
 sg13g2_fill_1 FILLER_80_1003 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_fill_2 FILLER_80_1022 ();
 sg13g2_fill_1 FILLER_80_1024 ();
 sg13g2_decap_8 FILLER_80_1055 ();
 sg13g2_decap_8 FILLER_80_1062 ();
 sg13g2_decap_8 FILLER_80_1069 ();
 sg13g2_fill_2 FILLER_80_1080 ();
 sg13g2_fill_2 FILLER_80_1108 ();
 sg13g2_fill_1 FILLER_80_1110 ();
 sg13g2_fill_2 FILLER_80_1115 ();
 sg13g2_fill_2 FILLER_80_1120 ();
 sg13g2_fill_1 FILLER_80_1122 ();
 sg13g2_decap_8 FILLER_80_1127 ();
 sg13g2_decap_8 FILLER_80_1134 ();
 sg13g2_fill_2 FILLER_80_1141 ();
 sg13g2_decap_4 FILLER_80_1147 ();
 sg13g2_fill_2 FILLER_80_1151 ();
 sg13g2_decap_4 FILLER_80_1157 ();
 sg13g2_fill_1 FILLER_80_1161 ();
 sg13g2_decap_8 FILLER_80_1166 ();
 sg13g2_decap_8 FILLER_80_1173 ();
 sg13g2_decap_8 FILLER_80_1180 ();
 sg13g2_decap_8 FILLER_80_1187 ();
 sg13g2_fill_2 FILLER_80_1194 ();
 sg13g2_decap_8 FILLER_80_1226 ();
 sg13g2_decap_8 FILLER_80_1233 ();
 sg13g2_decap_8 FILLER_80_1240 ();
 sg13g2_decap_4 FILLER_80_1260 ();
 sg13g2_fill_2 FILLER_80_1264 ();
 sg13g2_decap_8 FILLER_80_1270 ();
 sg13g2_fill_1 FILLER_80_1277 ();
 sg13g2_decap_8 FILLER_80_1281 ();
 sg13g2_decap_8 FILLER_80_1288 ();
 sg13g2_decap_8 FILLER_80_1295 ();
 sg13g2_decap_8 FILLER_80_1302 ();
 sg13g2_decap_4 FILLER_80_1309 ();
 sg13g2_decap_8 FILLER_80_1317 ();
 sg13g2_decap_4 FILLER_80_1324 ();
 sg13g2_fill_2 FILLER_80_1332 ();
 sg13g2_decap_8 FILLER_80_1338 ();
 sg13g2_decap_8 FILLER_80_1345 ();
 sg13g2_decap_8 FILLER_80_1352 ();
 sg13g2_decap_8 FILLER_80_1359 ();
 sg13g2_decap_8 FILLER_80_1366 ();
 sg13g2_decap_8 FILLER_80_1373 ();
 sg13g2_decap_8 FILLER_80_1380 ();
 sg13g2_decap_8 FILLER_80_1387 ();
 sg13g2_decap_8 FILLER_80_1394 ();
 sg13g2_decap_8 FILLER_80_1401 ();
 sg13g2_decap_8 FILLER_80_1408 ();
 sg13g2_decap_8 FILLER_80_1415 ();
 sg13g2_decap_8 FILLER_80_1422 ();
 sg13g2_decap_8 FILLER_80_1429 ();
 sg13g2_decap_8 FILLER_80_1436 ();
 sg13g2_decap_4 FILLER_80_1451 ();
 sg13g2_decap_8 FILLER_80_1459 ();
 sg13g2_decap_8 FILLER_80_1466 ();
 sg13g2_decap_8 FILLER_80_1473 ();
 sg13g2_decap_8 FILLER_80_1480 ();
 sg13g2_decap_8 FILLER_80_1487 ();
 sg13g2_decap_8 FILLER_80_1494 ();
 sg13g2_decap_8 FILLER_80_1501 ();
 sg13g2_decap_8 FILLER_80_1508 ();
 sg13g2_decap_8 FILLER_80_1515 ();
 sg13g2_decap_8 FILLER_80_1522 ();
 sg13g2_fill_2 FILLER_80_1529 ();
 sg13g2_fill_1 FILLER_80_1531 ();
 sg13g2_decap_8 FILLER_80_1543 ();
 sg13g2_decap_8 FILLER_80_1550 ();
 sg13g2_decap_8 FILLER_80_1557 ();
 sg13g2_decap_8 FILLER_80_1564 ();
 sg13g2_decap_8 FILLER_80_1571 ();
 sg13g2_decap_8 FILLER_80_1578 ();
 sg13g2_decap_8 FILLER_80_1585 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_fill_2 FILLER_80_1620 ();
 sg13g2_fill_1 FILLER_80_1622 ();
 sg13g2_decap_8 FILLER_80_1636 ();
 sg13g2_decap_8 FILLER_80_1643 ();
 sg13g2_decap_8 FILLER_80_1650 ();
 sg13g2_decap_4 FILLER_80_1657 ();
 sg13g2_fill_2 FILLER_80_1661 ();
 sg13g2_decap_8 FILLER_80_1667 ();
 sg13g2_decap_8 FILLER_80_1674 ();
 sg13g2_decap_8 FILLER_80_1681 ();
 sg13g2_decap_8 FILLER_80_1688 ();
 sg13g2_decap_8 FILLER_80_1695 ();
 sg13g2_decap_4 FILLER_80_1702 ();
 sg13g2_fill_2 FILLER_80_1721 ();
 sg13g2_fill_1 FILLER_80_1723 ();
 sg13g2_decap_8 FILLER_80_1728 ();
 sg13g2_decap_8 FILLER_80_1735 ();
 sg13g2_decap_8 FILLER_80_1742 ();
 sg13g2_decap_8 FILLER_80_1749 ();
 sg13g2_decap_4 FILLER_80_1756 ();
 sg13g2_fill_2 FILLER_80_1760 ();
 sg13g2_decap_4 FILLER_80_1766 ();
 sg13g2_decap_8 FILLER_80_1774 ();
 sg13g2_decap_8 FILLER_80_1781 ();
 sg13g2_decap_8 FILLER_80_1788 ();
 sg13g2_decap_8 FILLER_80_1795 ();
 sg13g2_decap_8 FILLER_80_1802 ();
 sg13g2_decap_8 FILLER_80_1809 ();
 sg13g2_decap_8 FILLER_80_1816 ();
 sg13g2_decap_8 FILLER_80_1823 ();
 sg13g2_decap_8 FILLER_80_1830 ();
 sg13g2_decap_8 FILLER_80_1841 ();
 sg13g2_decap_8 FILLER_80_1848 ();
 sg13g2_decap_8 FILLER_80_1855 ();
 sg13g2_fill_2 FILLER_80_1862 ();
 sg13g2_fill_1 FILLER_80_1864 ();
 sg13g2_decap_8 FILLER_80_1869 ();
 sg13g2_decap_8 FILLER_80_1876 ();
 sg13g2_decap_8 FILLER_80_1883 ();
 sg13g2_decap_4 FILLER_80_1890 ();
 sg13g2_fill_2 FILLER_80_1894 ();
 sg13g2_decap_4 FILLER_80_1922 ();
 sg13g2_decap_4 FILLER_80_1930 ();
 sg13g2_decap_8 FILLER_80_1938 ();
 sg13g2_decap_8 FILLER_80_1945 ();
 sg13g2_decap_8 FILLER_80_1952 ();
 sg13g2_fill_2 FILLER_80_1959 ();
 sg13g2_decap_8 FILLER_80_1969 ();
 sg13g2_decap_8 FILLER_80_1976 ();
 sg13g2_decap_8 FILLER_80_1983 ();
 sg13g2_decap_8 FILLER_80_1990 ();
 sg13g2_decap_8 FILLER_80_1997 ();
 sg13g2_decap_4 FILLER_80_2004 ();
 sg13g2_decap_8 FILLER_80_2038 ();
 sg13g2_fill_1 FILLER_80_2045 ();
 sg13g2_decap_4 FILLER_80_2060 ();
 sg13g2_fill_1 FILLER_80_2064 ();
 sg13g2_decap_8 FILLER_80_2073 ();
 sg13g2_decap_8 FILLER_80_2080 ();
 sg13g2_decap_8 FILLER_80_2087 ();
 sg13g2_fill_1 FILLER_80_2094 ();
 sg13g2_decap_8 FILLER_80_2099 ();
 sg13g2_decap_8 FILLER_80_2106 ();
 sg13g2_decap_8 FILLER_80_2113 ();
 sg13g2_decap_8 FILLER_80_2120 ();
 sg13g2_decap_8 FILLER_80_2131 ();
 sg13g2_decap_8 FILLER_80_2138 ();
 sg13g2_decap_8 FILLER_80_2145 ();
 sg13g2_decap_8 FILLER_80_2152 ();
 sg13g2_decap_8 FILLER_80_2159 ();
 sg13g2_decap_8 FILLER_80_2166 ();
 sg13g2_decap_8 FILLER_80_2173 ();
 sg13g2_decap_8 FILLER_80_2180 ();
 sg13g2_decap_8 FILLER_80_2187 ();
 sg13g2_decap_8 FILLER_80_2194 ();
 sg13g2_decap_8 FILLER_80_2201 ();
 sg13g2_decap_8 FILLER_80_2208 ();
 sg13g2_fill_2 FILLER_80_2245 ();
 sg13g2_fill_1 FILLER_80_2247 ();
 sg13g2_fill_1 FILLER_80_2252 ();
 sg13g2_decap_8 FILLER_80_2266 ();
 sg13g2_decap_8 FILLER_80_2273 ();
 sg13g2_fill_2 FILLER_80_2280 ();
 sg13g2_fill_1 FILLER_80_2282 ();
 sg13g2_decap_8 FILLER_80_2287 ();
 sg13g2_decap_8 FILLER_80_2294 ();
 sg13g2_decap_8 FILLER_80_2301 ();
 sg13g2_decap_8 FILLER_80_2308 ();
 sg13g2_fill_2 FILLER_80_2315 ();
 sg13g2_decap_8 FILLER_80_2321 ();
 sg13g2_decap_4 FILLER_80_2328 ();
 sg13g2_fill_2 FILLER_80_2332 ();
 sg13g2_decap_8 FILLER_80_2364 ();
 sg13g2_decap_4 FILLER_80_2381 ();
 sg13g2_fill_2 FILLER_80_2385 ();
 sg13g2_decap_8 FILLER_80_2391 ();
 sg13g2_decap_8 FILLER_80_2398 ();
 sg13g2_decap_8 FILLER_80_2405 ();
 sg13g2_decap_8 FILLER_80_2412 ();
 sg13g2_decap_8 FILLER_80_2445 ();
 sg13g2_decap_8 FILLER_80_2452 ();
 sg13g2_decap_8 FILLER_80_2459 ();
 sg13g2_decap_8 FILLER_80_2466 ();
 sg13g2_decap_4 FILLER_80_2473 ();
 sg13g2_fill_1 FILLER_80_2477 ();
 sg13g2_decap_8 FILLER_80_2482 ();
 sg13g2_decap_8 FILLER_80_2499 ();
 sg13g2_decap_4 FILLER_80_2506 ();
 sg13g2_fill_2 FILLER_80_2510 ();
 sg13g2_decap_4 FILLER_80_2522 ();
 sg13g2_decap_8 FILLER_80_2534 ();
 sg13g2_decap_8 FILLER_80_2541 ();
 sg13g2_decap_8 FILLER_80_2548 ();
 sg13g2_decap_8 FILLER_80_2555 ();
 sg13g2_decap_8 FILLER_80_2566 ();
 sg13g2_decap_8 FILLER_80_2573 ();
 sg13g2_decap_8 FILLER_80_2580 ();
 sg13g2_decap_8 FILLER_80_2587 ();
 sg13g2_decap_8 FILLER_80_2594 ();
 sg13g2_decap_8 FILLER_80_2601 ();
 sg13g2_decap_8 FILLER_80_2608 ();
 sg13g2_decap_8 FILLER_80_2615 ();
 sg13g2_decap_8 FILLER_80_2622 ();
 sg13g2_decap_8 FILLER_80_2629 ();
 sg13g2_decap_8 FILLER_80_2636 ();
 sg13g2_decap_8 FILLER_80_2643 ();
 sg13g2_decap_8 FILLER_80_2650 ();
 sg13g2_decap_8 FILLER_80_2657 ();
 sg13g2_decap_4 FILLER_80_2664 ();
 sg13g2_fill_2 FILLER_80_2668 ();
endmodule
