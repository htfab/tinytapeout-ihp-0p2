module tt_um_vga_glyph_mode (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire clknet_0_clk;
 wire net101;
 wire \a[0] ;
 wire \a[1] ;
 wire \b[0] ;
 wire \b[1] ;
 wire \b[2] ;
 wire \b[3] ;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \div3.in[0] ;
 wire \div3.in[1] ;
 wire \div3.in[2] ;
 wire \div3.in[3] ;
 wire \div3.in[4] ;
 wire \div3.in[5] ;
 wire \div3.in[6] ;
 wire \div3.out[0] ;
 wire \div3.out[1] ;
 wire \div3.out[2] ;
 wire \div3.out[3] ;
 wire \div3.out[4] ;
 wire \div3.out[5] ;
 wire \g_x[0] ;
 wire \g_x[1] ;
 wire \g_x[2] ;
 wire hsync;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 sg13g2_inv_1 _1698_ (.Y(_0109_),
    .A(net1));
 sg13g2_buf_8 _1699_ (.A(\a[1] ),
    .X(_0120_));
 sg13g2_inv_2 _1700_ (.Y(_0131_),
    .A(_0120_));
 sg13g2_buf_8 _1701_ (.A(\a[0] ),
    .X(_0142_));
 sg13g2_inv_1 _1702_ (.Y(_0153_),
    .A(_0142_));
 sg13g2_buf_1 _1703_ (.A(_0153_),
    .X(_0164_));
 sg13g2_buf_1 _1704_ (.A(\g_x[1] ),
    .X(_0175_));
 sg13g2_buf_1 _1705_ (.A(\g_x[0] ),
    .X(_0186_));
 sg13g2_nand2_1 _1706_ (.Y(_0197_),
    .A(_0175_),
    .B(_0186_));
 sg13g2_inv_1 _1707_ (.Y(_0208_),
    .A(_0197_));
 sg13g2_nand2_1 _1708_ (.Y(_0219_),
    .A(_0208_),
    .B(\g_x[2] ));
 sg13g2_nor2_1 _1709_ (.A(net76),
    .B(_0219_),
    .Y(_0230_));
 sg13g2_inv_1 _1710_ (.Y(_0241_),
    .A(_0230_));
 sg13g2_nor2_2 _1711_ (.A(_0131_),
    .B(_0241_),
    .Y(_0252_));
 sg13g2_buf_1 _1712_ (.A(\b[3] ),
    .X(_0263_));
 sg13g2_inv_1 _1713_ (.Y(_0274_),
    .A(net83));
 sg13g2_buf_2 _1714_ (.A(\hvsync_gen.hpos[9] ),
    .X(_0285_));
 sg13g2_inv_1 _1715_ (.Y(_0296_),
    .A(_0285_));
 sg13g2_buf_1 _1716_ (.A(\b[0] ),
    .X(_0307_));
 sg13g2_inv_1 _1717_ (.Y(_0318_),
    .A(net82));
 sg13g2_buf_1 _1718_ (.A(\b[2] ),
    .X(_0329_));
 sg13g2_inv_1 _1719_ (.Y(_0340_),
    .A(net81));
 sg13g2_buf_8 _1720_ (.A(\b[1] ),
    .X(_0351_));
 sg13g2_inv_1 _1721_ (.Y(_0362_),
    .A(_0351_));
 sg13g2_nand3_1 _1722_ (.B(_0340_),
    .C(_0362_),
    .A(_0318_),
    .Y(_0373_));
 sg13g2_nor3_1 _1723_ (.A(_0274_),
    .B(_0296_),
    .C(_0373_),
    .Y(_0384_));
 sg13g2_nand2_2 _1724_ (.Y(_0395_),
    .A(_0252_),
    .B(_0384_));
 sg13g2_inv_1 _1725_ (.Y(_0406_),
    .A(_0395_));
 sg13g2_nor2_2 _1726_ (.A(_0109_),
    .B(_0406_),
    .Y(_0417_));
 sg13g2_inv_1 _1727_ (.Y(_0428_),
    .A(_0417_));
 sg13g2_nor2_1 _1728_ (.A(_0008_),
    .B(_0428_),
    .Y(_0439_));
 sg13g2_inv_1 _1729_ (.Y(_0450_),
    .A(\div3.in[4] ));
 sg13g2_inv_1 _1730_ (.Y(_0461_),
    .A(\div3.in[5] ));
 sg13g2_inv_1 _1731_ (.Y(_0472_),
    .A(\div3.in[3] ));
 sg13g2_buf_1 _1732_ (.A(\hvsync_gen.vpos[1] ),
    .X(_0483_));
 sg13g2_buf_2 _1733_ (.A(\hvsync_gen.vpos[0] ),
    .X(_0494_));
 sg13g2_nand2_1 _1734_ (.Y(_0505_),
    .A(net80),
    .B(_0494_));
 sg13g2_buf_1 _1735_ (.A(_0505_),
    .X(_0516_));
 sg13g2_nand2_1 _1736_ (.Y(_0527_),
    .A(\div3.in[1] ),
    .B(\div3.in[0] ));
 sg13g2_nor2_1 _1737_ (.A(_0516_),
    .B(_0527_),
    .Y(_0538_));
 sg13g2_nand2_1 _1738_ (.Y(_0549_),
    .A(_0538_),
    .B(\div3.in[2] ));
 sg13g2_nor2_1 _1739_ (.A(_0472_),
    .B(_0549_),
    .Y(_0560_));
 sg13g2_inv_1 _1740_ (.Y(_0571_),
    .A(_0560_));
 sg13g2_nor3_1 _1741_ (.A(_0450_),
    .B(_0461_),
    .C(_0571_),
    .Y(_0582_));
 sg13g2_xnor2_1 _1742_ (.Y(_0593_),
    .A(_0008_),
    .B(_0582_));
 sg13g2_nand4_1 _1743_ (.B(_0362_),
    .C(net83),
    .A(_0340_),
    .Y(_0604_),
    .D(_0285_));
 sg13g2_nor4_1 _1744_ (.A(net82),
    .B(_0131_),
    .C(_0604_),
    .D(_0241_),
    .Y(_0615_));
 sg13g2_nor2_2 _1745_ (.A(net80),
    .B(_0494_),
    .Y(_0626_));
 sg13g2_inv_2 _1746_ (.Y(_0637_),
    .A(_0626_));
 sg13g2_nor4_1 _1747_ (.A(\div3.in[4] ),
    .B(\div3.in[3] ),
    .C(_0527_),
    .D(_0637_),
    .Y(_0648_));
 sg13g2_inv_1 _1748_ (.Y(_0659_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_nor4_1 _1749_ (.A(\div3.in[2] ),
    .B(\div3.in[5] ),
    .C(\div3.in[6] ),
    .D(_0659_),
    .Y(_0670_));
 sg13g2_nand2_1 _1750_ (.Y(_0681_),
    .A(_0648_),
    .B(_0670_));
 sg13g2_nand2_1 _1751_ (.Y(_0692_),
    .A(_0681_),
    .B(net1));
 sg13g2_inv_1 _1752_ (.Y(_0703_),
    .A(_0692_));
 sg13g2_nand3_1 _1753_ (.B(_0615_),
    .C(_0703_),
    .A(_0593_),
    .Y(_0714_));
 sg13g2_nor2b_1 _1754_ (.A(_0439_),
    .B_N(_0714_),
    .Y(_0725_));
 sg13g2_buf_2 _1755_ (.A(_0725_),
    .X(_0736_));
 sg13g2_nand3_1 _1756_ (.B(\div3.in[4] ),
    .C(_0560_),
    .A(_0428_),
    .Y(_0747_));
 sg13g2_nor2_1 _1757_ (.A(_0703_),
    .B(_0417_),
    .Y(_0758_));
 sg13g2_a21o_1 _1758_ (.A2(_0582_),
    .A1(_0428_),
    .B1(_0758_),
    .X(_0769_));
 sg13g2_a21oi_2 _1759_ (.B1(_0769_),
    .Y(_0056_),
    .A2(_0747_),
    .A1(_0461_));
 sg13g2_inv_1 _1760_ (.Y(_0790_),
    .A(_0056_));
 sg13g2_nor2_1 _1761_ (.A(_0736_),
    .B(_0790_),
    .Y(_0005_));
 sg13g2_inv_1 _1762_ (.Y(_0811_),
    .A(\div3.in[1] ));
 sg13g2_inv_1 _1763_ (.Y(_0822_),
    .A(\div3.in[0] ));
 sg13g2_nand3_1 _1764_ (.B(_0659_),
    .C(net80),
    .A(_0822_),
    .Y(_0833_));
 sg13g2_nand2_1 _1765_ (.Y(_0844_),
    .A(\div3.in[5] ),
    .B(\div3.in[6] ));
 sg13g2_nor3_1 _1766_ (.A(_0450_),
    .B(_0472_),
    .C(_0844_),
    .Y(_0855_));
 sg13g2_o21ai_1 _1767_ (.B1(_0855_),
    .Y(_0865_),
    .A1(_0494_),
    .A2(_0527_));
 sg13g2_nor4_1 _1768_ (.A(_0811_),
    .B(\div3.in[2] ),
    .C(_0833_),
    .D(_0865_),
    .Y(_0007_));
 sg13g2_nand2_1 _1769_ (.Y(_0883_),
    .A(_0131_),
    .B(_0362_));
 sg13g2_inv_1 _1770_ (.Y(_0891_),
    .A(_0883_));
 sg13g2_nor2_1 _1771_ (.A(net82),
    .B(net83),
    .Y(_0892_));
 sg13g2_nand2_1 _1772_ (.Y(_0893_),
    .A(_0120_),
    .B(_0351_));
 sg13g2_o21ai_1 _1773_ (.B1(_0274_),
    .Y(_0894_),
    .A1(_0318_),
    .A2(_0893_));
 sg13g2_inv_1 _1774_ (.Y(_0895_),
    .A(_0009_));
 sg13g2_o21ai_1 _1775_ (.B1(_0285_),
    .Y(_0896_),
    .A1(net81),
    .A2(net83));
 sg13g2_a221oi_1 _1776_ (.B2(_0895_),
    .C1(_0896_),
    .B1(_0894_),
    .A1(_0891_),
    .Y(_0006_),
    .A2(_0892_));
 sg13g2_nand2b_1 _1777_ (.Y(_0897_),
    .B(_0560_),
    .A_N(_0014_));
 sg13g2_nor2_2 _1778_ (.A(_0395_),
    .B(_0692_),
    .Y(_0898_));
 sg13g2_inv_1 _1779_ (.Y(_0899_),
    .A(_0898_));
 sg13g2_a21oi_1 _1780_ (.A1(_0014_),
    .A2(_0571_),
    .Y(_0900_),
    .B1(_0899_));
 sg13g2_a22oi_1 _1781_ (.Y(_0901_),
    .B1(_0897_),
    .B2(_0900_),
    .A2(_0417_),
    .A1(\div3.in[4] ));
 sg13g2_buf_2 _1782_ (.A(_0901_),
    .X(_0902_));
 sg13g2_xnor2_1 _1783_ (.Y(_0903_),
    .A(_0012_),
    .B(_0538_));
 sg13g2_a22oi_1 _1784_ (.Y(_0904_),
    .B1(_0903_),
    .B2(_0898_),
    .A2(\div3.in[2] ),
    .A1(_0417_));
 sg13g2_inv_1 _1785_ (.Y(_0053_),
    .A(_0904_));
 sg13g2_nor2_1 _1786_ (.A(_0822_),
    .B(net75),
    .Y(_0905_));
 sg13g2_xor2_1 _1787_ (.B(_0905_),
    .A(_0011_),
    .X(_0906_));
 sg13g2_inv_1 _1788_ (.Y(_0907_),
    .A(_0906_));
 sg13g2_a22oi_1 _1789_ (.Y(_0908_),
    .B1(_0907_),
    .B2(_0898_),
    .A2(\div3.in[1] ),
    .A1(_0417_));
 sg13g2_xnor2_1 _1790_ (.Y(_0909_),
    .A(_0010_),
    .B(net75));
 sg13g2_inv_1 _1791_ (.Y(_0910_),
    .A(_0909_));
 sg13g2_a22oi_1 _1792_ (.Y(_0911_),
    .B1(_0910_),
    .B2(_0898_),
    .A2(\div3.in[0] ),
    .A1(_0417_));
 sg13g2_nor2_1 _1793_ (.A(_0908_),
    .B(_0911_),
    .Y(_0912_));
 sg13g2_nor2_1 _1794_ (.A(_0053_),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_inv_1 _1795_ (.Y(_0914_),
    .A(_0913_));
 sg13g2_xor2_1 _1796_ (.B(_0549_),
    .A(_0013_),
    .X(_0915_));
 sg13g2_a22oi_1 _1797_ (.Y(_0916_),
    .B1(_0915_),
    .B2(_0898_),
    .A2(\div3.in[3] ),
    .A1(_0417_));
 sg13g2_buf_1 _1798_ (.A(_0916_),
    .X(_0917_));
 sg13g2_nor2_1 _1799_ (.A(_0908_),
    .B(_0904_),
    .Y(_0918_));
 sg13g2_nor2_1 _1800_ (.A(_0917_),
    .B(_0918_),
    .Y(_0919_));
 sg13g2_nand2_1 _1801_ (.Y(_0920_),
    .A(_0908_),
    .B(_0911_));
 sg13g2_inv_1 _1802_ (.Y(_0052_),
    .A(_0908_));
 sg13g2_nor2_1 _1803_ (.A(_0052_),
    .B(_0053_),
    .Y(_0921_));
 sg13g2_a21oi_1 _1804_ (.A1(_0920_),
    .A2(_0053_),
    .Y(_0922_),
    .B1(_0921_));
 sg13g2_inv_1 _1805_ (.Y(_0923_),
    .A(_0922_));
 sg13g2_a22oi_1 _1806_ (.Y(_0924_),
    .B1(_0917_),
    .B2(_0923_),
    .A2(_0919_),
    .A1(_0914_));
 sg13g2_nor2_1 _1807_ (.A(_0902_),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_inv_1 _1808_ (.Y(_0055_),
    .A(_0902_));
 sg13g2_inv_2 _1809_ (.Y(_0054_),
    .A(_0917_));
 sg13g2_nor2_1 _1810_ (.A(_0054_),
    .B(_0918_),
    .Y(_0926_));
 sg13g2_a21o_1 _1811_ (.A2(_0904_),
    .A1(_0920_),
    .B1(_0912_),
    .X(_0927_));
 sg13g2_a22oi_1 _1812_ (.Y(_0928_),
    .B1(_0054_),
    .B2(_0927_),
    .A2(_0926_),
    .A1(_0914_));
 sg13g2_nor2_1 _1813_ (.A(net71),
    .B(_0928_),
    .Y(_0929_));
 sg13g2_o21ai_1 _1814_ (.B1(_0790_),
    .Y(_0930_),
    .A1(_0925_),
    .A2(_0929_));
 sg13g2_nand2_1 _1815_ (.Y(_0931_),
    .A(_0922_),
    .B(_0054_));
 sg13g2_o21ai_1 _1816_ (.B1(_0931_),
    .Y(_0932_),
    .A1(_0054_),
    .A2(_0927_));
 sg13g2_inv_1 _1817_ (.Y(_0933_),
    .A(_0932_));
 sg13g2_nor2_1 _1818_ (.A(net71),
    .B(_0790_),
    .Y(_0934_));
 sg13g2_inv_1 _1819_ (.Y(_0935_),
    .A(_0928_));
 sg13g2_nor2_1 _1820_ (.A(_0902_),
    .B(_0790_),
    .Y(_0936_));
 sg13g2_a22oi_1 _1821_ (.Y(_0937_),
    .B1(_0935_),
    .B2(_0936_),
    .A2(_0934_),
    .A1(_0933_));
 sg13g2_inv_1 _1822_ (.Y(_0938_),
    .A(_0736_));
 sg13g2_a21oi_1 _1823_ (.A1(_0930_),
    .A2(_0937_),
    .Y(_0939_),
    .B1(_0938_));
 sg13g2_nand2_1 _1824_ (.Y(_0940_),
    .A(_0932_),
    .B(net71));
 sg13g2_nor2_1 _1825_ (.A(_0736_),
    .B(_0056_),
    .Y(_0941_));
 sg13g2_inv_1 _1826_ (.Y(_0942_),
    .A(_0941_));
 sg13g2_a21oi_1 _1827_ (.A1(_0924_),
    .A2(_0902_),
    .Y(_0943_),
    .B1(_0942_));
 sg13g2_a21o_1 _1828_ (.A2(_0923_),
    .A1(net71),
    .B1(_0929_),
    .X(_0944_));
 sg13g2_a22oi_1 _1829_ (.Y(_0945_),
    .B1(_0005_),
    .B2(_0944_),
    .A2(_0943_),
    .A1(_0940_));
 sg13g2_nand2b_1 _1830_ (.Y(_0000_),
    .B(_0945_),
    .A_N(_0939_));
 sg13g2_inv_1 _1831_ (.Y(_0946_),
    .A(_0921_));
 sg13g2_nor2_1 _1832_ (.A(_0054_),
    .B(_0053_),
    .Y(_0947_));
 sg13g2_a21oi_1 _1833_ (.A1(_0946_),
    .A2(_0054_),
    .Y(_0948_),
    .B1(_0947_));
 sg13g2_nor2b_1 _1834_ (.A(_0948_),
    .B_N(_0934_),
    .Y(_0949_));
 sg13g2_nor2_1 _1835_ (.A(_0921_),
    .B(_0902_),
    .Y(_0950_));
 sg13g2_nand2b_1 _1836_ (.Y(_0951_),
    .B(_0950_),
    .A_N(_0919_));
 sg13g2_nor2_1 _1837_ (.A(_0917_),
    .B(_0904_),
    .Y(_0952_));
 sg13g2_nor2_1 _1838_ (.A(_0952_),
    .B(net71),
    .Y(_0953_));
 sg13g2_inv_1 _1839_ (.Y(_0954_),
    .A(_0953_));
 sg13g2_nor2_1 _1840_ (.A(_0926_),
    .B(_0954_),
    .Y(_0955_));
 sg13g2_nor2_1 _1841_ (.A(_0056_),
    .B(_0955_),
    .Y(_0956_));
 sg13g2_inv_1 _1842_ (.Y(_0957_),
    .A(_0952_));
 sg13g2_a21oi_1 _1843_ (.A1(net71),
    .A2(_0957_),
    .Y(_0958_),
    .B1(_0790_));
 sg13g2_a221oi_1 _1844_ (.B2(_0956_),
    .C1(_0958_),
    .B1(_0951_),
    .A1(_0056_),
    .Y(_0959_),
    .A2(_0926_));
 sg13g2_o21ai_1 _1845_ (.B1(_0736_),
    .Y(_0960_),
    .A1(_0949_),
    .A2(_0959_));
 sg13g2_nand2_1 _1846_ (.Y(_0961_),
    .A(_0948_),
    .B(net71));
 sg13g2_o21ai_1 _1847_ (.B1(_0902_),
    .Y(_0962_),
    .A1(_0921_),
    .A2(_0919_));
 sg13g2_nand3_1 _1848_ (.B(_0941_),
    .C(_0962_),
    .A(_0961_),
    .Y(_0963_));
 sg13g2_o21ai_1 _1849_ (.B1(_0005_),
    .Y(_0964_),
    .A1(_0950_),
    .A2(_0955_));
 sg13g2_nand3_1 _1850_ (.B(_0963_),
    .C(_0964_),
    .A(_0960_),
    .Y(_0001_));
 sg13g2_a21oi_1 _1851_ (.A1(net71),
    .A2(_0054_),
    .Y(_0965_),
    .B1(_0056_));
 sg13g2_inv_1 _1852_ (.Y(_0966_),
    .A(_0947_));
 sg13g2_a22oi_1 _1853_ (.Y(_0967_),
    .B1(_0966_),
    .B2(_0958_),
    .A2(_0954_),
    .A1(_0965_));
 sg13g2_nand2_1 _1854_ (.Y(_0968_),
    .A(_0055_),
    .B(_0966_));
 sg13g2_a21oi_1 _1855_ (.A1(_0902_),
    .A2(_0917_),
    .Y(_0969_),
    .B1(_0056_));
 sg13g2_a22oi_1 _1856_ (.Y(_0970_),
    .B1(_0968_),
    .B2(_0969_),
    .A2(_0957_),
    .A1(_0934_));
 sg13g2_nor2_1 _1857_ (.A(_0736_),
    .B(_0970_),
    .Y(_0971_));
 sg13g2_a21oi_1 _1858_ (.A1(_0736_),
    .A2(_0967_),
    .Y(_0002_),
    .B1(_0971_));
 sg13g2_inv_1 _1859_ (.Y(_0972_),
    .A(_0936_));
 sg13g2_nand2_1 _1860_ (.Y(_0973_),
    .A(_0972_),
    .B(_0736_));
 sg13g2_nand2_1 _1861_ (.Y(_0974_),
    .A(_0969_),
    .B(_0938_));
 sg13g2_o21ai_1 _1862_ (.B1(_0974_),
    .Y(_0003_),
    .A1(_0965_),
    .A2(_0973_));
 sg13g2_a21oi_1 _1863_ (.A1(_0972_),
    .A2(_0736_),
    .Y(_0004_),
    .B1(_0005_));
 sg13g2_inv_1 _1864_ (.Y(_0975_),
    .A(_0494_));
 sg13g2_buf_1 _1865_ (.A(_0428_),
    .X(_0976_));
 sg13g2_nand2_1 _1866_ (.Y(_0977_),
    .A(_0898_),
    .B(_0026_));
 sg13g2_o21ai_1 _1867_ (.B1(_0977_),
    .Y(_0049_),
    .A1(_0975_),
    .A2(net72));
 sg13g2_inv_2 _1868_ (.Y(_0978_),
    .A(net80));
 sg13g2_nand2_1 _1869_ (.Y(_0979_),
    .A(_0637_),
    .B(net75));
 sg13g2_inv_1 _1870_ (.Y(_0980_),
    .A(_0979_));
 sg13g2_o21ai_1 _1871_ (.B1(net1),
    .Y(_0981_),
    .A1(_0980_),
    .A2(_0395_));
 sg13g2_a21oi_1 _1872_ (.A1(_0978_),
    .A2(_0395_),
    .Y(_0050_),
    .B1(_0981_));
 sg13g2_inv_1 _1873_ (.Y(_0051_),
    .A(_0911_));
 sg13g2_inv_1 _1874_ (.Y(_0982_),
    .A(\div3.in[6] ));
 sg13g2_o21ai_1 _1875_ (.B1(_0714_),
    .Y(_0057_),
    .A1(_0982_),
    .A2(net72));
 sg13g2_nor2_1 _1876_ (.A(_0844_),
    .B(_0747_),
    .Y(_0983_));
 sg13g2_xnor2_1 _1877_ (.Y(_0984_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_0983_));
 sg13g2_nor2_1 _1878_ (.A(_0758_),
    .B(_0984_),
    .Y(_0058_));
 sg13g2_nand2_1 _1879_ (.Y(_0985_),
    .A(net1),
    .B(_0027_));
 sg13g2_inv_1 _1880_ (.Y(_0029_),
    .A(_0985_));
 sg13g2_buf_1 _1881_ (.A(_0109_),
    .X(_0986_));
 sg13g2_nor2_1 _1882_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_0987_));
 sg13g2_nand2_1 _1883_ (.Y(_0988_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_inv_1 _1884_ (.Y(_0989_),
    .A(_0988_));
 sg13g2_nor3_1 _1885_ (.A(net79),
    .B(_0987_),
    .C(_0989_),
    .Y(_0030_));
 sg13g2_nor2_1 _1886_ (.A(\counter[2] ),
    .B(_0989_),
    .Y(_0990_));
 sg13g2_nand2_1 _1887_ (.Y(_0991_),
    .A(_0989_),
    .B(\counter[2] ));
 sg13g2_inv_1 _1888_ (.Y(_0992_),
    .A(_0991_));
 sg13g2_nor3_1 _1889_ (.A(net79),
    .B(_0990_),
    .C(_0992_),
    .Y(_0031_));
 sg13g2_inv_1 _1890_ (.Y(_0993_),
    .A(\counter[3] ));
 sg13g2_nor2_1 _1891_ (.A(_0993_),
    .B(_0991_),
    .Y(_0994_));
 sg13g2_nor2_1 _1892_ (.A(\counter[3] ),
    .B(_0992_),
    .Y(_0995_));
 sg13g2_nor3_1 _1893_ (.A(net79),
    .B(_0994_),
    .C(_0995_),
    .Y(_0032_));
 sg13g2_nor2_1 _1894_ (.A(\counter[4] ),
    .B(_0994_),
    .Y(_0996_));
 sg13g2_nand2_1 _1895_ (.Y(_0997_),
    .A(_0994_),
    .B(\counter[4] ));
 sg13g2_inv_1 _1896_ (.Y(_0998_),
    .A(_0997_));
 sg13g2_nor3_1 _1897_ (.A(net79),
    .B(_0996_),
    .C(_0998_),
    .Y(_0033_));
 sg13g2_nor2_1 _1898_ (.A(\counter[5] ),
    .B(_0998_),
    .Y(_0999_));
 sg13g2_nand2_1 _1899_ (.Y(_1000_),
    .A(_0998_),
    .B(\counter[5] ));
 sg13g2_inv_1 _1900_ (.Y(_1001_),
    .A(_1000_));
 sg13g2_nor3_1 _1901_ (.A(net79),
    .B(_0999_),
    .C(_1001_),
    .Y(_0034_));
 sg13g2_nor2_1 _1902_ (.A(\counter[6] ),
    .B(_1001_),
    .Y(_1002_));
 sg13g2_nand2_1 _1903_ (.Y(_1003_),
    .A(_1001_),
    .B(\counter[6] ));
 sg13g2_inv_1 _1904_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_nor3_1 _1905_ (.A(net79),
    .B(_1002_),
    .C(_1004_),
    .Y(_0035_));
 sg13g2_nor2_1 _1906_ (.A(\counter[7] ),
    .B(_1004_),
    .Y(_1005_));
 sg13g2_nand2_1 _1907_ (.Y(_1006_),
    .A(_1004_),
    .B(\counter[7] ));
 sg13g2_inv_1 _1908_ (.Y(_1007_),
    .A(_1006_));
 sg13g2_nor3_1 _1909_ (.A(net79),
    .B(_1005_),
    .C(_1007_),
    .Y(_0036_));
 sg13g2_inv_1 _1910_ (.Y(_1008_),
    .A(\counter[8] ));
 sg13g2_nor2_1 _1911_ (.A(_1008_),
    .B(_1006_),
    .Y(_1009_));
 sg13g2_nor2_1 _1912_ (.A(\counter[8] ),
    .B(_1007_),
    .Y(_1010_));
 sg13g2_nor3_1 _1913_ (.A(net79),
    .B(_1009_),
    .C(_1010_),
    .Y(_0037_));
 sg13g2_nor2_1 _1914_ (.A(\counter[9] ),
    .B(_1009_),
    .Y(_1011_));
 sg13g2_a21oi_1 _1915_ (.A1(_1009_),
    .A2(\counter[9] ),
    .Y(_1012_),
    .B1(_0109_));
 sg13g2_nor2b_1 _1916_ (.A(_1011_),
    .B_N(_1012_),
    .Y(_0038_));
 sg13g2_nor2b_1 _1917_ (.A(net72),
    .B_N(_0028_),
    .Y(_0039_));
 sg13g2_nor2_1 _1918_ (.A(_0175_),
    .B(_0186_),
    .Y(_1013_));
 sg13g2_nor3_1 _1919_ (.A(_0208_),
    .B(_1013_),
    .C(net72),
    .Y(_0040_));
 sg13g2_inv_1 _1920_ (.Y(_1014_),
    .A(_0219_));
 sg13g2_nor2_1 _1921_ (.A(\g_x[2] ),
    .B(_0208_),
    .Y(_1015_));
 sg13g2_nor3_1 _1922_ (.A(_1014_),
    .B(_1015_),
    .C(net72),
    .Y(_0041_));
 sg13g2_buf_1 _1923_ (.A(_0142_),
    .X(_1016_));
 sg13g2_nor2_1 _1924_ (.A(net78),
    .B(_1014_),
    .Y(_1017_));
 sg13g2_nor3_1 _1925_ (.A(_0986_),
    .B(_0230_),
    .C(_1017_),
    .Y(_0042_));
 sg13g2_buf_1 _1926_ (.A(_0120_),
    .X(_1018_));
 sg13g2_nor2_1 _1927_ (.A(_1018_),
    .B(_0230_),
    .Y(_1019_));
 sg13g2_nor3_1 _1928_ (.A(_0986_),
    .B(_1019_),
    .C(_0252_),
    .Y(_0043_));
 sg13g2_nor2_1 _1929_ (.A(net82),
    .B(_0252_),
    .Y(_1020_));
 sg13g2_nand2_1 _1930_ (.Y(_1021_),
    .A(_0252_),
    .B(net82));
 sg13g2_inv_1 _1931_ (.Y(_1022_),
    .A(_1021_));
 sg13g2_nor3_1 _1932_ (.A(_1020_),
    .B(_1022_),
    .C(_0976_),
    .Y(_0044_));
 sg13g2_nor2_1 _1933_ (.A(_0351_),
    .B(_1022_),
    .Y(_1023_));
 sg13g2_nor2_1 _1934_ (.A(_0362_),
    .B(_1021_),
    .Y(_1024_));
 sg13g2_nor3_1 _1935_ (.A(_1023_),
    .B(_1024_),
    .C(_0976_),
    .Y(_0045_));
 sg13g2_nor2_1 _1936_ (.A(net81),
    .B(_1024_),
    .Y(_1025_));
 sg13g2_nand2_1 _1937_ (.Y(_1026_),
    .A(_1024_),
    .B(net81));
 sg13g2_inv_1 _1938_ (.Y(_1027_),
    .A(_1026_));
 sg13g2_nor3_1 _1939_ (.A(net72),
    .B(_1025_),
    .C(_1027_),
    .Y(_0046_));
 sg13g2_nor2_1 _1940_ (.A(_0274_),
    .B(_1026_),
    .Y(_1028_));
 sg13g2_nor2_1 _1941_ (.A(net83),
    .B(_1027_),
    .Y(_1029_));
 sg13g2_nor3_1 _1942_ (.A(net72),
    .B(_1028_),
    .C(_1029_),
    .Y(_0047_));
 sg13g2_xnor2_1 _1943_ (.Y(_1030_),
    .A(_0285_),
    .B(_1028_));
 sg13g2_nor2_1 _1944_ (.A(net72),
    .B(_1030_),
    .Y(_0048_));
 sg13g2_buf_2 _1945_ (.A(\div3.out[0] ),
    .X(_1031_));
 sg13g2_xor2_1 _1946_ (.B(_1031_),
    .A(\div3.in[0] ),
    .X(_1032_));
 sg13g2_inv_1 _1947_ (.Y(_1033_),
    .A(_1032_));
 sg13g2_xor2_1 _1948_ (.B(\div3.out[1] ),
    .A(\div3.in[1] ),
    .X(_1034_));
 sg13g2_inv_1 _1949_ (.Y(_1035_),
    .A(_1034_));
 sg13g2_nor2_1 _1950_ (.A(_1033_),
    .B(_1035_),
    .Y(_1036_));
 sg13g2_buf_1 _1951_ (.A(_1036_),
    .X(_1037_));
 sg13g2_xor2_1 _1952_ (.B(_1031_),
    .A(net82),
    .X(_1038_));
 sg13g2_inv_1 _1953_ (.Y(_1039_),
    .A(_1038_));
 sg13g2_xnor2_1 _1954_ (.Y(_1040_),
    .A(_0142_),
    .B(\b[0] ));
 sg13g2_xnor2_1 _1955_ (.Y(_1041_),
    .A(_0329_),
    .B(net83));
 sg13g2_xnor2_1 _1956_ (.Y(_1042_),
    .A(_1040_),
    .B(_1041_));
 sg13g2_xnor2_1 _1957_ (.Y(_1043_),
    .A(_0120_),
    .B(_0351_));
 sg13g2_xnor2_1 _1958_ (.Y(_1044_),
    .A(_0895_),
    .B(_1043_));
 sg13g2_nand2_2 _1959_ (.Y(_1045_),
    .A(_1042_),
    .B(_1044_));
 sg13g2_xor2_1 _1960_ (.B(net83),
    .A(net81),
    .X(_1046_));
 sg13g2_nand2_1 _1961_ (.Y(_1047_),
    .A(_1046_),
    .B(_1040_));
 sg13g2_xor2_1 _1962_ (.B(net82),
    .A(_0142_),
    .X(_1048_));
 sg13g2_nand2_1 _1963_ (.Y(_1049_),
    .A(_1048_),
    .B(_1041_));
 sg13g2_nand2_1 _1964_ (.Y(_1050_),
    .A(_1047_),
    .B(_1049_));
 sg13g2_nand2_1 _1965_ (.Y(_1051_),
    .A(_1043_),
    .B(_0009_));
 sg13g2_nand3_1 _1966_ (.B(_0895_),
    .C(_0893_),
    .A(_0883_),
    .Y(_1052_));
 sg13g2_nand2_1 _1967_ (.Y(_1053_),
    .A(_1051_),
    .B(_1052_));
 sg13g2_nand2_2 _1968_ (.Y(_1054_),
    .A(_1050_),
    .B(_1053_));
 sg13g2_nand2_1 _1969_ (.Y(_1055_),
    .A(_1045_),
    .B(_1054_));
 sg13g2_nand2b_1 _1970_ (.Y(_1056_),
    .B(net73),
    .A_N(_0015_));
 sg13g2_inv_1 _1971_ (.Y(_1057_),
    .A(_0016_));
 sg13g2_nand3_1 _1972_ (.B(_1054_),
    .C(_1057_),
    .A(_1045_),
    .Y(_1058_));
 sg13g2_nand2_1 _1973_ (.Y(_1059_),
    .A(_1056_),
    .B(_1058_));
 sg13g2_nand2_1 _1974_ (.Y(_1060_),
    .A(_0285_),
    .B(\div3.out[2] ));
 sg13g2_nor2_1 _1975_ (.A(_0285_),
    .B(\div3.out[2] ),
    .Y(_1061_));
 sg13g2_a21oi_1 _1976_ (.A1(_1059_),
    .A2(_1060_),
    .Y(_1062_),
    .B1(_1061_));
 sg13g2_nand2_1 _1977_ (.Y(_1063_),
    .A(net73),
    .B(_1057_));
 sg13g2_inv_1 _1978_ (.Y(_1064_),
    .A(_0019_));
 sg13g2_nand3_1 _1979_ (.B(_1054_),
    .C(_1064_),
    .A(_1045_),
    .Y(_1065_));
 sg13g2_nand2_1 _1980_ (.Y(_1066_),
    .A(_1063_),
    .B(_1065_));
 sg13g2_nor2_1 _1981_ (.A(_0120_),
    .B(\div3.out[3] ),
    .Y(_1067_));
 sg13g2_inv_1 _1982_ (.Y(_1068_),
    .A(_1067_));
 sg13g2_nand2_1 _1983_ (.Y(_1069_),
    .A(_0120_),
    .B(\div3.out[3] ));
 sg13g2_nand2_1 _1984_ (.Y(_1070_),
    .A(_1068_),
    .B(_1069_));
 sg13g2_inv_1 _1985_ (.Y(_1071_),
    .A(_1070_));
 sg13g2_nand2_1 _1986_ (.Y(_1072_),
    .A(_1066_),
    .B(_1071_));
 sg13g2_nand3_1 _1987_ (.B(_1065_),
    .C(_1070_),
    .A(_1063_),
    .Y(_1073_));
 sg13g2_nand2_1 _1988_ (.Y(_1074_),
    .A(_1072_),
    .B(_1073_));
 sg13g2_nand2_1 _1989_ (.Y(_1075_),
    .A(_1062_),
    .B(_1074_));
 sg13g2_nand2_1 _1990_ (.Y(_1076_),
    .A(_0142_),
    .B(\div3.out[1] ));
 sg13g2_inv_1 _1991_ (.Y(_1077_),
    .A(_1076_));
 sg13g2_inv_1 _1992_ (.Y(_1078_),
    .A(_1061_));
 sg13g2_nand2_1 _1993_ (.Y(_1079_),
    .A(_1078_),
    .B(_1060_));
 sg13g2_inv_1 _1994_ (.Y(_1080_),
    .A(_1079_));
 sg13g2_nand2_1 _1995_ (.Y(_1081_),
    .A(_1059_),
    .B(_1080_));
 sg13g2_nand3_1 _1996_ (.B(_1058_),
    .C(_1079_),
    .A(_1056_),
    .Y(_1082_));
 sg13g2_nand2_1 _1997_ (.Y(_1083_),
    .A(_1081_),
    .B(_1082_));
 sg13g2_nor2_1 _1998_ (.A(_1077_),
    .B(_1083_),
    .Y(_1084_));
 sg13g2_xnor2_1 _1999_ (.Y(_1085_),
    .A(_1070_),
    .B(_1066_));
 sg13g2_nand2_1 _2000_ (.Y(_1086_),
    .A(_1081_),
    .B(_1078_));
 sg13g2_nand2_1 _2001_ (.Y(_1087_),
    .A(_1085_),
    .B(_1086_));
 sg13g2_inv_1 _2002_ (.Y(_1088_),
    .A(_1087_));
 sg13g2_a21oi_1 _2003_ (.A1(_1075_),
    .A2(_1084_),
    .Y(_1089_),
    .B1(_1088_));
 sg13g2_inv_1 _2004_ (.Y(_1090_),
    .A(_0020_));
 sg13g2_nand2_1 _2005_ (.Y(_1091_),
    .A(net73),
    .B(_1090_));
 sg13g2_inv_1 _2006_ (.Y(_1092_),
    .A(_0021_));
 sg13g2_nand3_1 _2007_ (.B(_1054_),
    .C(_1092_),
    .A(_1045_),
    .Y(_1093_));
 sg13g2_nand2_1 _2008_ (.Y(_1094_),
    .A(_1091_),
    .B(_1093_));
 sg13g2_xor2_1 _2009_ (.B(\div3.out[5] ),
    .A(_0120_),
    .X(_1095_));
 sg13g2_nand2_1 _2010_ (.Y(_1096_),
    .A(_1094_),
    .B(_1095_));
 sg13g2_inv_1 _2011_ (.Y(_1097_),
    .A(_1095_));
 sg13g2_nand3_1 _2012_ (.B(_1093_),
    .C(_1097_),
    .A(_1091_),
    .Y(_1098_));
 sg13g2_nand2_2 _2013_ (.Y(_1099_),
    .A(_1096_),
    .B(_1098_));
 sg13g2_nand2_1 _2014_ (.Y(_1100_),
    .A(net73),
    .B(_1064_));
 sg13g2_nand3_1 _2015_ (.B(_1054_),
    .C(_1090_),
    .A(_1045_),
    .Y(_1101_));
 sg13g2_nand2_1 _2016_ (.Y(_1102_),
    .A(_1100_),
    .B(_1101_));
 sg13g2_nand2_1 _2017_ (.Y(_1103_),
    .A(net81),
    .B(\div3.out[4] ));
 sg13g2_nor2_1 _2018_ (.A(net81),
    .B(\div3.out[4] ),
    .Y(_1104_));
 sg13g2_a21oi_2 _2019_ (.B1(_1104_),
    .Y(_1105_),
    .A2(_1103_),
    .A1(_1102_));
 sg13g2_xor2_1 _2020_ (.B(_1105_),
    .A(_1099_),
    .X(_1106_));
 sg13g2_nand2b_1 _2021_ (.Y(_1107_),
    .B(_1103_),
    .A_N(_1104_));
 sg13g2_xnor2_1 _2022_ (.Y(_1108_),
    .A(_1107_),
    .B(_1102_));
 sg13g2_a21oi_1 _2023_ (.A1(_1066_),
    .A2(_1069_),
    .Y(_1109_),
    .B1(_1067_));
 sg13g2_nand2_1 _2024_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nand2b_1 _2025_ (.Y(_1111_),
    .B(_1102_),
    .A_N(_1107_));
 sg13g2_nand3_1 _2026_ (.B(_1101_),
    .C(_1107_),
    .A(_1100_),
    .Y(_1112_));
 sg13g2_nand2_1 _2027_ (.Y(_1113_),
    .A(_1111_),
    .B(_1112_));
 sg13g2_nand2_1 _2028_ (.Y(_1114_),
    .A(_1072_),
    .B(_1068_));
 sg13g2_nand2_1 _2029_ (.Y(_1115_),
    .A(_1113_),
    .B(_1114_));
 sg13g2_nand2_1 _2030_ (.Y(_1116_),
    .A(_1110_),
    .B(_1115_));
 sg13g2_nand2_1 _2031_ (.Y(_1117_),
    .A(_1106_),
    .B(_1116_));
 sg13g2_nor2_1 _2032_ (.A(_1089_),
    .B(_1117_),
    .Y(_1118_));
 sg13g2_nand2_1 _2033_ (.Y(_1119_),
    .A(_1108_),
    .B(_1114_));
 sg13g2_inv_1 _2034_ (.Y(_1120_),
    .A(_1119_));
 sg13g2_nand2_1 _2035_ (.Y(_1121_),
    .A(_1105_),
    .B(_1099_));
 sg13g2_nor2_1 _2036_ (.A(_1099_),
    .B(_1105_),
    .Y(_1122_));
 sg13g2_a21oi_1 _2037_ (.A1(_1120_),
    .A2(_1121_),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_nor2b_1 _2038_ (.A(_1118_),
    .B_N(_1123_),
    .Y(_1124_));
 sg13g2_nand2_1 _2039_ (.Y(_1125_),
    .A(_1109_),
    .B(_1113_));
 sg13g2_nand2_1 _2040_ (.Y(_1126_),
    .A(_1119_),
    .B(_1125_));
 sg13g2_xnor2_1 _2041_ (.Y(_1127_),
    .A(_1099_),
    .B(_1105_));
 sg13g2_nor2_1 _2042_ (.A(_1126_),
    .B(_1127_),
    .Y(_1128_));
 sg13g2_nand2_1 _2043_ (.Y(_1129_),
    .A(_1083_),
    .B(_1077_));
 sg13g2_nand3_1 _2044_ (.B(_1082_),
    .C(_1076_),
    .A(_1081_),
    .Y(_1130_));
 sg13g2_nand2_1 _2045_ (.Y(_1131_),
    .A(_1129_),
    .B(_1130_));
 sg13g2_nand2_1 _2046_ (.Y(_1132_),
    .A(_1087_),
    .B(_1075_));
 sg13g2_nor2_1 _2047_ (.A(_1131_),
    .B(_1132_),
    .Y(_1133_));
 sg13g2_nor2_1 _2048_ (.A(_0993_),
    .B(net73),
    .Y(_1134_));
 sg13g2_nor2_1 _2049_ (.A(net82),
    .B(_1031_),
    .Y(_1135_));
 sg13g2_a21oi_1 _2050_ (.A1(_1134_),
    .A2(_1038_),
    .Y(_1136_),
    .B1(_1135_));
 sg13g2_xor2_1 _2051_ (.B(\div3.out[1] ),
    .A(_0142_),
    .X(_1137_));
 sg13g2_nand2_1 _2052_ (.Y(_1138_),
    .A(_1136_),
    .B(_1137_));
 sg13g2_nor2b_1 _2053_ (.A(net73),
    .B_N(_0015_),
    .Y(_1139_));
 sg13g2_a21oi_2 _2054_ (.B1(_1139_),
    .Y(_1140_),
    .A2(_1055_),
    .A1(_0017_));
 sg13g2_nor2_1 _2055_ (.A(_1137_),
    .B(_1136_),
    .Y(_1141_));
 sg13g2_a21oi_1 _2056_ (.A1(_1138_),
    .A2(_1140_),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_inv_2 _2057_ (.Y(_1143_),
    .A(_1142_));
 sg13g2_nand3_1 _2058_ (.B(_1133_),
    .C(_1143_),
    .A(_1128_),
    .Y(_1144_));
 sg13g2_nand2_1 _2059_ (.Y(_1145_),
    .A(_1124_),
    .B(_1144_));
 sg13g2_o21ai_1 _2060_ (.B1(_1096_),
    .Y(_1146_),
    .A1(_0120_),
    .A2(\div3.out[5] ));
 sg13g2_inv_1 _2061_ (.Y(_1147_),
    .A(_0023_));
 sg13g2_nor2_1 _2062_ (.A(\counter[9] ),
    .B(net73),
    .Y(_1148_));
 sg13g2_a21oi_1 _2063_ (.A1(_1008_),
    .A2(net73),
    .Y(_1149_),
    .B1(_1148_));
 sg13g2_xnor2_1 _2064_ (.Y(_1150_),
    .A(_1147_),
    .B(_1149_));
 sg13g2_xnor2_1 _2065_ (.Y(_1151_),
    .A(_1146_),
    .B(_1150_));
 sg13g2_inv_1 _2066_ (.Y(_1152_),
    .A(_1151_));
 sg13g2_nand2_1 _2067_ (.Y(_1153_),
    .A(_1145_),
    .B(_1152_));
 sg13g2_nand3_1 _2068_ (.B(_1144_),
    .C(_1151_),
    .A(_1124_),
    .Y(_1154_));
 sg13g2_nand2_1 _2069_ (.Y(_1155_),
    .A(_1153_),
    .B(_1154_));
 sg13g2_nand3_1 _2070_ (.B(net76),
    .C(_0018_),
    .A(_1155_),
    .Y(_1156_));
 sg13g2_inv_1 _2071_ (.Y(_1157_),
    .A(_1156_));
 sg13g2_xor2_1 _2072_ (.B(\div3.out[5] ),
    .A(_0263_),
    .X(_1158_));
 sg13g2_xnor2_1 _2073_ (.Y(_1159_),
    .A(_1137_),
    .B(_1156_));
 sg13g2_a22oi_1 _2074_ (.Y(_1160_),
    .B1(_1158_),
    .B2(_1159_),
    .A2(_1157_),
    .A1(\div3.out[1] ));
 sg13g2_nor2_1 _2075_ (.A(_1039_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_nand2_1 _2076_ (.Y(_1162_),
    .A(_1160_),
    .B(_1039_));
 sg13g2_inv_1 _2077_ (.Y(_1163_),
    .A(_1162_));
 sg13g2_nor2_1 _2078_ (.A(_1161_),
    .B(_1163_),
    .Y(_1164_));
 sg13g2_nand3_1 _2079_ (.B(_1154_),
    .C(net78),
    .A(_1153_),
    .Y(_1165_));
 sg13g2_a21oi_1 _2080_ (.A1(_1129_),
    .A2(_1141_),
    .Y(_1166_),
    .B1(_1084_));
 sg13g2_xnor2_1 _2081_ (.Y(_1167_),
    .A(_1086_),
    .B(_1074_));
 sg13g2_nand2_1 _2082_ (.Y(_1168_),
    .A(_1167_),
    .B(_1116_));
 sg13g2_nor2_1 _2083_ (.A(_1166_),
    .B(_1168_),
    .Y(_1169_));
 sg13g2_a21oi_1 _2084_ (.A1(_1088_),
    .A2(_1125_),
    .Y(_1170_),
    .B1(_1120_));
 sg13g2_nor2b_1 _2085_ (.A(_1169_),
    .B_N(_1170_),
    .Y(_1171_));
 sg13g2_nor2_1 _2086_ (.A(_1132_),
    .B(_1126_),
    .Y(_1172_));
 sg13g2_nand2b_1 _2087_ (.Y(_1173_),
    .B(_1138_),
    .A_N(_1141_));
 sg13g2_nor2_1 _2088_ (.A(_1173_),
    .B(_1131_),
    .Y(_1174_));
 sg13g2_nand3_1 _2089_ (.B(_1140_),
    .C(_1174_),
    .A(_1172_),
    .Y(_1175_));
 sg13g2_nand2_1 _2090_ (.Y(_1176_),
    .A(_1171_),
    .B(_1175_));
 sg13g2_nand2_1 _2091_ (.Y(_1177_),
    .A(_1176_),
    .B(_1127_));
 sg13g2_nand3_1 _2092_ (.B(_1175_),
    .C(_1106_),
    .A(_1171_),
    .Y(_1178_));
 sg13g2_nand3_1 _2093_ (.B(_1178_),
    .C(net76),
    .A(_1177_),
    .Y(_1179_));
 sg13g2_nand3_1 _2094_ (.B(_1179_),
    .C(_0018_),
    .A(_1165_),
    .Y(_1180_));
 sg13g2_xnor2_1 _2095_ (.Y(_1181_),
    .A(_1018_),
    .B(\div3.out[2] ));
 sg13g2_nand2_1 _2096_ (.Y(_1182_),
    .A(_1180_),
    .B(_1181_));
 sg13g2_xnor2_1 _2097_ (.Y(_1183_),
    .A(_0285_),
    .B(_1031_));
 sg13g2_inv_1 _2098_ (.Y(_1184_),
    .A(_1183_));
 sg13g2_nand2_1 _2099_ (.Y(_1185_),
    .A(_1145_),
    .B(_1151_));
 sg13g2_nand3_1 _2100_ (.B(_1144_),
    .C(_1152_),
    .A(_1124_),
    .Y(_1186_));
 sg13g2_nand3_1 _2101_ (.B(_1186_),
    .C(_1016_),
    .A(_1185_),
    .Y(_1187_));
 sg13g2_nand2_1 _2102_ (.Y(_1188_),
    .A(_1176_),
    .B(_1106_));
 sg13g2_nand3_1 _2103_ (.B(_1175_),
    .C(_1127_),
    .A(_1171_),
    .Y(_1189_));
 sg13g2_nand3_1 _2104_ (.B(_1189_),
    .C(_0153_),
    .A(_1188_),
    .Y(_1190_));
 sg13g2_nand2_1 _2105_ (.Y(_1191_),
    .A(_1187_),
    .B(_1190_));
 sg13g2_inv_1 _2106_ (.Y(_1192_),
    .A(_1181_));
 sg13g2_nand3_1 _2107_ (.B(_0018_),
    .C(_1192_),
    .A(_1191_),
    .Y(_1193_));
 sg13g2_inv_1 _2108_ (.Y(_1194_),
    .A(_1193_));
 sg13g2_a21oi_2 _2109_ (.B1(_1194_),
    .Y(_1195_),
    .A2(_1184_),
    .A1(_1182_));
 sg13g2_xnor2_1 _2110_ (.Y(_1196_),
    .A(_1158_),
    .B(_1159_));
 sg13g2_nor2_1 _2111_ (.A(_1195_),
    .B(_1196_),
    .Y(_1197_));
 sg13g2_xor2_1 _2112_ (.B(_1196_),
    .A(_1195_),
    .X(_1198_));
 sg13g2_nand3_1 _2113_ (.B(_1178_),
    .C(net78),
    .A(_1177_),
    .Y(_1199_));
 sg13g2_nand2_1 _2114_ (.Y(_1200_),
    .A(_1133_),
    .B(_1143_));
 sg13g2_nand2_1 _2115_ (.Y(_1201_),
    .A(_1200_),
    .B(_1089_));
 sg13g2_xnor2_1 _2116_ (.Y(_1202_),
    .A(_1116_),
    .B(_1201_));
 sg13g2_nand2_1 _2117_ (.Y(_1203_),
    .A(_1202_),
    .B(_0153_));
 sg13g2_nand3_1 _2118_ (.B(_0131_),
    .C(_1203_),
    .A(_1199_),
    .Y(_1204_));
 sg13g2_xnor2_1 _2119_ (.Y(_1205_),
    .A(net81),
    .B(\div3.out[3] ));
 sg13g2_nand3_1 _2120_ (.B(net76),
    .C(net77),
    .A(_1155_),
    .Y(_1206_));
 sg13g2_nand3_1 _2121_ (.B(_1205_),
    .C(_1206_),
    .A(_1204_),
    .Y(_1207_));
 sg13g2_a21oi_1 _2122_ (.A1(_1204_),
    .A2(_1206_),
    .Y(_1208_),
    .B1(_1205_));
 sg13g2_a21oi_2 _2123_ (.B1(_1208_),
    .Y(_1209_),
    .A2(_1137_),
    .A1(_1207_));
 sg13g2_nand3_1 _2124_ (.B(_1193_),
    .C(_1184_),
    .A(_1182_),
    .Y(_1210_));
 sg13g2_nand2_1 _2125_ (.Y(_1211_),
    .A(_1180_),
    .B(_1192_));
 sg13g2_nand3_1 _2126_ (.B(_0018_),
    .C(_1181_),
    .A(_1191_),
    .Y(_1212_));
 sg13g2_nand3_1 _2127_ (.B(_1212_),
    .C(_1183_),
    .A(_1211_),
    .Y(_1213_));
 sg13g2_nand2_1 _2128_ (.Y(_1214_),
    .A(_1210_),
    .B(_1213_));
 sg13g2_nor2_1 _2129_ (.A(_1209_),
    .B(_1214_),
    .Y(_1215_));
 sg13g2_nand2_1 _2130_ (.Y(_1216_),
    .A(_1198_),
    .B(_1215_));
 sg13g2_nand2b_1 _2131_ (.Y(_1217_),
    .B(_1216_),
    .A_N(_1197_));
 sg13g2_xnor2_1 _2132_ (.Y(_1218_),
    .A(_1195_),
    .B(_1196_));
 sg13g2_nand2_1 _2133_ (.Y(_1219_),
    .A(_1199_),
    .B(_1203_));
 sg13g2_nand2_1 _2134_ (.Y(_1220_),
    .A(_1219_),
    .B(_0131_));
 sg13g2_nand2_1 _2135_ (.Y(_1221_),
    .A(_1155_),
    .B(net76));
 sg13g2_nand2_1 _2136_ (.Y(_1222_),
    .A(_1221_),
    .B(net77));
 sg13g2_nand3_1 _2137_ (.B(_1205_),
    .C(_1222_),
    .A(_1220_),
    .Y(_1223_));
 sg13g2_inv_1 _2138_ (.Y(_1224_),
    .A(_1205_));
 sg13g2_nand3_1 _2139_ (.B(_1224_),
    .C(_1206_),
    .A(_1204_),
    .Y(_1225_));
 sg13g2_nand3_1 _2140_ (.B(_1225_),
    .C(_1137_),
    .A(_1223_),
    .Y(_1226_));
 sg13g2_nand3_1 _2141_ (.B(_1224_),
    .C(_1222_),
    .A(_1220_),
    .Y(_1227_));
 sg13g2_inv_1 _2142_ (.Y(_1228_),
    .A(_1137_));
 sg13g2_nand3_1 _2143_ (.B(_1207_),
    .C(_1228_),
    .A(_1227_),
    .Y(_1229_));
 sg13g2_nand2_1 _2144_ (.Y(_1230_),
    .A(_1226_),
    .B(_1229_));
 sg13g2_nand2_1 _2145_ (.Y(_1231_),
    .A(_1191_),
    .B(net77));
 sg13g2_xnor2_1 _2146_ (.Y(_1232_),
    .A(_0351_),
    .B(\div3.out[4] ));
 sg13g2_a21oi_1 _2147_ (.A1(_1143_),
    .A2(_1129_),
    .Y(_1233_),
    .B1(_1084_));
 sg13g2_xnor2_1 _2148_ (.Y(_1234_),
    .A(_1167_),
    .B(_1233_));
 sg13g2_nor2_1 _2149_ (.A(net78),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_a21oi_1 _2150_ (.A1(_1202_),
    .A2(net78),
    .Y(_1236_),
    .B1(_1235_));
 sg13g2_nand2_1 _2151_ (.Y(_1237_),
    .A(_1236_),
    .B(_0131_));
 sg13g2_nand3_1 _2152_ (.B(_1232_),
    .C(_1237_),
    .A(_1231_),
    .Y(_1238_));
 sg13g2_a21oi_1 _2153_ (.A1(_1231_),
    .A2(_1237_),
    .Y(_1239_),
    .B1(_1232_));
 sg13g2_a21oi_1 _2154_ (.A1(_1238_),
    .A2(_1192_),
    .Y(_1240_),
    .B1(_1239_));
 sg13g2_inv_1 _2155_ (.Y(_1241_),
    .A(_1240_));
 sg13g2_nand2_2 _2156_ (.Y(_1242_),
    .A(_1230_),
    .B(_1241_));
 sg13g2_nand2_1 _2157_ (.Y(_1243_),
    .A(_1182_),
    .B(_1193_));
 sg13g2_xnor2_1 _2158_ (.Y(_1244_),
    .A(_1184_),
    .B(_1243_));
 sg13g2_inv_2 _2159_ (.Y(_1245_),
    .A(_1209_));
 sg13g2_nand2_1 _2160_ (.Y(_1246_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_nand2_1 _2161_ (.Y(_1247_),
    .A(_1214_),
    .B(_1209_));
 sg13g2_nand2_1 _2162_ (.Y(_1248_),
    .A(_1246_),
    .B(_1247_));
 sg13g2_nor3_1 _2163_ (.A(_1218_),
    .B(_1242_),
    .C(_1248_),
    .Y(_1249_));
 sg13g2_nor3_1 _2164_ (.A(_1164_),
    .B(_1217_),
    .C(_1249_),
    .Y(_1250_));
 sg13g2_inv_1 _2165_ (.Y(_1251_),
    .A(_1217_));
 sg13g2_nor2_1 _2166_ (.A(_1245_),
    .B(_1244_),
    .Y(_1252_));
 sg13g2_nor2_1 _2167_ (.A(_1215_),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nand3_1 _2168_ (.B(_1207_),
    .C(_1137_),
    .A(_1227_),
    .Y(_1254_));
 sg13g2_nand3_1 _2169_ (.B(_1225_),
    .C(_1228_),
    .A(_1223_),
    .Y(_1255_));
 sg13g2_nand2_1 _2170_ (.Y(_1256_),
    .A(_1254_),
    .B(_1255_));
 sg13g2_nor2_1 _2171_ (.A(_1240_),
    .B(_1256_),
    .Y(_1257_));
 sg13g2_nand3_1 _2172_ (.B(_1198_),
    .C(_1257_),
    .A(_1253_),
    .Y(_1258_));
 sg13g2_nand2_1 _2173_ (.Y(_1259_),
    .A(_1251_),
    .B(_1258_));
 sg13g2_nand2_2 _2174_ (.Y(_1260_),
    .A(_1259_),
    .B(_1164_));
 sg13g2_inv_1 _2175_ (.Y(_1261_),
    .A(_1260_));
 sg13g2_a21oi_1 _2176_ (.A1(_1250_),
    .A2(_1161_),
    .Y(_1262_),
    .B1(_1261_));
 sg13g2_a21oi_1 _2177_ (.A1(_1257_),
    .A2(_1247_),
    .Y(_1263_),
    .B1(_1215_));
 sg13g2_xnor2_1 _2178_ (.Y(_1264_),
    .A(_1198_),
    .B(_1263_));
 sg13g2_nand2_1 _2179_ (.Y(_1265_),
    .A(_1262_),
    .B(_1264_));
 sg13g2_o21ai_1 _2180_ (.B1(_1246_),
    .Y(_1266_),
    .A1(_1252_),
    .A2(_1242_));
 sg13g2_nand2_1 _2181_ (.Y(_1267_),
    .A(_1266_),
    .B(_1198_));
 sg13g2_nand2_1 _2182_ (.Y(_1268_),
    .A(_1263_),
    .B(_1218_));
 sg13g2_nand2_1 _2183_ (.Y(_1269_),
    .A(_1253_),
    .B(_1242_));
 sg13g2_nand2_1 _2184_ (.Y(_1270_),
    .A(_1248_),
    .B(_1257_));
 sg13g2_nand2_1 _2185_ (.Y(_1271_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_nand3_1 _2186_ (.B(_1268_),
    .C(_1271_),
    .A(_1267_),
    .Y(_1272_));
 sg13g2_nand2_1 _2187_ (.Y(_1273_),
    .A(_1231_),
    .B(_1237_));
 sg13g2_xor2_1 _2188_ (.B(_1273_),
    .A(_1232_),
    .X(_1274_));
 sg13g2_xnor2_1 _2189_ (.Y(_1275_),
    .A(_1192_),
    .B(_1274_));
 sg13g2_nand2_1 _2190_ (.Y(_1276_),
    .A(_1256_),
    .B(_1240_));
 sg13g2_nand2_1 _2191_ (.Y(_1277_),
    .A(_1242_),
    .B(_1276_));
 sg13g2_inv_1 _2192_ (.Y(_1278_),
    .A(_1277_));
 sg13g2_a21oi_1 _2193_ (.A1(_1271_),
    .A2(_1275_),
    .Y(_1279_),
    .B1(_1278_));
 sg13g2_nor2_1 _2194_ (.A(_1271_),
    .B(_1264_),
    .Y(_1280_));
 sg13g2_a21oi_2 _2195_ (.B1(_1280_),
    .Y(_1281_),
    .A2(_1279_),
    .A1(_1272_));
 sg13g2_inv_2 _2196_ (.Y(_1282_),
    .A(_1281_));
 sg13g2_nand2_1 _2197_ (.Y(_1283_),
    .A(_1265_),
    .B(_1282_));
 sg13g2_nor2_1 _2198_ (.A(_1161_),
    .B(_1250_),
    .Y(_1284_));
 sg13g2_nand2_1 _2199_ (.Y(_1285_),
    .A(_1284_),
    .B(_1260_));
 sg13g2_nand2_1 _2200_ (.Y(_1286_),
    .A(_1262_),
    .B(_1285_));
 sg13g2_nand2_1 _2201_ (.Y(_1287_),
    .A(_1286_),
    .B(_1281_));
 sg13g2_nand2_1 _2202_ (.Y(_1288_),
    .A(_1283_),
    .B(_1287_));
 sg13g2_nand2_1 _2203_ (.Y(_1289_),
    .A(_1267_),
    .B(_1268_));
 sg13g2_nand3_1 _2204_ (.B(_1260_),
    .C(_1289_),
    .A(_1284_),
    .Y(_1290_));
 sg13g2_buf_8 _2205_ (.A(_1290_),
    .X(_1291_));
 sg13g2_nand2_1 _2206_ (.Y(_1292_),
    .A(_1288_),
    .B(_1291_));
 sg13g2_xnor2_1 _2207_ (.Y(_1293_),
    .A(net74),
    .B(_1292_));
 sg13g2_xnor2_1 _2208_ (.Y(_1294_),
    .A(_1242_),
    .B(_1248_));
 sg13g2_nand2_1 _2209_ (.Y(_1295_),
    .A(_1289_),
    .B(_1294_));
 sg13g2_nand2_1 _2210_ (.Y(_1296_),
    .A(_1295_),
    .B(_1272_));
 sg13g2_nand2b_1 _2211_ (.Y(_1297_),
    .B(_1296_),
    .A_N(_1279_));
 sg13g2_nand3_1 _2212_ (.B(_1272_),
    .C(_1279_),
    .A(_1295_),
    .Y(_1298_));
 sg13g2_nand2_1 _2213_ (.Y(_1299_),
    .A(_1297_),
    .B(_1298_));
 sg13g2_inv_1 _2214_ (.Y(_1300_),
    .A(_1036_));
 sg13g2_nand2_1 _2215_ (.Y(_1301_),
    .A(_1299_),
    .B(_1300_));
 sg13g2_nor2_1 _2216_ (.A(\div3.in[0] ),
    .B(_1031_),
    .Y(_1302_));
 sg13g2_xor2_1 _2217_ (.B(_1034_),
    .A(_1302_),
    .X(_1303_));
 sg13g2_inv_1 _2218_ (.Y(_1304_),
    .A(_1275_));
 sg13g2_nand2_1 _2219_ (.Y(_1305_),
    .A(_1277_),
    .B(_1304_));
 sg13g2_nand3_1 _2220_ (.B(_1276_),
    .C(_1275_),
    .A(_1242_),
    .Y(_1306_));
 sg13g2_nand2_1 _2221_ (.Y(_1307_),
    .A(_1305_),
    .B(_1306_));
 sg13g2_nand2b_1 _2222_ (.Y(_1308_),
    .B(_1307_),
    .A_N(_1303_));
 sg13g2_nor2_1 _2223_ (.A(_1033_),
    .B(_1275_),
    .Y(_1309_));
 sg13g2_nand3_1 _2224_ (.B(_1306_),
    .C(_1303_),
    .A(_1305_),
    .Y(_1310_));
 sg13g2_inv_1 _2225_ (.Y(_1311_),
    .A(_1310_));
 sg13g2_a21oi_1 _2226_ (.A1(_1308_),
    .A2(_1309_),
    .Y(_1312_),
    .B1(_1311_));
 sg13g2_nand3_1 _2227_ (.B(_1277_),
    .C(_1275_),
    .A(_1294_),
    .Y(_1313_));
 sg13g2_o21ai_1 _2228_ (.B1(_1271_),
    .Y(_1314_),
    .A1(_1278_),
    .A2(_1304_));
 sg13g2_a21oi_1 _2229_ (.A1(_1313_),
    .A2(_1314_),
    .Y(_1315_),
    .B1(net74));
 sg13g2_nand3_1 _2230_ (.B(_1314_),
    .C(net74),
    .A(_1313_),
    .Y(_1316_));
 sg13g2_o21ai_1 _2231_ (.B1(_1316_),
    .Y(_1317_),
    .A1(_1312_),
    .A2(_1315_));
 sg13g2_buf_2 _2232_ (.A(_1317_),
    .X(_1318_));
 sg13g2_nand3_1 _2233_ (.B(_1298_),
    .C(net74),
    .A(_1297_),
    .Y(_1319_));
 sg13g2_inv_1 _2234_ (.Y(_1320_),
    .A(_1319_));
 sg13g2_a21oi_1 _2235_ (.A1(_1301_),
    .A2(_1318_),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_nand2_1 _2236_ (.Y(_1322_),
    .A(_1285_),
    .B(_1264_));
 sg13g2_nand2_1 _2237_ (.Y(_1323_),
    .A(_1322_),
    .B(_1291_));
 sg13g2_nand2_1 _2238_ (.Y(_1324_),
    .A(_1323_),
    .B(_1282_));
 sg13g2_nand3_1 _2239_ (.B(_1291_),
    .C(_1281_),
    .A(_1322_),
    .Y(_1325_));
 sg13g2_nand2_1 _2240_ (.Y(_1326_),
    .A(_1324_),
    .B(_1325_));
 sg13g2_nor2_1 _2241_ (.A(net74),
    .B(_1326_),
    .Y(_1327_));
 sg13g2_nand2_1 _2242_ (.Y(_1328_),
    .A(_1326_),
    .B(net74));
 sg13g2_o21ai_1 _2243_ (.B1(_1328_),
    .Y(_1329_),
    .A1(_1321_),
    .A2(_1327_));
 sg13g2_nand2_1 _2244_ (.Y(_1330_),
    .A(_1282_),
    .B(_1322_));
 sg13g2_nand3_1 _2245_ (.B(_1262_),
    .C(_1291_),
    .A(_1330_),
    .Y(_1331_));
 sg13g2_nand2b_1 _2246_ (.Y(_1332_),
    .B(_1260_),
    .A_N(_1250_));
 sg13g2_nand2b_1 _2247_ (.Y(_1333_),
    .B(_1260_),
    .A_N(_1161_));
 sg13g2_nand4_1 _2248_ (.B(_1332_),
    .C(_1333_),
    .A(_1282_),
    .Y(_1334_),
    .D(_1289_));
 sg13g2_nand2_1 _2249_ (.Y(_1335_),
    .A(_1331_),
    .B(_1334_));
 sg13g2_nand2_1 _2250_ (.Y(_1336_),
    .A(_1335_),
    .B(net74));
 sg13g2_nand3_1 _2251_ (.B(_1334_),
    .C(_1300_),
    .A(_1331_),
    .Y(_1337_));
 sg13g2_nand2_2 _2252_ (.Y(_1338_),
    .A(_1336_),
    .B(_1337_));
 sg13g2_inv_1 _2253_ (.Y(_1339_),
    .A(_1338_));
 sg13g2_nand2_1 _2254_ (.Y(_1340_),
    .A(_1329_),
    .B(_1339_));
 sg13g2_nand2_1 _2255_ (.Y(_1341_),
    .A(_1340_),
    .B(_1336_));
 sg13g2_xor2_1 _2256_ (.B(_1341_),
    .A(_1293_),
    .X(_1342_));
 sg13g2_inv_1 _2257_ (.Y(_1343_),
    .A(_1312_));
 sg13g2_nand2_1 _2258_ (.Y(_1344_),
    .A(_1313_),
    .B(_1314_));
 sg13g2_nand2_1 _2259_ (.Y(_1345_),
    .A(_1344_),
    .B(_1300_));
 sg13g2_nand2_1 _2260_ (.Y(_1346_),
    .A(_1345_),
    .B(_1316_));
 sg13g2_xnor2_1 _2261_ (.Y(_1347_),
    .A(_1343_),
    .B(_1346_));
 sg13g2_buf_4 _2262_ (.X(_1348_),
    .A(_1347_));
 sg13g2_buf_8 _2263_ (.A(_1348_),
    .X(_1349_));
 sg13g2_buf_1 _2264_ (.A(net63),
    .X(_1350_));
 sg13g2_nand2_1 _2265_ (.Y(_1351_),
    .A(_1308_),
    .B(_1310_));
 sg13g2_inv_1 _2266_ (.Y(_1352_),
    .A(_1309_));
 sg13g2_nand2_1 _2267_ (.Y(_1353_),
    .A(_1351_),
    .B(_1352_));
 sg13g2_nand3_1 _2268_ (.B(_1310_),
    .C(_1309_),
    .A(_1308_),
    .Y(_1354_));
 sg13g2_nand2_2 _2269_ (.Y(_1355_),
    .A(_1353_),
    .B(_1354_));
 sg13g2_inv_2 _2270_ (.Y(_1356_),
    .A(_1355_));
 sg13g2_buf_8 _2271_ (.A(_1356_),
    .X(_1357_));
 sg13g2_buf_8 _2272_ (.A(net62),
    .X(_1358_));
 sg13g2_buf_1 _2273_ (.A(net49),
    .X(_1359_));
 sg13g2_nand2_1 _2274_ (.Y(_1360_),
    .A(_1275_),
    .B(_1033_));
 sg13g2_nand2_1 _2275_ (.Y(_1361_),
    .A(_1352_),
    .B(_1360_));
 sg13g2_buf_1 _2276_ (.A(_1361_),
    .X(_1362_));
 sg13g2_nor2_2 _2277_ (.A(net80),
    .B(net70),
    .Y(_1363_));
 sg13g2_inv_2 _2278_ (.Y(_1364_),
    .A(_1363_));
 sg13g2_nand2_2 _2279_ (.Y(_1365_),
    .A(net70),
    .B(net75));
 sg13g2_nand2_1 _2280_ (.Y(_1366_),
    .A(_1364_),
    .B(_1365_));
 sg13g2_nor2_2 _2281_ (.A(_0978_),
    .B(net70),
    .Y(_1367_));
 sg13g2_inv_4 _2282_ (.A(net70),
    .Y(_1368_));
 sg13g2_buf_1 _2283_ (.A(_1368_),
    .X(_1369_));
 sg13g2_nor2_1 _2284_ (.A(_0979_),
    .B(net67),
    .Y(_1370_));
 sg13g2_nor2_1 _2285_ (.A(_1367_),
    .B(_1370_),
    .Y(_1371_));
 sg13g2_inv_1 _2286_ (.Y(_1372_),
    .A(_1371_));
 sg13g2_nor2_2 _2287_ (.A(_1372_),
    .B(net62),
    .Y(_1373_));
 sg13g2_a21oi_1 _2288_ (.A1(net36),
    .A2(_1366_),
    .Y(_1374_),
    .B1(_1373_));
 sg13g2_inv_2 _2289_ (.Y(_1375_),
    .A(net75));
 sg13g2_nor2_2 _2290_ (.A(_1375_),
    .B(net70),
    .Y(_1376_));
 sg13g2_nor2_2 _2291_ (.A(_0626_),
    .B(_1368_),
    .Y(_1377_));
 sg13g2_nor2_1 _2292_ (.A(_1376_),
    .B(_1377_),
    .Y(_1378_));
 sg13g2_inv_1 _2293_ (.Y(_1379_),
    .A(_1378_));
 sg13g2_buf_8 _2294_ (.A(_1355_),
    .X(_1380_));
 sg13g2_buf_8 _2295_ (.A(net65),
    .X(_1381_));
 sg13g2_buf_1 _2296_ (.A(net61),
    .X(_1382_));
 sg13g2_nor2_1 _2297_ (.A(_1379_),
    .B(net48),
    .Y(_1383_));
 sg13g2_nand3_1 _2298_ (.B(_1345_),
    .C(_1316_),
    .A(_1343_),
    .Y(_1384_));
 sg13g2_nand2_1 _2299_ (.Y(_1385_),
    .A(_1346_),
    .B(_1312_));
 sg13g2_nand2_1 _2300_ (.Y(_1386_),
    .A(_1384_),
    .B(_1385_));
 sg13g2_buf_8 _2301_ (.A(_1386_),
    .X(_1387_));
 sg13g2_buf_8 _2302_ (.A(net60),
    .X(_1388_));
 sg13g2_nor2_1 _2303_ (.A(_1383_),
    .B(net47),
    .Y(_1389_));
 sg13g2_nor2_1 _2304_ (.A(_1376_),
    .B(net49),
    .Y(_1390_));
 sg13g2_nor2_1 _2305_ (.A(_0980_),
    .B(net67),
    .Y(_1391_));
 sg13g2_inv_1 _2306_ (.Y(_1392_),
    .A(_1391_));
 sg13g2_nand2_1 _2307_ (.Y(_1393_),
    .A(_1390_),
    .B(_1392_));
 sg13g2_nand2_1 _2308_ (.Y(_1394_),
    .A(_1389_),
    .B(_1393_));
 sg13g2_o21ai_1 _2309_ (.B1(_1394_),
    .Y(_1395_),
    .A1(net50),
    .A2(_1374_));
 sg13g2_nand2_1 _2310_ (.Y(_1396_),
    .A(_1301_),
    .B(_1319_));
 sg13g2_xnor2_1 _2311_ (.Y(_1397_),
    .A(_1318_),
    .B(_1396_));
 sg13g2_buf_1 _2312_ (.A(_1397_),
    .X(_1398_));
 sg13g2_buf_8 _2313_ (.A(net35),
    .X(_1399_));
 sg13g2_buf_8 _2314_ (.A(net30),
    .X(_1400_));
 sg13g2_nand2_1 _2315_ (.Y(_1401_),
    .A(_1395_),
    .B(net25));
 sg13g2_inv_1 _2316_ (.Y(_1402_),
    .A(_1318_));
 sg13g2_nand2_1 _2317_ (.Y(_1403_),
    .A(_1396_),
    .B(_1402_));
 sg13g2_nand3_1 _2318_ (.B(_1319_),
    .C(_1318_),
    .A(_1301_),
    .Y(_1404_));
 sg13g2_nand2_1 _2319_ (.Y(_1405_),
    .A(_1403_),
    .B(_1404_));
 sg13g2_buf_8 _2320_ (.A(_1405_),
    .X(_1406_));
 sg13g2_buf_1 _2321_ (.A(net29),
    .X(_1407_));
 sg13g2_buf_8 _2322_ (.A(net60),
    .X(_1408_));
 sg13g2_buf_1 _2323_ (.A(net46),
    .X(_1409_));
 sg13g2_nand2_2 _2324_ (.Y(_1410_),
    .A(net62),
    .B(_1379_));
 sg13g2_buf_8 _2325_ (.A(net65),
    .X(_1411_));
 sg13g2_nor2_2 _2326_ (.A(_0978_),
    .B(_1369_),
    .Y(_1412_));
 sg13g2_inv_2 _2327_ (.Y(_1413_),
    .A(_1412_));
 sg13g2_nor2_2 _2328_ (.A(net80),
    .B(_0975_),
    .Y(_1414_));
 sg13g2_nor2_2 _2329_ (.A(_1414_),
    .B(_1362_),
    .Y(_1415_));
 sg13g2_inv_1 _2330_ (.Y(_1416_),
    .A(_1415_));
 sg13g2_nand3_1 _2331_ (.B(_1413_),
    .C(_1416_),
    .A(net59),
    .Y(_1417_));
 sg13g2_nand3_1 _2332_ (.B(_1410_),
    .C(_1417_),
    .A(net34),
    .Y(_1418_));
 sg13g2_buf_1 _2333_ (.A(net60),
    .X(_1419_));
 sg13g2_nor2_1 _2334_ (.A(_1390_),
    .B(net45),
    .Y(_1420_));
 sg13g2_nor2_1 _2335_ (.A(_0626_),
    .B(net70),
    .Y(_1421_));
 sg13g2_buf_8 _2336_ (.A(_1355_),
    .X(_1422_));
 sg13g2_nor2_1 _2337_ (.A(net69),
    .B(net64),
    .Y(_1423_));
 sg13g2_inv_1 _2338_ (.Y(_1424_),
    .A(_1423_));
 sg13g2_nand2_1 _2339_ (.Y(_1425_),
    .A(_1420_),
    .B(_1424_));
 sg13g2_nand3_1 _2340_ (.B(_1418_),
    .C(_1425_),
    .A(net24),
    .Y(_1426_));
 sg13g2_nand2_1 _2341_ (.Y(_1427_),
    .A(_1401_),
    .B(_1426_));
 sg13g2_inv_1 _2342_ (.Y(_1428_),
    .A(_1321_));
 sg13g2_nand3_1 _2343_ (.B(_1325_),
    .C(_1300_),
    .A(_1324_),
    .Y(_1429_));
 sg13g2_nand3_1 _2344_ (.B(_1328_),
    .C(_1429_),
    .A(_1428_),
    .Y(_1430_));
 sg13g2_nand2_1 _2345_ (.Y(_1431_),
    .A(_1328_),
    .B(_1429_));
 sg13g2_nand2_1 _2346_ (.Y(_1432_),
    .A(_1431_),
    .B(_1321_));
 sg13g2_nand2_1 _2347_ (.Y(_1433_),
    .A(_1430_),
    .B(_1432_));
 sg13g2_buf_1 _2348_ (.A(_1433_),
    .X(_1434_));
 sg13g2_buf_1 _2349_ (.A(net17),
    .X(_1435_));
 sg13g2_nand2_1 _2350_ (.Y(_1436_),
    .A(_1427_),
    .B(_1435_));
 sg13g2_xnor2_1 _2351_ (.Y(_1437_),
    .A(_1338_),
    .B(_1329_));
 sg13g2_buf_8 _2352_ (.A(_1437_),
    .X(_1438_));
 sg13g2_xnor2_1 _2353_ (.Y(_1439_),
    .A(_1428_),
    .B(_1431_));
 sg13g2_buf_1 _2354_ (.A(_1439_),
    .X(_1440_));
 sg13g2_buf_1 _2355_ (.A(_1440_),
    .X(_1441_));
 sg13g2_nor2_2 _2356_ (.A(net75),
    .B(_1368_),
    .Y(_1442_));
 sg13g2_inv_1 _2357_ (.Y(_1443_),
    .A(_1442_));
 sg13g2_nand2_2 _2358_ (.Y(_1444_),
    .A(_1355_),
    .B(_1443_));
 sg13g2_inv_1 _2359_ (.Y(_1445_),
    .A(_1444_));
 sg13g2_nand2_1 _2360_ (.Y(_1446_),
    .A(net67),
    .B(_1414_));
 sg13g2_nand2_1 _2361_ (.Y(_1447_),
    .A(_1445_),
    .B(_1446_));
 sg13g2_nor2_2 _2362_ (.A(_1413_),
    .B(net64),
    .Y(_1448_));
 sg13g2_inv_1 _2363_ (.Y(_1449_),
    .A(_1448_));
 sg13g2_nand2_1 _2364_ (.Y(_1450_),
    .A(_1447_),
    .B(_1449_));
 sg13g2_buf_8 _2365_ (.A(_1348_),
    .X(_1451_));
 sg13g2_buf_1 _2366_ (.A(net58),
    .X(_1452_));
 sg13g2_nand2_1 _2367_ (.Y(_1453_),
    .A(_1450_),
    .B(_1452_));
 sg13g2_nor2_1 _2368_ (.A(_1413_),
    .B(net36),
    .Y(_1454_));
 sg13g2_nor2_2 _2369_ (.A(net80),
    .B(_1368_),
    .Y(_1455_));
 sg13g2_nor2_1 _2370_ (.A(_1367_),
    .B(_1455_),
    .Y(_1456_));
 sg13g2_buf_1 _2371_ (.A(net64),
    .X(_1457_));
 sg13g2_buf_1 _2372_ (.A(net57),
    .X(_1458_));
 sg13g2_nor3_1 _2373_ (.A(_1375_),
    .B(_1456_),
    .C(net43),
    .Y(_1459_));
 sg13g2_buf_1 _2374_ (.A(_1386_),
    .X(_1460_));
 sg13g2_buf_8 _2375_ (.A(net56),
    .X(_1461_));
 sg13g2_o21ai_1 _2376_ (.B1(net42),
    .Y(_1462_),
    .A1(_1454_),
    .A2(_1459_));
 sg13g2_nand2_1 _2377_ (.Y(_1463_),
    .A(_1453_),
    .B(_1462_));
 sg13g2_nand2_1 _2378_ (.Y(_1464_),
    .A(_1463_),
    .B(net24));
 sg13g2_buf_1 _2379_ (.A(net35),
    .X(_1465_));
 sg13g2_inv_2 _2380_ (.Y(_1466_),
    .A(_1414_));
 sg13g2_nor2_2 _2381_ (.A(_1466_),
    .B(net67),
    .Y(_1467_));
 sg13g2_nor2_2 _2382_ (.A(_1467_),
    .B(net61),
    .Y(_1468_));
 sg13g2_o21ai_1 _2383_ (.B1(_1387_),
    .Y(_1469_),
    .A1(_1468_),
    .A2(_1445_));
 sg13g2_nor2_2 _2384_ (.A(_0494_),
    .B(_0978_),
    .Y(_1470_));
 sg13g2_nor2_1 _2385_ (.A(_1470_),
    .B(net65),
    .Y(_1471_));
 sg13g2_nand2_1 _2386_ (.Y(_1472_),
    .A(_1471_),
    .B(_1446_));
 sg13g2_buf_1 _2387_ (.A(net61),
    .X(_1473_));
 sg13g2_nor2_1 _2388_ (.A(net69),
    .B(_1455_),
    .Y(_1474_));
 sg13g2_nand2_1 _2389_ (.Y(_1475_),
    .A(_1473_),
    .B(_1474_));
 sg13g2_nand2_1 _2390_ (.Y(_1476_),
    .A(_1472_),
    .B(_1475_));
 sg13g2_buf_1 _2391_ (.A(_1348_),
    .X(_1477_));
 sg13g2_nand2_1 _2392_ (.Y(_1478_),
    .A(_1476_),
    .B(_1477_));
 sg13g2_nand2_1 _2393_ (.Y(_1479_),
    .A(_1469_),
    .B(_1478_));
 sg13g2_nand2_1 _2394_ (.Y(_1480_),
    .A(net28),
    .B(_1479_));
 sg13g2_nand2_1 _2395_ (.Y(_1481_),
    .A(_1464_),
    .B(_1480_));
 sg13g2_nand2_1 _2396_ (.Y(_1482_),
    .A(net16),
    .B(_1481_));
 sg13g2_nand3_1 _2397_ (.B(net23),
    .C(_1482_),
    .A(_1436_),
    .Y(_1483_));
 sg13g2_inv_1 _2398_ (.Y(_1484_),
    .A(_1328_));
 sg13g2_a21oi_1 _2399_ (.A1(_1428_),
    .A2(_1429_),
    .Y(_1485_),
    .B1(_1484_));
 sg13g2_nand2_1 _2400_ (.Y(_1486_),
    .A(_1485_),
    .B(_1338_));
 sg13g2_nand2_2 _2401_ (.Y(_1487_),
    .A(_1340_),
    .B(_1486_));
 sg13g2_buf_1 _2402_ (.A(_1487_),
    .X(_1488_));
 sg13g2_buf_1 _2403_ (.A(net70),
    .X(_1489_));
 sg13g2_nor2_2 _2404_ (.A(_0979_),
    .B(net68),
    .Y(_1490_));
 sg13g2_nor3_1 _2405_ (.A(_1442_),
    .B(_1490_),
    .C(net59),
    .Y(_1491_));
 sg13g2_nand2_2 _2406_ (.Y(_1492_),
    .A(net59),
    .B(_1364_));
 sg13g2_inv_1 _2407_ (.Y(_1493_),
    .A(_1492_));
 sg13g2_buf_1 _2408_ (.A(net60),
    .X(_1494_));
 sg13g2_nor3_1 _2409_ (.A(_1491_),
    .B(_1493_),
    .C(net40),
    .Y(_1495_));
 sg13g2_nor2_1 _2410_ (.A(_1490_),
    .B(_1412_),
    .Y(_1496_));
 sg13g2_nand2_1 _2411_ (.Y(_1497_),
    .A(_1473_),
    .B(_1496_));
 sg13g2_inv_1 _2412_ (.Y(_1498_),
    .A(_1497_));
 sg13g2_nor2_1 _2413_ (.A(_1370_),
    .B(_1381_),
    .Y(_1499_));
 sg13g2_nand2b_1 _2414_ (.Y(_1500_),
    .B(net60),
    .A_N(_1499_));
 sg13g2_nor2_1 _2415_ (.A(_1498_),
    .B(_1500_),
    .Y(_1501_));
 sg13g2_nor2_1 _2416_ (.A(_1495_),
    .B(_1501_),
    .Y(_1502_));
 sg13g2_buf_1 _2417_ (.A(net29),
    .X(_1503_));
 sg13g2_nand2_1 _2418_ (.Y(_1504_),
    .A(_1502_),
    .B(net21));
 sg13g2_buf_8 _2419_ (.A(_1348_),
    .X(_1505_));
 sg13g2_buf_1 _2420_ (.A(net54),
    .X(_1506_));
 sg13g2_buf_8 _2421_ (.A(net48),
    .X(_1507_));
 sg13g2_nor2_2 _2422_ (.A(net80),
    .B(net65),
    .Y(_1508_));
 sg13g2_a21oi_1 _2423_ (.A1(net33),
    .A2(_1391_),
    .Y(_1509_),
    .B1(_1508_));
 sg13g2_nor2_1 _2424_ (.A(_1470_),
    .B(net67),
    .Y(_1510_));
 sg13g2_o21ai_1 _2425_ (.B1(net41),
    .Y(_1511_),
    .A1(_1510_),
    .A2(_1415_));
 sg13g2_nand2_1 _2426_ (.Y(_1512_),
    .A(_1511_),
    .B(_1410_));
 sg13g2_nand2_1 _2427_ (.Y(_1513_),
    .A(_1512_),
    .B(net44));
 sg13g2_o21ai_1 _2428_ (.B1(_1513_),
    .Y(_1514_),
    .A1(net39),
    .A2(_1509_));
 sg13g2_nand2_1 _2429_ (.Y(_1515_),
    .A(_1514_),
    .B(net28));
 sg13g2_nand2_1 _2430_ (.Y(_1516_),
    .A(_1504_),
    .B(_1515_));
 sg13g2_nand2_1 _2431_ (.Y(_1517_),
    .A(_1516_),
    .B(net16));
 sg13g2_nor2_1 _2432_ (.A(_1363_),
    .B(net65),
    .Y(_1518_));
 sg13g2_nand2_1 _2433_ (.Y(_1519_),
    .A(net68),
    .B(_1470_));
 sg13g2_nand2_1 _2434_ (.Y(_1520_),
    .A(_1518_),
    .B(_1519_));
 sg13g2_o21ai_1 _2435_ (.B1(net41),
    .Y(_1521_),
    .A1(_0980_),
    .A2(_1363_));
 sg13g2_nand2_1 _2436_ (.Y(_1522_),
    .A(_1520_),
    .B(_1521_));
 sg13g2_nand2_1 _2437_ (.Y(_1523_),
    .A(_1522_),
    .B(net44));
 sg13g2_nor2_1 _2438_ (.A(net75),
    .B(net70),
    .Y(_1524_));
 sg13g2_nor2_1 _2439_ (.A(_1524_),
    .B(_1455_),
    .Y(_1525_));
 sg13g2_nand2_1 _2440_ (.Y(_1526_),
    .A(net62),
    .B(_1525_));
 sg13g2_nand2_1 _2441_ (.Y(_1527_),
    .A(net41),
    .B(_1413_));
 sg13g2_nand2_1 _2442_ (.Y(_1528_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_nand2_1 _2443_ (.Y(_1529_),
    .A(net42),
    .B(_1528_));
 sg13g2_nand2_1 _2444_ (.Y(_1530_),
    .A(_1523_),
    .B(_1529_));
 sg13g2_nand2_1 _2445_ (.Y(_1531_),
    .A(net28),
    .B(_1530_));
 sg13g2_inv_1 _2446_ (.Y(_1532_),
    .A(_1455_));
 sg13g2_nor2_1 _2447_ (.A(_1532_),
    .B(net57),
    .Y(_1533_));
 sg13g2_nand2_1 _2448_ (.Y(_1534_),
    .A(net50),
    .B(_1533_));
 sg13g2_nand2_1 _2449_ (.Y(_1535_),
    .A(net24),
    .B(_1534_));
 sg13g2_nand2_1 _2450_ (.Y(_1536_),
    .A(_1531_),
    .B(_1535_));
 sg13g2_nand2_1 _2451_ (.Y(_1537_),
    .A(net12),
    .B(_1536_));
 sg13g2_nand3_1 _2452_ (.B(_1517_),
    .C(_1537_),
    .A(net11),
    .Y(_1538_));
 sg13g2_nand3_1 _2453_ (.B(_1483_),
    .C(_1538_),
    .A(_1342_),
    .Y(_1539_));
 sg13g2_xnor2_1 _2454_ (.Y(_1540_),
    .A(_1293_),
    .B(_1341_));
 sg13g2_inv_1 _2455_ (.Y(_1541_),
    .A(_1377_));
 sg13g2_nand2_1 _2456_ (.Y(_1542_),
    .A(net65),
    .B(_0978_));
 sg13g2_o21ai_1 _2457_ (.B1(_1542_),
    .Y(_1543_),
    .A1(net43),
    .A2(_1541_));
 sg13g2_nor2_1 _2458_ (.A(_0980_),
    .B(_1412_),
    .Y(_1544_));
 sg13g2_inv_1 _2459_ (.Y(_1545_),
    .A(_1544_));
 sg13g2_nand2_1 _2460_ (.Y(_1546_),
    .A(net57),
    .B(_1545_));
 sg13g2_nor2_1 _2461_ (.A(_1362_),
    .B(_1351_),
    .Y(_1547_));
 sg13g2_nand2_1 _2462_ (.Y(_1548_),
    .A(_1547_),
    .B(_1375_));
 sg13g2_nand2_1 _2463_ (.Y(_1549_),
    .A(_1546_),
    .B(_1548_));
 sg13g2_nor2_1 _2464_ (.A(_1549_),
    .B(net47),
    .Y(_1550_));
 sg13g2_a21oi_1 _2465_ (.A1(net40),
    .A2(_1543_),
    .Y(_1551_),
    .B1(_1550_));
 sg13g2_buf_8 _2466_ (.A(net35),
    .X(_1552_));
 sg13g2_nor2_1 _2467_ (.A(_1551_),
    .B(net27),
    .Y(_1553_));
 sg13g2_buf_8 _2468_ (.A(net29),
    .X(_1554_));
 sg13g2_nand2_2 _2469_ (.Y(_1555_),
    .A(net68),
    .B(_1466_));
 sg13g2_nand2_2 _2470_ (.Y(_1556_),
    .A(_1381_),
    .B(net75));
 sg13g2_o21ai_1 _2471_ (.B1(_1556_),
    .Y(_1557_),
    .A1(net43),
    .A2(_1555_));
 sg13g2_nand2_1 _2472_ (.Y(_1558_),
    .A(net49),
    .B(_1545_));
 sg13g2_a21oi_1 _2473_ (.A1(_1444_),
    .A2(_1558_),
    .Y(_1559_),
    .B1(net46));
 sg13g2_a21oi_1 _2474_ (.A1(net42),
    .A2(_1557_),
    .Y(_1560_),
    .B1(_1559_));
 sg13g2_nor2_1 _2475_ (.A(net20),
    .B(_1560_),
    .Y(_1561_));
 sg13g2_nor2_1 _2476_ (.A(_1553_),
    .B(_1561_),
    .Y(_1562_));
 sg13g2_buf_8 _2477_ (.A(net22),
    .X(_1563_));
 sg13g2_nand2_1 _2478_ (.Y(_1564_),
    .A(_1562_),
    .B(net15));
 sg13g2_nand2_1 _2479_ (.Y(_1565_),
    .A(_1541_),
    .B(_1416_));
 sg13g2_nor2b_1 _2480_ (.A(net65),
    .B_N(_1565_),
    .Y(_1566_));
 sg13g2_inv_1 _2481_ (.Y(_1567_),
    .A(_1542_));
 sg13g2_nor2_1 _2482_ (.A(_1566_),
    .B(_1567_),
    .Y(_1568_));
 sg13g2_nor2_1 _2483_ (.A(_1568_),
    .B(_1348_),
    .Y(_1569_));
 sg13g2_inv_1 _2484_ (.Y(_1570_),
    .A(_1367_));
 sg13g2_nand2_1 _2485_ (.Y(_1571_),
    .A(_1468_),
    .B(_1570_));
 sg13g2_inv_1 _2486_ (.Y(_1572_),
    .A(_1365_));
 sg13g2_nor2_1 _2487_ (.A(_1470_),
    .B(net68),
    .Y(_1573_));
 sg13g2_o21ai_1 _2488_ (.B1(net48),
    .Y(_1574_),
    .A1(_1572_),
    .A2(_1573_));
 sg13g2_a21oi_1 _2489_ (.A1(_1571_),
    .A2(_1574_),
    .Y(_1575_),
    .B1(net47));
 sg13g2_nor2_1 _2490_ (.A(_1569_),
    .B(_1575_),
    .Y(_1576_));
 sg13g2_nor2_1 _2491_ (.A(net20),
    .B(_1576_),
    .Y(_1577_));
 sg13g2_buf_1 _2492_ (.A(net64),
    .X(_1578_));
 sg13g2_nor2_1 _2493_ (.A(_1443_),
    .B(net53),
    .Y(_1579_));
 sg13g2_inv_1 _2494_ (.Y(_1580_),
    .A(_1470_));
 sg13g2_nor2_1 _2495_ (.A(_1580_),
    .B(net68),
    .Y(_1581_));
 sg13g2_nor2_1 _2496_ (.A(_1581_),
    .B(_1356_),
    .Y(_1582_));
 sg13g2_inv_1 _2497_ (.Y(_1583_),
    .A(_1582_));
 sg13g2_nand2b_1 _2498_ (.Y(_1584_),
    .B(_1583_),
    .A_N(_1579_));
 sg13g2_nand2_2 _2499_ (.Y(_1585_),
    .A(_1411_),
    .B(net67));
 sg13g2_inv_1 _2500_ (.Y(_1586_),
    .A(_1490_));
 sg13g2_nand2_1 _2501_ (.Y(_1587_),
    .A(_1585_),
    .B(_1586_));
 sg13g2_nor2_1 _2502_ (.A(_1587_),
    .B(net63),
    .Y(_1588_));
 sg13g2_a21oi_1 _2503_ (.A1(net55),
    .A2(_1584_),
    .Y(_1589_),
    .B1(_1588_));
 sg13g2_nor2_1 _2504_ (.A(_1589_),
    .B(net27),
    .Y(_1590_));
 sg13g2_nor2_1 _2505_ (.A(_1577_),
    .B(_1590_),
    .Y(_1591_));
 sg13g2_buf_1 _2506_ (.A(_1433_),
    .X(_1592_));
 sg13g2_nand2_1 _2507_ (.Y(_1593_),
    .A(_1591_),
    .B(net14));
 sg13g2_nand2_1 _2508_ (.Y(_1594_),
    .A(_1564_),
    .B(_1593_));
 sg13g2_nand2_1 _2509_ (.Y(_1595_),
    .A(_1594_),
    .B(net23));
 sg13g2_buf_1 _2510_ (.A(net62),
    .X(_1596_));
 sg13g2_nand2_1 _2511_ (.Y(_1597_),
    .A(net38),
    .B(_1490_));
 sg13g2_o21ai_1 _2512_ (.B1(net64),
    .Y(_1598_),
    .A1(_0626_),
    .A2(_1363_));
 sg13g2_nand3_1 _2513_ (.B(_1597_),
    .C(_1598_),
    .A(net44),
    .Y(_1599_));
 sg13g2_nor2_1 _2514_ (.A(_1367_),
    .B(net64),
    .Y(_1600_));
 sg13g2_inv_1 _2515_ (.Y(_1601_),
    .A(_1600_));
 sg13g2_inv_1 _2516_ (.Y(_1602_),
    .A(_1555_));
 sg13g2_nor2_1 _2517_ (.A(_1376_),
    .B(_1602_),
    .Y(_1603_));
 sg13g2_nand2b_1 _2518_ (.Y(_1604_),
    .B(net59),
    .A_N(_1603_));
 sg13g2_nand2_1 _2519_ (.Y(_1605_),
    .A(_1601_),
    .B(_1604_));
 sg13g2_nand2_1 _2520_ (.Y(_1606_),
    .A(net42),
    .B(_1605_));
 sg13g2_nand2_1 _2521_ (.Y(_1607_),
    .A(_1599_),
    .B(_1606_));
 sg13g2_nand2_1 _2522_ (.Y(_1608_),
    .A(_1607_),
    .B(net24));
 sg13g2_nor2_2 _2523_ (.A(_1364_),
    .B(_1351_),
    .Y(_1609_));
 sg13g2_nand2_1 _2524_ (.Y(_1610_),
    .A(_1609_),
    .B(_0975_));
 sg13g2_inv_1 _2525_ (.Y(_1611_),
    .A(net66));
 sg13g2_a21oi_1 _2526_ (.A1(_1382_),
    .A2(net68),
    .Y(_1612_),
    .B1(_1611_));
 sg13g2_nand2_1 _2527_ (.Y(_1613_),
    .A(net39),
    .B(_1612_));
 sg13g2_nand2_1 _2528_ (.Y(_1614_),
    .A(_1552_),
    .B(_1613_));
 sg13g2_nand2_1 _2529_ (.Y(_1615_),
    .A(_1608_),
    .B(_1614_));
 sg13g2_nand2_1 _2530_ (.Y(_1616_),
    .A(net16),
    .B(_1615_));
 sg13g2_buf_1 _2531_ (.A(net47),
    .X(_1617_));
 sg13g2_nor2_2 _2532_ (.A(_1367_),
    .B(net62),
    .Y(_1618_));
 sg13g2_nor2_1 _2533_ (.A(_1376_),
    .B(_1442_),
    .Y(_1619_));
 sg13g2_nand2_1 _2534_ (.Y(_1620_),
    .A(net62),
    .B(_1619_));
 sg13g2_inv_1 _2535_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_nor2_1 _2536_ (.A(_1618_),
    .B(_1621_),
    .Y(_1622_));
 sg13g2_nand2_1 _2537_ (.Y(_1623_),
    .A(_1570_),
    .B(_1555_));
 sg13g2_nand2_1 _2538_ (.Y(_1624_),
    .A(net49),
    .B(_1623_));
 sg13g2_nand2_1 _2539_ (.Y(_1625_),
    .A(_1624_),
    .B(_1585_));
 sg13g2_nand2_1 _2540_ (.Y(_1626_),
    .A(net40),
    .B(_1625_));
 sg13g2_o21ai_1 _2541_ (.B1(_1626_),
    .Y(_1627_),
    .A1(_1617_),
    .A2(_1622_));
 sg13g2_nand2_1 _2542_ (.Y(_1628_),
    .A(net28),
    .B(_1627_));
 sg13g2_nor2_1 _2543_ (.A(_1375_),
    .B(net65),
    .Y(_1629_));
 sg13g2_nor2_2 _2544_ (.A(_0637_),
    .B(net67),
    .Y(_1630_));
 sg13g2_inv_1 _2545_ (.Y(_1631_),
    .A(_1630_));
 sg13g2_nand2_1 _2546_ (.Y(_1632_),
    .A(_1629_),
    .B(_1631_));
 sg13g2_nand2_1 _2547_ (.Y(_1633_),
    .A(_1422_),
    .B(net68));
 sg13g2_nand2_1 _2548_ (.Y(_1634_),
    .A(_1632_),
    .B(_1633_));
 sg13g2_nand2_1 _2549_ (.Y(_1635_),
    .A(_1634_),
    .B(net55));
 sg13g2_nand2_1 _2550_ (.Y(_1636_),
    .A(net48),
    .B(_1379_));
 sg13g2_o21ai_1 _2551_ (.B1(_1636_),
    .Y(_1637_),
    .A1(net43),
    .A2(_1372_));
 sg13g2_nand2_1 _2552_ (.Y(_1638_),
    .A(_1637_),
    .B(net40));
 sg13g2_nand2_1 _2553_ (.Y(_1639_),
    .A(_1635_),
    .B(_1638_));
 sg13g2_nand2_1 _2554_ (.Y(_1640_),
    .A(_1407_),
    .B(_1639_));
 sg13g2_nand2_1 _2555_ (.Y(_1641_),
    .A(_1628_),
    .B(_1640_));
 sg13g2_nand2_1 _2556_ (.Y(_1642_),
    .A(_1592_),
    .B(_1641_));
 sg13g2_nand3_1 _2557_ (.B(_1616_),
    .C(_1642_),
    .A(net11),
    .Y(_1643_));
 sg13g2_nand3_1 _2558_ (.B(_1595_),
    .C(_1643_),
    .A(_1540_),
    .Y(_1644_));
 sg13g2_a21oi_1 _2559_ (.A1(_1330_),
    .A2(_1291_),
    .Y(_1645_),
    .B1(_1286_));
 sg13g2_xnor2_1 _2560_ (.Y(_1646_),
    .A(net74),
    .B(_1645_));
 sg13g2_inv_1 _2561_ (.Y(_1647_),
    .A(_1299_));
 sg13g2_o21ai_1 _2562_ (.B1(_1037_),
    .Y(_1648_),
    .A1(_1647_),
    .A2(_1326_));
 sg13g2_nor3_1 _2563_ (.A(_1293_),
    .B(_1648_),
    .C(_1338_),
    .Y(_1649_));
 sg13g2_o21ai_1 _2564_ (.B1(_1037_),
    .Y(_1650_),
    .A1(_1292_),
    .A2(_1335_));
 sg13g2_nor2b_1 _2565_ (.A(_1649_),
    .B_N(_1650_),
    .Y(_1651_));
 sg13g2_nor2_1 _2566_ (.A(_1293_),
    .B(_1338_),
    .Y(_1652_));
 sg13g2_nor2_1 _2567_ (.A(_1396_),
    .B(_1431_),
    .Y(_1653_));
 sg13g2_nand3_1 _2568_ (.B(_1318_),
    .C(_1653_),
    .A(_1652_),
    .Y(_1654_));
 sg13g2_nand2_1 _2569_ (.Y(_1655_),
    .A(_1651_),
    .B(_1654_));
 sg13g2_nand2b_1 _2570_ (.Y(_1656_),
    .B(_1655_),
    .A_N(_1646_));
 sg13g2_nand3_1 _2571_ (.B(_1654_),
    .C(_1646_),
    .A(_1651_),
    .Y(_1657_));
 sg13g2_nand2_2 _2572_ (.Y(_1658_),
    .A(_1656_),
    .B(_1657_));
 sg13g2_buf_8 _2573_ (.A(_1658_),
    .X(_1659_));
 sg13g2_nand3_1 _2574_ (.B(_1644_),
    .C(net10),
    .A(_1539_),
    .Y(_1660_));
 sg13g2_inv_1 _2575_ (.Y(_1661_),
    .A(_0186_));
 sg13g2_nor2_2 _2576_ (.A(_0637_),
    .B(_1489_),
    .Y(_1662_));
 sg13g2_nor2_1 _2577_ (.A(_1662_),
    .B(net57),
    .Y(_1663_));
 sg13g2_nand2_1 _2578_ (.Y(_1664_),
    .A(net50),
    .B(_1663_));
 sg13g2_buf_1 _2579_ (.A(net42),
    .X(_1665_));
 sg13g2_nor2_1 _2580_ (.A(_1442_),
    .B(net41),
    .Y(_1666_));
 sg13g2_a21oi_1 _2581_ (.A1(net33),
    .A2(_1379_),
    .Y(_1667_),
    .B1(_1666_));
 sg13g2_a21oi_2 _2582_ (.B1(net21),
    .Y(_1668_),
    .A2(_1667_),
    .A1(net31));
 sg13g2_nor2_1 _2583_ (.A(net48),
    .B(net60),
    .Y(_1669_));
 sg13g2_nand2_1 _2584_ (.Y(_1670_),
    .A(_1387_),
    .B(net53));
 sg13g2_inv_1 _2585_ (.Y(_1671_),
    .A(_1670_));
 sg13g2_inv_1 _2586_ (.Y(_1672_),
    .A(_1619_));
 sg13g2_a221oi_1 _2587_ (.B2(_1672_),
    .C1(net25),
    .B1(_1671_),
    .A1(_0483_),
    .Y(_1673_),
    .A2(_1669_));
 sg13g2_a21oi_1 _2588_ (.A1(_1664_),
    .A2(_1668_),
    .Y(_1674_),
    .B1(_1673_));
 sg13g2_nor2b_1 _2589_ (.A(net10),
    .B_N(_1674_),
    .Y(_1675_));
 sg13g2_nor2_1 _2590_ (.A(_1661_),
    .B(_1675_),
    .Y(_1676_));
 sg13g2_nand2_1 _2591_ (.Y(_1677_),
    .A(_1660_),
    .B(_1676_));
 sg13g2_inv_1 _2592_ (.Y(_1678_),
    .A(_1662_));
 sg13g2_nand2_1 _2593_ (.Y(_0059_),
    .A(net64),
    .B(_1678_));
 sg13g2_inv_1 _2594_ (.Y(_0060_),
    .A(_0059_));
 sg13g2_nor2_1 _2595_ (.A(_0060_),
    .B(net55),
    .Y(_0061_));
 sg13g2_a21oi_1 _2596_ (.A1(_0059_),
    .A2(net66),
    .Y(_0062_),
    .B1(net46));
 sg13g2_buf_1 _2597_ (.A(net29),
    .X(_0063_));
 sg13g2_o21ai_1 _2598_ (.B1(_0063_),
    .Y(_0064_),
    .A1(_0061_),
    .A2(_0062_));
 sg13g2_nand2_1 _2599_ (.Y(_0065_),
    .A(_1422_),
    .B(_1662_));
 sg13g2_inv_1 _2600_ (.Y(_0066_),
    .A(_0065_));
 sg13g2_o21ai_1 _2601_ (.B1(net54),
    .Y(_0067_),
    .A1(_1448_),
    .A2(_0066_));
 sg13g2_inv_1 _2602_ (.Y(_0068_),
    .A(_1456_));
 sg13g2_nand2_1 _2603_ (.Y(_0069_),
    .A(net59),
    .B(_0068_));
 sg13g2_o21ai_1 _2604_ (.B1(_0069_),
    .Y(_0070_),
    .A1(net48),
    .A2(_1525_));
 sg13g2_nand2_1 _2605_ (.Y(_0071_),
    .A(_0070_),
    .B(_1419_));
 sg13g2_nand2_1 _2606_ (.Y(_0072_),
    .A(_0067_),
    .B(_0071_));
 sg13g2_nand2_1 _2607_ (.Y(_0073_),
    .A(_1552_),
    .B(_0072_));
 sg13g2_nand2_1 _2608_ (.Y(_0074_),
    .A(_0064_),
    .B(_0073_));
 sg13g2_nand2_1 _2609_ (.Y(_0075_),
    .A(_0074_),
    .B(net15));
 sg13g2_nand2_1 _2610_ (.Y(_0076_),
    .A(_1472_),
    .B(_1585_));
 sg13g2_nand2_1 _2611_ (.Y(_0077_),
    .A(_0076_),
    .B(net54));
 sg13g2_nor2_1 _2612_ (.A(net69),
    .B(_1510_),
    .Y(_0078_));
 sg13g2_inv_1 _2613_ (.Y(_0079_),
    .A(_1547_));
 sg13g2_nor2_2 _2614_ (.A(_1375_),
    .B(_0079_),
    .Y(_0080_));
 sg13g2_inv_1 _2615_ (.Y(_0081_),
    .A(_0080_));
 sg13g2_o21ai_1 _2616_ (.B1(_0081_),
    .Y(_0082_),
    .A1(_0078_),
    .A2(net38));
 sg13g2_buf_1 _2617_ (.A(net60),
    .X(_0083_));
 sg13g2_nand2_1 _2618_ (.Y(_0084_),
    .A(_0082_),
    .B(net37));
 sg13g2_nand2_1 _2619_ (.Y(_0085_),
    .A(_0077_),
    .B(_0084_));
 sg13g2_nand2_1 _2620_ (.Y(_0086_),
    .A(_1399_),
    .B(_0085_));
 sg13g2_nand2_1 _2621_ (.Y(_0087_),
    .A(_1669_),
    .B(_1467_));
 sg13g2_nand2_1 _2622_ (.Y(_0088_),
    .A(_0063_),
    .B(_0087_));
 sg13g2_nand2_1 _2623_ (.Y(_0089_),
    .A(_0086_),
    .B(_0088_));
 sg13g2_nand2_1 _2624_ (.Y(_0090_),
    .A(net14),
    .B(_0089_));
 sg13g2_nand2_1 _2625_ (.Y(_0091_),
    .A(_0075_),
    .B(_0090_));
 sg13g2_nand2_1 _2626_ (.Y(_0092_),
    .A(_0091_),
    .B(net11));
 sg13g2_nand2_1 _2627_ (.Y(_0093_),
    .A(_1357_),
    .B(_1519_));
 sg13g2_nand2_1 _2628_ (.Y(_0094_),
    .A(_1380_),
    .B(_1466_));
 sg13g2_nand3_1 _2629_ (.B(_1633_),
    .C(_0094_),
    .A(_0093_),
    .Y(_0095_));
 sg13g2_nand2_1 _2630_ (.Y(_0096_),
    .A(_0095_),
    .B(_1348_));
 sg13g2_nand2_1 _2631_ (.Y(_0097_),
    .A(_1469_),
    .B(_0096_));
 sg13g2_nand2_1 _2632_ (.Y(_0098_),
    .A(net35),
    .B(_0097_));
 sg13g2_buf_1 _2633_ (.A(_1348_),
    .X(_0099_));
 sg13g2_o21ai_1 _2634_ (.B1(net52),
    .Y(_0100_),
    .A1(_0066_),
    .A2(_1663_));
 sg13g2_nor2_1 _2635_ (.A(_1541_),
    .B(net49),
    .Y(_0101_));
 sg13g2_o21ai_1 _2636_ (.B1(net56),
    .Y(_0102_),
    .A1(_1533_),
    .A2(_0101_));
 sg13g2_nand2_1 _2637_ (.Y(_0103_),
    .A(_0100_),
    .B(_0102_));
 sg13g2_buf_1 _2638_ (.A(net29),
    .X(_0104_));
 sg13g2_nand2_1 _2639_ (.Y(_0105_),
    .A(_0103_),
    .B(net18));
 sg13g2_nand2_1 _2640_ (.Y(_0106_),
    .A(_0098_),
    .B(_0105_));
 sg13g2_nand2_1 _2641_ (.Y(_0107_),
    .A(net15),
    .B(_0106_));
 sg13g2_a21oi_1 _2642_ (.A1(net41),
    .A2(_1630_),
    .Y(_0108_),
    .B1(_0080_));
 sg13g2_nand2_1 _2643_ (.Y(_0110_),
    .A(_1598_),
    .B(_1620_));
 sg13g2_nand2_1 _2644_ (.Y(_0111_),
    .A(_0110_),
    .B(net37));
 sg13g2_o21ai_1 _2645_ (.B1(_0111_),
    .Y(_0112_),
    .A1(net46),
    .A2(_0108_));
 sg13g2_buf_1 _2646_ (.A(net35),
    .X(_0113_));
 sg13g2_nand2_1 _2647_ (.Y(_0114_),
    .A(_0112_),
    .B(net26));
 sg13g2_o21ai_1 _2648_ (.B1(_1620_),
    .Y(_0115_),
    .A1(_1596_),
    .A2(_1415_));
 sg13g2_nand2_1 _2649_ (.Y(_0116_),
    .A(_0115_),
    .B(_0099_));
 sg13g2_nand2_1 _2650_ (.Y(_0117_),
    .A(_1417_),
    .B(_0081_));
 sg13g2_nand2_1 _2651_ (.Y(_0118_),
    .A(_0117_),
    .B(net56));
 sg13g2_nand2_1 _2652_ (.Y(_0119_),
    .A(_0116_),
    .B(_0118_));
 sg13g2_nand2_1 _2653_ (.Y(_0121_),
    .A(net19),
    .B(_0119_));
 sg13g2_nand2_1 _2654_ (.Y(_0122_),
    .A(_0114_),
    .B(_0121_));
 sg13g2_nand2_1 _2655_ (.Y(_0123_),
    .A(_0122_),
    .B(_1434_));
 sg13g2_nand2_1 _2656_ (.Y(_0124_),
    .A(_0107_),
    .B(_0123_));
 sg13g2_nand2_1 _2657_ (.Y(_0125_),
    .A(_0124_),
    .B(net23));
 sg13g2_nand2_1 _2658_ (.Y(_0126_),
    .A(_0092_),
    .B(_0125_));
 sg13g2_nand2_1 _2659_ (.Y(_0127_),
    .A(_0126_),
    .B(_1342_));
 sg13g2_buf_1 _2660_ (.A(_1386_),
    .X(_0128_));
 sg13g2_nand2_1 _2661_ (.Y(_0129_),
    .A(net51),
    .B(_1492_));
 sg13g2_o21ai_1 _2662_ (.B1(_0129_),
    .Y(_0130_),
    .A1(net47),
    .A2(_1612_));
 sg13g2_nand2_1 _2663_ (.Y(_0132_),
    .A(net30),
    .B(_0130_));
 sg13g2_a21oi_1 _2664_ (.A1(net41),
    .A2(_1623_),
    .Y(_0133_),
    .B1(_1508_));
 sg13g2_nor2_1 _2665_ (.A(net69),
    .B(_1630_),
    .Y(_0134_));
 sg13g2_inv_1 _2666_ (.Y(_0135_),
    .A(_0134_));
 sg13g2_a21oi_1 _2667_ (.A1(net57),
    .A2(_0135_),
    .Y(_0136_),
    .B1(_1609_));
 sg13g2_nand2_1 _2668_ (.Y(_0137_),
    .A(net52),
    .B(_0136_));
 sg13g2_o21ai_1 _2669_ (.B1(_0137_),
    .Y(_0138_),
    .A1(net63),
    .A2(_0133_));
 sg13g2_nand2_1 _2670_ (.Y(_0139_),
    .A(_0138_),
    .B(net18));
 sg13g2_nand2_1 _2671_ (.Y(_0140_),
    .A(_0132_),
    .B(_0139_));
 sg13g2_nand2_1 _2672_ (.Y(_0141_),
    .A(net22),
    .B(_0140_));
 sg13g2_nor2_2 _2673_ (.A(_1364_),
    .B(_1356_),
    .Y(_0143_));
 sg13g2_o21ai_1 _2674_ (.B1(net52),
    .Y(_0144_),
    .A1(_1611_),
    .A2(_0143_));
 sg13g2_o21ai_1 _2675_ (.B1(net56),
    .Y(_0145_),
    .A1(_1602_),
    .A2(_1424_));
 sg13g2_nand2_1 _2676_ (.Y(_0146_),
    .A(_0144_),
    .B(_0145_));
 sg13g2_nand2_1 _2677_ (.Y(_0147_),
    .A(net30),
    .B(_0146_));
 sg13g2_nand2_1 _2678_ (.Y(_0148_),
    .A(_1632_),
    .B(_0059_));
 sg13g2_nand2_1 _2679_ (.Y(_0149_),
    .A(_0148_),
    .B(_1348_));
 sg13g2_nand2_1 _2680_ (.Y(_0150_),
    .A(net49),
    .B(_0068_));
 sg13g2_nand2_1 _2681_ (.Y(_0151_),
    .A(net51),
    .B(_0150_));
 sg13g2_nand2_1 _2682_ (.Y(_0152_),
    .A(_0149_),
    .B(_0151_));
 sg13g2_nand2_1 _2683_ (.Y(_0154_),
    .A(_0104_),
    .B(_0152_));
 sg13g2_nand2_1 _2684_ (.Y(_0155_),
    .A(_0147_),
    .B(_0154_));
 sg13g2_nand2_1 _2685_ (.Y(_0156_),
    .A(_0155_),
    .B(net17));
 sg13g2_nand2_1 _2686_ (.Y(_0157_),
    .A(_0141_),
    .B(_0156_));
 sg13g2_nand2_1 _2687_ (.Y(_0158_),
    .A(_0157_),
    .B(_1487_));
 sg13g2_a21oi_1 _2688_ (.A1(net38),
    .A2(_1545_),
    .Y(_0159_),
    .B1(_0066_));
 sg13g2_nand2_1 _2689_ (.Y(_0160_),
    .A(_1624_),
    .B(_1444_));
 sg13g2_nand2_1 _2690_ (.Y(_0161_),
    .A(_0083_),
    .B(_0160_));
 sg13g2_o21ai_1 _2691_ (.B1(_0161_),
    .Y(_0162_),
    .A1(_1388_),
    .A2(_0159_));
 sg13g2_nand2_1 _2692_ (.Y(_0163_),
    .A(_0162_),
    .B(net35));
 sg13g2_o21ai_1 _2693_ (.B1(_1556_),
    .Y(_0165_),
    .A1(net57),
    .A2(_1662_));
 sg13g2_nand2_1 _2694_ (.Y(_0166_),
    .A(_0165_),
    .B(net51));
 sg13g2_nand2_1 _2695_ (.Y(_0167_),
    .A(_1570_),
    .B(_1365_));
 sg13g2_nand2_1 _2696_ (.Y(_0168_),
    .A(net64),
    .B(_0167_));
 sg13g2_nand2_1 _2697_ (.Y(_0169_),
    .A(_0168_),
    .B(_0081_));
 sg13g2_nand2_1 _2698_ (.Y(_0170_),
    .A(net58),
    .B(_0169_));
 sg13g2_nand2_1 _2699_ (.Y(_0171_),
    .A(_0166_),
    .B(_0170_));
 sg13g2_nand2_1 _2700_ (.Y(_0172_),
    .A(_1406_),
    .B(_0171_));
 sg13g2_nand2_1 _2701_ (.Y(_0173_),
    .A(_0163_),
    .B(_0172_));
 sg13g2_nand2_1 _2702_ (.Y(_0174_),
    .A(net22),
    .B(_0173_));
 sg13g2_inv_1 _2703_ (.Y(_0176_),
    .A(_1569_));
 sg13g2_nor2_2 _2704_ (.A(_1524_),
    .B(_1380_),
    .Y(_0177_));
 sg13g2_nand2_1 _2705_ (.Y(_0178_),
    .A(_0177_),
    .B(_1541_));
 sg13g2_nand2b_1 _2706_ (.Y(_0179_),
    .B(net58),
    .A_N(_0178_));
 sg13g2_nand2_1 _2707_ (.Y(_0180_),
    .A(_0176_),
    .B(_0179_));
 sg13g2_nand2_1 _2708_ (.Y(_0181_),
    .A(net35),
    .B(_0180_));
 sg13g2_inv_1 _2709_ (.Y(_0182_),
    .A(_0143_));
 sg13g2_nand2_1 _2710_ (.Y(_0183_),
    .A(_0182_),
    .B(_1449_));
 sg13g2_nand2_1 _2711_ (.Y(_0184_),
    .A(_0183_),
    .B(_1451_));
 sg13g2_inv_1 _2712_ (.Y(_0185_),
    .A(_1518_));
 sg13g2_nand2_1 _2713_ (.Y(_0187_),
    .A(_1457_),
    .B(_1586_));
 sg13g2_nand2_1 _2714_ (.Y(_0188_),
    .A(_0185_),
    .B(_0187_));
 sg13g2_nand2_1 _2715_ (.Y(_0189_),
    .A(net51),
    .B(_0188_));
 sg13g2_nand2_1 _2716_ (.Y(_0190_),
    .A(_0184_),
    .B(_0189_));
 sg13g2_nand2_1 _2717_ (.Y(_0191_),
    .A(net29),
    .B(_0190_));
 sg13g2_nand2_1 _2718_ (.Y(_0192_),
    .A(_0181_),
    .B(_0191_));
 sg13g2_nand2_1 _2719_ (.Y(_0193_),
    .A(net17),
    .B(_0192_));
 sg13g2_nand2_1 _2720_ (.Y(_0194_),
    .A(_0174_),
    .B(_0193_));
 sg13g2_nand2_1 _2721_ (.Y(_0195_),
    .A(_0194_),
    .B(_1437_));
 sg13g2_nand2_1 _2722_ (.Y(_0196_),
    .A(_0158_),
    .B(_0195_));
 sg13g2_nand2_1 _2723_ (.Y(_0198_),
    .A(_0196_),
    .B(_1540_));
 sg13g2_nand3_1 _2724_ (.B(_0198_),
    .C(net10),
    .A(_0127_),
    .Y(_0199_));
 sg13g2_buf_1 _2725_ (.A(net20),
    .X(_0200_));
 sg13g2_a21oi_1 _2726_ (.A1(net36),
    .A2(_1367_),
    .Y(_0201_),
    .B1(net34));
 sg13g2_inv_1 _2727_ (.Y(_0202_),
    .A(_1508_));
 sg13g2_nand2_1 _2728_ (.Y(_0203_),
    .A(_0202_),
    .B(_0168_));
 sg13g2_o21ai_1 _2729_ (.B1(_1665_),
    .Y(_0204_),
    .A1(_1547_),
    .A2(_0203_));
 sg13g2_nand2b_1 _2730_ (.Y(_0205_),
    .B(_0204_),
    .A_N(_0201_));
 sg13g2_nor2_1 _2731_ (.A(_1377_),
    .B(_1457_),
    .Y(_0206_));
 sg13g2_nor2_1 _2732_ (.A(_0206_),
    .B(net56),
    .Y(_0207_));
 sg13g2_nand2_1 _2733_ (.Y(_0209_),
    .A(_0207_),
    .B(_1633_));
 sg13g2_a22oi_1 _2734_ (.Y(_0210_),
    .B1(_0209_),
    .B2(_1668_),
    .A2(_0205_),
    .A1(net13));
 sg13g2_nor2b_1 _2735_ (.A(_1658_),
    .B_N(_0210_),
    .Y(_0211_));
 sg13g2_nor2_1 _2736_ (.A(_0186_),
    .B(_0211_),
    .Y(_0212_));
 sg13g2_nand2_1 _2737_ (.Y(_0213_),
    .A(_0199_),
    .B(_0212_));
 sg13g2_nand3_1 _2738_ (.B(_0213_),
    .C(_0175_),
    .A(_1677_),
    .Y(_0214_));
 sg13g2_o21ai_1 _2739_ (.B1(net59),
    .Y(_0215_),
    .A1(_1442_),
    .A2(_1581_));
 sg13g2_inv_1 _2740_ (.Y(_0216_),
    .A(_1376_));
 sg13g2_nand2_1 _2741_ (.Y(_0217_),
    .A(_1532_),
    .B(_0216_));
 sg13g2_nand2_2 _2742_ (.Y(_0218_),
    .A(net62),
    .B(_0217_));
 sg13g2_a21oi_1 _2743_ (.A1(_0215_),
    .A2(_0218_),
    .Y(_0220_),
    .B1(net34));
 sg13g2_o21ai_1 _2744_ (.B1(net32),
    .Y(_0221_),
    .A1(_1566_),
    .A2(_1618_));
 sg13g2_nor2b_1 _2745_ (.A(_0220_),
    .B_N(_0221_),
    .Y(_0222_));
 sg13g2_inv_1 _2746_ (.Y(_0223_),
    .A(_1609_));
 sg13g2_a22oi_1 _2747_ (.Y(_0224_),
    .B1(net66),
    .B2(net34),
    .A2(_0223_),
    .A1(_1492_));
 sg13g2_nand2b_1 _2748_ (.Y(_0225_),
    .B(_1503_),
    .A_N(_0224_));
 sg13g2_o21ai_1 _2749_ (.B1(_0225_),
    .Y(_0226_),
    .A1(net13),
    .A2(_0222_));
 sg13g2_nand2b_1 _2750_ (.Y(_0227_),
    .B(_1435_),
    .A_N(_0226_));
 sg13g2_o21ai_1 _2751_ (.B1(net61),
    .Y(_0228_),
    .A1(_1572_),
    .A2(_1421_));
 sg13g2_a21oi_1 _2752_ (.A1(_0228_),
    .A2(_0081_),
    .Y(_0229_),
    .B1(net31));
 sg13g2_inv_1 _2753_ (.Y(_0231_),
    .A(_0166_));
 sg13g2_o21ai_1 _2754_ (.B1(net13),
    .Y(_0232_),
    .A1(_0229_),
    .A2(_0231_));
 sg13g2_inv_1 _2755_ (.Y(_0233_),
    .A(_0228_));
 sg13g2_inv_1 _2756_ (.Y(_0234_),
    .A(_0093_));
 sg13g2_o21ai_1 _2757_ (.B1(net34),
    .Y(_0235_),
    .A1(_1445_),
    .A2(_0234_));
 sg13g2_o21ai_1 _2758_ (.B1(_0235_),
    .Y(_0236_),
    .A1(net31),
    .A2(_0233_));
 sg13g2_nand2_1 _2759_ (.Y(_0237_),
    .A(_0236_),
    .B(net25));
 sg13g2_nand3_1 _2760_ (.B(_0232_),
    .C(_0237_),
    .A(net16),
    .Y(_0238_));
 sg13g2_nand3_1 _2761_ (.B(net23),
    .C(_0238_),
    .A(_0227_),
    .Y(_0239_));
 sg13g2_nand2_2 _2762_ (.Y(_0240_),
    .A(_1357_),
    .B(_0167_));
 sg13g2_o21ai_1 _2763_ (.B1(_0240_),
    .Y(_0242_),
    .A1(_1359_),
    .A2(_1573_));
 sg13g2_nor2b_1 _2764_ (.A(net31),
    .B_N(_0242_),
    .Y(_0243_));
 sg13g2_nand3_1 _2765_ (.B(net36),
    .C(_1467_),
    .A(_1408_),
    .Y(_0244_));
 sg13g2_nand2_1 _2766_ (.Y(_0245_),
    .A(_1398_),
    .B(_0244_));
 sg13g2_nand2_1 _2767_ (.Y(_0246_),
    .A(net49),
    .B(_1489_));
 sg13g2_nand2_1 _2768_ (.Y(_0247_),
    .A(_1461_),
    .B(_0246_));
 sg13g2_nand2_1 _2769_ (.Y(_0248_),
    .A(_0149_),
    .B(_0247_));
 sg13g2_nand2_1 _2770_ (.Y(_0249_),
    .A(net21),
    .B(_0248_));
 sg13g2_o21ai_1 _2771_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_0243_),
    .A2(_0245_));
 sg13g2_nand2_1 _2772_ (.Y(_0251_),
    .A(_0250_),
    .B(net12));
 sg13g2_inv_1 _2773_ (.Y(_0253_),
    .A(_0129_));
 sg13g2_o21ai_1 _2774_ (.B1(_1465_),
    .Y(_0254_),
    .A1(_1389_),
    .A2(_0253_));
 sg13g2_nand2_1 _2775_ (.Y(_0255_),
    .A(_1582_),
    .B(_1466_));
 sg13g2_nand3_1 _2776_ (.B(_0255_),
    .C(_1601_),
    .A(net32),
    .Y(_0256_));
 sg13g2_nor2_1 _2777_ (.A(_1663_),
    .B(net47),
    .Y(_0257_));
 sg13g2_o21ai_1 _2778_ (.B1(net61),
    .Y(_0258_),
    .A1(_1377_),
    .A2(_1363_));
 sg13g2_nand2_1 _2779_ (.Y(_0259_),
    .A(_0257_),
    .B(_0258_));
 sg13g2_nand3_1 _2780_ (.B(_0256_),
    .C(_0259_),
    .A(net24),
    .Y(_0260_));
 sg13g2_nand2_1 _2781_ (.Y(_0261_),
    .A(_0254_),
    .B(_0260_));
 sg13g2_nand2_1 _2782_ (.Y(_0262_),
    .A(_0261_),
    .B(_1441_));
 sg13g2_nand2_1 _2783_ (.Y(_0264_),
    .A(_0251_),
    .B(_0262_));
 sg13g2_nand2_1 _2784_ (.Y(_0265_),
    .A(_0264_),
    .B(net11));
 sg13g2_nand3_1 _2785_ (.B(_0265_),
    .C(_1540_),
    .A(_0239_),
    .Y(_0266_));
 sg13g2_a21oi_1 _2786_ (.A1(net34),
    .A2(_0228_),
    .Y(_0267_),
    .B1(_0257_));
 sg13g2_nand2_1 _2787_ (.Y(_0268_),
    .A(_0267_),
    .B(_0200_));
 sg13g2_nand2_1 _2788_ (.Y(_0269_),
    .A(net51),
    .B(_0185_));
 sg13g2_nor2_1 _2789_ (.A(_1445_),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_a21oi_1 _2790_ (.A1(_1632_),
    .A2(_1492_),
    .Y(_0271_),
    .B1(_1409_));
 sg13g2_o21ai_1 _2791_ (.B1(net25),
    .Y(_0272_),
    .A1(_0270_),
    .A2(_0271_));
 sg13g2_nand3_1 _2792_ (.B(_0268_),
    .C(_0272_),
    .A(net16),
    .Y(_0273_));
 sg13g2_o21ai_1 _2793_ (.B1(_1461_),
    .Y(_0275_),
    .A1(_0206_),
    .A2(_0060_));
 sg13g2_nor2_1 _2794_ (.A(_1377_),
    .B(_1358_),
    .Y(_0276_));
 sg13g2_o21ai_1 _2795_ (.B1(net50),
    .Y(_0277_),
    .A1(_1471_),
    .A2(_0276_));
 sg13g2_nand3_1 _2796_ (.B(_0275_),
    .C(_0277_),
    .A(net25),
    .Y(_0278_));
 sg13g2_nand2_1 _2797_ (.Y(_0279_),
    .A(net12),
    .B(_0278_));
 sg13g2_nand2_1 _2798_ (.Y(_0280_),
    .A(_0273_),
    .B(_0279_));
 sg13g2_nand2_1 _2799_ (.Y(_0281_),
    .A(_0280_),
    .B(net11));
 sg13g2_nand3_1 _2800_ (.B(_0240_),
    .C(_1598_),
    .A(net32),
    .Y(_0282_));
 sg13g2_nor2_1 _2801_ (.A(_0080_),
    .B(_1494_),
    .Y(_0283_));
 sg13g2_nand2b_1 _2802_ (.Y(_0284_),
    .B(net61),
    .A_N(_1525_));
 sg13g2_nand2_1 _2803_ (.Y(_0286_),
    .A(_0283_),
    .B(_0284_));
 sg13g2_nand3_1 _2804_ (.B(_0282_),
    .C(_0286_),
    .A(net28),
    .Y(_0287_));
 sg13g2_nand4_1 _2805_ (.B(_1556_),
    .C(_1633_),
    .A(_1506_),
    .Y(_0288_),
    .D(_0240_));
 sg13g2_nor2_1 _2806_ (.A(_0080_),
    .B(net63),
    .Y(_0289_));
 sg13g2_nand2_1 _2807_ (.Y(_0290_),
    .A(_0289_),
    .B(_1542_));
 sg13g2_nand3_1 _2808_ (.B(_1554_),
    .C(_0290_),
    .A(_0288_),
    .Y(_0291_));
 sg13g2_nand2_1 _2809_ (.Y(_0292_),
    .A(_0287_),
    .B(_0291_));
 sg13g2_nand2_1 _2810_ (.Y(_0293_),
    .A(_0292_),
    .B(net12));
 sg13g2_nand2_1 _2811_ (.Y(_0294_),
    .A(_0257_),
    .B(_0182_));
 sg13g2_nand2_1 _2812_ (.Y(_0295_),
    .A(net38),
    .B(_0216_));
 sg13g2_nand2_1 _2813_ (.Y(_0297_),
    .A(net61),
    .B(_1532_));
 sg13g2_nand3_1 _2814_ (.B(_0295_),
    .C(_0297_),
    .A(net32),
    .Y(_0298_));
 sg13g2_nand3_1 _2815_ (.B(_0294_),
    .C(_0298_),
    .A(net24),
    .Y(_0299_));
 sg13g2_nand2_1 _2816_ (.Y(_0300_),
    .A(_0299_),
    .B(_0098_));
 sg13g2_nand2_1 _2817_ (.Y(_0301_),
    .A(_0300_),
    .B(_1441_));
 sg13g2_nand2_1 _2818_ (.Y(_0302_),
    .A(_0293_),
    .B(_0301_));
 sg13g2_nand2_1 _2819_ (.Y(_0303_),
    .A(_0302_),
    .B(_1438_));
 sg13g2_nand3_1 _2820_ (.B(_0303_),
    .C(_1342_),
    .A(_0281_),
    .Y(_0304_));
 sg13g2_nand3_1 _2821_ (.B(_0304_),
    .C(net10),
    .A(_0266_),
    .Y(_0305_));
 sg13g2_o21ai_1 _2822_ (.B1(_1668_),
    .Y(_0306_),
    .A1(net31),
    .A2(_1585_));
 sg13g2_nor2_1 _2823_ (.A(_1621_),
    .B(net50),
    .Y(_0308_));
 sg13g2_o21ai_1 _2824_ (.B1(_0200_),
    .Y(_0309_),
    .A1(_0308_),
    .A2(_0201_));
 sg13g2_a21oi_1 _2825_ (.A1(_0306_),
    .A2(_0309_),
    .Y(_0310_),
    .B1(net10));
 sg13g2_nor2_1 _2826_ (.A(_0175_),
    .B(_0028_),
    .Y(_0311_));
 sg13g2_nor2b_1 _2827_ (.A(_0310_),
    .B_N(_0311_),
    .Y(_0312_));
 sg13g2_a21oi_1 _2828_ (.A1(_0305_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(\g_x[2] ));
 sg13g2_inv_1 _2829_ (.Y(_0314_),
    .A(_0024_));
 sg13g2_o21ai_1 _2830_ (.B1(_0285_),
    .Y(_0315_),
    .A1(net83),
    .A2(_0314_));
 sg13g2_nand3b_1 _2831_ (.B(_0659_),
    .C(_0315_),
    .Y(_0316_),
    .A_N(_0855_));
 sg13g2_a21oi_1 _2832_ (.A1(_0214_),
    .A2(_0313_),
    .Y(_0317_),
    .B1(_0316_));
 sg13g2_a21oi_1 _2833_ (.A1(_1571_),
    .A2(_1521_),
    .Y(_0319_),
    .B1(net55));
 sg13g2_nor2_1 _2834_ (.A(_1545_),
    .B(net48),
    .Y(_0320_));
 sg13g2_nand3b_1 _2835_ (.B(net44),
    .C(_0284_),
    .Y(_0321_),
    .A_N(_0320_));
 sg13g2_nand2b_1 _2836_ (.Y(_0322_),
    .B(_0321_),
    .A_N(_0319_));
 sg13g2_nand2_1 _2837_ (.Y(_0323_),
    .A(_0322_),
    .B(net28));
 sg13g2_a21oi_1 _2838_ (.A1(_1580_),
    .A2(net33),
    .Y(_0324_),
    .B1(_1448_));
 sg13g2_nand2_1 _2839_ (.Y(_0325_),
    .A(_1598_),
    .B(_1424_));
 sg13g2_nand2_1 _2840_ (.Y(_0326_),
    .A(_0325_),
    .B(net44));
 sg13g2_o21ai_1 _2841_ (.B1(_0326_),
    .Y(_0327_),
    .A1(net39),
    .A2(_0324_));
 sg13g2_nand2_1 _2842_ (.Y(_0328_),
    .A(_0327_),
    .B(net21));
 sg13g2_nand2_1 _2843_ (.Y(_0330_),
    .A(_0323_),
    .B(_0328_));
 sg13g2_nand2_1 _2844_ (.Y(_0331_),
    .A(_0330_),
    .B(net16));
 sg13g2_nand2_1 _2845_ (.Y(_0332_),
    .A(net38),
    .B(_1366_));
 sg13g2_nand2_1 _2846_ (.Y(_0333_),
    .A(_0332_),
    .B(_1546_));
 sg13g2_nor2b_1 _2847_ (.A(net39),
    .B_N(_0333_),
    .Y(_0334_));
 sg13g2_a21oi_1 _2848_ (.A1(_1583_),
    .A2(_0150_),
    .Y(_0335_),
    .B1(net32));
 sg13g2_o21ai_1 _2849_ (.B1(net21),
    .Y(_0336_),
    .A1(_0334_),
    .A2(_0335_));
 sg13g2_nor2_1 _2850_ (.A(_1555_),
    .B(_1458_),
    .Y(_0337_));
 sg13g2_nand2_1 _2851_ (.Y(_0338_),
    .A(net53),
    .B(_1572_));
 sg13g2_nand2b_1 _2852_ (.Y(_0339_),
    .B(_0338_),
    .A_N(_1573_));
 sg13g2_o21ai_1 _2853_ (.B1(net44),
    .Y(_0341_),
    .A1(_0337_),
    .A2(_0339_));
 sg13g2_nor2_1 _2854_ (.A(net69),
    .B(net36),
    .Y(_0342_));
 sg13g2_o21ai_1 _2855_ (.B1(net42),
    .Y(_0343_),
    .A1(_1566_),
    .A2(_0342_));
 sg13g2_nand2_1 _2856_ (.Y(_0344_),
    .A(_0341_),
    .B(_0343_));
 sg13g2_nand2_1 _2857_ (.Y(_0345_),
    .A(_0344_),
    .B(net28));
 sg13g2_nand2_1 _2858_ (.Y(_0346_),
    .A(_0336_),
    .B(_0345_));
 sg13g2_nand2_1 _2859_ (.Y(_0347_),
    .A(_0346_),
    .B(net12));
 sg13g2_nand3_1 _2860_ (.B(_0331_),
    .C(_0347_),
    .A(_1438_),
    .Y(_0348_));
 sg13g2_inv_1 _2861_ (.Y(_0349_),
    .A(_0338_));
 sg13g2_nor3_1 _2862_ (.A(_0080_),
    .B(_0349_),
    .C(net40),
    .Y(_0350_));
 sg13g2_nor2b_1 _2863_ (.A(_0151_),
    .B_N(_1636_),
    .Y(_0352_));
 sg13g2_nor2_1 _2864_ (.A(_0350_),
    .B(_0352_),
    .Y(_0353_));
 sg13g2_nand2_1 _2865_ (.Y(_0354_),
    .A(_0353_),
    .B(_1407_));
 sg13g2_a21oi_1 _2866_ (.A1(_1359_),
    .A2(_1623_),
    .Y(_0355_),
    .B1(_0143_));
 sg13g2_nand2_1 _2867_ (.Y(_0356_),
    .A(_0240_),
    .B(_1542_));
 sg13g2_nand2_1 _2868_ (.Y(_0357_),
    .A(_1477_),
    .B(_0356_));
 sg13g2_o21ai_1 _2869_ (.B1(_0357_),
    .Y(_0358_),
    .A1(_1506_),
    .A2(_0355_));
 sg13g2_nand2_1 _2870_ (.Y(_0359_),
    .A(_0358_),
    .B(_1465_));
 sg13g2_nand2_1 _2871_ (.Y(_0360_),
    .A(_0354_),
    .B(_0359_));
 sg13g2_nand2_1 _2872_ (.Y(_0361_),
    .A(_0360_),
    .B(net12));
 sg13g2_nor2_1 _2873_ (.A(_0494_),
    .B(net67),
    .Y(_0363_));
 sg13g2_nand2b_1 _2874_ (.Y(_0364_),
    .B(_1629_),
    .A_N(_0363_));
 sg13g2_nand2_1 _2875_ (.Y(_0365_),
    .A(_1382_),
    .B(_0135_));
 sg13g2_nand2_1 _2876_ (.Y(_0366_),
    .A(_0364_),
    .B(_0365_));
 sg13g2_nand2_1 _2877_ (.Y(_0367_),
    .A(_0366_),
    .B(_1452_));
 sg13g2_nand2_1 _2878_ (.Y(_0368_),
    .A(_0367_),
    .B(_1670_));
 sg13g2_nand2_1 _2879_ (.Y(_0369_),
    .A(net28),
    .B(_0368_));
 sg13g2_o21ai_1 _2880_ (.B1(_0332_),
    .Y(_0370_),
    .A1(_0626_),
    .A2(net36));
 sg13g2_nand2_1 _2881_ (.Y(_0371_),
    .A(_0370_),
    .B(net55));
 sg13g2_o21ai_1 _2882_ (.B1(net66),
    .Y(_0372_),
    .A1(_1555_),
    .A2(net36));
 sg13g2_nand2_1 _2883_ (.Y(_0374_),
    .A(_0372_),
    .B(net40));
 sg13g2_nand2_1 _2884_ (.Y(_0375_),
    .A(_0371_),
    .B(_0374_));
 sg13g2_nand2_1 _2885_ (.Y(_0376_),
    .A(net24),
    .B(_0375_));
 sg13g2_nand2_1 _2886_ (.Y(_0377_),
    .A(_0369_),
    .B(_0376_));
 sg13g2_nand2_1 _2887_ (.Y(_0378_),
    .A(net16),
    .B(_0377_));
 sg13g2_nand3_1 _2888_ (.B(_0361_),
    .C(_0378_),
    .A(_1488_),
    .Y(_0379_));
 sg13g2_nand3_1 _2889_ (.B(_1540_),
    .C(_0379_),
    .A(_0348_),
    .Y(_0380_));
 sg13g2_nor2_1 _2890_ (.A(_1412_),
    .B(_0094_),
    .Y(_0381_));
 sg13g2_o21ai_1 _2891_ (.B1(net54),
    .Y(_0382_),
    .A1(_1579_),
    .A2(_0381_));
 sg13g2_nor2_1 _2892_ (.A(_0167_),
    .B(net38),
    .Y(_0383_));
 sg13g2_o21ai_1 _2893_ (.B1(net45),
    .Y(_0385_),
    .A1(_0177_),
    .A2(_0383_));
 sg13g2_nand2_1 _2894_ (.Y(_0386_),
    .A(_0382_),
    .B(_0385_));
 sg13g2_nand2_1 _2895_ (.Y(_0387_),
    .A(_0386_),
    .B(net19));
 sg13g2_o21ai_1 _2896_ (.B1(net59),
    .Y(_0388_),
    .A1(_1442_),
    .A2(_1662_));
 sg13g2_nand2_1 _2897_ (.Y(_0389_),
    .A(_1472_),
    .B(_0388_));
 sg13g2_nand2_1 _2898_ (.Y(_0390_),
    .A(_0389_),
    .B(_0099_));
 sg13g2_nand2b_1 _2899_ (.Y(_0391_),
    .B(net37),
    .A_N(_0136_));
 sg13g2_nand2_1 _2900_ (.Y(_0392_),
    .A(_0390_),
    .B(_0391_));
 sg13g2_nand2_1 _2901_ (.Y(_0393_),
    .A(net26),
    .B(_0392_));
 sg13g2_nand2_1 _2902_ (.Y(_0394_),
    .A(_0387_),
    .B(_0393_));
 sg13g2_nand2_1 _2903_ (.Y(_0396_),
    .A(net15),
    .B(_0394_));
 sg13g2_a21oi_1 _2904_ (.A1(_1629_),
    .A2(_1631_),
    .Y(_0397_),
    .B1(_1373_));
 sg13g2_nand2_1 _2905_ (.Y(_0398_),
    .A(_1410_),
    .B(_1604_));
 sg13g2_nand2_1 _2906_ (.Y(_0399_),
    .A(net54),
    .B(_0398_));
 sg13g2_o21ai_1 _2907_ (.B1(_0399_),
    .Y(_0400_),
    .A1(net63),
    .A2(_0397_));
 sg13g2_nand2_1 _2908_ (.Y(_0401_),
    .A(_0400_),
    .B(net26));
 sg13g2_o21ai_1 _2909_ (.B1(net54),
    .Y(_0402_),
    .A1(_1508_),
    .A2(_0101_));
 sg13g2_nand2_1 _2910_ (.Y(_0403_),
    .A(_1598_),
    .B(_1410_));
 sg13g2_nand2_1 _2911_ (.Y(_0404_),
    .A(_0403_),
    .B(net45));
 sg13g2_nand2_1 _2912_ (.Y(_0405_),
    .A(_0402_),
    .B(_0404_));
 sg13g2_nand2_1 _2913_ (.Y(_0407_),
    .A(_0405_),
    .B(net18));
 sg13g2_nand2_1 _2914_ (.Y(_0408_),
    .A(_0401_),
    .B(_0407_));
 sg13g2_nand2_1 _2915_ (.Y(_0409_),
    .A(_0408_),
    .B(net17));
 sg13g2_nand2_1 _2916_ (.Y(_0410_),
    .A(_0396_),
    .B(_0409_));
 sg13g2_nand2_1 _2917_ (.Y(_0411_),
    .A(_0410_),
    .B(net23));
 sg13g2_nor3_1 _2918_ (.A(_1491_),
    .B(_1390_),
    .C(net56),
    .Y(_0412_));
 sg13g2_nor2_1 _2919_ (.A(_1490_),
    .B(_1444_),
    .Y(_0413_));
 sg13g2_nor2_1 _2920_ (.A(_0413_),
    .B(_1500_),
    .Y(_0414_));
 sg13g2_nor2_1 _2921_ (.A(_0412_),
    .B(_0414_),
    .Y(_0415_));
 sg13g2_nand2_1 _2922_ (.Y(_0416_),
    .A(_0415_),
    .B(net19));
 sg13g2_nand2_1 _2923_ (.Y(_0418_),
    .A(_1447_),
    .B(_0079_));
 sg13g2_nand2_1 _2924_ (.Y(_0419_),
    .A(_0418_),
    .B(net58));
 sg13g2_o21ai_1 _2925_ (.B1(_0218_),
    .Y(_0420_),
    .A1(net38),
    .A2(_0068_));
 sg13g2_nand2_1 _2926_ (.Y(_0421_),
    .A(_0420_),
    .B(net37));
 sg13g2_nand2_1 _2927_ (.Y(_0422_),
    .A(_0419_),
    .B(_0421_));
 sg13g2_nand2_1 _2928_ (.Y(_0423_),
    .A(_0113_),
    .B(_0422_));
 sg13g2_nand2_1 _2929_ (.Y(_0424_),
    .A(_0416_),
    .B(_0423_));
 sg13g2_nand2_1 _2930_ (.Y(_0425_),
    .A(_0424_),
    .B(net22));
 sg13g2_o21ai_1 _2931_ (.B1(net60),
    .Y(_0426_),
    .A1(_1596_),
    .A2(_1443_));
 sg13g2_nand2_1 _2932_ (.Y(_0427_),
    .A(_1411_),
    .B(_1366_));
 sg13g2_nand2_1 _2933_ (.Y(_0429_),
    .A(_1520_),
    .B(_0427_));
 sg13g2_nand2_1 _2934_ (.Y(_0430_),
    .A(_0429_),
    .B(net58));
 sg13g2_nand2_1 _2935_ (.Y(_0431_),
    .A(_0426_),
    .B(_0430_));
 sg13g2_nand2_1 _2936_ (.Y(_0432_),
    .A(net35),
    .B(_0431_));
 sg13g2_nand2_1 _2937_ (.Y(_0433_),
    .A(net55),
    .B(_0320_));
 sg13g2_nand2_1 _2938_ (.Y(_0434_),
    .A(net29),
    .B(_0433_));
 sg13g2_nand2_1 _2939_ (.Y(_0435_),
    .A(_0432_),
    .B(_0434_));
 sg13g2_nand2_1 _2940_ (.Y(_0436_),
    .A(net17),
    .B(_0435_));
 sg13g2_nand2_1 _2941_ (.Y(_0437_),
    .A(_0425_),
    .B(_0436_));
 sg13g2_nand2_1 _2942_ (.Y(_0438_),
    .A(_0437_),
    .B(_1487_));
 sg13g2_nand2_1 _2943_ (.Y(_0440_),
    .A(_0411_),
    .B(_0438_));
 sg13g2_nand2_1 _2944_ (.Y(_0441_),
    .A(_0440_),
    .B(_1342_));
 sg13g2_nand3_1 _2945_ (.B(_0441_),
    .C(net10),
    .A(_0380_),
    .Y(_0442_));
 sg13g2_a221oi_1 _2946_ (.B2(_1378_),
    .C1(net13),
    .B1(_1671_),
    .A1(_1669_),
    .Y(_0443_),
    .A2(_0135_));
 sg13g2_o21ai_1 _2947_ (.B1(_1358_),
    .Y(_0444_),
    .A1(_1630_),
    .A2(_1363_));
 sg13g2_nor2_1 _2948_ (.A(_1455_),
    .B(_1578_),
    .Y(_0445_));
 sg13g2_nand2_1 _2949_ (.Y(_0446_),
    .A(_0445_),
    .B(_1586_));
 sg13g2_nand3_1 _2950_ (.B(_0065_),
    .C(_0338_),
    .A(_0446_),
    .Y(_0447_));
 sg13g2_o21ai_1 _2951_ (.B1(net13),
    .Y(_0448_),
    .A1(_1350_),
    .A2(_0447_));
 sg13g2_a21oi_1 _2952_ (.A1(_1350_),
    .A2(_0444_),
    .Y(_0449_),
    .B1(_0448_));
 sg13g2_nor2_1 _2953_ (.A(_0443_),
    .B(_0449_),
    .Y(_0451_));
 sg13g2_nor2b_1 _2954_ (.A(_1658_),
    .B_N(_0451_),
    .Y(_0452_));
 sg13g2_nor2_1 _2955_ (.A(_0186_),
    .B(_0452_),
    .Y(_0453_));
 sg13g2_a21oi_1 _2956_ (.A1(_0442_),
    .A2(_0453_),
    .Y(_0454_),
    .B1(_0175_));
 sg13g2_nor2_1 _2957_ (.A(_1365_),
    .B(net61),
    .Y(_0455_));
 sg13g2_nor2_1 _2958_ (.A(_0455_),
    .B(_1582_),
    .Y(_0456_));
 sg13g2_nor2_1 _2959_ (.A(net42),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_a21oi_1 _2960_ (.A1(_0218_),
    .A2(_0297_),
    .Y(_0458_),
    .B1(net44));
 sg13g2_nor3_1 _2961_ (.A(_0457_),
    .B(_0458_),
    .C(net27),
    .Y(_0459_));
 sg13g2_nand2_1 _2962_ (.Y(_0460_),
    .A(_0284_),
    .B(net66));
 sg13g2_nand2_1 _2963_ (.Y(_0462_),
    .A(net51),
    .B(_0460_));
 sg13g2_o21ai_1 _2964_ (.B1(_1466_),
    .Y(_0463_),
    .A1(_1580_),
    .A2(net68));
 sg13g2_o21ai_1 _2965_ (.B1(_1574_),
    .Y(_0464_),
    .A1(net33),
    .A2(_0463_));
 sg13g2_nand2_1 _2966_ (.Y(_0465_),
    .A(_0464_),
    .B(net39));
 sg13g2_nand3_1 _2967_ (.B(_0462_),
    .C(_0465_),
    .A(net27),
    .Y(_0466_));
 sg13g2_nand3b_1 _2968_ (.B(net14),
    .C(_0466_),
    .Y(_0467_),
    .A_N(_0459_));
 sg13g2_a21oi_1 _2969_ (.A1(net43),
    .A2(net69),
    .Y(_0468_),
    .B1(_0320_));
 sg13g2_nand2_1 _2970_ (.Y(_0469_),
    .A(_1364_),
    .B(_1519_));
 sg13g2_nor2_1 _2971_ (.A(_1603_),
    .B(net48),
    .Y(_0470_));
 sg13g2_a21oi_1 _2972_ (.A1(net43),
    .A2(_0469_),
    .Y(_0471_),
    .B1(_0470_));
 sg13g2_nor2_1 _2973_ (.A(net55),
    .B(_0471_),
    .Y(_0473_));
 sg13g2_a21oi_1 _2974_ (.A1(net39),
    .A2(_0468_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_a21oi_1 _2975_ (.A1(_1556_),
    .A2(_1424_),
    .Y(_0475_),
    .B1(net46));
 sg13g2_nand2_1 _2976_ (.Y(_0476_),
    .A(net53),
    .B(_0980_));
 sg13g2_nand2_1 _2977_ (.Y(_0477_),
    .A(net51),
    .B(_0476_));
 sg13g2_nand2_1 _2978_ (.Y(_0478_),
    .A(_1423_),
    .B(_1413_));
 sg13g2_nor2b_1 _2979_ (.A(_0477_),
    .B_N(_0478_),
    .Y(_0479_));
 sg13g2_o21ai_1 _2980_ (.B1(net20),
    .Y(_0480_),
    .A1(_0475_),
    .A2(_0479_));
 sg13g2_o21ai_1 _2981_ (.B1(_0480_),
    .Y(_0481_),
    .A1(net20),
    .A2(_0474_));
 sg13g2_nand2_1 _2982_ (.Y(_0482_),
    .A(_0481_),
    .B(net15));
 sg13g2_nand2_1 _2983_ (.Y(_0484_),
    .A(_0467_),
    .B(_0482_));
 sg13g2_nand2_1 _2984_ (.Y(_0485_),
    .A(_0484_),
    .B(net23));
 sg13g2_nand3_1 _2985_ (.B(_0364_),
    .C(_1585_),
    .A(_1494_),
    .Y(_0486_));
 sg13g2_a21oi_1 _2986_ (.A1(_0357_),
    .A2(_0486_),
    .Y(_0487_),
    .B1(_1554_));
 sg13g2_nand3_1 _2987_ (.B(_0388_),
    .C(_0185_),
    .A(net44),
    .Y(_0488_));
 sg13g2_a21oi_1 _2988_ (.A1(_1500_),
    .A2(_0488_),
    .Y(_0489_),
    .B1(net27));
 sg13g2_o21ai_1 _2989_ (.B1(net14),
    .Y(_0490_),
    .A1(_0487_),
    .A2(_0489_));
 sg13g2_nand2_1 _2990_ (.Y(_0491_),
    .A(net41),
    .B(_1631_));
 sg13g2_a21oi_1 _2991_ (.A1(_0218_),
    .A2(_0491_),
    .Y(_0492_),
    .B1(net47));
 sg13g2_o21ai_1 _2992_ (.B1(net57),
    .Y(_0493_),
    .A1(_1375_),
    .A2(_0363_));
 sg13g2_a21oi_1 _2993_ (.A1(net66),
    .A2(_0493_),
    .Y(_0495_),
    .B1(net63));
 sg13g2_nor2_1 _2994_ (.A(_0492_),
    .B(_0495_),
    .Y(_0496_));
 sg13g2_nor2_1 _2995_ (.A(_0496_),
    .B(net27),
    .Y(_0497_));
 sg13g2_a21oi_1 _2996_ (.A1(_1410_),
    .A2(_1420_),
    .Y(_0498_),
    .B1(net20));
 sg13g2_o21ai_1 _2997_ (.B1(net15),
    .Y(_0499_),
    .A1(_0497_),
    .A2(_0498_));
 sg13g2_nand2_1 _2998_ (.Y(_0500_),
    .A(_0490_),
    .B(_0499_));
 sg13g2_nand2_1 _2999_ (.Y(_0501_),
    .A(_0500_),
    .B(net11));
 sg13g2_nand2_1 _3000_ (.Y(_0502_),
    .A(_0485_),
    .B(_0501_));
 sg13g2_nand2_1 _3001_ (.Y(_0503_),
    .A(_0502_),
    .B(_1540_));
 sg13g2_a21oi_1 _3002_ (.A1(_1471_),
    .A2(_1446_),
    .Y(_0504_),
    .B1(_0413_));
 sg13g2_o21ai_1 _3003_ (.B1(_0275_),
    .Y(_0506_),
    .A1(_1409_),
    .A2(_0504_));
 sg13g2_nand2_1 _3004_ (.Y(_0507_),
    .A(_0506_),
    .B(net25));
 sg13g2_o21ai_1 _3005_ (.B1(net21),
    .Y(_0508_),
    .A1(_0079_),
    .A2(net31));
 sg13g2_a21oi_1 _3006_ (.A1(_0507_),
    .A2(_0508_),
    .Y(_0509_),
    .B1(net15));
 sg13g2_inv_1 _3007_ (.Y(_0510_),
    .A(_0218_));
 sg13g2_a21oi_1 _3008_ (.A1(net33),
    .A2(_1365_),
    .Y(_0511_),
    .B1(_0510_));
 sg13g2_o21ai_1 _3009_ (.B1(_0419_),
    .Y(_0512_),
    .A1(net50),
    .A2(_0511_));
 sg13g2_nand2_1 _3010_ (.Y(_0513_),
    .A(_0512_),
    .B(net25));
 sg13g2_nand2b_1 _3011_ (.Y(_0514_),
    .B(_1671_),
    .A_N(_1496_));
 sg13g2_o21ai_1 _3012_ (.B1(net39),
    .Y(_0515_),
    .A1(_1448_),
    .A2(net69));
 sg13g2_nand3_1 _3013_ (.B(_0514_),
    .C(_0515_),
    .A(net21),
    .Y(_0517_));
 sg13g2_nand2_1 _3014_ (.Y(_0518_),
    .A(_0513_),
    .B(_0517_));
 sg13g2_nand2_1 _3015_ (.Y(_0519_),
    .A(_0518_),
    .B(net16));
 sg13g2_nand3b_1 _3016_ (.B(_1488_),
    .C(_0519_),
    .Y(_0520_),
    .A_N(_0509_));
 sg13g2_nor2_1 _3017_ (.A(_1413_),
    .B(_0234_),
    .Y(_0521_));
 sg13g2_o21ai_1 _3018_ (.B1(net32),
    .Y(_0522_),
    .A1(_1468_),
    .A2(_0276_));
 sg13g2_o21ai_1 _3019_ (.B1(_0522_),
    .Y(_0523_),
    .A1(_0521_),
    .A2(_0096_));
 sg13g2_nand2_1 _3020_ (.Y(_0524_),
    .A(_0523_),
    .B(_1400_));
 sg13g2_nor2_1 _3021_ (.A(_1474_),
    .B(_1507_),
    .Y(_0525_));
 sg13g2_inv_1 _3022_ (.Y(_0526_),
    .A(_0026_));
 sg13g2_a21oi_1 _3023_ (.A1(_0526_),
    .A2(_1369_),
    .Y(_0528_),
    .B1(_0297_));
 sg13g2_o21ai_1 _3024_ (.B1(net39),
    .Y(_0529_),
    .A1(_0525_),
    .A2(_0528_));
 sg13g2_o21ai_1 _3025_ (.B1(_1617_),
    .Y(_0530_),
    .A1(_0177_),
    .A2(_1498_));
 sg13g2_nand2_1 _3026_ (.Y(_0531_),
    .A(_0529_),
    .B(_0530_));
 sg13g2_nand2_1 _3027_ (.Y(_0532_),
    .A(_0531_),
    .B(_1503_));
 sg13g2_a21oi_1 _3028_ (.A1(_0524_),
    .A2(_0532_),
    .Y(_0533_),
    .B1(net12));
 sg13g2_nand2b_1 _3029_ (.Y(_0534_),
    .B(_1420_),
    .A_N(_0177_));
 sg13g2_nand2_1 _3030_ (.Y(_0535_),
    .A(_1507_),
    .B(_1630_));
 sg13g2_nand3_1 _3031_ (.B(net66),
    .C(_0535_),
    .A(net32),
    .Y(_0536_));
 sg13g2_nand3_1 _3032_ (.B(_0534_),
    .C(_0536_),
    .A(net24),
    .Y(_0537_));
 sg13g2_a21oi_1 _3033_ (.A1(net33),
    .A2(_1623_),
    .Y(_0539_),
    .B1(_1609_));
 sg13g2_nor2_1 _3034_ (.A(_1510_),
    .B(_1458_),
    .Y(_0540_));
 sg13g2_o21ai_1 _3035_ (.B1(net40),
    .Y(_0541_),
    .A1(_0540_),
    .A2(_1373_));
 sg13g2_o21ai_1 _3036_ (.B1(_0541_),
    .Y(_0542_),
    .A1(net32),
    .A2(_0539_));
 sg13g2_nand2_1 _3037_ (.Y(_0543_),
    .A(_0542_),
    .B(net27));
 sg13g2_nand2_1 _3038_ (.Y(_0544_),
    .A(_0537_),
    .B(_0543_));
 sg13g2_a21oi_1 _3039_ (.A1(net12),
    .A2(_0544_),
    .Y(_0545_),
    .B1(_1487_));
 sg13g2_nand2b_1 _3040_ (.Y(_0546_),
    .B(_0545_),
    .A_N(_0533_));
 sg13g2_nand3_1 _3041_ (.B(_0546_),
    .C(_1342_),
    .A(_0520_),
    .Y(_0547_));
 sg13g2_nand3_1 _3042_ (.B(_0547_),
    .C(_1659_),
    .A(_0503_),
    .Y(_0548_));
 sg13g2_a21oi_1 _3043_ (.A1(_0446_),
    .A2(_0427_),
    .Y(_0550_),
    .B1(net50));
 sg13g2_a21oi_1 _3044_ (.A1(_0626_),
    .A2(_1669_),
    .Y(_0551_),
    .B1(_0550_));
 sg13g2_nor2_1 _3045_ (.A(_1400_),
    .B(_0551_),
    .Y(_0552_));
 sg13g2_nor3_1 _3046_ (.A(_0552_),
    .B(_1668_),
    .C(_1658_),
    .Y(_0553_));
 sg13g2_nor2_1 _3047_ (.A(_1661_),
    .B(_0553_),
    .Y(_0554_));
 sg13g2_nand2_1 _3048_ (.Y(_0555_),
    .A(_0548_),
    .B(_0554_));
 sg13g2_nand2_1 _3049_ (.Y(_0556_),
    .A(_0454_),
    .B(_0555_));
 sg13g2_nor2_1 _3050_ (.A(_0143_),
    .B(_1491_),
    .Y(_0557_));
 sg13g2_nor2_1 _3051_ (.A(net40),
    .B(_0557_),
    .Y(_0558_));
 sg13g2_o21ai_1 _3052_ (.B1(net19),
    .Y(_0559_),
    .A1(_0289_),
    .A2(_0558_));
 sg13g2_nand2_1 _3053_ (.Y(_0561_),
    .A(_0559_),
    .B(_0245_));
 sg13g2_nor2_1 _3054_ (.A(_1592_),
    .B(_0561_),
    .Y(_0562_));
 sg13g2_nor2_1 _3055_ (.A(_1487_),
    .B(_0562_),
    .Y(_0563_));
 sg13g2_nor2_1 _3056_ (.A(_1524_),
    .B(net38),
    .Y(_0564_));
 sg13g2_nor2_1 _3057_ (.A(_1666_),
    .B(_0564_),
    .Y(_0565_));
 sg13g2_nor2_1 _3058_ (.A(net34),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_a21oi_1 _3059_ (.A1(_1410_),
    .A2(_1527_),
    .Y(_0567_),
    .B1(net50));
 sg13g2_o21ai_1 _3060_ (.B1(net21),
    .Y(_0568_),
    .A1(_0566_),
    .A2(_0567_));
 sg13g2_nand2b_1 _3061_ (.Y(_0569_),
    .B(_0216_),
    .A_N(_1510_));
 sg13g2_inv_1 _3062_ (.Y(_0570_),
    .A(_1410_));
 sg13g2_a21oi_1 _3063_ (.A1(net33),
    .A2(_0569_),
    .Y(_0572_),
    .B1(_0570_));
 sg13g2_a21oi_1 _3064_ (.A1(net33),
    .A2(_1370_),
    .Y(_0573_),
    .B1(_1448_));
 sg13g2_nand2_1 _3065_ (.Y(_0574_),
    .A(_0573_),
    .B(net42));
 sg13g2_o21ai_1 _3066_ (.B1(_0574_),
    .Y(_0575_),
    .A1(net34),
    .A2(_0572_));
 sg13g2_nand2_1 _3067_ (.Y(_0576_),
    .A(_0575_),
    .B(net25));
 sg13g2_nand3_1 _3068_ (.B(_0568_),
    .C(_0576_),
    .A(net14),
    .Y(_0577_));
 sg13g2_nand2_1 _3069_ (.Y(_0578_),
    .A(_0563_),
    .B(_0577_));
 sg13g2_nor3_1 _3070_ (.A(_0564_),
    .B(_0445_),
    .C(_1419_),
    .Y(_0579_));
 sg13g2_nor2_1 _3071_ (.A(_1586_),
    .B(_1670_),
    .Y(_0580_));
 sg13g2_nor2_1 _3072_ (.A(_0579_),
    .B(_0580_),
    .Y(_0581_));
 sg13g2_nand2_1 _3073_ (.Y(_0583_),
    .A(_0581_),
    .B(net20));
 sg13g2_o21ai_1 _3074_ (.B1(net54),
    .Y(_0584_),
    .A1(_1468_),
    .A2(_0383_));
 sg13g2_nand2_1 _3075_ (.Y(_0585_),
    .A(_0584_),
    .B(_0426_));
 sg13g2_nand2_1 _3076_ (.Y(_0586_),
    .A(net27),
    .B(_0585_));
 sg13g2_nand2_1 _3077_ (.Y(_0587_),
    .A(_0583_),
    .B(_0586_));
 sg13g2_nand2_1 _3078_ (.Y(_0588_),
    .A(_0587_),
    .B(net15));
 sg13g2_o21ai_1 _3079_ (.B1(net63),
    .Y(_0589_),
    .A1(_0510_),
    .A2(_0233_));
 sg13g2_o21ai_1 _3080_ (.B1(net45),
    .Y(_0590_),
    .A1(_1412_),
    .A2(_0295_));
 sg13g2_nand2_1 _3081_ (.Y(_0591_),
    .A(_0589_),
    .B(_0590_));
 sg13g2_nand2_1 _3082_ (.Y(_0592_),
    .A(_0591_),
    .B(net30));
 sg13g2_nor2_1 _3083_ (.A(net69),
    .B(_1391_),
    .Y(_0594_));
 sg13g2_nor2_1 _3084_ (.A(_0594_),
    .B(net36),
    .Y(_0595_));
 sg13g2_nand2_1 _3085_ (.Y(_0596_),
    .A(net45),
    .B(_0079_));
 sg13g2_o21ai_1 _3086_ (.B1(_0596_),
    .Y(_0597_),
    .A1(_1408_),
    .A2(_0595_));
 sg13g2_nand2_1 _3087_ (.Y(_0598_),
    .A(_0597_),
    .B(net19));
 sg13g2_nand2_1 _3088_ (.Y(_0599_),
    .A(_0592_),
    .B(_0598_));
 sg13g2_nand2_1 _3089_ (.Y(_0600_),
    .A(_0599_),
    .B(net14));
 sg13g2_nand2_1 _3090_ (.Y(_0601_),
    .A(_0588_),
    .B(_0600_));
 sg13g2_nand2_1 _3091_ (.Y(_0602_),
    .A(_0601_),
    .B(net11));
 sg13g2_nand2_1 _3092_ (.Y(_0603_),
    .A(_0578_),
    .B(_0602_));
 sg13g2_nand2_1 _3093_ (.Y(_0605_),
    .A(_0603_),
    .B(_1342_));
 sg13g2_nand2_1 _3094_ (.Y(_0606_),
    .A(net57),
    .B(_1378_));
 sg13g2_nor2b_1 _3095_ (.A(net52),
    .B_N(_0606_),
    .Y(_0607_));
 sg13g2_a21oi_1 _3096_ (.A1(_0607_),
    .A2(_0202_),
    .Y(_0608_),
    .B1(_0207_));
 sg13g2_nand2_1 _3097_ (.Y(_0609_),
    .A(_0608_),
    .B(net20));
 sg13g2_nand2_1 _3098_ (.Y(_0610_),
    .A(_0128_),
    .B(_0168_));
 sg13g2_o21ai_1 _3099_ (.B1(_0610_),
    .Y(_0611_),
    .A1(net46),
    .A2(_1383_));
 sg13g2_nand2_1 _3100_ (.Y(_0612_),
    .A(net30),
    .B(_0611_));
 sg13g2_nand2_1 _3101_ (.Y(_0613_),
    .A(_0609_),
    .B(_0612_));
 sg13g2_nand2_1 _3102_ (.Y(_0614_),
    .A(_0613_),
    .B(_1563_));
 sg13g2_nor2b_1 _3103_ (.A(net43),
    .B_N(_0469_),
    .Y(_0616_));
 sg13g2_nor2_1 _3104_ (.A(_1541_),
    .B(net53),
    .Y(_0617_));
 sg13g2_nand2b_1 _3105_ (.Y(_0618_),
    .B(_0128_),
    .A_N(_0617_));
 sg13g2_o21ai_1 _3106_ (.B1(_0618_),
    .Y(_0619_),
    .A1(net47),
    .A2(_0616_));
 sg13g2_nand2_1 _3107_ (.Y(_0620_),
    .A(net30),
    .B(_0619_));
 sg13g2_nand2_1 _3108_ (.Y(_0621_),
    .A(_0149_),
    .B(_0618_));
 sg13g2_nand2_1 _3109_ (.Y(_0622_),
    .A(net19),
    .B(_0621_));
 sg13g2_nand2_1 _3110_ (.Y(_0623_),
    .A(_0620_),
    .B(_0622_));
 sg13g2_nand2_1 _3111_ (.Y(_0624_),
    .A(net14),
    .B(_0623_));
 sg13g2_nand2_1 _3112_ (.Y(_0625_),
    .A(_0614_),
    .B(_0624_));
 sg13g2_nand2_1 _3113_ (.Y(_0627_),
    .A(_0625_),
    .B(net11));
 sg13g2_o21ai_1 _3114_ (.B1(net45),
    .Y(_0628_),
    .A1(_1508_),
    .A2(_0068_));
 sg13g2_nand2_1 _3115_ (.Y(_0629_),
    .A(_1505_),
    .B(_0365_));
 sg13g2_nand2_1 _3116_ (.Y(_0630_),
    .A(_0628_),
    .B(_0629_));
 sg13g2_nand2_1 _3117_ (.Y(_0631_),
    .A(net30),
    .B(_0630_));
 sg13g2_o21ai_1 _3118_ (.B1(_0094_),
    .Y(_0632_),
    .A1(_1578_),
    .A2(_0078_));
 sg13g2_nand2_1 _3119_ (.Y(_0633_),
    .A(_0632_),
    .B(net37));
 sg13g2_nand2_1 _3120_ (.Y(_0634_),
    .A(_1526_),
    .B(_1444_));
 sg13g2_nand2_1 _3121_ (.Y(_0635_),
    .A(net52),
    .B(_0634_));
 sg13g2_nand2_1 _3122_ (.Y(_0636_),
    .A(_0633_),
    .B(_0635_));
 sg13g2_nand2_1 _3123_ (.Y(_0638_),
    .A(net18),
    .B(_0636_));
 sg13g2_nand2_1 _3124_ (.Y(_0639_),
    .A(_0631_),
    .B(_0638_));
 sg13g2_nand2_1 _3125_ (.Y(_0640_),
    .A(net22),
    .B(_0639_));
 sg13g2_o21ai_1 _3126_ (.B1(net56),
    .Y(_0641_),
    .A1(net43),
    .A2(_1565_));
 sg13g2_nor2_1 _3127_ (.A(_1415_),
    .B(_1455_),
    .Y(_0642_));
 sg13g2_inv_1 _3128_ (.Y(_0643_),
    .A(_0642_));
 sg13g2_nand2_1 _3129_ (.Y(_0644_),
    .A(net49),
    .B(_0643_));
 sg13g2_nand2_1 _3130_ (.Y(_0645_),
    .A(_0215_),
    .B(_0644_));
 sg13g2_nand2_1 _3131_ (.Y(_0646_),
    .A(_0645_),
    .B(net52));
 sg13g2_nand2_1 _3132_ (.Y(_0647_),
    .A(_0641_),
    .B(_0646_));
 sg13g2_nand2_1 _3133_ (.Y(_0649_),
    .A(net26),
    .B(_0647_));
 sg13g2_nand3_1 _3134_ (.B(_0185_),
    .C(_0258_),
    .A(_1349_),
    .Y(_0650_));
 sg13g2_nand2_1 _3135_ (.Y(_0651_),
    .A(net18),
    .B(_0650_));
 sg13g2_nand2_1 _3136_ (.Y(_0652_),
    .A(_0649_),
    .B(_0651_));
 sg13g2_nand2_1 _3137_ (.Y(_0653_),
    .A(net17),
    .B(_0652_));
 sg13g2_nand2_1 _3138_ (.Y(_0654_),
    .A(_0640_),
    .B(_0653_));
 sg13g2_nand2_1 _3139_ (.Y(_0655_),
    .A(_0654_),
    .B(net23));
 sg13g2_nand2_1 _3140_ (.Y(_0656_),
    .A(_0627_),
    .B(_0655_));
 sg13g2_nand2_1 _3141_ (.Y(_0657_),
    .A(_0656_),
    .B(_1540_));
 sg13g2_nand3_1 _3142_ (.B(_0657_),
    .C(net10),
    .A(_0605_),
    .Y(_0658_));
 sg13g2_inv_1 _3143_ (.Y(_0660_),
    .A(_0446_));
 sg13g2_o21ai_1 _3144_ (.B1(net31),
    .Y(_0661_),
    .A1(_1618_),
    .A2(_0660_));
 sg13g2_o21ai_1 _3145_ (.B1(_0661_),
    .Y(_0662_),
    .A1(_1665_),
    .A2(_1609_));
 sg13g2_nand2_1 _3146_ (.Y(_0663_),
    .A(_1420_),
    .B(net66));
 sg13g2_nor2_1 _3147_ (.A(_1666_),
    .B(_0066_),
    .Y(_0664_));
 sg13g2_a21oi_1 _3148_ (.A1(net31),
    .A2(_0664_),
    .Y(_0665_),
    .B1(net13));
 sg13g2_a22oi_1 _3149_ (.Y(_0666_),
    .B1(_0663_),
    .B2(_0665_),
    .A2(net13),
    .A1(_0662_));
 sg13g2_nor2b_1 _3150_ (.A(net10),
    .B_N(_0666_),
    .Y(_0667_));
 sg13g2_nor2_1 _3151_ (.A(_1661_),
    .B(_0667_),
    .Y(_0668_));
 sg13g2_nand2_1 _3152_ (.Y(_0669_),
    .A(_0658_),
    .B(_0668_));
 sg13g2_nand2_1 _3153_ (.Y(_0671_),
    .A(_1447_),
    .B(_0093_));
 sg13g2_nand2_1 _3154_ (.Y(_0672_),
    .A(_0671_),
    .B(net63));
 sg13g2_nand2_1 _3155_ (.Y(_0673_),
    .A(_0672_),
    .B(_1469_));
 sg13g2_nand2_1 _3156_ (.Y(_0674_),
    .A(net30),
    .B(_0673_));
 sg13g2_nand2_1 _3157_ (.Y(_0675_),
    .A(_0240_),
    .B(_0065_));
 sg13g2_nand2_1 _3158_ (.Y(_0676_),
    .A(_1349_),
    .B(_0675_));
 sg13g2_nand2_1 _3159_ (.Y(_0677_),
    .A(_0246_),
    .B(_0168_));
 sg13g2_nand2_1 _3160_ (.Y(_0678_),
    .A(net45),
    .B(_0677_));
 sg13g2_nand2_1 _3161_ (.Y(_0679_),
    .A(_0676_),
    .B(_0678_));
 sg13g2_nand2_1 _3162_ (.Y(_0680_),
    .A(net19),
    .B(_0679_));
 sg13g2_nand2_1 _3163_ (.Y(_0682_),
    .A(_0674_),
    .B(_0680_));
 sg13g2_nand2_1 _3164_ (.Y(_0683_),
    .A(_1563_),
    .B(_0682_));
 sg13g2_o21ai_1 _3165_ (.B1(net45),
    .Y(_0684_),
    .A1(_0206_),
    .A2(_1373_));
 sg13g2_nand2_1 _3166_ (.Y(_0685_),
    .A(_0493_),
    .B(_0223_));
 sg13g2_nand2_1 _3167_ (.Y(_0686_),
    .A(_0685_),
    .B(_1505_));
 sg13g2_nand2_1 _3168_ (.Y(_0687_),
    .A(_0684_),
    .B(_0686_));
 sg13g2_nand2_1 _3169_ (.Y(_0688_),
    .A(_1399_),
    .B(_0687_));
 sg13g2_a21oi_1 _3170_ (.A1(net41),
    .A2(_1416_),
    .Y(_0689_),
    .B1(_1629_));
 sg13g2_o21ai_1 _3171_ (.B1(_0462_),
    .Y(_0690_),
    .A1(net46),
    .A2(_0689_));
 sg13g2_nand2_1 _3172_ (.Y(_0691_),
    .A(_0690_),
    .B(net19));
 sg13g2_nand2_1 _3173_ (.Y(_0693_),
    .A(_0688_),
    .B(_0691_));
 sg13g2_nand2_1 _3174_ (.Y(_0694_),
    .A(_0693_),
    .B(net14));
 sg13g2_nand2_1 _3175_ (.Y(_0695_),
    .A(_0683_),
    .B(_0694_));
 sg13g2_nand2_1 _3176_ (.Y(_0696_),
    .A(_0695_),
    .B(net23));
 sg13g2_o21ai_1 _3177_ (.B1(net54),
    .Y(_0697_),
    .A1(_1468_),
    .A2(_0066_));
 sg13g2_nand3_1 _3178_ (.B(_1413_),
    .C(_1548_),
    .A(net37),
    .Y(_0698_));
 sg13g2_nand2_1 _3179_ (.Y(_0699_),
    .A(_0697_),
    .B(_0698_));
 sg13g2_nand2_1 _3180_ (.Y(_0700_),
    .A(_0699_),
    .B(net26));
 sg13g2_nor2_1 _3181_ (.A(_0134_),
    .B(_1567_),
    .Y(_0701_));
 sg13g2_o21ai_1 _3182_ (.B1(_0477_),
    .Y(_0702_),
    .A1(net46),
    .A2(_0701_));
 sg13g2_nand2_1 _3183_ (.Y(_0704_),
    .A(_0702_),
    .B(net18));
 sg13g2_nand2_1 _3184_ (.Y(_0705_),
    .A(_0700_),
    .B(_0704_));
 sg13g2_nand2_1 _3185_ (.Y(_0706_),
    .A(net22),
    .B(_0705_));
 sg13g2_o21ai_1 _3186_ (.B1(_1460_),
    .Y(_0707_),
    .A1(_0080_),
    .A2(_0060_));
 sg13g2_nand2_1 _3187_ (.Y(_0708_),
    .A(net52),
    .B(_0203_));
 sg13g2_nand2_1 _3188_ (.Y(_0709_),
    .A(_0707_),
    .B(_0708_));
 sg13g2_nand2_1 _3189_ (.Y(_0710_),
    .A(net26),
    .B(_0709_));
 sg13g2_nand2b_1 _3190_ (.Y(_0711_),
    .B(net55),
    .A_N(_1597_));
 sg13g2_nand2_1 _3191_ (.Y(_0712_),
    .A(net18),
    .B(_0711_));
 sg13g2_nand2_1 _3192_ (.Y(_0713_),
    .A(_0710_),
    .B(_0712_));
 sg13g2_nand2_1 _3193_ (.Y(_0715_),
    .A(net17),
    .B(_0713_));
 sg13g2_nand2_1 _3194_ (.Y(_0716_),
    .A(_0706_),
    .B(_0715_));
 sg13g2_nand2_1 _3195_ (.Y(_0717_),
    .A(_0716_),
    .B(_1487_));
 sg13g2_nand2_1 _3196_ (.Y(_0718_),
    .A(_0696_),
    .B(_0717_));
 sg13g2_nand2_1 _3197_ (.Y(_0719_),
    .A(_0718_),
    .B(_1342_));
 sg13g2_nor2_1 _3198_ (.A(_1618_),
    .B(_0570_),
    .Y(_0720_));
 sg13g2_o21ai_1 _3199_ (.B1(_0610_),
    .Y(_0721_),
    .A1(_1388_),
    .A2(_0720_));
 sg13g2_nand2_1 _3200_ (.Y(_0722_),
    .A(net26),
    .B(_0721_));
 sg13g2_o21ai_1 _3201_ (.B1(net37),
    .Y(_0723_),
    .A1(_1600_),
    .A2(_0276_));
 sg13g2_nand2_1 _3202_ (.Y(_0724_),
    .A(_0723_),
    .B(_0179_));
 sg13g2_nand2_1 _3203_ (.Y(_0726_),
    .A(_0724_),
    .B(net18));
 sg13g2_nand2_1 _3204_ (.Y(_0727_),
    .A(_0722_),
    .B(_0726_));
 sg13g2_nand2_1 _3205_ (.Y(_0728_),
    .A(net22),
    .B(_0727_));
 sg13g2_nand2_1 _3206_ (.Y(_0729_),
    .A(_0444_),
    .B(_1492_));
 sg13g2_nand2_1 _3207_ (.Y(_0730_),
    .A(_0729_),
    .B(_0083_));
 sg13g2_nand2_1 _3208_ (.Y(_0731_),
    .A(_1583_),
    .B(_0240_));
 sg13g2_nand2_1 _3209_ (.Y(_0732_),
    .A(_0731_),
    .B(_1451_));
 sg13g2_nand2_1 _3210_ (.Y(_0733_),
    .A(_0730_),
    .B(_0732_));
 sg13g2_nand2_1 _3211_ (.Y(_0734_),
    .A(_0113_),
    .B(_0733_));
 sg13g2_nand2_1 _3212_ (.Y(_0735_),
    .A(_1600_),
    .B(_1392_));
 sg13g2_nand2_1 _3213_ (.Y(_0737_),
    .A(_0735_),
    .B(_0059_));
 sg13g2_nand2_1 _3214_ (.Y(_0738_),
    .A(_0737_),
    .B(net58));
 sg13g2_nand2_1 _3215_ (.Y(_0739_),
    .A(_0738_),
    .B(_0269_));
 sg13g2_nand2_1 _3216_ (.Y(_0740_),
    .A(_0104_),
    .B(_0739_));
 sg13g2_nand2_1 _3217_ (.Y(_0741_),
    .A(_0734_),
    .B(_0740_));
 sg13g2_nand2_1 _3218_ (.Y(_0742_),
    .A(net17),
    .B(_0741_));
 sg13g2_nand2_1 _3219_ (.Y(_0743_),
    .A(_0728_),
    .B(_0742_));
 sg13g2_nand2_1 _3220_ (.Y(_0744_),
    .A(_0743_),
    .B(_1487_));
 sg13g2_nand2_1 _3221_ (.Y(_0745_),
    .A(_0178_),
    .B(_0606_));
 sg13g2_nand2_1 _3222_ (.Y(_0746_),
    .A(_0745_),
    .B(net37));
 sg13g2_nand2_1 _3223_ (.Y(_0748_),
    .A(_1558_),
    .B(_0297_));
 sg13g2_nand2_1 _3224_ (.Y(_0749_),
    .A(net52),
    .B(_0748_));
 sg13g2_nand2_1 _3225_ (.Y(_0750_),
    .A(_0746_),
    .B(_0749_));
 sg13g2_nand2_1 _3226_ (.Y(_0751_),
    .A(net26),
    .B(_0750_));
 sg13g2_o21ai_1 _3227_ (.B1(_0094_),
    .Y(_0752_),
    .A1(net53),
    .A2(_0594_));
 sg13g2_nand2_1 _3228_ (.Y(_0753_),
    .A(_0752_),
    .B(net56));
 sg13g2_nand2_1 _3229_ (.Y(_0754_),
    .A(_1526_),
    .B(_1556_));
 sg13g2_nand2_1 _3230_ (.Y(_0755_),
    .A(net58),
    .B(_0754_));
 sg13g2_nand2_1 _3231_ (.Y(_0756_),
    .A(_0753_),
    .B(_0755_));
 sg13g2_nand2_1 _3232_ (.Y(_0757_),
    .A(net29),
    .B(_0756_));
 sg13g2_nand2_1 _3233_ (.Y(_0759_),
    .A(_0751_),
    .B(_0757_));
 sg13g2_nand2_1 _3234_ (.Y(_0760_),
    .A(net22),
    .B(_0759_));
 sg13g2_nand2_1 _3235_ (.Y(_0761_),
    .A(_0069_),
    .B(_1610_));
 sg13g2_nand2_1 _3236_ (.Y(_0762_),
    .A(_1460_),
    .B(_0761_));
 sg13g2_nand2_1 _3237_ (.Y(_0763_),
    .A(_1570_),
    .B(_0637_));
 sg13g2_nor2b_1 _3238_ (.A(net53),
    .B_N(_0763_),
    .Y(_0764_));
 sg13g2_nand3_1 _3239_ (.B(_1385_),
    .C(_0764_),
    .A(_1384_),
    .Y(_0765_));
 sg13g2_nand2_1 _3240_ (.Y(_0766_),
    .A(_0762_),
    .B(_0765_));
 sg13g2_nand3_1 _3241_ (.B(_1404_),
    .C(_1403_),
    .A(_0766_),
    .Y(_0767_));
 sg13g2_nand2b_1 _3242_ (.Y(_0768_),
    .B(_0258_),
    .A_N(_0455_));
 sg13g2_nand2_1 _3243_ (.Y(_0770_),
    .A(_0768_),
    .B(net58));
 sg13g2_nor2_1 _3244_ (.A(_0569_),
    .B(net59),
    .Y(_0771_));
 sg13g2_a21oi_1 _3245_ (.A1(net53),
    .A2(_1467_),
    .Y(_0772_),
    .B1(_0771_));
 sg13g2_nand2_1 _3246_ (.Y(_0773_),
    .A(_0772_),
    .B(net51));
 sg13g2_nand2_1 _3247_ (.Y(_0774_),
    .A(_0770_),
    .B(_0773_));
 sg13g2_nand2_1 _3248_ (.Y(_0775_),
    .A(_1406_),
    .B(_0774_));
 sg13g2_nand2_1 _3249_ (.Y(_0776_),
    .A(_0767_),
    .B(_0775_));
 sg13g2_nand2_1 _3250_ (.Y(_0777_),
    .A(_1434_),
    .B(_0776_));
 sg13g2_nand2_1 _3251_ (.Y(_0778_),
    .A(_0760_),
    .B(_0777_));
 sg13g2_nand2_1 _3252_ (.Y(_0779_),
    .A(_0778_),
    .B(_1437_));
 sg13g2_nand2_1 _3253_ (.Y(_0780_),
    .A(_0744_),
    .B(_0779_));
 sg13g2_nand2_1 _3254_ (.Y(_0781_),
    .A(_0780_),
    .B(_1540_));
 sg13g2_nand3_1 _3255_ (.B(_0781_),
    .C(_1659_),
    .A(_0719_),
    .Y(_0782_));
 sg13g2_or2_1 _3256_ (.X(_0783_),
    .B(_0550_),
    .A(_0283_));
 sg13g2_a22oi_1 _3257_ (.Y(_0784_),
    .B1(_1664_),
    .B2(_0665_),
    .A2(_0783_),
    .A1(net13));
 sg13g2_nor2b_1 _3258_ (.A(_1658_),
    .B_N(_0784_),
    .Y(_0785_));
 sg13g2_nor2_1 _3259_ (.A(_0186_),
    .B(_0785_),
    .Y(_0786_));
 sg13g2_nand2_1 _3260_ (.Y(_0787_),
    .A(_0782_),
    .B(_0786_));
 sg13g2_nand3_1 _3261_ (.B(_0787_),
    .C(_0175_),
    .A(_0669_),
    .Y(_0788_));
 sg13g2_nand3_1 _3262_ (.B(_0788_),
    .C(\g_x[2] ),
    .A(_0556_),
    .Y(_0789_));
 sg13g2_nand2_2 _3263_ (.Y(_0791_),
    .A(_0317_),
    .B(_0789_));
 sg13g2_xor2_1 _3264_ (.B(_1043_),
    .A(_0025_),
    .X(_0792_));
 sg13g2_nor2_2 _3265_ (.A(net78),
    .B(_0307_),
    .Y(_0793_));
 sg13g2_o21ai_1 _3266_ (.B1(_0793_),
    .Y(_0794_),
    .A1(_0025_),
    .A2(_1043_));
 sg13g2_nor2_1 _3267_ (.A(_0314_),
    .B(_1040_),
    .Y(_0795_));
 sg13g2_a21oi_1 _3268_ (.A1(_0023_),
    .A2(_1040_),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_o21ai_1 _3269_ (.B1(_0891_),
    .Y(_0797_),
    .A1(_0794_),
    .A2(_0796_));
 sg13g2_nor3_1 _3270_ (.A(net78),
    .B(_0797_),
    .C(_1202_),
    .Y(_0798_));
 sg13g2_nand2_1 _3271_ (.Y(_0799_),
    .A(_0891_),
    .B(_0793_));
 sg13g2_inv_1 _3272_ (.Y(_0800_),
    .A(_0799_));
 sg13g2_nor2_1 _3273_ (.A(_1147_),
    .B(_1040_),
    .Y(_0801_));
 sg13g2_a21oi_1 _3274_ (.A1(_0022_),
    .A2(_1040_),
    .Y(_0802_),
    .B1(_0801_));
 sg13g2_and3_1 _3275_ (.X(_0803_),
    .A(_1234_),
    .B(_0800_),
    .C(_0802_));
 sg13g2_nor3_1 _3276_ (.A(_0792_),
    .B(_0798_),
    .C(_0803_),
    .Y(_0804_));
 sg13g2_nor2_1 _3277_ (.A(_0893_),
    .B(_0793_),
    .Y(_0805_));
 sg13g2_a21oi_1 _3278_ (.A1(_0800_),
    .A2(_0025_),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_xor2_1 _3279_ (.B(_1043_),
    .A(_0793_),
    .X(_0807_));
 sg13g2_a21oi_1 _3280_ (.A1(net76),
    .A2(_0307_),
    .Y(_0808_),
    .B1(_0807_));
 sg13g2_nor2b_1 _3281_ (.A(_0796_),
    .B_N(_0807_),
    .Y(_0809_));
 sg13g2_o21ai_1 _3282_ (.B1(_0799_),
    .Y(_0810_),
    .A1(_0808_),
    .A2(_0809_));
 sg13g2_nand3_1 _3283_ (.B(_0806_),
    .C(_0810_),
    .A(_1155_),
    .Y(_0812_));
 sg13g2_a22oi_1 _3284_ (.Y(_0813_),
    .B1(_0807_),
    .B2(_0802_),
    .A2(_0800_),
    .A1(_0314_));
 sg13g2_nor2_1 _3285_ (.A(_0805_),
    .B(_0813_),
    .Y(_0814_));
 sg13g2_nand3_1 _3286_ (.B(_1189_),
    .C(_0814_),
    .A(_1188_),
    .Y(_0815_));
 sg13g2_nand3_1 _3287_ (.B(_0812_),
    .C(_0815_),
    .A(_0804_),
    .Y(_0816_));
 sg13g2_buf_1 _3288_ (.A(_0816_),
    .X(_0817_));
 sg13g2_buf_2 _3289_ (.A(ui_in[1]),
    .X(_0818_));
 sg13g2_xnor2_1 _3290_ (.Y(_0819_),
    .A(_1131_),
    .B(_1142_));
 sg13g2_nor2_1 _3291_ (.A(net76),
    .B(_1234_),
    .Y(_0820_));
 sg13g2_a21oi_1 _3292_ (.A1(net76),
    .A2(_0819_),
    .Y(_0821_),
    .B1(_0820_));
 sg13g2_nor2_1 _3293_ (.A(net77),
    .B(_0821_),
    .Y(_0823_));
 sg13g2_a21oi_2 _3294_ (.B1(_0823_),
    .Y(_0824_),
    .A2(net77),
    .A1(_1219_));
 sg13g2_nand2_1 _3295_ (.Y(_0825_),
    .A(_1236_),
    .B(net77));
 sg13g2_nand2_1 _3296_ (.Y(_0826_),
    .A(_0819_),
    .B(net78));
 sg13g2_xor2_1 _3297_ (.B(_1173_),
    .A(_1140_),
    .X(_0827_));
 sg13g2_nand2_1 _3298_ (.Y(_0828_),
    .A(_0827_),
    .B(_0164_));
 sg13g2_nand3_1 _3299_ (.B(_0828_),
    .C(_0131_),
    .A(_0826_),
    .Y(_0829_));
 sg13g2_nand2_1 _3300_ (.Y(_0830_),
    .A(_0825_),
    .B(_0829_));
 sg13g2_nand2_1 _3301_ (.Y(_0831_),
    .A(_0824_),
    .B(_0830_));
 sg13g2_buf_1 _3302_ (.A(ui_in[0]),
    .X(_0832_));
 sg13g2_nand2_1 _3303_ (.Y(_0834_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_nor2_1 _3304_ (.A(_0818_),
    .B(_0834_),
    .Y(_0835_));
 sg13g2_inv_1 _3305_ (.Y(_0836_),
    .A(_0832_));
 sg13g2_inv_1 _3306_ (.Y(_0837_),
    .A(_0818_));
 sg13g2_nand2_1 _3307_ (.Y(_0838_),
    .A(_0827_),
    .B(_1016_));
 sg13g2_xnor2_1 _3308_ (.Y(_0839_),
    .A(_1038_),
    .B(_1134_));
 sg13g2_a21oi_1 _3309_ (.A1(_0839_),
    .A2(_0164_),
    .Y(_0840_),
    .B1(net77));
 sg13g2_a22oi_1 _3310_ (.Y(_0841_),
    .B1(net77),
    .B2(_0821_),
    .A2(_0840_),
    .A1(_0838_));
 sg13g2_inv_1 _3311_ (.Y(_0842_),
    .A(_0830_));
 sg13g2_nor2_1 _3312_ (.A(_0841_),
    .B(_0842_),
    .Y(_0843_));
 sg13g2_nor2_1 _3313_ (.A(_0842_),
    .B(_0824_),
    .Y(_0845_));
 sg13g2_nor4_1 _3314_ (.A(_0836_),
    .B(_0837_),
    .C(_0843_),
    .D(_0845_),
    .Y(_0846_));
 sg13g2_nand3_1 _3315_ (.B(_0827_),
    .C(_0839_),
    .A(_0819_),
    .Y(_0847_));
 sg13g2_inv_1 _3316_ (.Y(_0848_),
    .A(_0841_));
 sg13g2_nor2_1 _3317_ (.A(_0830_),
    .B(_0848_),
    .Y(_0849_));
 sg13g2_inv_1 _3318_ (.Y(_0850_),
    .A(_0849_));
 sg13g2_nor2_1 _3319_ (.A(_0824_),
    .B(_0850_),
    .Y(_0851_));
 sg13g2_inv_1 _3320_ (.Y(_0852_),
    .A(_0851_));
 sg13g2_a21oi_1 _3321_ (.A1(_0832_),
    .A2(_0847_),
    .Y(_0853_),
    .B1(_0852_));
 sg13g2_nor3_1 _3322_ (.A(_0835_),
    .B(_0846_),
    .C(_0853_),
    .Y(_0854_));
 sg13g2_nor2_1 _3323_ (.A(_0817_),
    .B(_0854_),
    .Y(_0856_));
 sg13g2_nor2b_1 _3324_ (.A(_0791_),
    .B_N(_0856_),
    .Y(net2));
 sg13g2_nor2_1 _3325_ (.A(_0824_),
    .B(_0843_),
    .Y(_0857_));
 sg13g2_nor2_1 _3326_ (.A(_0830_),
    .B(_0824_),
    .Y(_0858_));
 sg13g2_nand2_1 _3327_ (.Y(_0859_),
    .A(_0858_),
    .B(_0836_));
 sg13g2_o21ai_1 _3328_ (.B1(_0859_),
    .Y(_0860_),
    .A1(_0857_),
    .A2(_0834_));
 sg13g2_nor2_2 _3329_ (.A(_0847_),
    .B(_0852_),
    .Y(_0861_));
 sg13g2_a21oi_1 _3330_ (.A1(_0860_),
    .A2(_0818_),
    .Y(_0862_),
    .B1(_0861_));
 sg13g2_nand2_1 _3331_ (.Y(_0863_),
    .A(_0831_),
    .B(_0836_));
 sg13g2_inv_1 _3332_ (.Y(_0864_),
    .A(_0863_));
 sg13g2_o21ai_1 _3333_ (.B1(_0837_),
    .Y(_0866_),
    .A1(_0864_),
    .A2(_0851_));
 sg13g2_a21oi_1 _3334_ (.A1(_0862_),
    .A2(_0866_),
    .Y(_0867_),
    .B1(_0817_));
 sg13g2_nor2b_1 _3335_ (.A(_0791_),
    .B_N(_0867_),
    .Y(net3));
 sg13g2_o21ai_1 _3336_ (.B1(_0818_),
    .Y(_0868_),
    .A1(_0857_),
    .A2(_0864_));
 sg13g2_nand2_1 _3337_ (.Y(_0869_),
    .A(_0858_),
    .B(_0837_));
 sg13g2_a21oi_1 _3338_ (.A1(_0868_),
    .A2(_0869_),
    .Y(_0870_),
    .B1(_0817_));
 sg13g2_nor2b_1 _3339_ (.A(_0791_),
    .B_N(_0870_),
    .Y(net4));
 sg13g2_nand2_1 _3340_ (.Y(_0871_),
    .A(_0824_),
    .B(_0848_));
 sg13g2_inv_1 _3341_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_nand2_1 _3342_ (.Y(_0873_),
    .A(_0842_),
    .B(_0818_));
 sg13g2_nor2_1 _3343_ (.A(_0837_),
    .B(_0824_),
    .Y(_0874_));
 sg13g2_a21oi_1 _3344_ (.A1(_0872_),
    .A2(_0873_),
    .Y(_0875_),
    .B1(_0874_));
 sg13g2_o21ai_1 _3345_ (.B1(_0832_),
    .Y(_0876_),
    .A1(_0849_),
    .A2(_0875_));
 sg13g2_nor3_1 _3346_ (.A(_0824_),
    .B(_0843_),
    .C(_0849_),
    .Y(_0877_));
 sg13g2_a21oi_1 _3347_ (.A1(_0836_),
    .A2(_0877_),
    .Y(_0878_),
    .B1(_0861_));
 sg13g2_a21oi_1 _3348_ (.A1(_0876_),
    .A2(_0878_),
    .Y(_0879_),
    .B1(_0817_));
 sg13g2_nor2b_1 _3349_ (.A(_0791_),
    .B_N(_0879_),
    .Y(net6));
 sg13g2_nor2_1 _3350_ (.A(_0858_),
    .B(_0834_),
    .Y(_0880_));
 sg13g2_a22oi_1 _3351_ (.Y(_0881_),
    .B1(_0841_),
    .B2(_0880_),
    .A2(_0845_),
    .A1(_0836_));
 sg13g2_nor2_1 _3352_ (.A(_0837_),
    .B(_0861_),
    .Y(_0882_));
 sg13g2_nor2_1 _3353_ (.A(_0832_),
    .B(_0872_),
    .Y(_0884_));
 sg13g2_nor3_1 _3354_ (.A(_0818_),
    .B(_0884_),
    .C(_0861_),
    .Y(_0885_));
 sg13g2_nand2_1 _3355_ (.Y(_0886_),
    .A(_0877_),
    .B(_0832_));
 sg13g2_a221oi_1 _3356_ (.B2(_0886_),
    .C1(_0817_),
    .B1(_0885_),
    .A1(_0881_),
    .Y(_0887_),
    .A2(_0882_));
 sg13g2_nor2b_1 _3357_ (.A(_0791_),
    .B_N(_0887_),
    .Y(net7));
 sg13g2_a221oi_1 _3358_ (.B2(_0874_),
    .C1(_0861_),
    .B1(_0841_),
    .A1(_0845_),
    .Y(_0888_),
    .A2(_0837_));
 sg13g2_nand2_1 _3359_ (.Y(_0889_),
    .A(_0884_),
    .B(_0818_));
 sg13g2_a21oi_1 _3360_ (.A1(_0888_),
    .A2(_0889_),
    .Y(_0890_),
    .B1(_0817_));
 sg13g2_nor2b_1 _3361_ (.A(_0791_),
    .B_N(_0890_),
    .Y(net8));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_buf_1 _3364_ (.A(net85),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3365_ (.A(net86),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3366_ (.A(net87),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3367_ (.A(net88),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3368_ (.A(net89),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3369_ (.A(net90),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3370_ (.A(net91),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3371_ (.A(net92),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3372_ (.A(net93),
    .X(uio_out[0]));
 sg13g2_buf_1 _3373_ (.A(net94),
    .X(uio_out[1]));
 sg13g2_buf_1 _3374_ (.A(net95),
    .X(uio_out[2]));
 sg13g2_buf_1 _3375_ (.A(net96),
    .X(uio_out[3]));
 sg13g2_buf_1 _3376_ (.A(net97),
    .X(uio_out[4]));
 sg13g2_buf_1 _3377_ (.A(net98),
    .X(uio_out[5]));
 sg13g2_buf_1 _3378_ (.A(net99),
    .X(uio_out[6]));
 sg13g2_buf_1 _3379_ (.A(net100),
    .X(uio_out[7]));
 sg13g2_buf_1 _3380_ (.A(\hvsync_gen.vsync ),
    .X(net5));
 sg13g2_buf_1 _3381_ (.A(hsync),
    .X(net9));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net101),
    .D(_0029_),
    .Q_N(_0027_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net102),
    .D(_0030_),
    .Q_N(_1689_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net103),
    .D(_0031_),
    .Q_N(_1688_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net104),
    .D(_0032_),
    .Q_N(_0017_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(\hvsync_gen.vsync ),
    .RESET_B(net105),
    .D(_0033_),
    .Q_N(_0015_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net106),
    .D(_0034_),
    .Q_N(_0016_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net107),
    .D(_0035_),
    .Q_N(_0019_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net108),
    .D(_0036_),
    .Q_N(_0020_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net109),
    .D(_0037_),
    .Q_N(_0021_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(net84),
    .RESET_B(net110),
    .D(_0038_),
    .Q_N(_1687_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net111),
    .D(_0039_),
    .Q_N(_0028_),
    .Q(\g_x[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net112),
    .D(_0040_),
    .Q_N(_1686_),
    .Q(\g_x[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net113),
    .D(_0041_),
    .Q_N(_1685_),
    .Q(\g_x[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net114),
    .D(_0042_),
    .Q_N(_1684_),
    .Q(\a[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net115),
    .D(_0043_),
    .Q_N(_0018_),
    .Q(\a[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net116),
    .D(_0044_),
    .Q_N(_0022_),
    .Q(\b[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PN0_  (.CLK(clknet_2_2__leaf_clk),
    .RESET_B(net117),
    .D(_0045_),
    .Q_N(_0023_),
    .Q(\b[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net118),
    .D(_0046_),
    .Q_N(_0024_),
    .Q(\b[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net119),
    .D(_0047_),
    .Q_N(_0025_),
    .Q(\b[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PN0_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net120),
    .D(_0048_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net121),
    .D(_0006_),
    .Q_N(_1683_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net122),
    .D(_0049_),
    .Q_N(_0026_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0N_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net123),
    .D(_0050_),
    .Q_N(_1682_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net124),
    .D(_0051_),
    .Q_N(_0010_),
    .Q(\div3.in[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net125),
    .D(_0052_),
    .Q_N(_0011_),
    .Q(\div3.in[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net126),
    .D(_0053_),
    .Q_N(_0012_),
    .Q(\div3.in[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net127),
    .D(_0054_),
    .Q_N(_0013_),
    .Q(\div3.in[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net128),
    .D(_0055_),
    .Q_N(_0014_),
    .Q(\div3.in[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0N_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net129),
    .D(_0056_),
    .Q_N(_1681_),
    .Q(\div3.in[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0N_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net130),
    .D(_0057_),
    .Q_N(_0008_),
    .Q(\div3.in[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0N_  (.CLK(clknet_2_0__leaf_clk),
    .RESET_B(net131),
    .D(_0058_),
    .Q_N(_1690_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net132),
    .D(_0007_),
    .Q_N(_1691_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \yb[0]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net133),
    .D(_0000_),
    .Q_N(_1692_),
    .Q(\div3.out[0] ));
 sg13g2_dfrbp_1 \yb[1]$_DFF_P_  (.CLK(clknet_2_3__leaf_clk),
    .RESET_B(net134),
    .D(_0001_),
    .Q_N(_1693_),
    .Q(\div3.out[1] ));
 sg13g2_dfrbp_1 \yb[2]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net135),
    .D(_0002_),
    .Q_N(_1694_),
    .Q(\div3.out[2] ));
 sg13g2_dfrbp_1 \yb[3]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net136),
    .D(_0003_),
    .Q_N(_1695_),
    .Q(\div3.out[3] ));
 sg13g2_dfrbp_1 \yb[4]$_DFF_P_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net137),
    .D(_0004_),
    .Q_N(_1680_),
    .Q(\div3.out[4] ));
 sg13g2_dfrbp_1 \yb[5]$_SDFF_PN0_  (.CLK(clknet_2_1__leaf_clk),
    .RESET_B(net138),
    .D(_0005_),
    .Q_N(_1679_),
    .Q(\div3.out[5] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uo_out[0]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[1]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[2]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[3]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[4]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[5]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[6]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout10 (.A(_1659_),
    .X(net10));
 sg13g2_buf_2 fanout11 (.A(_1488_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_1435_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_0200_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_1592_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1563_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_1441_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1434_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0104_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0063_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_1554_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1503_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_1440_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_1438_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_1407_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1400_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0113_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1552_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1465_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1406_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1399_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1665_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1617_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1507_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1409_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1398_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1359_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0083_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1596_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1506_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1494_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1473_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1461_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1458_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1452_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1419_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1408_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1388_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1382_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1358_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1350_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0128_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0099_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1578_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1505_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1477_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1460_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1457_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1451_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1411_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1387_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1381_),
    .X(net61));
 sg13g2_buf_4 fanout62 (.X(net62),
    .A(_1357_));
 sg13g2_buf_2 fanout63 (.A(_1349_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1422_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_1380_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_1610_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1369_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1489_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1421_),
    .X(net69));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_1362_));
 sg13g2_buf_2 fanout71 (.A(_0055_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0976_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1055_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1037_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_0516_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0164_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_1018_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_1016_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0986_),
    .X(net79));
 sg13g2_buf_4 fanout80 (.X(net80),
    .A(_0483_));
 sg13g2_buf_2 fanout81 (.A(_0329_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0307_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_0263_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(\hvsync_gen.vsync ),
    .X(net84));
 sg13g2_tielo _3364__85 (.L_LO(net85));
 sg13g2_tielo _3365__86 (.L_LO(net86));
 sg13g2_tielo _3366__87 (.L_LO(net87));
 sg13g2_tielo _3367__88 (.L_LO(net88));
 sg13g2_tielo _3368__89 (.L_LO(net89));
 sg13g2_tielo _3369__90 (.L_LO(net90));
 sg13g2_tielo _3370__91 (.L_LO(net91));
 sg13g2_tielo _3371__92 (.L_LO(net92));
 sg13g2_tielo _3372__93 (.L_LO(net93));
 sg13g2_tielo _3373__94 (.L_LO(net94));
 sg13g2_tielo _3374__95 (.L_LO(net95));
 sg13g2_tielo _3375__96 (.L_LO(net96));
 sg13g2_tielo _3376__97 (.L_LO(net97));
 sg13g2_tielo _3377__98 (.L_LO(net98));
 sg13g2_tielo _3378__99 (.L_LO(net99));
 sg13g2_tielo _3379__100 (.L_LO(net100));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__121  (.L_HI(net121));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0N__122  (.L_HI(net122));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0N__123  (.L_HI(net123));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0N__124  (.L_HI(net124));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0N__125  (.L_HI(net125));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0N__126  (.L_HI(net126));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0N__127  (.L_HI(net127));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0N__128  (.L_HI(net128));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0N__129  (.L_HI(net129));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0N__130  (.L_HI(net130));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0N__131  (.L_HI(net131));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__132  (.L_HI(net132));
 sg13g2_tiehi \yb[0]$_DFF_P__133  (.L_HI(net133));
 sg13g2_tiehi \yb[1]$_DFF_P__134  (.L_HI(net134));
 sg13g2_tiehi \yb[2]$_DFF_P__135  (.L_HI(net135));
 sg13g2_tiehi \yb[3]$_DFF_P__136  (.L_HI(net136));
 sg13g2_tiehi \yb[4]$_DFF_P__137  (.L_HI(net137));
 sg13g2_tiehi \yb[5]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_buf_1 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sg13g2_buf_1 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sg13g2_buf_1 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sg13g2_buf_1 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_fill_2 FILLER_0_105 ();
 sg13g2_fill_1 FILLER_0_107 ();
 sg13g2_decap_8 FILLER_0_116 ();
 sg13g2_decap_8 FILLER_0_123 ();
 sg13g2_decap_8 FILLER_0_130 ();
 sg13g2_decap_8 FILLER_0_137 ();
 sg13g2_decap_8 FILLER_0_144 ();
 sg13g2_decap_8 FILLER_0_151 ();
 sg13g2_decap_8 FILLER_0_158 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_4 FILLER_0_172 ();
 sg13g2_fill_2 FILLER_0_176 ();
 sg13g2_decap_4 FILLER_0_182 ();
 sg13g2_fill_2 FILLER_0_186 ();
 sg13g2_fill_1 FILLER_0_192 ();
 sg13g2_decap_8 FILLER_0_197 ();
 sg13g2_decap_8 FILLER_0_204 ();
 sg13g2_decap_4 FILLER_0_215 ();
 sg13g2_fill_1 FILLER_0_232 ();
 sg13g2_decap_8 FILLER_0_250 ();
 sg13g2_decap_8 FILLER_0_257 ();
 sg13g2_decap_8 FILLER_0_264 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_278 ();
 sg13g2_decap_8 FILLER_0_285 ();
 sg13g2_decap_8 FILLER_0_292 ();
 sg13g2_decap_8 FILLER_0_299 ();
 sg13g2_decap_8 FILLER_0_306 ();
 sg13g2_decap_8 FILLER_0_313 ();
 sg13g2_decap_8 FILLER_0_320 ();
 sg13g2_decap_8 FILLER_0_327 ();
 sg13g2_decap_8 FILLER_0_334 ();
 sg13g2_decap_8 FILLER_0_341 ();
 sg13g2_decap_8 FILLER_0_348 ();
 sg13g2_decap_8 FILLER_0_355 ();
 sg13g2_decap_8 FILLER_0_362 ();
 sg13g2_decap_8 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_376 ();
 sg13g2_decap_8 FILLER_0_383 ();
 sg13g2_decap_8 FILLER_0_390 ();
 sg13g2_decap_8 FILLER_0_397 ();
 sg13g2_decap_8 FILLER_0_404 ();
 sg13g2_decap_8 FILLER_0_411 ();
 sg13g2_decap_8 FILLER_0_418 ();
 sg13g2_decap_4 FILLER_0_425 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_4 FILLER_1_77 ();
 sg13g2_fill_2 FILLER_1_81 ();
 sg13g2_decap_8 FILLER_1_117 ();
 sg13g2_decap_4 FILLER_1_124 ();
 sg13g2_fill_2 FILLER_1_132 ();
 sg13g2_fill_1 FILLER_1_134 ();
 sg13g2_fill_2 FILLER_1_140 ();
 sg13g2_fill_1 FILLER_1_142 ();
 sg13g2_decap_8 FILLER_1_160 ();
 sg13g2_decap_4 FILLER_1_167 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_2 FILLER_1_193 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_fill_1 FILLER_1_224 ();
 sg13g2_decap_4 FILLER_1_245 ();
 sg13g2_fill_1 FILLER_1_249 ();
 sg13g2_fill_2 FILLER_1_263 ();
 sg13g2_fill_1 FILLER_1_265 ();
 sg13g2_decap_4 FILLER_1_283 ();
 sg13g2_fill_1 FILLER_1_287 ();
 sg13g2_decap_4 FILLER_1_296 ();
 sg13g2_fill_2 FILLER_1_300 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_decap_4 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_341 ();
 sg13g2_decap_8 FILLER_1_348 ();
 sg13g2_decap_8 FILLER_1_355 ();
 sg13g2_decap_8 FILLER_1_362 ();
 sg13g2_decap_8 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_376 ();
 sg13g2_decap_8 FILLER_1_383 ();
 sg13g2_decap_8 FILLER_1_390 ();
 sg13g2_decap_8 FILLER_1_397 ();
 sg13g2_decap_8 FILLER_1_404 ();
 sg13g2_decap_8 FILLER_1_411 ();
 sg13g2_decap_8 FILLER_1_418 ();
 sg13g2_decap_4 FILLER_1_425 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_fill_1 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_73 ();
 sg13g2_decap_8 FILLER_2_80 ();
 sg13g2_fill_2 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_89 ();
 sg13g2_fill_1 FILLER_2_95 ();
 sg13g2_fill_1 FILLER_2_104 ();
 sg13g2_decap_4 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_117 ();
 sg13g2_decap_4 FILLER_2_128 ();
 sg13g2_fill_2 FILLER_2_136 ();
 sg13g2_fill_1 FILLER_2_138 ();
 sg13g2_decap_4 FILLER_2_153 ();
 sg13g2_fill_1 FILLER_2_157 ();
 sg13g2_fill_1 FILLER_2_163 ();
 sg13g2_fill_2 FILLER_2_179 ();
 sg13g2_fill_1 FILLER_2_181 ();
 sg13g2_fill_1 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_205 ();
 sg13g2_fill_2 FILLER_2_212 ();
 sg13g2_fill_1 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_239 ();
 sg13g2_fill_1 FILLER_2_245 ();
 sg13g2_fill_1 FILLER_2_258 ();
 sg13g2_decap_8 FILLER_2_276 ();
 sg13g2_decap_4 FILLER_2_283 ();
 sg13g2_fill_2 FILLER_2_287 ();
 sg13g2_fill_2 FILLER_2_301 ();
 sg13g2_fill_1 FILLER_2_303 ();
 sg13g2_decap_8 FILLER_2_316 ();
 sg13g2_decap_4 FILLER_2_323 ();
 sg13g2_fill_2 FILLER_2_327 ();
 sg13g2_decap_8 FILLER_2_337 ();
 sg13g2_fill_2 FILLER_2_344 ();
 sg13g2_decap_8 FILLER_2_359 ();
 sg13g2_decap_8 FILLER_2_366 ();
 sg13g2_decap_8 FILLER_2_373 ();
 sg13g2_decap_8 FILLER_2_380 ();
 sg13g2_decap_8 FILLER_2_387 ();
 sg13g2_decap_8 FILLER_2_394 ();
 sg13g2_decap_8 FILLER_2_401 ();
 sg13g2_decap_8 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_422 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_2 FILLER_3_57 ();
 sg13g2_fill_1 FILLER_3_59 ();
 sg13g2_fill_1 FILLER_3_64 ();
 sg13g2_fill_1 FILLER_3_68 ();
 sg13g2_decap_8 FILLER_3_79 ();
 sg13g2_decap_4 FILLER_3_86 ();
 sg13g2_fill_1 FILLER_3_90 ();
 sg13g2_decap_4 FILLER_3_95 ();
 sg13g2_fill_2 FILLER_3_99 ();
 sg13g2_fill_2 FILLER_3_110 ();
 sg13g2_fill_1 FILLER_3_112 ();
 sg13g2_fill_2 FILLER_3_117 ();
 sg13g2_fill_1 FILLER_3_139 ();
 sg13g2_fill_1 FILLER_3_154 ();
 sg13g2_fill_2 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_fill_1 FILLER_3_184 ();
 sg13g2_decap_4 FILLER_3_197 ();
 sg13g2_fill_2 FILLER_3_201 ();
 sg13g2_decap_4 FILLER_3_211 ();
 sg13g2_fill_1 FILLER_3_215 ();
 sg13g2_fill_2 FILLER_3_221 ();
 sg13g2_fill_1 FILLER_3_248 ();
 sg13g2_fill_1 FILLER_3_258 ();
 sg13g2_fill_1 FILLER_3_275 ();
 sg13g2_fill_2 FILLER_3_281 ();
 sg13g2_fill_1 FILLER_3_283 ();
 sg13g2_decap_4 FILLER_3_293 ();
 sg13g2_fill_1 FILLER_3_321 ();
 sg13g2_fill_1 FILLER_3_335 ();
 sg13g2_fill_2 FILLER_3_340 ();
 sg13g2_fill_1 FILLER_3_342 ();
 sg13g2_fill_2 FILLER_3_355 ();
 sg13g2_fill_1 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_60 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_132 ();
 sg13g2_fill_1 FILLER_4_137 ();
 sg13g2_fill_2 FILLER_4_142 ();
 sg13g2_fill_1 FILLER_4_152 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_decap_4 FILLER_4_165 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_183 ();
 sg13g2_fill_2 FILLER_4_190 ();
 sg13g2_decap_4 FILLER_4_196 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_215 ();
 sg13g2_decap_4 FILLER_4_261 ();
 sg13g2_decap_8 FILLER_4_269 ();
 sg13g2_decap_4 FILLER_4_276 ();
 sg13g2_fill_1 FILLER_4_280 ();
 sg13g2_fill_1 FILLER_4_286 ();
 sg13g2_decap_8 FILLER_4_299 ();
 sg13g2_decap_8 FILLER_4_306 ();
 sg13g2_decap_8 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_320 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_4 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_fill_2 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_108 ();
 sg13g2_decap_4 FILLER_5_120 ();
 sg13g2_fill_2 FILLER_5_133 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_2 FILLER_5_145 ();
 sg13g2_decap_4 FILLER_5_156 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_fill_1 FILLER_5_184 ();
 sg13g2_fill_1 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_194 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_209 ();
 sg13g2_decap_4 FILLER_5_216 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_8 FILLER_5_230 ();
 sg13g2_decap_4 FILLER_5_237 ();
 sg13g2_fill_2 FILLER_5_249 ();
 sg13g2_fill_1 FILLER_5_251 ();
 sg13g2_fill_1 FILLER_5_268 ();
 sg13g2_fill_2 FILLER_5_276 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_4 FILLER_5_325 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_decap_4 FILLER_5_350 ();
 sg13g2_fill_1 FILLER_5_354 ();
 sg13g2_fill_1 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_372 ();
 sg13g2_decap_8 FILLER_5_379 ();
 sg13g2_decap_8 FILLER_5_386 ();
 sg13g2_decap_8 FILLER_5_393 ();
 sg13g2_decap_8 FILLER_5_400 ();
 sg13g2_decap_8 FILLER_5_407 ();
 sg13g2_decap_8 FILLER_5_414 ();
 sg13g2_decap_8 FILLER_5_421 ();
 sg13g2_fill_2 FILLER_5_428 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_fill_2 FILLER_6_49 ();
 sg13g2_fill_2 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_57 ();
 sg13g2_fill_2 FILLER_6_68 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_2 FILLER_6_78 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_106 ();
 sg13g2_fill_1 FILLER_6_108 ();
 sg13g2_fill_2 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_135 ();
 sg13g2_fill_1 FILLER_6_146 ();
 sg13g2_decap_8 FILLER_6_156 ();
 sg13g2_fill_2 FILLER_6_163 ();
 sg13g2_fill_2 FILLER_6_173 ();
 sg13g2_fill_1 FILLER_6_184 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_fill_2 FILLER_6_204 ();
 sg13g2_decap_8 FILLER_6_215 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_1 FILLER_6_227 ();
 sg13g2_decap_8 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_239 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_262 ();
 sg13g2_fill_1 FILLER_6_273 ();
 sg13g2_fill_1 FILLER_6_278 ();
 sg13g2_fill_1 FILLER_6_283 ();
 sg13g2_fill_2 FILLER_6_288 ();
 sg13g2_fill_2 FILLER_6_302 ();
 sg13g2_fill_1 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_313 ();
 sg13g2_fill_2 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_4 FILLER_6_351 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_6_361 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_fill_2 FILLER_7_76 ();
 sg13g2_fill_1 FILLER_7_82 ();
 sg13g2_fill_2 FILLER_7_90 ();
 sg13g2_fill_2 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_127 ();
 sg13g2_fill_1 FILLER_7_129 ();
 sg13g2_fill_1 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_138 ();
 sg13g2_fill_1 FILLER_7_145 ();
 sg13g2_fill_1 FILLER_7_151 ();
 sg13g2_fill_2 FILLER_7_168 ();
 sg13g2_decap_8 FILLER_7_176 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_fill_1 FILLER_7_221 ();
 sg13g2_fill_2 FILLER_7_227 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_238 ();
 sg13g2_fill_2 FILLER_7_244 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_fill_2 FILLER_7_260 ();
 sg13g2_fill_2 FILLER_7_266 ();
 sg13g2_fill_1 FILLER_7_272 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_288 ();
 sg13g2_decap_4 FILLER_7_294 ();
 sg13g2_fill_2 FILLER_7_302 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_fill_2 FILLER_7_315 ();
 sg13g2_fill_1 FILLER_7_317 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_fill_2 FILLER_7_329 ();
 sg13g2_fill_1 FILLER_7_331 ();
 sg13g2_decap_4 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_349 ();
 sg13g2_fill_1 FILLER_7_356 ();
 sg13g2_fill_2 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_8 FILLER_7_404 ();
 sg13g2_decap_8 FILLER_7_411 ();
 sg13g2_decap_8 FILLER_7_418 ();
 sg13g2_decap_4 FILLER_7_425 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_fill_2 FILLER_8_60 ();
 sg13g2_fill_1 FILLER_8_62 ();
 sg13g2_fill_1 FILLER_8_72 ();
 sg13g2_fill_2 FILLER_8_85 ();
 sg13g2_fill_2 FILLER_8_92 ();
 sg13g2_decap_4 FILLER_8_103 ();
 sg13g2_fill_1 FILLER_8_107 ();
 sg13g2_fill_1 FILLER_8_116 ();
 sg13g2_fill_2 FILLER_8_121 ();
 sg13g2_fill_1 FILLER_8_123 ();
 sg13g2_decap_4 FILLER_8_136 ();
 sg13g2_fill_1 FILLER_8_140 ();
 sg13g2_decap_4 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_161 ();
 sg13g2_fill_1 FILLER_8_169 ();
 sg13g2_decap_8 FILLER_8_179 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_fill_1 FILLER_8_188 ();
 sg13g2_fill_1 FILLER_8_194 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_fill_2 FILLER_8_209 ();
 sg13g2_fill_2 FILLER_8_242 ();
 sg13g2_decap_4 FILLER_8_261 ();
 sg13g2_fill_1 FILLER_8_265 ();
 sg13g2_fill_2 FILLER_8_270 ();
 sg13g2_fill_1 FILLER_8_272 ();
 sg13g2_fill_2 FILLER_8_277 ();
 sg13g2_fill_2 FILLER_8_284 ();
 sg13g2_fill_2 FILLER_8_290 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_302 ();
 sg13g2_fill_1 FILLER_8_304 ();
 sg13g2_decap_4 FILLER_8_313 ();
 sg13g2_fill_2 FILLER_8_333 ();
 sg13g2_fill_1 FILLER_8_335 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_4 FILLER_9_28 ();
 sg13g2_fill_1 FILLER_9_32 ();
 sg13g2_fill_1 FILLER_9_59 ();
 sg13g2_fill_1 FILLER_9_64 ();
 sg13g2_fill_2 FILLER_9_82 ();
 sg13g2_fill_2 FILLER_9_89 ();
 sg13g2_fill_2 FILLER_9_95 ();
 sg13g2_decap_8 FILLER_9_106 ();
 sg13g2_decap_4 FILLER_9_118 ();
 sg13g2_fill_2 FILLER_9_122 ();
 sg13g2_decap_8 FILLER_9_130 ();
 sg13g2_decap_4 FILLER_9_137 ();
 sg13g2_decap_8 FILLER_9_145 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_fill_1 FILLER_9_154 ();
 sg13g2_fill_2 FILLER_9_160 ();
 sg13g2_decap_4 FILLER_9_174 ();
 sg13g2_decap_4 FILLER_9_193 ();
 sg13g2_fill_1 FILLER_9_210 ();
 sg13g2_fill_2 FILLER_9_215 ();
 sg13g2_decap_8 FILLER_9_237 ();
 sg13g2_fill_1 FILLER_9_244 ();
 sg13g2_decap_4 FILLER_9_260 ();
 sg13g2_fill_1 FILLER_9_264 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_1 FILLER_9_289 ();
 sg13g2_decap_4 FILLER_9_299 ();
 sg13g2_fill_1 FILLER_9_303 ();
 sg13g2_decap_8 FILLER_9_312 ();
 sg13g2_fill_2 FILLER_9_319 ();
 sg13g2_fill_1 FILLER_9_321 ();
 sg13g2_decap_4 FILLER_9_330 ();
 sg13g2_fill_2 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_fill_2 FILLER_9_384 ();
 sg13g2_fill_1 FILLER_9_386 ();
 sg13g2_decap_8 FILLER_9_400 ();
 sg13g2_decap_8 FILLER_9_407 ();
 sg13g2_decap_8 FILLER_9_414 ();
 sg13g2_decap_8 FILLER_9_421 ();
 sg13g2_fill_2 FILLER_9_428 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_4 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_39 ();
 sg13g2_decap_4 FILLER_10_45 ();
 sg13g2_fill_2 FILLER_10_68 ();
 sg13g2_fill_2 FILLER_10_84 ();
 sg13g2_fill_2 FILLER_10_96 ();
 sg13g2_fill_1 FILLER_10_101 ();
 sg13g2_decap_4 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_110 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_1 FILLER_10_123 ();
 sg13g2_fill_2 FILLER_10_128 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_fill_1 FILLER_10_157 ();
 sg13g2_decap_4 FILLER_10_162 ();
 sg13g2_decap_8 FILLER_10_183 ();
 sg13g2_decap_8 FILLER_10_201 ();
 sg13g2_decap_8 FILLER_10_211 ();
 sg13g2_fill_1 FILLER_10_218 ();
 sg13g2_fill_2 FILLER_10_232 ();
 sg13g2_decap_4 FILLER_10_238 ();
 sg13g2_fill_1 FILLER_10_251 ();
 sg13g2_fill_2 FILLER_10_263 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_fill_1 FILLER_10_270 ();
 sg13g2_fill_1 FILLER_10_275 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_fill_1 FILLER_10_285 ();
 sg13g2_fill_2 FILLER_10_302 ();
 sg13g2_fill_1 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_316 ();
 sg13g2_fill_1 FILLER_10_327 ();
 sg13g2_fill_1 FILLER_10_332 ();
 sg13g2_fill_2 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_339 ();
 sg13g2_decap_4 FILLER_10_344 ();
 sg13g2_fill_2 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_375 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_1 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_10_409 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_fill_2 FILLER_11_60 ();
 sg13g2_fill_1 FILLER_11_69 ();
 sg13g2_decap_4 FILLER_11_80 ();
 sg13g2_fill_2 FILLER_11_84 ();
 sg13g2_fill_2 FILLER_11_94 ();
 sg13g2_fill_1 FILLER_11_96 ();
 sg13g2_fill_2 FILLER_11_106 ();
 sg13g2_fill_2 FILLER_11_118 ();
 sg13g2_decap_8 FILLER_11_136 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_decap_4 FILLER_11_154 ();
 sg13g2_fill_2 FILLER_11_162 ();
 sg13g2_fill_1 FILLER_11_164 ();
 sg13g2_fill_2 FILLER_11_169 ();
 sg13g2_fill_1 FILLER_11_171 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_1 FILLER_11_182 ();
 sg13g2_fill_2 FILLER_11_188 ();
 sg13g2_decap_4 FILLER_11_214 ();
 sg13g2_decap_4 FILLER_11_222 ();
 sg13g2_decap_4 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_247 ();
 sg13g2_decap_4 FILLER_11_252 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_decap_4 FILLER_11_295 ();
 sg13g2_decap_4 FILLER_11_303 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_decap_8 FILLER_11_317 ();
 sg13g2_fill_2 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_348 ();
 sg13g2_decap_8 FILLER_11_355 ();
 sg13g2_decap_8 FILLER_11_362 ();
 sg13g2_decap_8 FILLER_11_369 ();
 sg13g2_decap_8 FILLER_11_376 ();
 sg13g2_fill_1 FILLER_11_383 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_8 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_11_412 ();
 sg13g2_decap_8 FILLER_11_419 ();
 sg13g2_decap_4 FILLER_11_426 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_4 FILLER_12_28 ();
 sg13g2_fill_2 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_71 ();
 sg13g2_fill_2 FILLER_12_77 ();
 sg13g2_fill_2 FILLER_12_89 ();
 sg13g2_fill_1 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_101 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_fill_2 FILLER_12_113 ();
 sg13g2_fill_2 FILLER_12_136 ();
 sg13g2_fill_1 FILLER_12_157 ();
 sg13g2_fill_1 FILLER_12_184 ();
 sg13g2_fill_1 FILLER_12_193 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_214 ();
 sg13g2_fill_2 FILLER_12_219 ();
 sg13g2_decap_8 FILLER_12_231 ();
 sg13g2_decap_8 FILLER_12_238 ();
 sg13g2_fill_2 FILLER_12_245 ();
 sg13g2_fill_1 FILLER_12_247 ();
 sg13g2_fill_2 FILLER_12_252 ();
 sg13g2_fill_1 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_270 ();
 sg13g2_fill_1 FILLER_12_276 ();
 sg13g2_decap_8 FILLER_12_282 ();
 sg13g2_fill_2 FILLER_12_289 ();
 sg13g2_fill_1 FILLER_12_291 ();
 sg13g2_fill_1 FILLER_12_301 ();
 sg13g2_fill_2 FILLER_12_315 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_331 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_fill_2 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_345 ();
 sg13g2_fill_1 FILLER_12_359 ();
 sg13g2_fill_2 FILLER_12_368 ();
 sg13g2_decap_4 FILLER_12_374 ();
 sg13g2_fill_1 FILLER_12_378 ();
 sg13g2_decap_4 FILLER_12_387 ();
 sg13g2_fill_2 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_397 ();
 sg13g2_decap_8 FILLER_12_404 ();
 sg13g2_decap_8 FILLER_12_411 ();
 sg13g2_decap_8 FILLER_12_418 ();
 sg13g2_decap_4 FILLER_12_425 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_50 ();
 sg13g2_fill_1 FILLER_13_52 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_fill_1 FILLER_13_64 ();
 sg13g2_fill_2 FILLER_13_79 ();
 sg13g2_fill_2 FILLER_13_84 ();
 sg13g2_fill_1 FILLER_13_86 ();
 sg13g2_decap_4 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_118 ();
 sg13g2_decap_4 FILLER_13_123 ();
 sg13g2_fill_2 FILLER_13_131 ();
 sg13g2_fill_1 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_2 FILLER_13_171 ();
 sg13g2_fill_1 FILLER_13_173 ();
 sg13g2_decap_4 FILLER_13_179 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_fill_1 FILLER_13_197 ();
 sg13g2_fill_1 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_208 ();
 sg13g2_fill_1 FILLER_13_215 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_238 ();
 sg13g2_fill_2 FILLER_13_244 ();
 sg13g2_fill_1 FILLER_13_246 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_2 FILLER_13_265 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_294 ();
 sg13g2_fill_1 FILLER_13_300 ();
 sg13g2_fill_2 FILLER_13_310 ();
 sg13g2_fill_1 FILLER_13_312 ();
 sg13g2_fill_1 FILLER_13_321 ();
 sg13g2_fill_2 FILLER_13_326 ();
 sg13g2_fill_1 FILLER_13_328 ();
 sg13g2_fill_1 FILLER_13_333 ();
 sg13g2_decap_4 FILLER_13_338 ();
 sg13g2_fill_2 FILLER_13_342 ();
 sg13g2_decap_8 FILLER_13_348 ();
 sg13g2_decap_8 FILLER_13_355 ();
 sg13g2_fill_1 FILLER_13_362 ();
 sg13g2_decap_8 FILLER_13_376 ();
 sg13g2_fill_2 FILLER_13_383 ();
 sg13g2_decap_8 FILLER_13_418 ();
 sg13g2_decap_4 FILLER_13_425 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_4 FILLER_14_35 ();
 sg13g2_fill_2 FILLER_14_39 ();
 sg13g2_decap_4 FILLER_14_55 ();
 sg13g2_fill_1 FILLER_14_59 ();
 sg13g2_fill_1 FILLER_14_65 ();
 sg13g2_decap_4 FILLER_14_111 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_decap_4 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_136 ();
 sg13g2_fill_2 FILLER_14_142 ();
 sg13g2_fill_2 FILLER_14_153 ();
 sg13g2_fill_1 FILLER_14_155 ();
 sg13g2_decap_4 FILLER_14_161 ();
 sg13g2_fill_1 FILLER_14_165 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_fill_2 FILLER_14_191 ();
 sg13g2_decap_4 FILLER_14_198 ();
 sg13g2_fill_2 FILLER_14_219 ();
 sg13g2_fill_1 FILLER_14_221 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_244 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_2 FILLER_14_269 ();
 sg13g2_fill_2 FILLER_14_276 ();
 sg13g2_fill_1 FILLER_14_278 ();
 sg13g2_fill_2 FILLER_14_284 ();
 sg13g2_fill_1 FILLER_14_286 ();
 sg13g2_fill_2 FILLER_14_299 ();
 sg13g2_fill_2 FILLER_14_306 ();
 sg13g2_fill_1 FILLER_14_308 ();
 sg13g2_fill_2 FILLER_14_314 ();
 sg13g2_fill_2 FILLER_14_321 ();
 sg13g2_decap_4 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_344 ();
 sg13g2_decap_8 FILLER_14_351 ();
 sg13g2_decap_4 FILLER_14_358 ();
 sg13g2_fill_1 FILLER_14_362 ();
 sg13g2_fill_1 FILLER_14_370 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_fill_2 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_4 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_419 ();
 sg13g2_decap_4 FILLER_14_426 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_42 ();
 sg13g2_fill_2 FILLER_15_49 ();
 sg13g2_fill_1 FILLER_15_51 ();
 sg13g2_fill_1 FILLER_15_56 ();
 sg13g2_fill_2 FILLER_15_65 ();
 sg13g2_fill_1 FILLER_15_71 ();
 sg13g2_decap_4 FILLER_15_86 ();
 sg13g2_fill_2 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_102 ();
 sg13g2_fill_1 FILLER_15_110 ();
 sg13g2_fill_1 FILLER_15_120 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_decap_8 FILLER_15_162 ();
 sg13g2_fill_2 FILLER_15_185 ();
 sg13g2_fill_2 FILLER_15_209 ();
 sg13g2_fill_2 FILLER_15_215 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_242 ();
 sg13g2_fill_1 FILLER_15_271 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_292 ();
 sg13g2_fill_2 FILLER_15_297 ();
 sg13g2_fill_1 FILLER_15_308 ();
 sg13g2_fill_2 FILLER_15_319 ();
 sg13g2_fill_1 FILLER_15_321 ();
 sg13g2_fill_1 FILLER_15_342 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_4 FILLER_15_361 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_2 FILLER_15_376 ();
 sg13g2_decap_4 FILLER_15_383 ();
 sg13g2_decap_4 FILLER_15_391 ();
 sg13g2_fill_1 FILLER_15_395 ();
 sg13g2_fill_2 FILLER_15_412 ();
 sg13g2_fill_1 FILLER_15_414 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_fill_1 FILLER_16_56 ();
 sg13g2_fill_2 FILLER_16_61 ();
 sg13g2_fill_1 FILLER_16_63 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_fill_1 FILLER_16_71 ();
 sg13g2_fill_1 FILLER_16_94 ();
 sg13g2_fill_1 FILLER_16_120 ();
 sg13g2_fill_2 FILLER_16_126 ();
 sg13g2_fill_1 FILLER_16_128 ();
 sg13g2_fill_1 FILLER_16_134 ();
 sg13g2_fill_1 FILLER_16_157 ();
 sg13g2_decap_8 FILLER_16_170 ();
 sg13g2_decap_4 FILLER_16_181 ();
 sg13g2_decap_4 FILLER_16_197 ();
 sg13g2_fill_1 FILLER_16_213 ();
 sg13g2_decap_8 FILLER_16_227 ();
 sg13g2_decap_8 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_241 ();
 sg13g2_fill_1 FILLER_16_253 ();
 sg13g2_decap_4 FILLER_16_273 ();
 sg13g2_fill_2 FILLER_16_277 ();
 sg13g2_decap_8 FILLER_16_288 ();
 sg13g2_decap_4 FILLER_16_295 ();
 sg13g2_fill_1 FILLER_16_299 ();
 sg13g2_decap_4 FILLER_16_309 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_fill_2 FILLER_16_333 ();
 sg13g2_fill_1 FILLER_16_347 ();
 sg13g2_decap_8 FILLER_16_352 ();
 sg13g2_decap_8 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_decap_8 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_fill_1 FILLER_16_409 ();
 sg13g2_decap_8 FILLER_16_418 ();
 sg13g2_decap_4 FILLER_16_425 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_78 ();
 sg13g2_fill_2 FILLER_17_95 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_1 FILLER_17_102 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_decap_4 FILLER_17_122 ();
 sg13g2_decap_4 FILLER_17_134 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_2 FILLER_17_145 ();
 sg13g2_decap_4 FILLER_17_151 ();
 sg13g2_decap_4 FILLER_17_159 ();
 sg13g2_fill_1 FILLER_17_167 ();
 sg13g2_fill_1 FILLER_17_172 ();
 sg13g2_fill_1 FILLER_17_178 ();
 sg13g2_fill_2 FILLER_17_204 ();
 sg13g2_fill_1 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_4 FILLER_17_235 ();
 sg13g2_fill_1 FILLER_17_239 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_fill_1 FILLER_17_282 ();
 sg13g2_fill_1 FILLER_17_294 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_fill_1 FILLER_17_302 ();
 sg13g2_fill_2 FILLER_17_322 ();
 sg13g2_fill_2 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_fill_1 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_17_404 ();
 sg13g2_fill_1 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_4 FILLER_18_49 ();
 sg13g2_fill_2 FILLER_18_53 ();
 sg13g2_fill_2 FILLER_18_69 ();
 sg13g2_fill_1 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_77 ();
 sg13g2_fill_1 FILLER_18_85 ();
 sg13g2_fill_2 FILLER_18_90 ();
 sg13g2_fill_2 FILLER_18_103 ();
 sg13g2_fill_2 FILLER_18_125 ();
 sg13g2_fill_1 FILLER_18_133 ();
 sg13g2_fill_2 FILLER_18_138 ();
 sg13g2_decap_4 FILLER_18_150 ();
 sg13g2_fill_2 FILLER_18_154 ();
 sg13g2_fill_1 FILLER_18_182 ();
 sg13g2_fill_1 FILLER_18_186 ();
 sg13g2_decap_4 FILLER_18_198 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_213 ();
 sg13g2_fill_1 FILLER_18_215 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_244 ();
 sg13g2_decap_4 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_4 FILLER_18_273 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_decap_8 FILLER_18_282 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_decap_8 FILLER_18_296 ();
 sg13g2_fill_2 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_325 ();
 sg13g2_fill_2 FILLER_18_332 ();
 sg13g2_fill_1 FILLER_18_334 ();
 sg13g2_decap_4 FILLER_18_340 ();
 sg13g2_fill_2 FILLER_18_344 ();
 sg13g2_decap_8 FILLER_18_351 ();
 sg13g2_decap_8 FILLER_18_358 ();
 sg13g2_fill_2 FILLER_18_365 ();
 sg13g2_fill_1 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_fill_2 FILLER_18_385 ();
 sg13g2_fill_2 FILLER_18_405 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_fill_2 FILLER_18_428 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_53 ();
 sg13g2_fill_1 FILLER_19_83 ();
 sg13g2_fill_1 FILLER_19_102 ();
 sg13g2_fill_1 FILLER_19_109 ();
 sg13g2_fill_2 FILLER_19_120 ();
 sg13g2_decap_4 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_158 ();
 sg13g2_fill_1 FILLER_19_166 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_217 ();
 sg13g2_decap_4 FILLER_19_222 ();
 sg13g2_decap_4 FILLER_19_231 ();
 sg13g2_decap_4 FILLER_19_239 ();
 sg13g2_fill_1 FILLER_19_243 ();
 sg13g2_decap_4 FILLER_19_249 ();
 sg13g2_fill_1 FILLER_19_253 ();
 sg13g2_decap_4 FILLER_19_260 ();
 sg13g2_decap_4 FILLER_19_269 ();
 sg13g2_fill_1 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_296 ();
 sg13g2_decap_8 FILLER_19_302 ();
 sg13g2_decap_4 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_decap_8 FILLER_19_345 ();
 sg13g2_decap_8 FILLER_19_352 ();
 sg13g2_decap_8 FILLER_19_359 ();
 sg13g2_fill_1 FILLER_19_366 ();
 sg13g2_fill_1 FILLER_19_376 ();
 sg13g2_decap_8 FILLER_19_391 ();
 sg13g2_fill_1 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_4 FILLER_19_410 ();
 sg13g2_fill_1 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_42 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_fill_1 FILLER_20_102 ();
 sg13g2_decap_4 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_124 ();
 sg13g2_decap_4 FILLER_20_132 ();
 sg13g2_fill_2 FILLER_20_136 ();
 sg13g2_fill_2 FILLER_20_141 ();
 sg13g2_decap_8 FILLER_20_147 ();
 sg13g2_decap_8 FILLER_20_154 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_decap_4 FILLER_20_182 ();
 sg13g2_fill_2 FILLER_20_186 ();
 sg13g2_decap_4 FILLER_20_196 ();
 sg13g2_fill_1 FILLER_20_200 ();
 sg13g2_decap_4 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_decap_4 FILLER_20_226 ();
 sg13g2_fill_1 FILLER_20_230 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_fill_1 FILLER_20_257 ();
 sg13g2_fill_1 FILLER_20_272 ();
 sg13g2_fill_2 FILLER_20_283 ();
 sg13g2_fill_2 FILLER_20_290 ();
 sg13g2_fill_2 FILLER_20_322 ();
 sg13g2_fill_1 FILLER_20_324 ();
 sg13g2_decap_8 FILLER_20_334 ();
 sg13g2_decap_8 FILLER_20_341 ();
 sg13g2_decap_8 FILLER_20_348 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_8 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_1 FILLER_20_418 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_fill_2 FILLER_21_35 ();
 sg13g2_fill_1 FILLER_21_37 ();
 sg13g2_fill_1 FILLER_21_41 ();
 sg13g2_decap_8 FILLER_21_68 ();
 sg13g2_decap_8 FILLER_21_75 ();
 sg13g2_decap_8 FILLER_21_82 ();
 sg13g2_decap_8 FILLER_21_89 ();
 sg13g2_decap_4 FILLER_21_96 ();
 sg13g2_fill_2 FILLER_21_100 ();
 sg13g2_decap_8 FILLER_21_110 ();
 sg13g2_decap_8 FILLER_21_117 ();
 sg13g2_decap_8 FILLER_21_124 ();
 sg13g2_fill_1 FILLER_21_131 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_147 ();
 sg13g2_fill_2 FILLER_21_153 ();
 sg13g2_decap_8 FILLER_21_160 ();
 sg13g2_decap_4 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_8 FILLER_21_184 ();
 sg13g2_decap_8 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_198 ();
 sg13g2_decap_8 FILLER_21_205 ();
 sg13g2_decap_8 FILLER_21_212 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_decap_8 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_233 ();
 sg13g2_decap_8 FILLER_21_240 ();
 sg13g2_decap_8 FILLER_21_247 ();
 sg13g2_decap_8 FILLER_21_254 ();
 sg13g2_decap_8 FILLER_21_261 ();
 sg13g2_decap_8 FILLER_21_268 ();
 sg13g2_decap_4 FILLER_21_275 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_4 FILLER_21_291 ();
 sg13g2_decap_4 FILLER_21_305 ();
 sg13g2_fill_2 FILLER_21_309 ();
 sg13g2_fill_2 FILLER_21_316 ();
 sg13g2_fill_1 FILLER_21_318 ();
 sg13g2_decap_4 FILLER_21_323 ();
 sg13g2_fill_1 FILLER_21_327 ();
 sg13g2_fill_2 FILLER_21_345 ();
 sg13g2_fill_1 FILLER_21_356 ();
 sg13g2_fill_2 FILLER_21_360 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_decap_8 FILLER_21_368 ();
 sg13g2_decap_4 FILLER_21_375 ();
 sg13g2_decap_8 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_391 ();
 sg13g2_fill_2 FILLER_21_398 ();
 sg13g2_fill_1 FILLER_21_412 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_4 FILLER_22_28 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_78 ();
 sg13g2_decap_4 FILLER_22_91 ();
 sg13g2_fill_1 FILLER_22_95 ();
 sg13g2_fill_1 FILLER_22_108 ();
 sg13g2_fill_1 FILLER_22_116 ();
 sg13g2_decap_4 FILLER_22_122 ();
 sg13g2_fill_2 FILLER_22_126 ();
 sg13g2_fill_1 FILLER_22_132 ();
 sg13g2_fill_2 FILLER_22_159 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_decap_8 FILLER_22_196 ();
 sg13g2_decap_8 FILLER_22_203 ();
 sg13g2_decap_8 FILLER_22_210 ();
 sg13g2_fill_2 FILLER_22_217 ();
 sg13g2_fill_2 FILLER_22_234 ();
 sg13g2_fill_1 FILLER_22_236 ();
 sg13g2_fill_2 FILLER_22_244 ();
 sg13g2_fill_2 FILLER_22_285 ();
 sg13g2_fill_2 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_299 ();
 sg13g2_decap_8 FILLER_22_306 ();
 sg13g2_decap_8 FILLER_22_313 ();
 sg13g2_decap_8 FILLER_22_320 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_338 ();
 sg13g2_decap_8 FILLER_22_345 ();
 sg13g2_decap_8 FILLER_22_352 ();
 sg13g2_decap_4 FILLER_22_359 ();
 sg13g2_fill_2 FILLER_22_363 ();
 sg13g2_fill_2 FILLER_22_395 ();
 sg13g2_fill_1 FILLER_22_397 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_fill_2 FILLER_22_412 ();
 sg13g2_decap_8 FILLER_22_420 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_4 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_18 ();
 sg13g2_fill_2 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_30 ();
 sg13g2_fill_1 FILLER_23_64 ();
 sg13g2_decap_8 FILLER_23_88 ();
 sg13g2_decap_4 FILLER_23_99 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_121 ();
 sg13g2_decap_8 FILLER_23_128 ();
 sg13g2_decap_4 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_139 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_191 ();
 sg13g2_fill_1 FILLER_23_226 ();
 sg13g2_decap_8 FILLER_23_235 ();
 sg13g2_fill_1 FILLER_23_242 ();
 sg13g2_decap_8 FILLER_23_247 ();
 sg13g2_decap_4 FILLER_23_254 ();
 sg13g2_decap_8 FILLER_23_262 ();
 sg13g2_decap_8 FILLER_23_269 ();
 sg13g2_decap_8 FILLER_23_276 ();
 sg13g2_decap_4 FILLER_23_283 ();
 sg13g2_decap_8 FILLER_23_299 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_2 FILLER_23_372 ();
 sg13g2_decap_4 FILLER_23_379 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_4 FILLER_23_395 ();
 sg13g2_fill_2 FILLER_23_399 ();
 sg13g2_fill_1 FILLER_23_414 ();
 sg13g2_decap_4 FILLER_23_425 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_22 ();
 sg13g2_fill_2 FILLER_24_27 ();
 sg13g2_fill_1 FILLER_24_29 ();
 sg13g2_decap_8 FILLER_24_37 ();
 sg13g2_fill_2 FILLER_24_44 ();
 sg13g2_fill_1 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_51 ();
 sg13g2_decap_4 FILLER_24_58 ();
 sg13g2_fill_1 FILLER_24_66 ();
 sg13g2_decap_4 FILLER_24_75 ();
 sg13g2_decap_8 FILLER_24_93 ();
 sg13g2_fill_1 FILLER_24_100 ();
 sg13g2_fill_1 FILLER_24_108 ();
 sg13g2_fill_1 FILLER_24_112 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_fill_1 FILLER_24_126 ();
 sg13g2_fill_2 FILLER_24_131 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_170 ();
 sg13g2_decap_8 FILLER_24_177 ();
 sg13g2_decap_4 FILLER_24_184 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_202 ();
 sg13g2_fill_1 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_212 ();
 sg13g2_fill_1 FILLER_24_216 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_4 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_fill_2 FILLER_24_284 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_8 FILLER_24_324 ();
 sg13g2_decap_8 FILLER_24_331 ();
 sg13g2_decap_8 FILLER_24_338 ();
 sg13g2_decap_8 FILLER_24_345 ();
 sg13g2_decap_8 FILLER_24_352 ();
 sg13g2_decap_8 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_366 ();
 sg13g2_decap_8 FILLER_24_394 ();
 sg13g2_decap_8 FILLER_24_401 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_9 ();
 sg13g2_fill_2 FILLER_25_33 ();
 sg13g2_decap_8 FILLER_25_50 ();
 sg13g2_decap_4 FILLER_25_57 ();
 sg13g2_fill_1 FILLER_25_61 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_4 FILLER_25_95 ();
 sg13g2_decap_4 FILLER_25_102 ();
 sg13g2_decap_4 FILLER_25_109 ();
 sg13g2_fill_2 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_149 ();
 sg13g2_fill_1 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_159 ();
 sg13g2_decap_8 FILLER_25_166 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_decap_4 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_205 ();
 sg13g2_fill_1 FILLER_25_212 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_2 FILLER_25_228 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_decap_8 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_248 ();
 sg13g2_fill_1 FILLER_25_255 ();
 sg13g2_decap_4 FILLER_25_260 ();
 sg13g2_decap_4 FILLER_25_277 ();
 sg13g2_decap_4 FILLER_25_301 ();
 sg13g2_fill_1 FILLER_25_305 ();
 sg13g2_decap_8 FILLER_25_310 ();
 sg13g2_fill_2 FILLER_25_317 ();
 sg13g2_decap_8 FILLER_25_332 ();
 sg13g2_decap_8 FILLER_25_339 ();
 sg13g2_decap_4 FILLER_25_346 ();
 sg13g2_fill_2 FILLER_25_364 ();
 sg13g2_fill_2 FILLER_25_370 ();
 sg13g2_fill_1 FILLER_25_372 ();
 sg13g2_fill_1 FILLER_25_381 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_399 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_fill_2 FILLER_26_29 ();
 sg13g2_fill_2 FILLER_26_40 ();
 sg13g2_fill_2 FILLER_26_47 ();
 sg13g2_decap_8 FILLER_26_58 ();
 sg13g2_decap_8 FILLER_26_65 ();
 sg13g2_decap_8 FILLER_26_72 ();
 sg13g2_fill_2 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_137 ();
 sg13g2_fill_1 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_173 ();
 sg13g2_fill_2 FILLER_26_178 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_fill_1 FILLER_26_216 ();
 sg13g2_fill_2 FILLER_26_233 ();
 sg13g2_decap_4 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_248 ();
 sg13g2_decap_8 FILLER_26_326 ();
 sg13g2_fill_2 FILLER_26_333 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_fill_2 FILLER_26_378 ();
 sg13g2_fill_1 FILLER_26_388 ();
 sg13g2_fill_2 FILLER_26_397 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_26_409 ();
 sg13g2_decap_8 FILLER_26_421 ();
 sg13g2_fill_2 FILLER_26_428 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_31 ();
 sg13g2_fill_1 FILLER_27_38 ();
 sg13g2_decap_8 FILLER_27_65 ();
 sg13g2_decap_8 FILLER_27_98 ();
 sg13g2_decap_8 FILLER_27_105 ();
 sg13g2_decap_8 FILLER_27_112 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_fill_1 FILLER_27_132 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_decap_4 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_176 ();
 sg13g2_decap_8 FILLER_27_183 ();
 sg13g2_fill_2 FILLER_27_190 ();
 sg13g2_decap_4 FILLER_27_197 ();
 sg13g2_fill_1 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_246 ();
 sg13g2_decap_4 FILLER_27_253 ();
 sg13g2_fill_1 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_272 ();
 sg13g2_decap_8 FILLER_27_281 ();
 sg13g2_decap_4 FILLER_27_288 ();
 sg13g2_decap_8 FILLER_27_336 ();
 sg13g2_decap_4 FILLER_27_343 ();
 sg13g2_fill_2 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_355 ();
 sg13g2_decap_4 FILLER_27_365 ();
 sg13g2_fill_2 FILLER_27_369 ();
 sg13g2_decap_8 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_27_386 ();
 sg13g2_fill_1 FILLER_27_393 ();
 sg13g2_decap_8 FILLER_27_420 ();
 sg13g2_fill_2 FILLER_27_427 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_11 ();
 sg13g2_fill_2 FILLER_28_47 ();
 sg13g2_fill_2 FILLER_28_54 ();
 sg13g2_fill_1 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_62 ();
 sg13g2_decap_8 FILLER_28_69 ();
 sg13g2_decap_4 FILLER_28_76 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_fill_2 FILLER_28_91 ();
 sg13g2_decap_4 FILLER_28_123 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_fill_1 FILLER_28_161 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_decap_8 FILLER_28_197 ();
 sg13g2_fill_1 FILLER_28_229 ();
 sg13g2_decap_8 FILLER_28_241 ();
 sg13g2_decap_8 FILLER_28_248 ();
 sg13g2_decap_8 FILLER_28_255 ();
 sg13g2_fill_2 FILLER_28_262 ();
 sg13g2_decap_4 FILLER_28_273 ();
 sg13g2_fill_2 FILLER_28_277 ();
 sg13g2_decap_8 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_304 ();
 sg13g2_fill_2 FILLER_28_309 ();
 sg13g2_fill_2 FILLER_28_324 ();
 sg13g2_decap_4 FILLER_28_334 ();
 sg13g2_fill_2 FILLER_28_357 ();
 sg13g2_fill_1 FILLER_28_362 ();
 sg13g2_fill_1 FILLER_28_367 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_387 ();
 sg13g2_decap_4 FILLER_28_394 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_fill_1 FILLER_29_9 ();
 sg13g2_fill_2 FILLER_29_13 ();
 sg13g2_fill_1 FILLER_29_19 ();
 sg13g2_fill_1 FILLER_29_30 ();
 sg13g2_fill_1 FILLER_29_38 ();
 sg13g2_decap_4 FILLER_29_104 ();
 sg13g2_fill_2 FILLER_29_108 ();
 sg13g2_decap_8 FILLER_29_114 ();
 sg13g2_decap_8 FILLER_29_121 ();
 sg13g2_fill_1 FILLER_29_128 ();
 sg13g2_fill_1 FILLER_29_133 ();
 sg13g2_decap_8 FILLER_29_138 ();
 sg13g2_decap_4 FILLER_29_145 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_160 ();
 sg13g2_decap_8 FILLER_29_167 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_207 ();
 sg13g2_fill_1 FILLER_29_234 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_282 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_4 FILLER_29_322 ();
 sg13g2_decap_8 FILLER_29_329 ();
 sg13g2_fill_1 FILLER_29_336 ();
 sg13g2_decap_8 FILLER_29_341 ();
 sg13g2_fill_2 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_350 ();
 sg13g2_decap_4 FILLER_29_377 ();
 sg13g2_fill_2 FILLER_29_381 ();
 sg13g2_decap_8 FILLER_29_391 ();
 sg13g2_fill_2 FILLER_29_398 ();
 sg13g2_decap_8 FILLER_29_421 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_4 FILLER_30_14 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_28 ();
 sg13g2_fill_2 FILLER_30_43 ();
 sg13g2_fill_1 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_50 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_84 ();
 sg13g2_fill_2 FILLER_30_118 ();
 sg13g2_fill_2 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_148 ();
 sg13g2_fill_1 FILLER_30_154 ();
 sg13g2_fill_2 FILLER_30_181 ();
 sg13g2_fill_1 FILLER_30_183 ();
 sg13g2_decap_8 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_195 ();
 sg13g2_decap_8 FILLER_30_201 ();
 sg13g2_fill_2 FILLER_30_208 ();
 sg13g2_fill_1 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_fill_2 FILLER_30_252 ();
 sg13g2_fill_1 FILLER_30_254 ();
 sg13g2_decap_8 FILLER_30_263 ();
 sg13g2_fill_1 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_284 ();
 sg13g2_fill_2 FILLER_30_290 ();
 sg13g2_fill_2 FILLER_30_299 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_312 ();
 sg13g2_fill_1 FILLER_30_319 ();
 sg13g2_decap_4 FILLER_30_350 ();
 sg13g2_fill_2 FILLER_30_354 ();
 sg13g2_decap_4 FILLER_30_360 ();
 sg13g2_decap_4 FILLER_30_368 ();
 sg13g2_decap_8 FILLER_30_395 ();
 sg13g2_decap_4 FILLER_30_402 ();
 sg13g2_fill_2 FILLER_30_406 ();
 sg13g2_fill_1 FILLER_30_416 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_51 ();
 sg13g2_decap_8 FILLER_31_58 ();
 sg13g2_decap_8 FILLER_31_65 ();
 sg13g2_decap_8 FILLER_31_76 ();
 sg13g2_decap_8 FILLER_31_109 ();
 sg13g2_decap_8 FILLER_31_116 ();
 sg13g2_decap_8 FILLER_31_123 ();
 sg13g2_decap_8 FILLER_31_130 ();
 sg13g2_decap_8 FILLER_31_137 ();
 sg13g2_fill_2 FILLER_31_144 ();
 sg13g2_fill_1 FILLER_31_173 ();
 sg13g2_fill_1 FILLER_31_181 ();
 sg13g2_decap_4 FILLER_31_185 ();
 sg13g2_fill_1 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_199 ();
 sg13g2_fill_2 FILLER_31_206 ();
 sg13g2_fill_1 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_230 ();
 sg13g2_decap_8 FILLER_31_236 ();
 sg13g2_decap_8 FILLER_31_243 ();
 sg13g2_fill_2 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_decap_8 FILLER_31_276 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_1 FILLER_31_285 ();
 sg13g2_decap_4 FILLER_31_296 ();
 sg13g2_fill_2 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_346 ();
 sg13g2_fill_2 FILLER_31_353 ();
 sg13g2_decap_4 FILLER_31_359 ();
 sg13g2_fill_1 FILLER_31_363 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_fill_2 FILLER_31_380 ();
 sg13g2_fill_1 FILLER_31_382 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_4 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_417 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_4 FILLER_32_35 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_4 FILLER_32_102 ();
 sg13g2_fill_2 FILLER_32_106 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_152 ();
 sg13g2_decap_8 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_191 ();
 sg13g2_decap_8 FILLER_32_198 ();
 sg13g2_decap_4 FILLER_32_205 ();
 sg13g2_decap_4 FILLER_32_221 ();
 sg13g2_decap_4 FILLER_32_239 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_fill_2 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_fill_1 FILLER_32_276 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_decap_8 FILLER_32_292 ();
 sg13g2_decap_4 FILLER_32_299 ();
 sg13g2_fill_2 FILLER_32_303 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_decap_4 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_332 ();
 sg13g2_decap_4 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_362 ();
 sg13g2_fill_1 FILLER_32_373 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_1 FILLER_32_392 ();
 sg13g2_decap_8 FILLER_32_398 ();
 sg13g2_decap_4 FILLER_32_425 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_4 FILLER_33_91 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_128 ();
 sg13g2_decap_4 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_159 ();
 sg13g2_decap_4 FILLER_33_166 ();
 sg13g2_fill_2 FILLER_33_170 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_4 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_204 ();
 sg13g2_fill_1 FILLER_33_208 ();
 sg13g2_decap_8 FILLER_33_214 ();
 sg13g2_fill_1 FILLER_33_221 ();
 sg13g2_fill_1 FILLER_33_227 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_decap_8 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_fill_1 FILLER_33_274 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_1 FILLER_33_288 ();
 sg13g2_fill_1 FILLER_33_293 ();
 sg13g2_decap_4 FILLER_33_306 ();
 sg13g2_decap_8 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_338 ();
 sg13g2_fill_1 FILLER_33_358 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_377 ();
 sg13g2_fill_2 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_400 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_decap_8 FILLER_34_77 ();
 sg13g2_decap_8 FILLER_34_84 ();
 sg13g2_decap_8 FILLER_34_91 ();
 sg13g2_decap_8 FILLER_34_98 ();
 sg13g2_decap_8 FILLER_34_109 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_fill_1 FILLER_34_120 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_fill_2 FILLER_34_137 ();
 sg13g2_decap_4 FILLER_34_201 ();
 sg13g2_fill_1 FILLER_34_205 ();
 sg13g2_fill_1 FILLER_34_217 ();
 sg13g2_fill_2 FILLER_34_223 ();
 sg13g2_fill_2 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_239 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_decap_4 FILLER_34_250 ();
 sg13g2_fill_1 FILLER_34_277 ();
 sg13g2_decap_4 FILLER_34_287 ();
 sg13g2_fill_2 FILLER_34_291 ();
 sg13g2_fill_2 FILLER_34_306 ();
 sg13g2_decap_4 FILLER_34_321 ();
 sg13g2_fill_2 FILLER_34_334 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_fill_2 FILLER_34_345 ();
 sg13g2_fill_1 FILLER_34_347 ();
 sg13g2_decap_4 FILLER_34_352 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_decap_8 FILLER_34_379 ();
 sg13g2_decap_8 FILLER_34_386 ();
 sg13g2_decap_8 FILLER_34_393 ();
 sg13g2_decap_8 FILLER_34_400 ();
 sg13g2_decap_8 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_4 FILLER_35_91 ();
 sg13g2_fill_1 FILLER_35_95 ();
 sg13g2_decap_8 FILLER_35_130 ();
 sg13g2_decap_8 FILLER_35_137 ();
 sg13g2_fill_1 FILLER_35_148 ();
 sg13g2_decap_8 FILLER_35_153 ();
 sg13g2_decap_8 FILLER_35_160 ();
 sg13g2_fill_2 FILLER_35_167 ();
 sg13g2_decap_8 FILLER_35_173 ();
 sg13g2_decap_4 FILLER_35_180 ();
 sg13g2_decap_4 FILLER_35_188 ();
 sg13g2_fill_2 FILLER_35_192 ();
 sg13g2_fill_2 FILLER_35_207 ();
 sg13g2_fill_1 FILLER_35_209 ();
 sg13g2_decap_8 FILLER_35_219 ();
 sg13g2_decap_8 FILLER_35_226 ();
 sg13g2_decap_8 FILLER_35_233 ();
 sg13g2_decap_4 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_244 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_257 ();
 sg13g2_decap_8 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_282 ();
 sg13g2_decap_4 FILLER_35_295 ();
 sg13g2_fill_1 FILLER_35_307 ();
 sg13g2_decap_4 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_326 ();
 sg13g2_decap_8 FILLER_35_341 ();
 sg13g2_decap_8 FILLER_35_348 ();
 sg13g2_decap_4 FILLER_35_355 ();
 sg13g2_fill_1 FILLER_35_359 ();
 sg13g2_decap_8 FILLER_35_363 ();
 sg13g2_fill_1 FILLER_35_370 ();
 sg13g2_decap_4 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_35_390 ();
 sg13g2_fill_1 FILLER_35_392 ();
 sg13g2_fill_1 FILLER_35_403 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_415 ();
 sg13g2_decap_8 FILLER_35_422 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_fill_2 FILLER_36_98 ();
 sg13g2_fill_1 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_fill_2 FILLER_36_112 ();
 sg13g2_fill_2 FILLER_36_117 ();
 sg13g2_decap_8 FILLER_36_131 ();
 sg13g2_decap_8 FILLER_36_138 ();
 sg13g2_fill_2 FILLER_36_145 ();
 sg13g2_fill_1 FILLER_36_179 ();
 sg13g2_decap_8 FILLER_36_184 ();
 sg13g2_decap_4 FILLER_36_194 ();
 sg13g2_fill_2 FILLER_36_198 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_fill_1 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_221 ();
 sg13g2_fill_2 FILLER_36_228 ();
 sg13g2_fill_1 FILLER_36_230 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_4 FILLER_36_266 ();
 sg13g2_fill_1 FILLER_36_270 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_fill_1 FILLER_36_282 ();
 sg13g2_decap_4 FILLER_36_299 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_fill_2 FILLER_36_343 ();
 sg13g2_fill_1 FILLER_36_345 ();
 sg13g2_fill_1 FILLER_36_363 ();
 sg13g2_fill_2 FILLER_36_385 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_2 FILLER_36_398 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_decap_8 FILLER_36_412 ();
 sg13g2_decap_8 FILLER_36_419 ();
 sg13g2_decap_4 FILLER_36_426 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_8 FILLER_37_28 ();
 sg13g2_decap_8 FILLER_37_35 ();
 sg13g2_decap_8 FILLER_37_42 ();
 sg13g2_decap_8 FILLER_37_49 ();
 sg13g2_decap_8 FILLER_37_56 ();
 sg13g2_decap_8 FILLER_37_63 ();
 sg13g2_decap_8 FILLER_37_70 ();
 sg13g2_decap_8 FILLER_37_77 ();
 sg13g2_decap_8 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_91 ();
 sg13g2_fill_2 FILLER_37_97 ();
 sg13g2_decap_4 FILLER_37_129 ();
 sg13g2_decap_4 FILLER_37_163 ();
 sg13g2_fill_2 FILLER_37_167 ();
 sg13g2_decap_4 FILLER_37_195 ();
 sg13g2_fill_2 FILLER_37_199 ();
 sg13g2_fill_2 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_220 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_decap_8 FILLER_37_234 ();
 sg13g2_decap_8 FILLER_37_241 ();
 sg13g2_decap_8 FILLER_37_248 ();
 sg13g2_decap_8 FILLER_37_255 ();
 sg13g2_decap_8 FILLER_37_262 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_300 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_2 FILLER_37_324 ();
 sg13g2_decap_8 FILLER_37_330 ();
 sg13g2_fill_2 FILLER_37_337 ();
 sg13g2_fill_1 FILLER_37_339 ();
 sg13g2_fill_2 FILLER_37_345 ();
 sg13g2_fill_1 FILLER_37_352 ();
 sg13g2_fill_2 FILLER_37_371 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_392 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_72 ();
 sg13g2_fill_1 FILLER_38_197 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_242 ();
 sg13g2_fill_2 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_299 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_decap_8 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_320 ();
 sg13g2_decap_8 FILLER_38_327 ();
 sg13g2_decap_8 FILLER_38_334 ();
 sg13g2_decap_4 FILLER_38_351 ();
 sg13g2_fill_2 FILLER_38_363 ();
 sg13g2_fill_2 FILLER_38_412 ();
 sg13g2_fill_1 FILLER_38_414 ();
 sg13g2_decap_8 FILLER_38_419 ();
 sg13g2_decap_4 FILLER_38_426 ();
endmodule
