module tt_um_dvxf_dj8v (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire \DJ8.ACC[0] ;
 wire \DJ8.ACC[1] ;
 wire \DJ8.ACC[2] ;
 wire \DJ8.ACC[3] ;
 wire \DJ8.ACC[4] ;
 wire \DJ8.ACC[5] ;
 wire \DJ8.ACC[6] ;
 wire \DJ8.ACC[7] ;
 wire \DJ8.ALU.c_in ;
 wire \DJ8.ALU.opalu[0] ;
 wire \DJ8.ALU.opalu[1] ;
 wire \DJ8.ALU.opalu[2] ;
 wire \DJ8.EF[0] ;
 wire \DJ8.EF[10] ;
 wire \DJ8.EF[11] ;
 wire \DJ8.EF[12] ;
 wire \DJ8.EF[13] ;
 wire \DJ8.EF[14] ;
 wire \DJ8.EF[15] ;
 wire \DJ8.EF[1] ;
 wire \DJ8.EF[2] ;
 wire \DJ8.EF[3] ;
 wire \DJ8.EF[4] ;
 wire \DJ8.EF[5] ;
 wire \DJ8.EF[6] ;
 wire \DJ8.EF[7] ;
 wire \DJ8.EF[8] ;
 wire \DJ8.EF[9] ;
 wire \DJ8.GH[0] ;
 wire \DJ8.GH[10] ;
 wire \DJ8.GH[11] ;
 wire \DJ8.GH[12] ;
 wire \DJ8.GH[13] ;
 wire \DJ8.GH[14] ;
 wire \DJ8.GH[15] ;
 wire \DJ8.GH[1] ;
 wire \DJ8.GH[2] ;
 wire \DJ8.GH[3] ;
 wire \DJ8.GH[4] ;
 wire \DJ8.GH[5] ;
 wire \DJ8.GH[6] ;
 wire \DJ8.GH[7] ;
 wire \DJ8.GH[8] ;
 wire \DJ8.GH[9] ;
 wire \DJ8.REGS.regs[1][0] ;
 wire \DJ8.REGS.regs[1][1] ;
 wire \DJ8.REGS.regs[1][2] ;
 wire \DJ8.REGS.regs[1][3] ;
 wire \DJ8.REGS.regs[1][4] ;
 wire \DJ8.REGS.regs[1][5] ;
 wire \DJ8.REGS.regs[1][6] ;
 wire \DJ8.REGS.regs[1][7] ;
 wire \DJ8.REGS.regs[2][0] ;
 wire \DJ8.REGS.regs[2][1] ;
 wire \DJ8.REGS.regs[2][2] ;
 wire \DJ8.REGS.regs[2][3] ;
 wire \DJ8.REGS.regs[2][4] ;
 wire \DJ8.REGS.regs[2][5] ;
 wire \DJ8.REGS.regs[2][6] ;
 wire \DJ8.REGS.regs[2][7] ;
 wire \DJ8.REGS.regs[3][0] ;
 wire \DJ8.REGS.regs[3][1] ;
 wire \DJ8.REGS.regs[3][2] ;
 wire \DJ8.REGS.regs[3][3] ;
 wire \DJ8.REGS.regs[3][4] ;
 wire \DJ8.REGS.regs[3][5] ;
 wire \DJ8.REGS.regs[3][6] ;
 wire \DJ8.REGS.regs[3][7] ;
 wire \DJ8.REGS.write_addr[0] ;
 wire \DJ8.REGS.write_addr[1] ;
 wire \DJ8.REGS.write_addr[2] ;
 wire \DJ8.flag_Z ;
 wire \DJ8.ir[0] ;
 wire \DJ8.ir[14] ;
 wire \DJ8.ir[15] ;
 wire \DJ8.ir[1] ;
 wire \DJ8.ir[2] ;
 wire \DJ8.ir[3] ;
 wire \DJ8.ir[4] ;
 wire \DJ8.ir[5] ;
 wire \DJ8.ir[6] ;
 wire \DJ8.ir[7] ;
 wire \DJ8.pc[0] ;
 wire \DJ8.pc[10] ;
 wire \DJ8.pc[11] ;
 wire \DJ8.pc[12] ;
 wire \DJ8.pc[13] ;
 wire \DJ8.pc[14] ;
 wire \DJ8.pc[1] ;
 wire \DJ8.pc[2] ;
 wire \DJ8.pc[3] ;
 wire \DJ8.pc[4] ;
 wire \DJ8.pc[5] ;
 wire \DJ8.pc[6] ;
 wire \DJ8.pc[7] ;
 wire \DJ8.pc[8] ;
 wire \DJ8.pc[9] ;
 wire \DJ8.state[0] ;
 wire \DJ8.state[1] ;
 wire \DJ8.state[2] ;
 wire \DJ8.state[3] ;
 wire \DJ8.we ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire clknet_0_clk;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire net115;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][0]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net103),
    .D(_0038_),
    .Q_N(_1549_),
    .Q(\DJ8.ACC[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][1]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net103),
    .D(_0039_),
    .Q_N(_0015_),
    .Q(\DJ8.ACC[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net103),
    .D(_0040_),
    .Q_N(_0017_),
    .Q(\DJ8.ACC[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][3]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net103),
    .D(_0041_),
    .Q_N(_0019_),
    .Q(\DJ8.ACC[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][4]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0042_),
    .Q_N(_0020_),
    .Q(\DJ8.ACC[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][5]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net103),
    .D(_0043_),
    .Q_N(_0022_),
    .Q(\DJ8.ACC[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][6]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0044_),
    .Q_N(_0024_),
    .Q(\DJ8.ACC[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[0][7]$_DFFE_PN1P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0045_),
    .Q_N(\DJ8.ACC[7] ),
    .Q(_0026_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][0]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net95),
    .D(_0046_),
    .Q_N(_1548_),
    .Q(\DJ8.REGS.regs[1][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][1]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0047_),
    .Q_N(_1547_),
    .Q(\DJ8.REGS.regs[1][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][2]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net94),
    .D(_0048_),
    .Q_N(_1546_),
    .Q(\DJ8.REGS.regs[1][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][3]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(_0049_),
    .Q_N(_1545_),
    .Q(\DJ8.REGS.regs[1][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][4]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(_0050_),
    .Q_N(_1544_),
    .Q(\DJ8.REGS.regs[1][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][5]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_0051_),
    .Q_N(_1543_),
    .Q(\DJ8.REGS.regs[1][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][6]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0052_),
    .Q_N(_1542_),
    .Q(\DJ8.REGS.regs[1][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[1][7]$_DFFE_PN1P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0053_),
    .Q_N(\DJ8.REGS.regs[1][7] ),
    .Q(_0027_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][0]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net95),
    .D(_0054_),
    .Q_N(_1541_),
    .Q(\DJ8.REGS.regs[2][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][1]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_0055_),
    .Q_N(_1540_),
    .Q(\DJ8.REGS.regs[2][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net95),
    .D(_0056_),
    .Q_N(_1539_),
    .Q(\DJ8.REGS.regs[2][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][3]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net90),
    .D(_0057_),
    .Q_N(_1538_),
    .Q(\DJ8.REGS.regs[2][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][4]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0058_),
    .Q_N(_1537_),
    .Q(\DJ8.REGS.regs[2][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][5]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0059_),
    .Q_N(_1536_),
    .Q(\DJ8.REGS.regs[2][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][6]$_DFFE_PN0P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net94),
    .D(_0060_),
    .Q_N(_1535_),
    .Q(\DJ8.REGS.regs[2][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[2][7]$_DFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0061_),
    .Q_N(\DJ8.REGS.regs[2][7] ),
    .Q(_0028_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][0]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net95),
    .D(_0062_),
    .Q_N(_1534_),
    .Q(\DJ8.REGS.regs[3][0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][1]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0063_),
    .Q_N(_1533_),
    .Q(\DJ8.REGS.regs[3][1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][2]$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net103),
    .D(_0064_),
    .Q_N(_1532_),
    .Q(\DJ8.REGS.regs[3][2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][3]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(_0065_),
    .Q_N(_1531_),
    .Q(\DJ8.REGS.regs[3][3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][4]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(_0066_),
    .Q_N(_1530_),
    .Q(\DJ8.REGS.regs[3][4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][5]$_DFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net89),
    .D(_0067_),
    .Q_N(_1529_),
    .Q(\DJ8.REGS.regs[3][5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][6]$_DFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net94),
    .D(_0068_),
    .Q_N(_1528_),
    .Q(\DJ8.REGS.regs[3][6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[3][7]$_DFFE_PN1P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net90),
    .D(_0069_),
    .Q_N(\DJ8.REGS.regs[3][7] ),
    .Q(_0029_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][0]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0070_),
    .Q_N(_1527_),
    .Q(\DJ8.EF[8] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][1]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net89),
    .D(_0071_),
    .Q_N(_1526_),
    .Q(\DJ8.EF[9] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][2]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0072_),
    .Q_N(_1525_),
    .Q(\DJ8.EF[10] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][3]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net93),
    .D(_0073_),
    .Q_N(_1524_),
    .Q(\DJ8.EF[11] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][4]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net93),
    .D(_0074_),
    .Q_N(_1523_),
    .Q(\DJ8.EF[12] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][5]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net91),
    .D(_0075_),
    .Q_N(_1522_),
    .Q(\DJ8.EF[13] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][6]$_DFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net90),
    .D(_0076_),
    .Q_N(_1521_),
    .Q(\DJ8.EF[14] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[4][7]$_DFFE_PN1P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0077_),
    .Q_N(\DJ8.EF[15] ),
    .Q(_0030_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][0]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net96),
    .D(_0078_),
    .Q_N(_1520_),
    .Q(\DJ8.EF[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][1]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(_0079_),
    .Q_N(_0008_),
    .Q(\DJ8.EF[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][2]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net96),
    .D(_0080_),
    .Q_N(_0011_),
    .Q(\DJ8.EF[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][3]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0081_),
    .Q_N(_1519_),
    .Q(\DJ8.EF[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][4]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0082_),
    .Q_N(_1518_),
    .Q(\DJ8.EF[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][5]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net91),
    .D(_0083_),
    .Q_N(_1517_),
    .Q(\DJ8.EF[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][6]$_DFFE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net92),
    .D(_0084_),
    .Q_N(_1516_),
    .Q(\DJ8.EF[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[5][7]$_DFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net91),
    .D(_0085_),
    .Q_N(\DJ8.EF[7] ),
    .Q(_0031_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][0]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net92),
    .D(_0086_),
    .Q_N(_1515_),
    .Q(\DJ8.GH[8] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][1]$_DFFE_PN0P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net91),
    .D(_0087_),
    .Q_N(_1514_),
    .Q(\DJ8.GH[9] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][2]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net100),
    .D(_0088_),
    .Q_N(_1513_),
    .Q(\DJ8.GH[10] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][3]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0089_),
    .Q_N(_1512_),
    .Q(\DJ8.GH[11] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][4]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0090_),
    .Q_N(_1511_),
    .Q(\DJ8.GH[12] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][5]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0091_),
    .Q_N(_1510_),
    .Q(\DJ8.GH[13] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][6]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net99),
    .D(_0092_),
    .Q_N(_1509_),
    .Q(\DJ8.GH[14] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[6][7]$_DFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net91),
    .D(_0093_),
    .Q_N(\DJ8.GH[15] ),
    .Q(_0032_));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][0]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0094_),
    .Q_N(_1508_),
    .Q(\DJ8.GH[0] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][1]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net96),
    .D(_0095_),
    .Q_N(_0007_),
    .Q(\DJ8.GH[1] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][2]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net100),
    .D(_0096_),
    .Q_N(_0010_),
    .Q(\DJ8.GH[2] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][3]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net100),
    .D(_0097_),
    .Q_N(_1507_),
    .Q(\DJ8.GH[3] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][4]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0098_),
    .Q_N(_1506_),
    .Q(\DJ8.GH[4] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][5]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0099_),
    .Q_N(_1505_),
    .Q(\DJ8.GH[5] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][6]$_DFFE_PN0P_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net99),
    .D(_0100_),
    .Q_N(_1504_),
    .Q(\DJ8.GH[6] ));
 sg13g2_dfrbp_1 \DJ8.REGS.regs[7][7]$_DFFE_PN1P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net92),
    .D(_0101_),
    .Q_N(\DJ8.GH[7] ),
    .Q(_0033_));
 sg13g2_dfrbp_1 \DJ8.flag_C$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net103),
    .D(_0102_),
    .Q_N(_1503_),
    .Q(\DJ8.ALU.c_in ));
 sg13g2_dfrbp_1 \DJ8.flag_Z$_DFFE_PN0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net103),
    .D(_0103_),
    .Q_N(_1502_),
    .Q(\DJ8.flag_Z ));
 sg13g2_dfrbp_1 \DJ8.ir[0]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net106),
    .D(_0104_),
    .Q_N(_1501_),
    .Q(\DJ8.ir[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[10]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0105_),
    .Q_N(_0001_),
    .Q(\DJ8.REGS.write_addr[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[11]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net105),
    .D(_0106_),
    .Q_N(_1500_),
    .Q(\DJ8.ALU.opalu[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[12]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net105),
    .D(_0107_),
    .Q_N(_1499_),
    .Q(\DJ8.ALU.opalu[1] ));
 sg13g2_dfrbp_1 \DJ8.ir[13]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net105),
    .D(_0108_),
    .Q_N(_0013_),
    .Q(\DJ8.ALU.opalu[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[14]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net104),
    .D(_0109_),
    .Q_N(_1498_),
    .Q(\DJ8.ir[14] ));
 sg13g2_dfrbp_1 \DJ8.ir[15]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net100),
    .D(_0110_),
    .Q_N(_1497_),
    .Q(\DJ8.ir[15] ));
 sg13g2_dfrbp_1 \DJ8.ir[1]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net104),
    .D(_0111_),
    .Q_N(_0014_),
    .Q(\DJ8.ir[1] ));
 sg13g2_dfrbp_1 \DJ8.ir[2]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net104),
    .D(_0112_),
    .Q_N(_0016_),
    .Q(\DJ8.ir[2] ));
 sg13g2_dfrbp_1 \DJ8.ir[3]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net104),
    .D(_0113_),
    .Q_N(_0018_),
    .Q(\DJ8.ir[3] ));
 sg13g2_dfrbp_1 \DJ8.ir[4]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net100),
    .D(_0114_),
    .Q_N(_0005_),
    .Q(\DJ8.ir[4] ));
 sg13g2_dfrbp_1 \DJ8.ir[5]$_DFFE_PN0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net104),
    .D(_0115_),
    .Q_N(_0021_),
    .Q(\DJ8.ir[5] ));
 sg13g2_dfrbp_1 \DJ8.ir[6]$_DFFE_PN0P_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net96),
    .D(_0116_),
    .Q_N(_0023_),
    .Q(\DJ8.ir[6] ));
 sg13g2_dfrbp_1 \DJ8.ir[7]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net106),
    .D(_0117_),
    .Q_N(_0003_),
    .Q(\DJ8.ir[7] ));
 sg13g2_dfrbp_1 \DJ8.ir[8]$_DFFE_PN0P_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net105),
    .D(_0118_),
    .Q_N(_1496_),
    .Q(\DJ8.REGS.write_addr[0] ));
 sg13g2_dfrbp_1 \DJ8.ir[9]$_DFFE_PN0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net97),
    .D(_0119_),
    .Q_N(_1495_),
    .Q(\DJ8.REGS.write_addr[1] ));
 sg13g2_dfrbp_1 \DJ8.pc[0]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net100),
    .D(_0120_),
    .Q_N(_0006_),
    .Q(\DJ8.pc[0] ));
 sg13g2_dfrbp_1 \DJ8.pc[10]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0121_),
    .Q_N(_1494_),
    .Q(\DJ8.pc[10] ));
 sg13g2_dfrbp_1 \DJ8.pc[11]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0122_),
    .Q_N(_1493_),
    .Q(\DJ8.pc[11] ));
 sg13g2_dfrbp_1 \DJ8.pc[12]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0123_),
    .Q_N(_1492_),
    .Q(\DJ8.pc[12] ));
 sg13g2_dfrbp_1 \DJ8.pc[13]$_DFFE_PN1P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0124_),
    .Q_N(\DJ8.pc[13] ),
    .Q(_0034_));
 sg13g2_dfrbp_1 \DJ8.pc[14]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0125_),
    .Q_N(_0004_),
    .Q(\DJ8.pc[14] ));
 sg13g2_dfrbp_1 \DJ8.pc[1]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net100),
    .D(_0126_),
    .Q_N(_0009_),
    .Q(\DJ8.pc[1] ));
 sg13g2_dfrbp_1 \DJ8.pc[2]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net100),
    .D(_0127_),
    .Q_N(_1491_),
    .Q(\DJ8.pc[2] ));
 sg13g2_dfrbp_1 \DJ8.pc[3]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_0128_),
    .Q_N(_1490_),
    .Q(\DJ8.pc[3] ));
 sg13g2_dfrbp_1 \DJ8.pc[4]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net98),
    .D(_0129_),
    .Q_N(_0012_),
    .Q(\DJ8.pc[4] ));
 sg13g2_dfrbp_1 \DJ8.pc[5]$_DFFE_PN0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net98),
    .D(_0130_),
    .Q_N(_1489_),
    .Q(\DJ8.pc[5] ));
 sg13g2_dfrbp_1 \DJ8.pc[6]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net99),
    .D(_0131_),
    .Q_N(_1488_),
    .Q(\DJ8.pc[6] ));
 sg13g2_dfrbp_1 \DJ8.pc[7]$_DFFE_PN0P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net101),
    .D(_0132_),
    .Q_N(_1487_),
    .Q(\DJ8.pc[7] ));
 sg13g2_dfrbp_1 \DJ8.pc[8]$_DFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net98),
    .D(_0133_),
    .Q_N(_1486_),
    .Q(\DJ8.pc[8] ));
 sg13g2_dfrbp_1 \DJ8.pc[9]$_DFFE_PN0P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_0134_),
    .Q_N(_1485_),
    .Q(\DJ8.pc[9] ));
 sg13g2_dfrbp_1 \DJ8.state[0]$_DFF_PN1_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_0036_),
    .Q_N(\DJ8.state[0] ),
    .Q(_1551_));
 sg13g2_dfrbp_1 \DJ8.state[1]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(\DJ8.state[2] ),
    .Q_N(_0002_),
    .Q(\DJ8.state[1] ));
 sg13g2_dfrbp_1 \DJ8.state[2]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(\DJ8.state[0] ),
    .Q_N(_1550_),
    .Q(\DJ8.state[2] ));
 sg13g2_dfrbp_1 \DJ8.state[3]$_DFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net101),
    .D(_0000_),
    .Q_N(_0025_),
    .Q(\DJ8.state[3] ));
 sg13g2_dfrbp_1 \DJ8.we$_DFFE_NN1P_  (.CLK(net115),
    .RESET_B(net101),
    .D(_0135_),
    .Q_N(\DJ8.we ),
    .Q(_0035_));
 sg13g2_buf_8 _1553_ (.A(\DJ8.ir[0] ),
    .X(_0752_));
 sg13g2_inv_1 _1554_ (.Y(_0753_),
    .A(_0752_));
 sg13g2_buf_8 _1555_ (.A(\DJ8.ir[14] ),
    .X(_0754_));
 sg13g2_inv_8 _1556_ (.Y(_0755_),
    .A(_0754_));
 sg13g2_nand2_1 _1557_ (.Y(_0756_),
    .A(_0755_),
    .B(\DJ8.ir[15] ));
 sg13g2_nor2_1 _1558_ (.A(_0753_),
    .B(_0756_),
    .Y(_0757_));
 sg13g2_inv_1 _1559_ (.Y(_0758_),
    .A(_0757_));
 sg13g2_nor2_1 _1560_ (.A(_0002_),
    .B(_0758_),
    .Y(_0000_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_inv_1 _1562_ (.Y(_0759_),
    .A(\DJ8.ACC[0] ));
 sg13g2_buf_2 _1563_ (.A(\DJ8.REGS.write_addr[1] ),
    .X(_0760_));
 sg13g2_buf_2 _1564_ (.A(\DJ8.REGS.write_addr[0] ),
    .X(_0761_));
 sg13g2_buf_1 _1565_ (.A(\DJ8.state[1] ),
    .X(_0762_));
 sg13g2_nand2_1 _1566_ (.Y(_0763_),
    .A(\DJ8.ir[15] ),
    .B(_0762_));
 sg13g2_a21oi_1 _1567_ (.A1(_0752_),
    .A2(_0755_),
    .Y(_0764_),
    .B1(_0763_));
 sg13g2_inv_1 _1568_ (.Y(_0765_),
    .A(_0764_));
 sg13g2_nor2_1 _1569_ (.A(\DJ8.REGS.write_addr[2] ),
    .B(_0765_),
    .Y(_0766_));
 sg13g2_inv_2 _1570_ (.Y(_0767_),
    .A(_0766_));
 sg13g2_nor3_2 _1571_ (.A(_0760_),
    .B(_0761_),
    .C(_0767_),
    .Y(_0768_));
 sg13g2_buf_1 _1572_ (.A(_0768_),
    .X(_0769_));
 sg13g2_nor2_1 _1573_ (.A(_0752_),
    .B(\DJ8.ir[1] ),
    .Y(_0770_));
 sg13g2_nor2_1 _1574_ (.A(_0770_),
    .B(_0756_),
    .Y(_0771_));
 sg13g2_buf_1 _1575_ (.A(\DJ8.state[2] ),
    .X(_0772_));
 sg13g2_buf_1 _1576_ (.A(\DJ8.state[0] ),
    .X(_0773_));
 sg13g2_nor2_1 _1577_ (.A(_0772_),
    .B(_0773_),
    .Y(_0774_));
 sg13g2_nand2_2 _1578_ (.Y(_0775_),
    .A(_0771_),
    .B(_0774_));
 sg13g2_buf_1 _1579_ (.A(_0775_),
    .X(_0776_));
 sg13g2_buf_1 _1580_ (.A(\DJ8.ir[4] ),
    .X(_0777_));
 sg13g2_buf_1 _1581_ (.A(_0777_),
    .X(_0778_));
 sg13g2_buf_1 _1582_ (.A(net87),
    .X(_0779_));
 sg13g2_inv_1 _1583_ (.Y(_0780_),
    .A(\DJ8.GH[7] ));
 sg13g2_nor2_1 _1584_ (.A(net87),
    .B(_0780_),
    .Y(_0781_));
 sg13g2_a21oi_1 _1585_ (.A1(net84),
    .A2(\DJ8.EF[7] ),
    .Y(_0782_),
    .B1(_0781_));
 sg13g2_nor2_1 _1586_ (.A(_0782_),
    .B(net74),
    .Y(_0783_));
 sg13g2_a21oi_2 _1587_ (.B1(_0783_),
    .Y(_0784_),
    .A2(net74),
    .A1(\DJ8.pc[6] ));
 sg13g2_inv_1 _1588_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_nor2b_1 _1589_ (.A(_0770_),
    .B_N(_0755_),
    .Y(_0786_));
 sg13g2_inv_1 _1590_ (.Y(_0787_),
    .A(\DJ8.ir[15] ));
 sg13g2_nor2_1 _1591_ (.A(net88),
    .B(_0787_),
    .Y(_0788_));
 sg13g2_nand2_2 _1592_ (.Y(_0789_),
    .A(_0786_),
    .B(_0788_));
 sg13g2_inv_1 _1593_ (.Y(_0790_),
    .A(_0010_));
 sg13g2_nand2_1 _1594_ (.Y(_0791_),
    .A(_0777_),
    .B(_0011_));
 sg13g2_o21ai_1 _1595_ (.B1(_0791_),
    .Y(_0792_),
    .A1(_0778_),
    .A2(_0790_));
 sg13g2_nor2b_2 _1596_ (.A(_0789_),
    .B_N(_0792_),
    .Y(_0793_));
 sg13g2_nand2_1 _1597_ (.Y(_0794_),
    .A(_0789_),
    .B(_0009_));
 sg13g2_inv_2 _1598_ (.Y(_0795_),
    .A(_0773_));
 sg13g2_nand2_1 _1599_ (.Y(_0796_),
    .A(_0794_),
    .B(_0795_));
 sg13g2_nor2_1 _1600_ (.A(_0793_),
    .B(_0796_),
    .Y(_0797_));
 sg13g2_buf_1 _1601_ (.A(_0773_),
    .X(_0798_));
 sg13g2_nand2b_1 _1602_ (.Y(_0799_),
    .B(net86),
    .A_N(_0009_));
 sg13g2_nor2b_1 _1603_ (.A(_0797_),
    .B_N(_0799_),
    .Y(_0800_));
 sg13g2_buf_2 _1604_ (.A(_0800_),
    .X(_0801_));
 sg13g2_inv_1 _1605_ (.Y(_0802_),
    .A(_0777_));
 sg13g2_nand2_1 _1606_ (.Y(_0803_),
    .A(_0802_),
    .B(_0007_));
 sg13g2_nand2_1 _1607_ (.Y(_0804_),
    .A(_0777_),
    .B(_0008_));
 sg13g2_nand2_1 _1608_ (.Y(_0805_),
    .A(_0803_),
    .B(_0804_));
 sg13g2_nand3_1 _1609_ (.B(_0786_),
    .C(_0788_),
    .A(_0805_),
    .Y(_0806_));
 sg13g2_nand2_1 _1610_ (.Y(_0807_),
    .A(_0789_),
    .B(_0006_));
 sg13g2_nand3_1 _1611_ (.B(_0807_),
    .C(_0795_),
    .A(_0806_),
    .Y(_0808_));
 sg13g2_buf_1 _1612_ (.A(_0808_),
    .X(_0809_));
 sg13g2_inv_1 _1613_ (.Y(_0810_),
    .A(\DJ8.GH[0] ));
 sg13g2_nand2_1 _1614_ (.Y(_0811_),
    .A(_0810_),
    .B(_0802_));
 sg13g2_inv_1 _1615_ (.Y(_0812_),
    .A(\DJ8.EF[0] ));
 sg13g2_nand2_1 _1616_ (.Y(_0813_),
    .A(_0812_),
    .B(_0777_));
 sg13g2_nand2_1 _1617_ (.Y(_0814_),
    .A(_0811_),
    .B(_0813_));
 sg13g2_nor2b_2 _1618_ (.A(_0789_),
    .B_N(_0814_),
    .Y(_0815_));
 sg13g2_nor2_2 _1619_ (.A(_0773_),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_inv_4 _1620_ (.A(_0816_),
    .Y(_0817_));
 sg13g2_nor2_1 _1621_ (.A(_0006_),
    .B(_0795_),
    .Y(_0818_));
 sg13g2_inv_1 _1622_ (.Y(_0819_),
    .A(_0818_));
 sg13g2_nand3_1 _1623_ (.B(_0817_),
    .C(_0819_),
    .A(net71),
    .Y(_0820_));
 sg13g2_buf_2 _1624_ (.A(_0820_),
    .X(_0821_));
 sg13g2_nor2_1 _1625_ (.A(_0801_),
    .B(_0821_),
    .Y(_0822_));
 sg13g2_inv_1 _1626_ (.Y(_0823_),
    .A(_0775_));
 sg13g2_mux2_1 _1627_ (.A0(\DJ8.GH[3] ),
    .A1(\DJ8.EF[3] ),
    .S(net87),
    .X(_0824_));
 sg13g2_nand2_1 _1628_ (.Y(_0825_),
    .A(_0823_),
    .B(_0824_));
 sg13g2_nand2_1 _1629_ (.Y(_0826_),
    .A(_0775_),
    .B(\DJ8.pc[2] ));
 sg13g2_nand2_2 _1630_ (.Y(_0827_),
    .A(_0825_),
    .B(_0826_));
 sg13g2_inv_1 _1631_ (.Y(_0828_),
    .A(\DJ8.GH[4] ));
 sg13g2_nand2_1 _1632_ (.Y(_0829_),
    .A(net87),
    .B(\DJ8.EF[4] ));
 sg13g2_o21ai_1 _1633_ (.B1(_0829_),
    .Y(_0830_),
    .A1(_0778_),
    .A2(_0828_));
 sg13g2_nand2_1 _1634_ (.Y(_0831_),
    .A(_0823_),
    .B(_0830_));
 sg13g2_nand2_1 _1635_ (.Y(_0832_),
    .A(_0775_),
    .B(\DJ8.pc[3] ));
 sg13g2_nand2_1 _1636_ (.Y(_0833_),
    .A(_0831_),
    .B(_0832_));
 sg13g2_buf_2 _1637_ (.A(_0833_),
    .X(_0834_));
 sg13g2_nand2_1 _1638_ (.Y(_0835_),
    .A(_0827_),
    .B(_0834_));
 sg13g2_inv_2 _1639_ (.Y(_0836_),
    .A(_0835_));
 sg13g2_inv_1 _1640_ (.Y(_0837_),
    .A(_0012_));
 sg13g2_inv_1 _1641_ (.Y(_0838_),
    .A(\DJ8.GH[5] ));
 sg13g2_nor2_1 _1642_ (.A(net87),
    .B(_0838_),
    .Y(_0839_));
 sg13g2_a21oi_1 _1643_ (.A1(net87),
    .A2(\DJ8.EF[5] ),
    .Y(_0840_),
    .B1(_0839_));
 sg13g2_nor2_1 _1644_ (.A(_0840_),
    .B(_0775_),
    .Y(_0841_));
 sg13g2_a21oi_2 _1645_ (.B1(_0841_),
    .Y(_0842_),
    .A2(_0775_),
    .A1(_0837_));
 sg13g2_inv_1 _1646_ (.Y(_0843_),
    .A(_0842_));
 sg13g2_buf_1 _1647_ (.A(_0843_),
    .X(_0844_));
 sg13g2_a21oi_1 _1648_ (.A1(_0822_),
    .A2(net39),
    .Y(_0845_),
    .B1(net54));
 sg13g2_inv_1 _1649_ (.Y(_0846_),
    .A(_0845_));
 sg13g2_buf_8 _1650_ (.A(_0801_),
    .X(_0847_));
 sg13g2_nand2_1 _1651_ (.Y(_0848_),
    .A(_0807_),
    .B(_0795_));
 sg13g2_nor2b_1 _1652_ (.A(_0848_),
    .B_N(_0806_),
    .Y(_0849_));
 sg13g2_buf_2 _1653_ (.A(_0849_),
    .X(_0850_));
 sg13g2_nand2_1 _1654_ (.Y(_0851_),
    .A(_0850_),
    .B(_0816_));
 sg13g2_nor2_1 _1655_ (.A(_0834_),
    .B(_0827_),
    .Y(_0852_));
 sg13g2_buf_1 _1656_ (.A(_0852_),
    .X(_0853_));
 sg13g2_nand4_1 _1657_ (.B(net46),
    .C(_0851_),
    .A(_0821_),
    .Y(_0854_),
    .D(net38));
 sg13g2_inv_4 _1658_ (.A(_0827_),
    .Y(_0855_));
 sg13g2_a21oi_1 _1659_ (.A1(_0789_),
    .A2(_0009_),
    .Y(_0856_),
    .B1(net86));
 sg13g2_inv_2 _1660_ (.Y(_0857_),
    .A(_0793_));
 sg13g2_nand2_1 _1661_ (.Y(_0858_),
    .A(_0856_),
    .B(_0857_));
 sg13g2_nand2_2 _1662_ (.Y(_0859_),
    .A(_0858_),
    .B(_0799_));
 sg13g2_nand2_2 _1663_ (.Y(_0860_),
    .A(net71),
    .B(_0819_));
 sg13g2_nand2_1 _1664_ (.Y(_0861_),
    .A(_0859_),
    .B(_0860_));
 sg13g2_nor2_1 _1665_ (.A(_0855_),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_buf_8 _1666_ (.A(_0816_),
    .X(_0863_));
 sg13g2_buf_8 _1667_ (.A(_0834_),
    .X(_0864_));
 sg13g2_nor2_2 _1668_ (.A(net70),
    .B(net45),
    .Y(_0865_));
 sg13g2_nand2_1 _1669_ (.Y(_0866_),
    .A(_0862_),
    .B(_0865_));
 sg13g2_nand2_1 _1670_ (.Y(_0867_),
    .A(_0854_),
    .B(_0866_));
 sg13g2_nor2_1 _1671_ (.A(_0846_),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_buf_8 _1672_ (.A(_0817_),
    .X(_0869_));
 sg13g2_nor2_2 _1673_ (.A(net65),
    .B(_0797_),
    .Y(_0870_));
 sg13g2_buf_1 _1674_ (.A(_0827_),
    .X(_0871_));
 sg13g2_nand4_1 _1675_ (.B(net53),
    .C(net71),
    .A(_0870_),
    .Y(_0872_),
    .D(net45));
 sg13g2_inv_1 _1676_ (.Y(_0873_),
    .A(\DJ8.GH[6] ));
 sg13g2_nor2_1 _1677_ (.A(net87),
    .B(_0873_),
    .Y(_0874_));
 sg13g2_a21oi_1 _1678_ (.A1(net87),
    .A2(\DJ8.EF[6] ),
    .Y(_0875_),
    .B1(_0874_));
 sg13g2_nor2_1 _1679_ (.A(_0875_),
    .B(_0775_),
    .Y(_0876_));
 sg13g2_a21oi_1 _1680_ (.A1(\DJ8.pc[5] ),
    .A2(net74),
    .Y(_0877_),
    .B1(_0876_));
 sg13g2_buf_1 _1681_ (.A(_0877_),
    .X(_0878_));
 sg13g2_inv_1 _1682_ (.Y(_0879_),
    .A(net64));
 sg13g2_a21oi_1 _1683_ (.A1(_0872_),
    .A2(net54),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_nor2b_1 _1684_ (.A(_0868_),
    .B_N(_0880_),
    .Y(_0881_));
 sg13g2_nor2_1 _1685_ (.A(net55),
    .B(_0881_),
    .Y(_0882_));
 sg13g2_nor3_1 _1686_ (.A(_0818_),
    .B(net70),
    .C(_0850_),
    .Y(_0883_));
 sg13g2_nand2_1 _1687_ (.Y(_0884_),
    .A(_0883_),
    .B(_0801_));
 sg13g2_nor3_2 _1688_ (.A(_0793_),
    .B(_0815_),
    .C(_0796_),
    .Y(_0885_));
 sg13g2_nand2_1 _1689_ (.Y(_0886_),
    .A(_0885_),
    .B(net71));
 sg13g2_nand2_1 _1690_ (.Y(_0887_),
    .A(_0884_),
    .B(_0886_));
 sg13g2_nand2_2 _1691_ (.Y(_0888_),
    .A(_0855_),
    .B(_0834_));
 sg13g2_inv_2 _1692_ (.Y(_0889_),
    .A(_0888_));
 sg13g2_nand2_1 _1693_ (.Y(_0890_),
    .A(_0887_),
    .B(_0889_));
 sg13g2_nor2_1 _1694_ (.A(_0834_),
    .B(_0855_),
    .Y(_0891_));
 sg13g2_buf_1 _1695_ (.A(_0891_),
    .X(_0892_));
 sg13g2_nand2_1 _1696_ (.Y(_0893_),
    .A(net37),
    .B(_0885_));
 sg13g2_nor2_1 _1697_ (.A(net65),
    .B(_0850_),
    .Y(_0894_));
 sg13g2_nand2_1 _1698_ (.Y(_0895_),
    .A(_0894_),
    .B(net38));
 sg13g2_nand2_1 _1699_ (.Y(_0896_),
    .A(_0893_),
    .B(_0895_));
 sg13g2_nor2_1 _1700_ (.A(_0842_),
    .B(_0896_),
    .Y(_0897_));
 sg13g2_a21oi_1 _1701_ (.A1(_0890_),
    .A2(_0897_),
    .Y(_0898_),
    .B1(net64));
 sg13g2_nor2_2 _1702_ (.A(net65),
    .B(_0809_),
    .Y(_0899_));
 sg13g2_nor2_1 _1703_ (.A(net53),
    .B(_0899_),
    .Y(_0900_));
 sg13g2_nand2_1 _1704_ (.Y(_0901_),
    .A(_0821_),
    .B(_0834_));
 sg13g2_o21ai_1 _1705_ (.B1(_0842_),
    .Y(_0902_),
    .A1(_0900_),
    .A2(_0901_));
 sg13g2_a21oi_2 _1706_ (.B1(net70),
    .Y(_0903_),
    .A2(_0819_),
    .A1(net71));
 sg13g2_a21oi_1 _1707_ (.A1(net86),
    .A2(\DJ8.pc[1] ),
    .Y(_0904_),
    .B1(_0797_));
 sg13g2_buf_1 _1708_ (.A(_0904_),
    .X(_0905_));
 sg13g2_nand2_1 _1709_ (.Y(_0906_),
    .A(_0903_),
    .B(net52));
 sg13g2_nand2_2 _1710_ (.Y(_0907_),
    .A(net71),
    .B(_0816_));
 sg13g2_nand2_1 _1711_ (.Y(_0908_),
    .A(_0906_),
    .B(_0907_));
 sg13g2_nand3_1 _1712_ (.B(net71),
    .C(net70),
    .A(_0858_),
    .Y(_0909_));
 sg13g2_buf_1 _1713_ (.A(_0909_),
    .X(_0910_));
 sg13g2_buf_8 _1714_ (.A(_0855_),
    .X(_0911_));
 sg13g2_nand2_1 _1715_ (.Y(_0912_),
    .A(_0910_),
    .B(net44));
 sg13g2_inv_2 _1716_ (.Y(_0913_),
    .A(_0834_));
 sg13g2_buf_1 _1717_ (.A(_0913_),
    .X(_0914_));
 sg13g2_nand3_1 _1718_ (.B(_0912_),
    .C(net36),
    .A(_0908_),
    .Y(_0915_));
 sg13g2_nand2b_1 _1719_ (.Y(_0916_),
    .B(_0915_),
    .A_N(_0902_));
 sg13g2_nand2_1 _1720_ (.Y(_0917_),
    .A(_0898_),
    .B(_0916_));
 sg13g2_nand2_1 _1721_ (.Y(_0918_),
    .A(_0882_),
    .B(_0917_));
 sg13g2_nor2_1 _1722_ (.A(_0855_),
    .B(_0859_),
    .Y(_0919_));
 sg13g2_nand2_1 _1723_ (.Y(_0920_),
    .A(_0919_),
    .B(_0903_));
 sg13g2_nand2_1 _1724_ (.Y(_0921_),
    .A(_0920_),
    .B(net45));
 sg13g2_nor2_1 _1725_ (.A(net64),
    .B(net54),
    .Y(_0922_));
 sg13g2_nand2_1 _1726_ (.Y(_0923_),
    .A(_0921_),
    .B(_0922_));
 sg13g2_nor2_1 _1727_ (.A(_0827_),
    .B(_0907_),
    .Y(_0924_));
 sg13g2_nor2_1 _1728_ (.A(net45),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nand2_1 _1729_ (.Y(_0926_),
    .A(_0919_),
    .B(_0899_));
 sg13g2_nand2_1 _1730_ (.Y(_0927_),
    .A(_0925_),
    .B(_0926_));
 sg13g2_nor2b_1 _1731_ (.A(_0923_),
    .B_N(_0927_),
    .Y(_0928_));
 sg13g2_buf_8 _1732_ (.A(_0859_),
    .X(_0929_));
 sg13g2_buf_1 _1733_ (.A(_0860_),
    .X(_0930_));
 sg13g2_nor2_2 _1734_ (.A(net70),
    .B(_0827_),
    .Y(_0931_));
 sg13g2_nand3_1 _1735_ (.B(net50),
    .C(_0931_),
    .A(net51),
    .Y(_0932_));
 sg13g2_nand2_1 _1736_ (.Y(_0933_),
    .A(_0932_),
    .B(net36));
 sg13g2_nand2_2 _1737_ (.Y(_0934_),
    .A(_0827_),
    .B(_0869_));
 sg13g2_inv_2 _1738_ (.Y(_0935_),
    .A(_0934_));
 sg13g2_nand3_1 _1739_ (.B(_0930_),
    .C(_0935_),
    .A(net52),
    .Y(_0936_));
 sg13g2_nor2b_1 _1740_ (.A(_0933_),
    .B_N(_0936_),
    .Y(_0937_));
 sg13g2_nor2_1 _1741_ (.A(net46),
    .B(_0894_),
    .Y(_0938_));
 sg13g2_nand2_2 _1742_ (.Y(_0939_),
    .A(_0860_),
    .B(net65));
 sg13g2_nand2_1 _1743_ (.Y(_0940_),
    .A(_0938_),
    .B(_0939_));
 sg13g2_nand2_1 _1744_ (.Y(_0941_),
    .A(_0940_),
    .B(net45));
 sg13g2_nand2_1 _1745_ (.Y(_0942_),
    .A(_0844_),
    .B(_0879_));
 sg13g2_nor2_1 _1746_ (.A(_0942_),
    .B(_0889_),
    .Y(_0943_));
 sg13g2_nand2_1 _1747_ (.Y(_0944_),
    .A(_0941_),
    .B(_0943_));
 sg13g2_nor2_1 _1748_ (.A(_0937_),
    .B(_0944_),
    .Y(_0945_));
 sg13g2_nor3_1 _1749_ (.A(_0784_),
    .B(_0928_),
    .C(_0945_),
    .Y(_0946_));
 sg13g2_nand2_1 _1750_ (.Y(_0947_),
    .A(_0821_),
    .B(_0851_));
 sg13g2_nor2_1 _1751_ (.A(net51),
    .B(_0947_),
    .Y(_0948_));
 sg13g2_inv_2 _1752_ (.Y(_0949_),
    .A(_0948_));
 sg13g2_nor2_1 _1753_ (.A(_0863_),
    .B(_0801_),
    .Y(_0950_));
 sg13g2_inv_1 _1754_ (.Y(_0951_),
    .A(_0950_));
 sg13g2_nand2_1 _1755_ (.Y(_0952_),
    .A(_0949_),
    .B(_0951_));
 sg13g2_nand2_1 _1756_ (.Y(_0953_),
    .A(_0952_),
    .B(net38));
 sg13g2_inv_1 _1757_ (.Y(_0954_),
    .A(net37));
 sg13g2_nand2_1 _1758_ (.Y(_0955_),
    .A(_0939_),
    .B(net46));
 sg13g2_nand2_1 _1759_ (.Y(_0956_),
    .A(_0821_),
    .B(_0859_));
 sg13g2_nand2_1 _1760_ (.Y(_0957_),
    .A(_0955_),
    .B(_0956_));
 sg13g2_nor2_1 _1761_ (.A(_0954_),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_nand2_1 _1762_ (.Y(_0959_),
    .A(_0801_),
    .B(_0899_));
 sg13g2_nand2_1 _1763_ (.Y(_0960_),
    .A(_0959_),
    .B(_0886_));
 sg13g2_nand2_1 _1764_ (.Y(_0961_),
    .A(_0960_),
    .B(net39));
 sg13g2_nand2_1 _1765_ (.Y(_0962_),
    .A(_0961_),
    .B(net54));
 sg13g2_nor2_1 _1766_ (.A(_0958_),
    .B(_0962_),
    .Y(_0963_));
 sg13g2_nand2_1 _1767_ (.Y(_0964_),
    .A(_0953_),
    .B(_0963_));
 sg13g2_buf_1 _1768_ (.A(_0879_),
    .X(_0965_));
 sg13g2_nand2_1 _1769_ (.Y(_0966_),
    .A(net46),
    .B(_0907_));
 sg13g2_nand2_1 _1770_ (.Y(_0967_),
    .A(_0956_),
    .B(_0966_));
 sg13g2_nor2_1 _1771_ (.A(_0954_),
    .B(_0967_),
    .Y(_0968_));
 sg13g2_a21oi_1 _1772_ (.A1(_0929_),
    .A2(net70),
    .Y(_0969_),
    .B1(net50));
 sg13g2_nand2_1 _1773_ (.Y(_0970_),
    .A(_0969_),
    .B(_0889_));
 sg13g2_inv_1 _1774_ (.Y(_0971_),
    .A(_0815_));
 sg13g2_nand3_1 _1775_ (.B(_0857_),
    .C(_0971_),
    .A(_0856_),
    .Y(_0972_));
 sg13g2_nor2_1 _1776_ (.A(net71),
    .B(_0972_),
    .Y(_0973_));
 sg13g2_a21oi_1 _1777_ (.A1(_0973_),
    .A2(net39),
    .Y(_0974_),
    .B1(net54));
 sg13g2_nand2_1 _1778_ (.Y(_0975_),
    .A(_0970_),
    .B(_0974_));
 sg13g2_nor2_1 _1779_ (.A(_0968_),
    .B(_0975_),
    .Y(_0976_));
 sg13g2_nor2_1 _1780_ (.A(net43),
    .B(_0976_),
    .Y(_0977_));
 sg13g2_nand2_1 _1781_ (.Y(_0978_),
    .A(_0964_),
    .B(_0977_));
 sg13g2_nand2_1 _1782_ (.Y(_0979_),
    .A(_0946_),
    .B(_0978_));
 sg13g2_inv_1 _1783_ (.Y(_0980_),
    .A(\DJ8.GH[15] ));
 sg13g2_nand2_1 _1784_ (.Y(_0981_),
    .A(\DJ8.EF[15] ),
    .B(net84));
 sg13g2_o21ai_1 _1785_ (.B1(_0981_),
    .Y(_0982_),
    .A1(net84),
    .A2(_0980_));
 sg13g2_nor2_1 _1786_ (.A(_0982_),
    .B(net74),
    .Y(_0983_));
 sg13g2_a21oi_1 _1787_ (.A1(_0004_),
    .A2(net74),
    .Y(_0984_),
    .B1(_0983_));
 sg13g2_nand3_1 _1788_ (.B(_0979_),
    .C(_0984_),
    .A(_0918_),
    .Y(_0985_));
 sg13g2_buf_1 _1789_ (.A(_0754_),
    .X(_0986_));
 sg13g2_inv_1 _1790_ (.Y(_0987_),
    .A(\DJ8.ir[1] ));
 sg13g2_nor2_1 _1791_ (.A(_0986_),
    .B(_0987_),
    .Y(_0988_));
 sg13g2_inv_2 _1792_ (.Y(_0989_),
    .A(_0984_));
 sg13g2_nand2_1 _1793_ (.Y(_0990_),
    .A(_0989_),
    .B(net2));
 sg13g2_nand3_1 _1794_ (.B(_0988_),
    .C(_0990_),
    .A(_0985_),
    .Y(_0991_));
 sg13g2_inv_1 _1795_ (.Y(_0992_),
    .A(\DJ8.ir[6] ));
 sg13g2_nand2_1 _1796_ (.Y(_0993_),
    .A(_0754_),
    .B(_0760_));
 sg13g2_o21ai_1 _1797_ (.B1(_0993_),
    .Y(_0994_),
    .A1(_0754_),
    .A2(_0992_));
 sg13g2_inv_2 _1798_ (.Y(_0995_),
    .A(_0761_));
 sg13g2_nor2_1 _1799_ (.A(_0754_),
    .B(\DJ8.ir[5] ),
    .Y(_0996_));
 sg13g2_a21oi_1 _1800_ (.A1(_0754_),
    .A2(_0995_),
    .Y(_0997_),
    .B1(_0996_));
 sg13g2_nor2_1 _1801_ (.A(_0994_),
    .B(_0997_),
    .Y(_0998_));
 sg13g2_inv_1 _1802_ (.Y(_0999_),
    .A(_0001_));
 sg13g2_nor2_1 _1803_ (.A(_0754_),
    .B(_0003_),
    .Y(_1000_));
 sg13g2_a21o_1 _1804_ (.A2(_0999_),
    .A1(_0754_),
    .B1(_1000_),
    .X(_1001_));
 sg13g2_buf_1 _1805_ (.A(_1001_),
    .X(_1002_));
 sg13g2_nand2_1 _1806_ (.Y(_1003_),
    .A(_0998_),
    .B(_1002_));
 sg13g2_inv_2 _1807_ (.Y(_1004_),
    .A(_1003_));
 sg13g2_nor2b_1 _1808_ (.A(_0994_),
    .B_N(_0997_),
    .Y(_1005_));
 sg13g2_nand2_1 _1809_ (.Y(_1006_),
    .A(_1005_),
    .B(_1002_));
 sg13g2_inv_2 _1810_ (.Y(_1007_),
    .A(_1006_));
 sg13g2_inv_1 _1811_ (.Y(_1008_),
    .A(\DJ8.GH[8] ));
 sg13g2_nor2b_1 _1812_ (.A(_0997_),
    .B_N(_0994_),
    .Y(_1009_));
 sg13g2_nand2_2 _1813_ (.Y(_1010_),
    .A(_1009_),
    .B(_1002_));
 sg13g2_nand2_1 _1814_ (.Y(_1011_),
    .A(_0997_),
    .B(_0994_));
 sg13g2_inv_1 _1815_ (.Y(_1012_),
    .A(_1002_));
 sg13g2_nor2_2 _1816_ (.A(_1011_),
    .B(_1012_),
    .Y(_1013_));
 sg13g2_nand2_1 _1817_ (.Y(_1014_),
    .A(_1013_),
    .B(\DJ8.GH[0] ));
 sg13g2_o21ai_1 _1818_ (.B1(_1014_),
    .Y(_1015_),
    .A1(_1008_),
    .A2(_1010_));
 sg13g2_a221oi_1 _1819_ (.B2(_1007_),
    .C1(_1015_),
    .B1(\DJ8.EF[0] ),
    .A1(\DJ8.EF[8] ),
    .Y(_1016_),
    .A2(_1004_));
 sg13g2_nand2_1 _1820_ (.Y(_1017_),
    .A(_1005_),
    .B(_1012_));
 sg13g2_inv_2 _1821_ (.Y(_1018_),
    .A(_1017_));
 sg13g2_nand2_1 _1822_ (.Y(_1019_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][0] ));
 sg13g2_nor2_2 _1823_ (.A(_1002_),
    .B(_1011_),
    .Y(_1020_));
 sg13g2_nand2_1 _1824_ (.Y(_1021_),
    .A(_1009_),
    .B(_1012_));
 sg13g2_inv_2 _1825_ (.Y(_1022_),
    .A(_1021_));
 sg13g2_a22oi_1 _1826_ (.Y(_1023_),
    .B1(\DJ8.REGS.regs[2][0] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][0] ));
 sg13g2_nand2_1 _1827_ (.Y(_1024_),
    .A(_1012_),
    .B(_0998_));
 sg13g2_inv_1 _1828_ (.Y(_1025_),
    .A(_1024_));
 sg13g2_nand2_1 _1829_ (.Y(_1026_),
    .A(net69),
    .B(\DJ8.ACC[0] ));
 sg13g2_nand4_1 _1830_ (.B(_1019_),
    .C(_1023_),
    .A(_1016_),
    .Y(_1027_),
    .D(_1026_));
 sg13g2_nor2_1 _1831_ (.A(_0988_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_inv_1 _1832_ (.Y(_1029_),
    .A(_1028_));
 sg13g2_nand2_1 _1833_ (.Y(_1030_),
    .A(_0752_),
    .B(_0986_));
 sg13g2_o21ai_1 _1834_ (.B1(_1030_),
    .Y(_1031_),
    .A1(net85),
    .A2(_0759_));
 sg13g2_nand3_1 _1835_ (.B(_1029_),
    .C(_1031_),
    .A(_0991_),
    .Y(_1032_));
 sg13g2_inv_4 _1836_ (.A(_1032_),
    .Y(_1033_));
 sg13g2_nor2_1 _1837_ (.A(net85),
    .B(_0015_),
    .Y(_1034_));
 sg13g2_nand2b_1 _1838_ (.Y(_1035_),
    .B(net85),
    .A_N(_0014_));
 sg13g2_nand2b_2 _1839_ (.Y(_1036_),
    .B(_1035_),
    .A_N(_1034_));
 sg13g2_nand2_1 _1840_ (.Y(_1037_),
    .A(_0887_),
    .B(net37));
 sg13g2_nand2_1 _1841_ (.Y(_1038_),
    .A(_0859_),
    .B(_0907_));
 sg13g2_nor2_1 _1842_ (.A(_0888_),
    .B(_0870_),
    .Y(_1039_));
 sg13g2_a22oi_1 _1843_ (.Y(_1040_),
    .B1(_1038_),
    .B2(_1039_),
    .A2(net38),
    .A1(_0863_));
 sg13g2_nand2_1 _1844_ (.Y(_1041_),
    .A(_1037_),
    .B(_1040_));
 sg13g2_buf_1 _1845_ (.A(net54),
    .X(_1042_));
 sg13g2_nand2_1 _1846_ (.Y(_1043_),
    .A(_1041_),
    .B(net42));
 sg13g2_nand2_1 _1847_ (.Y(_1044_),
    .A(_0885_),
    .B(net53));
 sg13g2_nand2_2 _1848_ (.Y(_1045_),
    .A(_0885_),
    .B(_0850_));
 sg13g2_nand2_1 _1849_ (.Y(_1046_),
    .A(_1044_),
    .B(_1045_));
 sg13g2_nor2_2 _1850_ (.A(_0913_),
    .B(_0843_),
    .Y(_1047_));
 sg13g2_a21oi_1 _1851_ (.A1(_1046_),
    .A2(_1047_),
    .Y(_1048_),
    .B1(net64));
 sg13g2_nand2_1 _1852_ (.Y(_1049_),
    .A(_1043_),
    .B(_1048_));
 sg13g2_nand2_1 _1853_ (.Y(_1050_),
    .A(_0910_),
    .B(_1045_));
 sg13g2_buf_1 _1854_ (.A(net44),
    .X(_1051_));
 sg13g2_nand3_1 _1855_ (.B(net35),
    .C(net54),
    .A(_1050_),
    .Y(_1052_));
 sg13g2_nor2_1 _1856_ (.A(_0911_),
    .B(_0910_),
    .Y(_1053_));
 sg13g2_inv_1 _1857_ (.Y(_1054_),
    .A(_1053_));
 sg13g2_nand2_1 _1858_ (.Y(_1055_),
    .A(_1052_),
    .B(_1054_));
 sg13g2_nand2_1 _1859_ (.Y(_1056_),
    .A(_1055_),
    .B(net36));
 sg13g2_o21ai_1 _1860_ (.B1(_0895_),
    .Y(_1057_),
    .A1(_0835_),
    .A2(_1045_));
 sg13g2_buf_1 _1861_ (.A(_0842_),
    .X(_1058_));
 sg13g2_a21oi_1 _1862_ (.A1(_1057_),
    .A2(net63),
    .Y(_1059_),
    .B1(net43));
 sg13g2_nand2_1 _1863_ (.Y(_1060_),
    .A(_1056_),
    .B(_1059_));
 sg13g2_nand2_1 _1864_ (.Y(_1061_),
    .A(_1049_),
    .B(_1060_));
 sg13g2_buf_1 _1865_ (.A(_0784_),
    .X(_1062_));
 sg13g2_a21oi_1 _1866_ (.A1(_1061_),
    .A2(net49),
    .Y(_1063_),
    .B1(_0989_));
 sg13g2_nand3_1 _1867_ (.B(_0799_),
    .C(net65),
    .A(_0858_),
    .Y(_1064_));
 sg13g2_buf_2 _1868_ (.A(_1064_),
    .X(_1065_));
 sg13g2_a21oi_1 _1869_ (.A1(_1045_),
    .A2(_1065_),
    .Y(_1066_),
    .B1(net53));
 sg13g2_buf_1 _1870_ (.A(_0864_),
    .X(_1067_));
 sg13g2_nand2b_1 _1871_ (.Y(_1068_),
    .B(net34),
    .A_N(_1066_));
 sg13g2_inv_1 _1872_ (.Y(_1069_),
    .A(_0886_));
 sg13g2_a21oi_1 _1873_ (.A1(_1069_),
    .A2(net53),
    .Y(_1070_),
    .B1(net34));
 sg13g2_nand2_1 _1874_ (.Y(_1071_),
    .A(_0907_),
    .B(_0855_));
 sg13g2_nor2_2 _1875_ (.A(_0859_),
    .B(_0903_),
    .Y(_1072_));
 sg13g2_nand2b_1 _1876_ (.Y(_1073_),
    .B(_1072_),
    .A_N(_1071_));
 sg13g2_nand2_1 _1877_ (.Y(_1074_),
    .A(_1070_),
    .B(_1073_));
 sg13g2_nand3_1 _1878_ (.B(net63),
    .C(_1074_),
    .A(_1068_),
    .Y(_1075_));
 sg13g2_nor2_1 _1879_ (.A(net36),
    .B(_1052_),
    .Y(_1076_));
 sg13g2_nor2_1 _1880_ (.A(_0834_),
    .B(_0934_),
    .Y(_1077_));
 sg13g2_nand2_1 _1881_ (.Y(_1078_),
    .A(_1077_),
    .B(_0801_));
 sg13g2_inv_1 _1882_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_nor2_1 _1883_ (.A(_1079_),
    .B(_0896_),
    .Y(_1080_));
 sg13g2_inv_1 _1884_ (.Y(_1081_),
    .A(_0870_));
 sg13g2_nand2_1 _1885_ (.Y(_1082_),
    .A(_1045_),
    .B(_1081_));
 sg13g2_nand2_1 _1886_ (.Y(_1083_),
    .A(_1082_),
    .B(net39));
 sg13g2_a21oi_1 _1887_ (.A1(_1080_),
    .A2(_1083_),
    .Y(_1084_),
    .B1(net63));
 sg13g2_nor2_1 _1888_ (.A(_1076_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nand2_1 _1889_ (.Y(_1086_),
    .A(_1075_),
    .B(_1085_));
 sg13g2_nand2_1 _1890_ (.Y(_1087_),
    .A(_1086_),
    .B(net64));
 sg13g2_nor2b_1 _1891_ (.A(_0895_),
    .B_N(_0922_),
    .Y(_1088_));
 sg13g2_nor2_1 _1892_ (.A(net49),
    .B(_1088_),
    .Y(_1089_));
 sg13g2_nand2_1 _1893_ (.Y(_1090_),
    .A(_1087_),
    .B(_1089_));
 sg13g2_nand2_1 _1894_ (.Y(_1091_),
    .A(_1063_),
    .B(_1090_));
 sg13g2_buf_1 _1895_ (.A(_0988_),
    .X(_1092_));
 sg13g2_nand2_1 _1896_ (.Y(_1093_),
    .A(_0989_),
    .B(net3));
 sg13g2_nand3_1 _1897_ (.B(net79),
    .C(_1093_),
    .A(_1091_),
    .Y(_1094_));
 sg13g2_a22oi_1 _1898_ (.Y(_1095_),
    .B1(\DJ8.EF[1] ),
    .B2(_1007_),
    .A2(_1013_),
    .A1(\DJ8.GH[1] ));
 sg13g2_a22oi_1 _1899_ (.Y(_1096_),
    .B1(\DJ8.REGS.regs[2][1] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][1] ));
 sg13g2_inv_1 _1900_ (.Y(_1097_),
    .A(\DJ8.GH[9] ));
 sg13g2_nor2_1 _1901_ (.A(_1097_),
    .B(_1010_),
    .Y(_1098_));
 sg13g2_a21oi_1 _1902_ (.A1(\DJ8.EF[9] ),
    .A2(_1004_),
    .Y(_1099_),
    .B1(_1098_));
 sg13g2_nand2_1 _1903_ (.Y(_1100_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][1] ));
 sg13g2_nand4_1 _1904_ (.B(_1096_),
    .C(_1099_),
    .A(_1095_),
    .Y(_1101_),
    .D(_1100_));
 sg13g2_a21oi_1 _1905_ (.A1(\DJ8.ACC[1] ),
    .A2(net69),
    .Y(_1102_),
    .B1(_1101_));
 sg13g2_inv_1 _1906_ (.Y(_1103_),
    .A(_0988_));
 sg13g2_nand2_1 _1907_ (.Y(_1104_),
    .A(_1102_),
    .B(_1103_));
 sg13g2_nand2_2 _1908_ (.Y(_1105_),
    .A(_1094_),
    .B(_1104_));
 sg13g2_xnor2_1 _1909_ (.Y(_1106_),
    .A(_1036_),
    .B(_1105_));
 sg13g2_xnor2_1 _1910_ (.Y(_1107_),
    .A(_1033_),
    .B(_1106_));
 sg13g2_nand2_1 _1911_ (.Y(_1108_),
    .A(_0991_),
    .B(_1029_));
 sg13g2_inv_1 _1912_ (.Y(_1109_),
    .A(_1031_));
 sg13g2_nand2_1 _1913_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nand3_1 _1914_ (.B(_1032_),
    .C(\DJ8.ALU.c_in ),
    .A(_1110_),
    .Y(_1111_));
 sg13g2_nand2_1 _1915_ (.Y(_1112_),
    .A(_1107_),
    .B(_1111_));
 sg13g2_inv_1 _1916_ (.Y(_1113_),
    .A(_1106_));
 sg13g2_nor2_1 _1917_ (.A(_1111_),
    .B(_1113_),
    .Y(_1114_));
 sg13g2_buf_2 _1918_ (.A(\DJ8.ALU.opalu[1] ),
    .X(_1115_));
 sg13g2_buf_2 _1919_ (.A(\DJ8.ALU.opalu[0] ),
    .X(_1116_));
 sg13g2_inv_2 _1920_ (.Y(_1117_),
    .A(_1116_));
 sg13g2_inv_1 _1921_ (.Y(_1118_),
    .A(_0013_));
 sg13g2_nor3_2 _1922_ (.A(_1115_),
    .B(_1117_),
    .C(_1118_),
    .Y(_1119_));
 sg13g2_nor2b_1 _1923_ (.A(_1114_),
    .B_N(_1119_),
    .Y(_1120_));
 sg13g2_inv_1 _1924_ (.Y(_1121_),
    .A(\DJ8.ALU.opalu[2] ));
 sg13g2_inv_1 _1925_ (.Y(_1122_),
    .A(_1115_));
 sg13g2_nor3_2 _1926_ (.A(_1116_),
    .B(_1121_),
    .C(_1122_),
    .Y(_1123_));
 sg13g2_inv_1 _1927_ (.Y(_1124_),
    .A(_1036_));
 sg13g2_nor2_1 _1928_ (.A(_1124_),
    .B(_1105_),
    .Y(_1125_));
 sg13g2_nand2_2 _1929_ (.Y(_1126_),
    .A(_1115_),
    .B(_1116_));
 sg13g2_nor2_2 _1930_ (.A(_1118_),
    .B(_1126_),
    .Y(_1127_));
 sg13g2_inv_1 _1931_ (.Y(_1128_),
    .A(_1127_));
 sg13g2_nor2_2 _1932_ (.A(_0013_),
    .B(_1126_),
    .Y(_1129_));
 sg13g2_inv_1 _1933_ (.Y(_1130_),
    .A(_1126_));
 sg13g2_a21oi_1 _1934_ (.A1(_1122_),
    .A2(_1117_),
    .Y(_1131_),
    .B1(_1118_));
 sg13g2_nor3_2 _1935_ (.A(\DJ8.ALU.opalu[2] ),
    .B(_1130_),
    .C(_1131_),
    .Y(_1132_));
 sg13g2_a21oi_1 _1936_ (.A1(_1129_),
    .A2(_1036_),
    .Y(_1133_),
    .B1(_1132_));
 sg13g2_o21ai_1 _1937_ (.B1(_1133_),
    .Y(_1134_),
    .A1(_1128_),
    .A2(_1105_));
 sg13g2_a21oi_1 _1938_ (.A1(_1123_),
    .A2(_1125_),
    .Y(_1135_),
    .B1(_1134_));
 sg13g2_nor3_2 _1939_ (.A(_1115_),
    .B(_1116_),
    .C(_1121_),
    .Y(_1136_));
 sg13g2_nand2_1 _1940_ (.Y(_1137_),
    .A(_1106_),
    .B(_1136_));
 sg13g2_nand2_1 _1941_ (.Y(_1138_),
    .A(_1105_),
    .B(_1124_));
 sg13g2_nor3_2 _1942_ (.A(_1115_),
    .B(_1121_),
    .C(_1117_),
    .Y(_1139_));
 sg13g2_nand2_1 _1943_ (.Y(_1140_),
    .A(_1138_),
    .B(_1139_));
 sg13g2_nand3_1 _1944_ (.B(_1137_),
    .C(_1140_),
    .A(_1135_),
    .Y(_1141_));
 sg13g2_a21oi_1 _1945_ (.A1(_1112_),
    .A2(_1120_),
    .Y(_1142_),
    .B1(_1141_));
 sg13g2_inv_1 _1946_ (.Y(_1143_),
    .A(\DJ8.ALU.c_in ));
 sg13g2_xnor2_1 _1947_ (.Y(_1144_),
    .A(_1143_),
    .B(_1031_));
 sg13g2_nand3_1 _1948_ (.B(_1029_),
    .C(_1144_),
    .A(_0991_),
    .Y(_1145_));
 sg13g2_nand2_1 _1949_ (.Y(_1146_),
    .A(_1109_),
    .B(_1143_));
 sg13g2_a21oi_1 _1950_ (.A1(_1145_),
    .A2(_1146_),
    .Y(_1147_),
    .B1(_1036_));
 sg13g2_inv_1 _1951_ (.Y(_1148_),
    .A(_1147_));
 sg13g2_nand3_1 _1952_ (.B(_1036_),
    .C(_1146_),
    .A(_1145_),
    .Y(_1149_));
 sg13g2_inv_1 _1953_ (.Y(_1150_),
    .A(_1105_));
 sg13g2_a21oi_1 _1954_ (.A1(_1148_),
    .A2(_1149_),
    .Y(_1151_),
    .B1(_1150_));
 sg13g2_nor3_2 _1955_ (.A(_1116_),
    .B(_1122_),
    .C(_1118_),
    .Y(_1152_));
 sg13g2_nand3_1 _1956_ (.B(_1149_),
    .C(_1150_),
    .A(_1148_),
    .Y(_1153_));
 sg13g2_nand3b_1 _1957_ (.B(_1152_),
    .C(_1153_),
    .Y(_1154_),
    .A_N(_1151_));
 sg13g2_nand2_1 _1958_ (.Y(_1155_),
    .A(_1142_),
    .B(_1154_));
 sg13g2_buf_1 _1959_ (.A(net85),
    .X(_1156_));
 sg13g2_inv_1 _1960_ (.Y(_1157_),
    .A(\DJ8.ir[2] ));
 sg13g2_nor3_1 _1961_ (.A(net83),
    .B(\DJ8.ir[3] ),
    .C(_1157_),
    .Y(_1158_));
 sg13g2_inv_1 _1962_ (.Y(_1159_),
    .A(\DJ8.ir[3] ));
 sg13g2_nor3_1 _1963_ (.A(net83),
    .B(\DJ8.ir[2] ),
    .C(_1159_),
    .Y(_1160_));
 sg13g2_nor2_2 _1964_ (.A(_1158_),
    .B(_1160_),
    .Y(_1161_));
 sg13g2_inv_2 _1965_ (.Y(_1162_),
    .A(_1161_));
 sg13g2_buf_1 _1966_ (.A(_1132_),
    .X(_1163_));
 sg13g2_nand2_1 _1967_ (.Y(_1164_),
    .A(_1107_),
    .B(net75));
 sg13g2_nand3_1 _1968_ (.B(_1162_),
    .C(_1164_),
    .A(_1155_),
    .Y(_1165_));
 sg13g2_inv_1 _1969_ (.Y(_1166_),
    .A(_1144_));
 sg13g2_nand3_1 _1970_ (.B(_1126_),
    .C(_1131_),
    .A(_1145_),
    .Y(_1167_));
 sg13g2_a21oi_1 _1971_ (.A1(_1108_),
    .A2(_1166_),
    .Y(_1168_),
    .B1(_1167_));
 sg13g2_a221oi_1 _1972_ (.B2(_1110_),
    .C1(_1168_),
    .B1(_1139_),
    .A1(_1129_),
    .Y(_1169_),
    .A2(_1031_));
 sg13g2_nor2b_1 _1973_ (.A(_1032_),
    .B_N(_1123_),
    .Y(_1170_));
 sg13g2_nor2_1 _1974_ (.A(_1128_),
    .B(_1108_),
    .Y(_1171_));
 sg13g2_nand2_1 _1975_ (.Y(_1172_),
    .A(_1110_),
    .B(_1032_));
 sg13g2_nor2b_1 _1976_ (.A(_1172_),
    .B_N(_1136_),
    .Y(_1173_));
 sg13g2_nor4_1 _1977_ (.A(_1132_),
    .B(_1170_),
    .C(_1171_),
    .D(_1173_),
    .Y(_1174_));
 sg13g2_nand2_1 _1978_ (.Y(_1175_),
    .A(_1169_),
    .B(_1174_));
 sg13g2_nand2_1 _1979_ (.Y(_1176_),
    .A(_1172_),
    .B(_1163_));
 sg13g2_nand3_1 _1980_ (.B(_1161_),
    .C(_1176_),
    .A(_1175_),
    .Y(_1177_));
 sg13g2_nand2_2 _1981_ (.Y(_1178_),
    .A(_1165_),
    .B(_1177_));
 sg13g2_nand2_1 _1982_ (.Y(_1179_),
    .A(_1178_),
    .B(_0768_));
 sg13g2_o21ai_1 _1983_ (.B1(_1179_),
    .Y(_0038_),
    .A1(_0759_),
    .A2(net66));
 sg13g2_a21oi_1 _1984_ (.A1(net52),
    .A2(net65),
    .Y(_1180_),
    .B1(_1071_));
 sg13g2_nor2_1 _1985_ (.A(net36),
    .B(_1180_),
    .Y(_1181_));
 sg13g2_nand2_1 _1986_ (.Y(_1182_),
    .A(_0956_),
    .B(_1065_));
 sg13g2_nand2_1 _1987_ (.Y(_1183_),
    .A(_1182_),
    .B(net53));
 sg13g2_nand2_1 _1988_ (.Y(_1184_),
    .A(_1181_),
    .B(_1183_));
 sg13g2_a21oi_1 _1989_ (.A1(_0907_),
    .A2(net44),
    .Y(_1185_),
    .B1(net54));
 sg13g2_nand2_1 _1990_ (.Y(_1186_),
    .A(_0948_),
    .B(_1185_));
 sg13g2_inv_1 _1991_ (.Y(_1187_),
    .A(_1047_));
 sg13g2_nand2_1 _1992_ (.Y(_1188_),
    .A(_1186_),
    .B(_1187_));
 sg13g2_nand2_1 _1993_ (.Y(_1189_),
    .A(_1184_),
    .B(_1188_));
 sg13g2_nand2_1 _1994_ (.Y(_1190_),
    .A(_1065_),
    .B(net38));
 sg13g2_nand2_1 _1995_ (.Y(_1191_),
    .A(_1190_),
    .B(_1078_));
 sg13g2_nor2_2 _1996_ (.A(_0818_),
    .B(_0850_),
    .Y(_1192_));
 sg13g2_nand2_1 _1997_ (.Y(_1193_),
    .A(_1191_),
    .B(_1192_));
 sg13g2_nand3_1 _1998_ (.B(net51),
    .C(net45),
    .A(_0924_),
    .Y(_1194_));
 sg13g2_nand2_1 _1999_ (.Y(_1195_),
    .A(_1193_),
    .B(_1194_));
 sg13g2_nand2_1 _2000_ (.Y(_1196_),
    .A(_1195_),
    .B(net42));
 sg13g2_a21oi_1 _2001_ (.A1(_1189_),
    .A2(_1196_),
    .Y(_1197_),
    .B1(net64));
 sg13g2_a21oi_1 _2002_ (.A1(_0861_),
    .A2(net65),
    .Y(_1198_),
    .B1(_0954_));
 sg13g2_nand2_1 _2003_ (.Y(_1199_),
    .A(_1038_),
    .B(net38));
 sg13g2_nor2_1 _2004_ (.A(_1199_),
    .B(_1072_),
    .Y(_1200_));
 sg13g2_nor2_1 _2005_ (.A(_1198_),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_nand2_1 _2006_ (.Y(_1202_),
    .A(_1201_),
    .B(_0845_));
 sg13g2_nand2_1 _2007_ (.Y(_1203_),
    .A(_0822_),
    .B(net38));
 sg13g2_a21oi_1 _2008_ (.A1(_0889_),
    .A2(_0870_),
    .Y(_1204_),
    .B1(_0842_));
 sg13g2_nand3_1 _2009_ (.B(_0893_),
    .C(_1204_),
    .A(_1203_),
    .Y(_1205_));
 sg13g2_nand3_1 _2010_ (.B(net64),
    .C(_1205_),
    .A(_1202_),
    .Y(_1206_));
 sg13g2_nand2_1 _2011_ (.Y(_1207_),
    .A(_1206_),
    .B(_0784_));
 sg13g2_nor2_1 _2012_ (.A(_1197_),
    .B(_1207_),
    .Y(_1208_));
 sg13g2_nor2_1 _2013_ (.A(_0989_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_buf_8 _2014_ (.A(_0847_),
    .X(_1210_));
 sg13g2_nor2_1 _2015_ (.A(net33),
    .B(_0901_),
    .Y(_1211_));
 sg13g2_nand2_1 _2016_ (.Y(_1212_),
    .A(_0939_),
    .B(net51));
 sg13g2_nand2_1 _2017_ (.Y(_1213_),
    .A(_0907_),
    .B(_0913_));
 sg13g2_nor2_1 _2018_ (.A(_0859_),
    .B(_0899_),
    .Y(_1214_));
 sg13g2_nor3_1 _2019_ (.A(net53),
    .B(_0842_),
    .C(_1214_),
    .Y(_1215_));
 sg13g2_o21ai_1 _2020_ (.B1(_1215_),
    .Y(_1216_),
    .A1(_1212_),
    .A2(_1213_));
 sg13g2_nor2_1 _2021_ (.A(_1211_),
    .B(_1216_),
    .Y(_1217_));
 sg13g2_nor2_1 _2022_ (.A(_0879_),
    .B(_1217_),
    .Y(_1218_));
 sg13g2_nor2_1 _2023_ (.A(net44),
    .B(_1045_),
    .Y(_1219_));
 sg13g2_nand2_1 _2024_ (.Y(_1220_),
    .A(net46),
    .B(_0935_));
 sg13g2_nor2_1 _2025_ (.A(_1192_),
    .B(_1220_),
    .Y(_1221_));
 sg13g2_nor3_1 _2026_ (.A(net45),
    .B(_1219_),
    .C(_1221_),
    .Y(_1222_));
 sg13g2_nand2_1 _2027_ (.Y(_1223_),
    .A(_0884_),
    .B(_1045_));
 sg13g2_nand2_1 _2028_ (.Y(_1224_),
    .A(_1223_),
    .B(net44));
 sg13g2_nand2_1 _2029_ (.Y(_1225_),
    .A(_1222_),
    .B(_1224_));
 sg13g2_nor2_1 _2030_ (.A(net44),
    .B(_0950_),
    .Y(_1226_));
 sg13g2_nand2_1 _2031_ (.Y(_1227_),
    .A(_1226_),
    .B(_0955_));
 sg13g2_nand2_1 _2032_ (.Y(_1228_),
    .A(_0973_),
    .B(_0911_));
 sg13g2_nand3_1 _2033_ (.B(net45),
    .C(_1228_),
    .A(_1227_),
    .Y(_1229_));
 sg13g2_nand3_1 _2034_ (.B(_1229_),
    .C(net63),
    .A(_1225_),
    .Y(_1230_));
 sg13g2_nand2_1 _2035_ (.Y(_1231_),
    .A(_1218_),
    .B(_1230_));
 sg13g2_inv_1 _2036_ (.Y(_1232_),
    .A(net52));
 sg13g2_o21ai_1 _2037_ (.B1(_0888_),
    .Y(_1233_),
    .A1(_1232_),
    .A2(_0901_));
 sg13g2_nand2_1 _2038_ (.Y(_1234_),
    .A(_0847_),
    .B(_0860_));
 sg13g2_nand2_1 _2039_ (.Y(_1235_),
    .A(_1234_),
    .B(_0931_));
 sg13g2_nand2_1 _2040_ (.Y(_1236_),
    .A(_1233_),
    .B(_1235_));
 sg13g2_nor2_1 _2041_ (.A(_0950_),
    .B(_1214_),
    .Y(_1237_));
 sg13g2_a21oi_1 _2042_ (.A1(_1237_),
    .A2(net37),
    .Y(_1238_),
    .B1(_0844_));
 sg13g2_nand2_1 _2043_ (.Y(_1239_),
    .A(_1236_),
    .B(_1238_));
 sg13g2_nor2_1 _2044_ (.A(_0899_),
    .B(net46),
    .Y(_1240_));
 sg13g2_nand2_1 _2045_ (.Y(_1241_),
    .A(net46),
    .B(net44));
 sg13g2_nor2_1 _2046_ (.A(_0864_),
    .B(_0939_),
    .Y(_1242_));
 sg13g2_a22oi_1 _2047_ (.Y(_1243_),
    .B1(_1241_),
    .B2(_1242_),
    .A2(_1240_),
    .A1(net39));
 sg13g2_nand2_1 _2048_ (.Y(_1244_),
    .A(_1243_),
    .B(net42));
 sg13g2_nand2_1 _2049_ (.Y(_1245_),
    .A(_1239_),
    .B(_1244_));
 sg13g2_nand2_1 _2050_ (.Y(_1246_),
    .A(_1245_),
    .B(net43));
 sg13g2_nand2_1 _2051_ (.Y(_1247_),
    .A(_1231_),
    .B(_1246_));
 sg13g2_nand2_1 _2052_ (.Y(_1248_),
    .A(_1247_),
    .B(net55));
 sg13g2_nand2_1 _2053_ (.Y(_1249_),
    .A(_1209_),
    .B(_1248_));
 sg13g2_nand2_1 _2054_ (.Y(_1250_),
    .A(_0989_),
    .B(net4));
 sg13g2_nand3_1 _2055_ (.B(net79),
    .C(_1250_),
    .A(_1249_),
    .Y(_1251_));
 sg13g2_inv_1 _2056_ (.Y(_1252_),
    .A(\DJ8.EF[10] ));
 sg13g2_nor2_1 _2057_ (.A(_1252_),
    .B(_1003_),
    .Y(_1253_));
 sg13g2_inv_1 _2058_ (.Y(_1254_),
    .A(\DJ8.GH[10] ));
 sg13g2_nor2_1 _2059_ (.A(_1254_),
    .B(_1010_),
    .Y(_1255_));
 sg13g2_inv_1 _2060_ (.Y(_1256_),
    .A(\DJ8.EF[2] ));
 sg13g2_nor2_1 _2061_ (.A(_1256_),
    .B(_1006_),
    .Y(_1257_));
 sg13g2_inv_1 _2062_ (.Y(_1258_),
    .A(\DJ8.GH[2] ));
 sg13g2_inv_1 _2063_ (.Y(_1259_),
    .A(_1013_));
 sg13g2_nor2_1 _2064_ (.A(_1258_),
    .B(_1259_),
    .Y(_1260_));
 sg13g2_nor4_1 _2065_ (.A(_1253_),
    .B(_1255_),
    .C(_1257_),
    .D(_1260_),
    .Y(_1261_));
 sg13g2_nand2_1 _2066_ (.Y(_1262_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][2] ));
 sg13g2_a22oi_1 _2067_ (.Y(_1263_),
    .B1(\DJ8.REGS.regs[2][2] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][2] ));
 sg13g2_nand2_1 _2068_ (.Y(_1264_),
    .A(net69),
    .B(\DJ8.ACC[2] ));
 sg13g2_nand4_1 _2069_ (.B(_1262_),
    .C(_1263_),
    .A(_1261_),
    .Y(_1265_),
    .D(_1264_));
 sg13g2_nand2b_1 _2070_ (.Y(_1266_),
    .B(_1103_),
    .A_N(_1265_));
 sg13g2_nand2_1 _2071_ (.Y(_1267_),
    .A(_1251_),
    .B(_1266_));
 sg13g2_nor2_1 _2072_ (.A(net85),
    .B(_0017_),
    .Y(_1268_));
 sg13g2_nand2b_1 _2073_ (.Y(_1269_),
    .B(net85),
    .A_N(_0016_));
 sg13g2_nand2b_1 _2074_ (.Y(_1270_),
    .B(_1269_),
    .A_N(_1268_));
 sg13g2_inv_1 _2075_ (.Y(_1271_),
    .A(_1270_));
 sg13g2_nand2_1 _2076_ (.Y(_1272_),
    .A(_1267_),
    .B(_1271_));
 sg13g2_nand3_1 _2077_ (.B(_1266_),
    .C(_1270_),
    .A(_1251_),
    .Y(_1273_));
 sg13g2_nand2_2 _2078_ (.Y(_1274_),
    .A(_1272_),
    .B(_1273_));
 sg13g2_a21oi_2 _2079_ (.B1(_1147_),
    .Y(_1275_),
    .A2(_1150_),
    .A1(_1149_));
 sg13g2_xnor2_1 _2080_ (.Y(_1276_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_nand2_1 _2081_ (.Y(_1277_),
    .A(_1267_),
    .B(_1270_));
 sg13g2_nand3_1 _2082_ (.B(_1266_),
    .C(_1271_),
    .A(_1251_),
    .Y(_1278_));
 sg13g2_nand2_1 _2083_ (.Y(_1279_),
    .A(_1277_),
    .B(_1278_));
 sg13g2_nand2_1 _2084_ (.Y(_1280_),
    .A(_1279_),
    .B(_1136_));
 sg13g2_nor2_1 _2085_ (.A(_1271_),
    .B(_1267_),
    .Y(_1281_));
 sg13g2_nand2_1 _2086_ (.Y(_1282_),
    .A(_1281_),
    .B(_1123_));
 sg13g2_nand2_1 _2087_ (.Y(_1283_),
    .A(_1272_),
    .B(_1139_));
 sg13g2_inv_1 _2088_ (.Y(_1284_),
    .A(_1129_));
 sg13g2_inv_1 _2089_ (.Y(_1285_),
    .A(_1132_));
 sg13g2_o21ai_1 _2090_ (.B1(_1285_),
    .Y(_1286_),
    .A1(_1284_),
    .A2(_1271_));
 sg13g2_nor2_1 _2091_ (.A(_1128_),
    .B(_1267_),
    .Y(_1287_));
 sg13g2_nor2_1 _2092_ (.A(_1286_),
    .B(_1287_),
    .Y(_1288_));
 sg13g2_nand4_1 _2093_ (.B(_1282_),
    .C(_1283_),
    .A(_1280_),
    .Y(_1289_),
    .D(_1288_));
 sg13g2_a21oi_1 _2094_ (.A1(_1276_),
    .A2(_1152_),
    .Y(_1290_),
    .B1(_1289_));
 sg13g2_a21oi_1 _2095_ (.A1(_1138_),
    .A2(_1033_),
    .Y(_1291_),
    .B1(_1125_));
 sg13g2_inv_1 _2096_ (.Y(_1292_),
    .A(_1291_));
 sg13g2_nand2_1 _2097_ (.Y(_1293_),
    .A(_1292_),
    .B(_1279_));
 sg13g2_nand2_1 _2098_ (.Y(_1294_),
    .A(_1291_),
    .B(_1274_));
 sg13g2_nand2_1 _2099_ (.Y(_1295_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_inv_1 _2100_ (.Y(_1296_),
    .A(_1114_));
 sg13g2_nand2_1 _2101_ (.Y(_1297_),
    .A(_1295_),
    .B(_1296_));
 sg13g2_nand3_1 _2102_ (.B(_1114_),
    .C(_1294_),
    .A(_1293_),
    .Y(_1298_));
 sg13g2_nand3_1 _2103_ (.B(_1298_),
    .C(_1119_),
    .A(_1297_),
    .Y(_1299_));
 sg13g2_nand2_1 _2104_ (.Y(_1300_),
    .A(_1290_),
    .B(_1299_));
 sg13g2_nand2_1 _2105_ (.Y(_1301_),
    .A(_1295_),
    .B(net75));
 sg13g2_nand3_1 _2106_ (.B(_1162_),
    .C(_1301_),
    .A(_1300_),
    .Y(_1302_));
 sg13g2_nand3_1 _2107_ (.B(_1161_),
    .C(_1164_),
    .A(_1155_),
    .Y(_1303_));
 sg13g2_nand2_1 _2108_ (.Y(_1304_),
    .A(_1302_),
    .B(_1303_));
 sg13g2_inv_2 _2109_ (.Y(_1305_),
    .A(_1304_));
 sg13g2_nor2_1 _2110_ (.A(\DJ8.ACC[1] ),
    .B(_0769_),
    .Y(_1306_));
 sg13g2_a21oi_1 _2111_ (.A1(_1305_),
    .A2(_0769_),
    .Y(_0039_),
    .B1(_1306_));
 sg13g2_nand3_1 _2112_ (.B(_1106_),
    .C(_1033_),
    .A(_1279_),
    .Y(_1307_));
 sg13g2_a21oi_2 _2113_ (.B1(_1281_),
    .Y(_1308_),
    .A2(_1125_),
    .A1(_1272_));
 sg13g2_nand2_1 _2114_ (.Y(_1309_),
    .A(_1307_),
    .B(_1308_));
 sg13g2_nor2_1 _2115_ (.A(net85),
    .B(_0019_),
    .Y(_1310_));
 sg13g2_nand2b_1 _2116_ (.Y(_1311_),
    .B(net85),
    .A_N(_0018_));
 sg13g2_nand2b_1 _2117_ (.Y(_1312_),
    .B(_1311_),
    .A_N(_1310_));
 sg13g2_nand2_1 _2118_ (.Y(_1313_),
    .A(_1192_),
    .B(net46));
 sg13g2_nand2_1 _2119_ (.Y(_1314_),
    .A(_1313_),
    .B(_0886_));
 sg13g2_a21oi_1 _2120_ (.A1(_1314_),
    .A2(_0853_),
    .Y(_1315_),
    .B1(_1079_));
 sg13g2_nor2_1 _2121_ (.A(_0888_),
    .B(_1065_),
    .Y(_1316_));
 sg13g2_a21oi_1 _2122_ (.A1(_1316_),
    .A2(net50),
    .Y(_1317_),
    .B1(net63));
 sg13g2_nand2_1 _2123_ (.Y(_1318_),
    .A(_1315_),
    .B(_1317_));
 sg13g2_o21ai_1 _2124_ (.B1(net34),
    .Y(_1319_),
    .A1(_0871_),
    .A2(_0907_));
 sg13g2_a21oi_1 _2125_ (.A1(_1313_),
    .A2(_0865_),
    .Y(_1320_),
    .B1(net42));
 sg13g2_o21ai_1 _2126_ (.B1(_1320_),
    .Y(_1321_),
    .A1(_1212_),
    .A2(_1319_));
 sg13g2_nand2_1 _2127_ (.Y(_1322_),
    .A(_1318_),
    .B(_1321_));
 sg13g2_nand2_1 _2128_ (.Y(_1323_),
    .A(_1322_),
    .B(net49));
 sg13g2_a21oi_1 _2129_ (.A1(net33),
    .A2(net50),
    .Y(_1324_),
    .B1(_0934_));
 sg13g2_nand3_1 _2130_ (.B(_0930_),
    .C(_0931_),
    .A(net52),
    .Y(_1325_));
 sg13g2_nand2_1 _2131_ (.Y(_1326_),
    .A(_1325_),
    .B(net63));
 sg13g2_nor2_1 _2132_ (.A(_0842_),
    .B(_0935_),
    .Y(_1327_));
 sg13g2_buf_1 _2133_ (.A(net34),
    .X(_1328_));
 sg13g2_a21oi_1 _2134_ (.A1(_0932_),
    .A2(_1327_),
    .Y(_1329_),
    .B1(_1328_));
 sg13g2_o21ai_1 _2135_ (.B1(_1329_),
    .Y(_1330_),
    .A1(_1324_),
    .A2(_1326_));
 sg13g2_nor2_1 _2136_ (.A(net70),
    .B(_0913_),
    .Y(_1331_));
 sg13g2_nor2b_1 _2137_ (.A(_0862_),
    .B_N(_1331_),
    .Y(_1332_));
 sg13g2_nor2_1 _2138_ (.A(net49),
    .B(_1332_),
    .Y(_1333_));
 sg13g2_nand2_1 _2139_ (.Y(_1334_),
    .A(_1330_),
    .B(_1333_));
 sg13g2_nand2_1 _2140_ (.Y(_1335_),
    .A(_1323_),
    .B(_1334_));
 sg13g2_a21oi_1 _2141_ (.A1(_1335_),
    .A2(net43),
    .Y(_1336_),
    .B1(_0989_));
 sg13g2_nand2_1 _2142_ (.Y(_1337_),
    .A(_0935_),
    .B(net51));
 sg13g2_inv_1 _2143_ (.Y(_1338_),
    .A(_1337_));
 sg13g2_nor3_1 _2144_ (.A(net34),
    .B(_1338_),
    .C(_1053_),
    .Y(_1339_));
 sg13g2_nand2_1 _2145_ (.Y(_1340_),
    .A(_0903_),
    .B(_0929_));
 sg13g2_nand2_1 _2146_ (.Y(_1341_),
    .A(_1340_),
    .B(_0910_));
 sg13g2_nand2_1 _2147_ (.Y(_1342_),
    .A(_1341_),
    .B(net35));
 sg13g2_nand2_1 _2148_ (.Y(_1343_),
    .A(_1339_),
    .B(_1342_));
 sg13g2_nand2_1 _2149_ (.Y(_1344_),
    .A(_1192_),
    .B(net51));
 sg13g2_a21oi_1 _2150_ (.A1(_1344_),
    .A2(_0931_),
    .Y(_1345_),
    .B1(net36));
 sg13g2_nand2_1 _2151_ (.Y(_1346_),
    .A(_1345_),
    .B(_0936_));
 sg13g2_nand2_1 _2152_ (.Y(_1347_),
    .A(_1343_),
    .B(_1346_));
 sg13g2_buf_1 _2153_ (.A(net42),
    .X(_1348_));
 sg13g2_nand2_1 _2154_ (.Y(_1349_),
    .A(_1347_),
    .B(net32));
 sg13g2_nor2_1 _2155_ (.A(net50),
    .B(net51),
    .Y(_1350_));
 sg13g2_nand3_1 _2156_ (.B(_1067_),
    .C(_0931_),
    .A(_1350_),
    .Y(_1351_));
 sg13g2_nand2_1 _2157_ (.Y(_1352_),
    .A(_1351_),
    .B(_1058_));
 sg13g2_nor3_1 _2158_ (.A(_1242_),
    .B(_1338_),
    .C(_1352_),
    .Y(_1353_));
 sg13g2_nor2_1 _2159_ (.A(net55),
    .B(_1353_),
    .Y(_1354_));
 sg13g2_nand2_1 _2160_ (.Y(_1355_),
    .A(_1349_),
    .B(_1354_));
 sg13g2_a21oi_1 _2161_ (.A1(net33),
    .A2(_0865_),
    .Y(_1356_),
    .B1(_0892_));
 sg13g2_a21oi_1 _2162_ (.A1(_0940_),
    .A2(_1065_),
    .Y(_1357_),
    .B1(_1356_));
 sg13g2_nor2_1 _2163_ (.A(_0888_),
    .B(_0957_),
    .Y(_1358_));
 sg13g2_nor2_1 _2164_ (.A(net42),
    .B(_1358_),
    .Y(_1359_));
 sg13g2_nand2b_1 _2165_ (.Y(_1360_),
    .B(_1359_),
    .A_N(_1357_));
 sg13g2_a21oi_1 _2166_ (.A1(net33),
    .A2(_0869_),
    .Y(_1361_),
    .B1(_0888_));
 sg13g2_nor2_1 _2167_ (.A(_0842_),
    .B(_1077_),
    .Y(_1362_));
 sg13g2_inv_1 _2168_ (.Y(_1363_),
    .A(_1362_));
 sg13g2_a21oi_1 _2169_ (.A1(_1361_),
    .A2(_1212_),
    .Y(_1364_),
    .B1(_1363_));
 sg13g2_buf_1 _2170_ (.A(net36),
    .X(_1365_));
 sg13g2_nand2_1 _2171_ (.Y(_1366_),
    .A(_1066_),
    .B(net30));
 sg13g2_nand2_1 _2172_ (.Y(_1367_),
    .A(_1341_),
    .B(_0836_));
 sg13g2_nand3_1 _2173_ (.B(_1366_),
    .C(_1367_),
    .A(_1364_),
    .Y(_1368_));
 sg13g2_nand3_1 _2174_ (.B(_1368_),
    .C(net55),
    .A(_1360_),
    .Y(_1369_));
 sg13g2_buf_1 _2175_ (.A(net64),
    .X(_1370_));
 sg13g2_nand3_1 _2176_ (.B(_1369_),
    .C(net48),
    .A(_1355_),
    .Y(_1371_));
 sg13g2_nand2_1 _2177_ (.Y(_1372_),
    .A(_1336_),
    .B(_1371_));
 sg13g2_buf_1 _2178_ (.A(_0989_),
    .X(_1373_));
 sg13g2_nand2_1 _2179_ (.Y(_1374_),
    .A(net41),
    .B(net5));
 sg13g2_nand3_1 _2180_ (.B(net79),
    .C(_1374_),
    .A(_1372_),
    .Y(_1375_));
 sg13g2_inv_1 _2181_ (.Y(_1376_),
    .A(\DJ8.GH[11] ));
 sg13g2_nand2_1 _2182_ (.Y(_1377_),
    .A(_1013_),
    .B(\DJ8.GH[3] ));
 sg13g2_o21ai_1 _2183_ (.B1(_1377_),
    .Y(_1378_),
    .A1(_1376_),
    .A2(_1010_));
 sg13g2_a221oi_1 _2184_ (.B2(_1007_),
    .C1(_1378_),
    .B1(\DJ8.EF[3] ),
    .A1(\DJ8.EF[11] ),
    .Y(_1379_),
    .A2(_1004_));
 sg13g2_nand2_1 _2185_ (.Y(_1380_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][3] ));
 sg13g2_a22oi_1 _2186_ (.Y(_1381_),
    .B1(\DJ8.REGS.regs[2][3] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][3] ));
 sg13g2_nand2_1 _2187_ (.Y(_1382_),
    .A(net69),
    .B(\DJ8.ACC[3] ));
 sg13g2_nand4_1 _2188_ (.B(_1380_),
    .C(_1381_),
    .A(_1379_),
    .Y(_1383_),
    .D(_1382_));
 sg13g2_nand2b_1 _2189_ (.Y(_1384_),
    .B(_1103_),
    .A_N(_1383_));
 sg13g2_nand2_1 _2190_ (.Y(_1385_),
    .A(_1375_),
    .B(_1384_));
 sg13g2_xnor2_1 _2191_ (.Y(_1386_),
    .A(_1312_),
    .B(_1385_));
 sg13g2_nand2_1 _2192_ (.Y(_1387_),
    .A(_1309_),
    .B(_1386_));
 sg13g2_inv_1 _2193_ (.Y(_1388_),
    .A(_1312_));
 sg13g2_nand2_1 _2194_ (.Y(_1389_),
    .A(_1385_),
    .B(_1388_));
 sg13g2_nand3_1 _2195_ (.B(_1312_),
    .C(_1384_),
    .A(_1375_),
    .Y(_1390_));
 sg13g2_nand2_2 _2196_ (.Y(_1391_),
    .A(_1389_),
    .B(_1390_));
 sg13g2_nand3_1 _2197_ (.B(_1391_),
    .C(_1308_),
    .A(_1307_),
    .Y(_1392_));
 sg13g2_nand2_1 _2198_ (.Y(_1393_),
    .A(_1387_),
    .B(_1392_));
 sg13g2_nand2_1 _2199_ (.Y(_1394_),
    .A(_1393_),
    .B(_1298_));
 sg13g2_nand2_1 _2200_ (.Y(_1395_),
    .A(_1309_),
    .B(_1391_));
 sg13g2_nand3_1 _2201_ (.B(_1386_),
    .C(_1308_),
    .A(_1307_),
    .Y(_1396_));
 sg13g2_nand2_1 _2202_ (.Y(_1397_),
    .A(_1395_),
    .B(_1396_));
 sg13g2_inv_2 _2203_ (.Y(_1398_),
    .A(_1298_));
 sg13g2_nand2_1 _2204_ (.Y(_1399_),
    .A(_1397_),
    .B(_1398_));
 sg13g2_nand3_1 _2205_ (.B(_1399_),
    .C(_1119_),
    .A(_1394_),
    .Y(_1400_));
 sg13g2_xor2_1 _2206_ (.B(_1391_),
    .A(_1277_),
    .X(_1401_));
 sg13g2_nand2_1 _2207_ (.Y(_1402_),
    .A(_1275_),
    .B(_1274_));
 sg13g2_xnor2_1 _2208_ (.Y(_1403_),
    .A(_1401_),
    .B(_1402_));
 sg13g2_nand2_1 _2209_ (.Y(_1404_),
    .A(_1372_),
    .B(_1374_));
 sg13g2_nand2_1 _2210_ (.Y(_1405_),
    .A(_1404_),
    .B(net79));
 sg13g2_nand2_1 _2211_ (.Y(_1406_),
    .A(_1383_),
    .B(_1103_));
 sg13g2_nand2_1 _2212_ (.Y(_1407_),
    .A(_1405_),
    .B(_1406_));
 sg13g2_o21ai_1 _2213_ (.B1(_1285_),
    .Y(_1408_),
    .A1(_1284_),
    .A2(_1388_));
 sg13g2_a221oi_1 _2214_ (.B2(_1139_),
    .C1(_1408_),
    .B1(_1389_),
    .A1(_1127_),
    .Y(_1409_),
    .A2(_1407_));
 sg13g2_nand2_1 _2215_ (.Y(_1410_),
    .A(_1386_),
    .B(_1136_));
 sg13g2_nor2_1 _2216_ (.A(_1388_),
    .B(_1385_),
    .Y(_1411_));
 sg13g2_nand2_1 _2217_ (.Y(_1412_),
    .A(_1411_),
    .B(_1123_));
 sg13g2_nand3_1 _2218_ (.B(_1410_),
    .C(_1412_),
    .A(_1409_),
    .Y(_1413_));
 sg13g2_a21oi_1 _2219_ (.A1(_1403_),
    .A2(_1152_),
    .Y(_1414_),
    .B1(_1413_));
 sg13g2_nand2_1 _2220_ (.Y(_1415_),
    .A(_1400_),
    .B(_1414_));
 sg13g2_nand2_1 _2221_ (.Y(_1416_),
    .A(_1393_),
    .B(net75));
 sg13g2_nand3_1 _2222_ (.B(_1162_),
    .C(_1416_),
    .A(_1415_),
    .Y(_1417_));
 sg13g2_nand3_1 _2223_ (.B(_1161_),
    .C(_1301_),
    .A(_1300_),
    .Y(_1418_));
 sg13g2_nand2_2 _2224_ (.Y(_1419_),
    .A(_1417_),
    .B(_1418_));
 sg13g2_mux2_1 _2225_ (.A0(\DJ8.ACC[2] ),
    .A1(_1419_),
    .S(_0768_),
    .X(_0040_));
 sg13g2_nor2_1 _2226_ (.A(_1298_),
    .B(_1393_),
    .Y(_1420_));
 sg13g2_nor2_1 _2227_ (.A(net83),
    .B(_0020_),
    .Y(_1421_));
 sg13g2_nand2b_1 _2228_ (.Y(_1422_),
    .B(net83),
    .A_N(_0005_));
 sg13g2_nand2b_2 _2229_ (.Y(_1423_),
    .B(_1422_),
    .A_N(_1421_));
 sg13g2_nand2_1 _2230_ (.Y(_1424_),
    .A(_0862_),
    .B(_1331_));
 sg13g2_nand3_1 _2231_ (.B(net50),
    .C(net35),
    .A(_1210_),
    .Y(_1425_));
 sg13g2_nand2_1 _2232_ (.Y(_1426_),
    .A(_1425_),
    .B(_0865_));
 sg13g2_nand2_1 _2233_ (.Y(_1427_),
    .A(_1424_),
    .B(_1426_));
 sg13g2_nor2_1 _2234_ (.A(_1352_),
    .B(_1427_),
    .Y(_1428_));
 sg13g2_nor2_1 _2235_ (.A(net55),
    .B(_1428_),
    .Y(_1429_));
 sg13g2_inv_1 _2236_ (.Y(_1430_),
    .A(_0931_));
 sg13g2_nor2_1 _2237_ (.A(_1210_),
    .B(_1430_),
    .Y(_1431_));
 sg13g2_nand2_1 _2238_ (.Y(_1432_),
    .A(net86),
    .B(\DJ8.pc[0] ));
 sg13g2_nor2b_1 _2239_ (.A(_0850_),
    .B_N(_1432_),
    .Y(_1433_));
 sg13g2_nor2_1 _2240_ (.A(_1433_),
    .B(_1241_),
    .Y(_1434_));
 sg13g2_nor2_1 _2241_ (.A(_1431_),
    .B(_1434_),
    .Y(_1435_));
 sg13g2_nand2_1 _2242_ (.Y(_1436_),
    .A(_1313_),
    .B(_0935_));
 sg13g2_nand2_1 _2243_ (.Y(_1437_),
    .A(_1435_),
    .B(_1436_));
 sg13g2_nand2_1 _2244_ (.Y(_1438_),
    .A(_1437_),
    .B(net30));
 sg13g2_buf_1 _2245_ (.A(net63),
    .X(_1439_));
 sg13g2_nand2_1 _2246_ (.Y(_1440_),
    .A(_1192_),
    .B(_0931_));
 sg13g2_a21oi_1 _2247_ (.A1(_1440_),
    .A2(_1065_),
    .Y(_1441_),
    .B1(_0914_));
 sg13g2_nor2_1 _2248_ (.A(net47),
    .B(_1441_),
    .Y(_1442_));
 sg13g2_nand2_1 _2249_ (.Y(_1443_),
    .A(_1438_),
    .B(_1442_));
 sg13g2_a21oi_1 _2250_ (.A1(_1429_),
    .A2(_1443_),
    .Y(_1444_),
    .B1(_0965_));
 sg13g2_buf_1 _2251_ (.A(_0871_),
    .X(_1445_));
 sg13g2_a21oi_1 _2252_ (.A1(_0940_),
    .A2(_1065_),
    .Y(_1446_),
    .B1(net40));
 sg13g2_nor2_1 _2253_ (.A(net35),
    .B(_1082_),
    .Y(_1447_));
 sg13g2_nor3_1 _2254_ (.A(net31),
    .B(net32),
    .C(_1447_),
    .Y(_1448_));
 sg13g2_nand2b_1 _2255_ (.Y(_1449_),
    .B(_1448_),
    .A_N(_1446_));
 sg13g2_nand2_1 _2256_ (.Y(_1450_),
    .A(_0939_),
    .B(_1430_));
 sg13g2_nand3_1 _2257_ (.B(_1450_),
    .C(net31),
    .A(_0955_),
    .Y(_1451_));
 sg13g2_inv_1 _2258_ (.Y(_1452_),
    .A(_0853_));
 sg13g2_nor2_1 _2259_ (.A(_0972_),
    .B(_1452_),
    .Y(_1453_));
 sg13g2_nor2_1 _2260_ (.A(_1453_),
    .B(_1363_),
    .Y(_1454_));
 sg13g2_nand2_1 _2261_ (.Y(_1455_),
    .A(_1451_),
    .B(_1454_));
 sg13g2_a21oi_1 _2262_ (.A1(_1436_),
    .A2(_1047_),
    .Y(_1456_),
    .B1(net49));
 sg13g2_nand3_1 _2263_ (.B(_1455_),
    .C(_1456_),
    .A(_1449_),
    .Y(_1457_));
 sg13g2_a21oi_1 _2264_ (.A1(_1444_),
    .A2(_1457_),
    .Y(_1458_),
    .B1(net41));
 sg13g2_nor2_1 _2265_ (.A(net40),
    .B(_1344_),
    .Y(_1459_));
 sg13g2_o21ai_1 _2266_ (.B1(net32),
    .Y(_1460_),
    .A1(net30),
    .A2(_1459_));
 sg13g2_a21oi_1 _2267_ (.A1(_0972_),
    .A2(net38),
    .Y(_1461_),
    .B1(_1198_));
 sg13g2_nor2_1 _2268_ (.A(_1434_),
    .B(_1461_),
    .Y(_1462_));
 sg13g2_nand2_1 _2269_ (.Y(_1463_),
    .A(_0939_),
    .B(_1047_));
 sg13g2_a21oi_1 _2270_ (.A1(_1038_),
    .A2(_1241_),
    .Y(_1464_),
    .B1(_1463_));
 sg13g2_o21ai_1 _2271_ (.B1(_0865_),
    .Y(_1465_),
    .A1(net35),
    .A2(_1234_));
 sg13g2_nor2_1 _2272_ (.A(net42),
    .B(_1465_),
    .Y(_1466_));
 sg13g2_nor3_1 _2273_ (.A(net55),
    .B(_1464_),
    .C(_1466_),
    .Y(_1467_));
 sg13g2_o21ai_1 _2274_ (.B1(_1467_),
    .Y(_1468_),
    .A1(_1460_),
    .A2(_1462_));
 sg13g2_nor2_1 _2275_ (.A(_0934_),
    .B(net50),
    .Y(_1469_));
 sg13g2_nor3_1 _2276_ (.A(_1058_),
    .B(_1331_),
    .C(_1469_),
    .Y(_1470_));
 sg13g2_nand2_1 _2277_ (.Y(_1471_),
    .A(_1073_),
    .B(_0951_));
 sg13g2_nand2_1 _2278_ (.Y(_1472_),
    .A(_1471_),
    .B(_0914_));
 sg13g2_nor2_1 _2279_ (.A(net42),
    .B(_1332_),
    .Y(_1473_));
 sg13g2_nand2_1 _2280_ (.Y(_1474_),
    .A(_1472_),
    .B(_1473_));
 sg13g2_nand2b_1 _2281_ (.Y(_1475_),
    .B(_1474_),
    .A_N(_1470_));
 sg13g2_nand2_1 _2282_ (.Y(_1476_),
    .A(_1475_),
    .B(net55));
 sg13g2_nand2_1 _2283_ (.Y(_1477_),
    .A(_1468_),
    .B(_1476_));
 sg13g2_nand2_1 _2284_ (.Y(_1478_),
    .A(_1477_),
    .B(net43));
 sg13g2_nand2_1 _2285_ (.Y(_1479_),
    .A(_1458_),
    .B(_1478_));
 sg13g2_nand2_1 _2286_ (.Y(_1480_),
    .A(net41),
    .B(net6));
 sg13g2_nand3_1 _2287_ (.B(_1092_),
    .C(_1480_),
    .A(_1479_),
    .Y(_1481_));
 sg13g2_inv_1 _2288_ (.Y(_1482_),
    .A(\DJ8.ACC[4] ));
 sg13g2_a221oi_1 _2289_ (.B2(\DJ8.EF[12] ),
    .C1(net69),
    .B1(_1004_),
    .A1(_1020_),
    .Y(_1483_),
    .A2(\DJ8.REGS.regs[3][4] ));
 sg13g2_inv_1 _2290_ (.Y(_1484_),
    .A(\DJ8.GH[12] ));
 sg13g2_a22oi_1 _2291_ (.Y(_0136_),
    .B1(\DJ8.EF[4] ),
    .B2(_1007_),
    .A2(_1013_),
    .A1(\DJ8.GH[4] ));
 sg13g2_o21ai_1 _2292_ (.B1(_0136_),
    .Y(_0137_),
    .A1(_1484_),
    .A2(_1010_));
 sg13g2_a221oi_1 _2293_ (.B2(_1018_),
    .C1(_0137_),
    .B1(\DJ8.REGS.regs[1][4] ),
    .A1(\DJ8.REGS.regs[2][4] ),
    .Y(_0138_),
    .A2(_1022_));
 sg13g2_a22oi_1 _2294_ (.Y(_0139_),
    .B1(_1483_),
    .B2(_0138_),
    .A2(net69),
    .A1(_1482_));
 sg13g2_nor2_1 _2295_ (.A(net79),
    .B(_0139_),
    .Y(_0140_));
 sg13g2_inv_1 _2296_ (.Y(_0141_),
    .A(_0140_));
 sg13g2_nand2_1 _2297_ (.Y(_0142_),
    .A(_1481_),
    .B(_0141_));
 sg13g2_xnor2_1 _2298_ (.Y(_0143_),
    .A(_1423_),
    .B(_0142_));
 sg13g2_nand2_1 _2299_ (.Y(_0144_),
    .A(_1281_),
    .B(_1389_));
 sg13g2_nand2_1 _2300_ (.Y(_0145_),
    .A(_0144_),
    .B(_1390_));
 sg13g2_nor2_1 _2301_ (.A(_1391_),
    .B(_1274_),
    .Y(_0146_));
 sg13g2_nand2_1 _2302_ (.Y(_0147_),
    .A(_0146_),
    .B(_1292_));
 sg13g2_nand2b_1 _2303_ (.Y(_0148_),
    .B(_0147_),
    .A_N(_0145_));
 sg13g2_xnor2_1 _2304_ (.Y(_0149_),
    .A(_0143_),
    .B(_0148_));
 sg13g2_inv_1 _2305_ (.Y(_0150_),
    .A(_0149_));
 sg13g2_nand2_1 _2306_ (.Y(_0151_),
    .A(_1420_),
    .B(_0150_));
 sg13g2_nand2_1 _2307_ (.Y(_0152_),
    .A(_1399_),
    .B(_0149_));
 sg13g2_nand3_1 _2308_ (.B(_0152_),
    .C(_1119_),
    .A(_0151_),
    .Y(_0153_));
 sg13g2_nor2_1 _2309_ (.A(_1388_),
    .B(_1407_),
    .Y(_0154_));
 sg13g2_nand2b_1 _2310_ (.Y(_0155_),
    .B(_0143_),
    .A_N(_0154_));
 sg13g2_inv_1 _2311_ (.Y(_0156_),
    .A(_1423_));
 sg13g2_nand2_1 _2312_ (.Y(_0157_),
    .A(_0142_),
    .B(_0156_));
 sg13g2_nand3_1 _2313_ (.B(_1423_),
    .C(_0141_),
    .A(_1481_),
    .Y(_0158_));
 sg13g2_nand2_1 _2314_ (.Y(_0159_),
    .A(_0157_),
    .B(_0158_));
 sg13g2_nand2_1 _2315_ (.Y(_0160_),
    .A(_0159_),
    .B(_0154_));
 sg13g2_nand2_1 _2316_ (.Y(_0161_),
    .A(_0155_),
    .B(_0160_));
 sg13g2_nor2_1 _2317_ (.A(_1279_),
    .B(_1275_),
    .Y(_0162_));
 sg13g2_nor2b_1 _2318_ (.A(_1386_),
    .B_N(_1278_),
    .Y(_0163_));
 sg13g2_nor2b_1 _2319_ (.A(_0162_),
    .B_N(_0163_),
    .Y(_0164_));
 sg13g2_nor2_1 _2320_ (.A(_0161_),
    .B(_0164_),
    .Y(_0165_));
 sg13g2_nor2b_1 _2321_ (.A(_0165_),
    .B_N(_1152_),
    .Y(_0166_));
 sg13g2_nand2_1 _2322_ (.Y(_0167_),
    .A(_0164_),
    .B(_0161_));
 sg13g2_inv_1 _2323_ (.Y(_0168_),
    .A(_0142_));
 sg13g2_o21ai_1 _2324_ (.B1(_1285_),
    .Y(_0169_),
    .A1(_1284_),
    .A2(_0156_));
 sg13g2_a221oi_1 _2325_ (.B2(_1139_),
    .C1(_0169_),
    .B1(_0157_),
    .A1(_0168_),
    .Y(_0170_),
    .A2(_1127_));
 sg13g2_nand2_1 _2326_ (.Y(_0171_),
    .A(_0143_),
    .B(_1136_));
 sg13g2_inv_1 _2327_ (.Y(_0172_),
    .A(_0158_));
 sg13g2_nand2_1 _2328_ (.Y(_0173_),
    .A(_0172_),
    .B(_1123_));
 sg13g2_nand3_1 _2329_ (.B(_0171_),
    .C(_0173_),
    .A(_0170_),
    .Y(_0174_));
 sg13g2_a21oi_1 _2330_ (.A1(_0166_),
    .A2(_0167_),
    .Y(_0175_),
    .B1(_0174_));
 sg13g2_nand2_1 _2331_ (.Y(_0176_),
    .A(_0153_),
    .B(_0175_));
 sg13g2_nand2_1 _2332_ (.Y(_0177_),
    .A(_0149_),
    .B(net75));
 sg13g2_nand3_1 _2333_ (.B(_1162_),
    .C(_0177_),
    .A(_0176_),
    .Y(_0178_));
 sg13g2_nand3_1 _2334_ (.B(_1161_),
    .C(_1416_),
    .A(_1415_),
    .Y(_0179_));
 sg13g2_nand2_1 _2335_ (.Y(_0180_),
    .A(_0178_),
    .B(_0179_));
 sg13g2_inv_2 _2336_ (.Y(_0181_),
    .A(_0180_));
 sg13g2_nor2_1 _2337_ (.A(\DJ8.ACC[3] ),
    .B(net66),
    .Y(_0182_));
 sg13g2_a21oi_1 _2338_ (.A1(_0181_),
    .A2(net66),
    .Y(_0041_),
    .B1(_0182_));
 sg13g2_a21oi_1 _2339_ (.A1(_0176_),
    .A2(_0177_),
    .Y(_0183_),
    .B1(_1162_));
 sg13g2_nor3_1 _2340_ (.A(_0835_),
    .B(net52),
    .C(_0939_),
    .Y(_0184_));
 sg13g2_nand2_1 _2341_ (.Y(_0185_),
    .A(_0900_),
    .B(net51));
 sg13g2_a21oi_1 _2342_ (.A1(_0185_),
    .A2(_0884_),
    .Y(_0186_),
    .B1(net31));
 sg13g2_o21ai_1 _2343_ (.B1(net47),
    .Y(_0187_),
    .A1(_0184_),
    .A2(_0186_));
 sg13g2_a21oi_1 _2344_ (.A1(_0926_),
    .A2(_0932_),
    .Y(_0188_),
    .B1(_1187_));
 sg13g2_nand2_1 _2345_ (.Y(_0189_),
    .A(_0851_),
    .B(net34));
 sg13g2_nor2_1 _2346_ (.A(_1433_),
    .B(net33),
    .Y(_0190_));
 sg13g2_nor2_1 _2347_ (.A(_0189_),
    .B(_0190_),
    .Y(_0191_));
 sg13g2_nand2_1 _2348_ (.Y(_0192_),
    .A(_0851_),
    .B(net44));
 sg13g2_a21oi_1 _2349_ (.A1(_0192_),
    .A2(_1065_),
    .Y(_0193_),
    .B1(net34));
 sg13g2_nor2_1 _2350_ (.A(_0191_),
    .B(_0193_),
    .Y(_0194_));
 sg13g2_nor2_1 _2351_ (.A(net63),
    .B(_0194_),
    .Y(_0195_));
 sg13g2_nor2_1 _2352_ (.A(_0188_),
    .B(_0195_),
    .Y(_0196_));
 sg13g2_nand3_1 _2353_ (.B(_0196_),
    .C(net48),
    .A(_0187_),
    .Y(_0197_));
 sg13g2_inv_1 _2354_ (.Y(_0198_),
    .A(_1433_));
 sg13g2_nor2_1 _2355_ (.A(net35),
    .B(_0885_),
    .Y(_0199_));
 sg13g2_o21ai_1 _2356_ (.B1(_0199_),
    .Y(_0200_),
    .A1(net70),
    .A2(_0198_));
 sg13g2_inv_1 _2357_ (.Y(_0201_),
    .A(_0861_));
 sg13g2_nand2_1 _2358_ (.Y(_0202_),
    .A(_0201_),
    .B(_1051_));
 sg13g2_nand2_1 _2359_ (.Y(_0203_),
    .A(_0200_),
    .B(_0202_));
 sg13g2_a21oi_1 _2360_ (.A1(_0203_),
    .A2(net30),
    .Y(_0204_),
    .B1(_0942_));
 sg13g2_nor2_1 _2361_ (.A(net33),
    .B(_0947_),
    .Y(_0205_));
 sg13g2_nand2_1 _2362_ (.Y(_0206_),
    .A(_0205_),
    .B(net39));
 sg13g2_nand2_1 _2363_ (.Y(_0207_),
    .A(_1194_),
    .B(_0922_));
 sg13g2_o21ai_1 _2364_ (.B1(net55),
    .Y(_0208_),
    .A1(_0193_),
    .A2(_0207_));
 sg13g2_a21oi_1 _2365_ (.A1(_0204_),
    .A2(_0206_),
    .Y(_0209_),
    .B1(_0208_));
 sg13g2_a21oi_1 _2366_ (.A1(_0197_),
    .A2(_0209_),
    .Y(_0210_),
    .B1(_1373_));
 sg13g2_inv_1 _2367_ (.Y(_0211_),
    .A(_1344_));
 sg13g2_a22oi_1 _2368_ (.Y(_0212_),
    .B1(_0892_),
    .B2(_1072_),
    .A2(net39),
    .A1(_0211_));
 sg13g2_nor2_1 _2369_ (.A(net32),
    .B(_0212_),
    .Y(_0213_));
 sg13g2_nor2_1 _2370_ (.A(_1042_),
    .B(_1452_),
    .Y(_0214_));
 sg13g2_inv_1 _2371_ (.Y(_0215_),
    .A(_0214_));
 sg13g2_nor2_1 _2372_ (.A(net50),
    .B(_0905_),
    .Y(_0216_));
 sg13g2_a21oi_1 _2373_ (.A1(_0905_),
    .A2(_0903_),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_o21ai_1 _2374_ (.B1(_0878_),
    .Y(_0218_),
    .A1(_0215_),
    .A2(_0217_));
 sg13g2_nor2_1 _2375_ (.A(_0213_),
    .B(_0218_),
    .Y(_0219_));
 sg13g2_a21oi_1 _2376_ (.A1(net40),
    .A2(_0870_),
    .Y(_0220_),
    .B1(_1431_));
 sg13g2_nor2_1 _2377_ (.A(net30),
    .B(_0220_),
    .Y(_0221_));
 sg13g2_nor2_1 _2378_ (.A(_1051_),
    .B(_1214_),
    .Y(_0222_));
 sg13g2_nor3_1 _2379_ (.A(net31),
    .B(_0201_),
    .C(_0222_),
    .Y(_0223_));
 sg13g2_o21ai_1 _2380_ (.B1(_1348_),
    .Y(_0224_),
    .A1(_0221_),
    .A2(_0223_));
 sg13g2_a21oi_1 _2381_ (.A1(_0219_),
    .A2(_0224_),
    .Y(_0225_),
    .B1(_0785_));
 sg13g2_nor2_1 _2382_ (.A(net53),
    .B(_0967_),
    .Y(_0226_));
 sg13g2_nor2_1 _2383_ (.A(net36),
    .B(_0226_),
    .Y(_0227_));
 sg13g2_nand2_1 _2384_ (.Y(_0228_),
    .A(_1212_),
    .B(net40));
 sg13g2_nand2_1 _2385_ (.Y(_0229_),
    .A(_0227_),
    .B(_0228_));
 sg13g2_nor2_1 _2386_ (.A(net34),
    .B(_0950_),
    .Y(_0230_));
 sg13g2_o21ai_1 _2387_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_1445_),
    .A2(_1072_));
 sg13g2_nand2_1 _2388_ (.Y(_0232_),
    .A(_0229_),
    .B(_0231_));
 sg13g2_nand2_1 _2389_ (.Y(_0233_),
    .A(_0232_),
    .B(_1439_));
 sg13g2_nor2_1 _2390_ (.A(net40),
    .B(_0822_),
    .Y(_0234_));
 sg13g2_nor2_1 _2391_ (.A(_1067_),
    .B(_1469_),
    .Y(_0235_));
 sg13g2_nand2_1 _2392_ (.Y(_0236_),
    .A(_0235_),
    .B(_0926_));
 sg13g2_o21ai_1 _2393_ (.B1(_1042_),
    .Y(_0237_),
    .A1(_0234_),
    .A2(_0236_));
 sg13g2_nor2_1 _2394_ (.A(_0227_),
    .B(_0237_),
    .Y(_0238_));
 sg13g2_nor2_1 _2395_ (.A(net48),
    .B(_0238_),
    .Y(_0239_));
 sg13g2_nand2_1 _2396_ (.Y(_0240_),
    .A(_0233_),
    .B(_0239_));
 sg13g2_nand2_1 _2397_ (.Y(_0241_),
    .A(_0225_),
    .B(_0240_));
 sg13g2_nand2_1 _2398_ (.Y(_0242_),
    .A(_0210_),
    .B(_0241_));
 sg13g2_nand2b_1 _2399_ (.Y(_0243_),
    .B(net41),
    .A_N(net7));
 sg13g2_nand3_1 _2400_ (.B(_1092_),
    .C(_0243_),
    .A(_0242_),
    .Y(_0244_));
 sg13g2_a22oi_1 _2401_ (.Y(_0245_),
    .B1(\DJ8.EF[5] ),
    .B2(_1007_),
    .A2(\DJ8.EF[13] ),
    .A1(_1004_));
 sg13g2_a22oi_1 _2402_ (.Y(_0246_),
    .B1(\DJ8.REGS.regs[2][5] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][5] ));
 sg13g2_inv_1 _2403_ (.Y(_0247_),
    .A(\DJ8.GH[13] ));
 sg13g2_nor2_1 _2404_ (.A(_0247_),
    .B(_1010_),
    .Y(_0248_));
 sg13g2_a21oi_1 _2405_ (.A1(\DJ8.GH[5] ),
    .A2(_1013_),
    .Y(_0249_),
    .B1(_0248_));
 sg13g2_nand2_1 _2406_ (.Y(_0250_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][5] ));
 sg13g2_nand4_1 _2407_ (.B(_0246_),
    .C(_0249_),
    .A(_0245_),
    .Y(_0251_),
    .D(_0250_));
 sg13g2_a21oi_1 _2408_ (.A1(\DJ8.ACC[5] ),
    .A2(_1025_),
    .Y(_0252_),
    .B1(_0251_));
 sg13g2_nand2b_1 _2409_ (.Y(_0253_),
    .B(_1103_),
    .A_N(_0252_));
 sg13g2_nand2_1 _2410_ (.Y(_0254_),
    .A(_0244_),
    .B(_0253_));
 sg13g2_nor2_1 _2411_ (.A(_1156_),
    .B(_0022_),
    .Y(_0255_));
 sg13g2_nand2b_1 _2412_ (.Y(_0256_),
    .B(_1156_),
    .A_N(_0021_));
 sg13g2_nand2b_1 _2413_ (.Y(_0257_),
    .B(_0256_),
    .A_N(_0255_));
 sg13g2_nand2_1 _2414_ (.Y(_0258_),
    .A(_0254_),
    .B(_0257_));
 sg13g2_inv_1 _2415_ (.Y(_0259_),
    .A(_0257_));
 sg13g2_nand3_1 _2416_ (.B(_0253_),
    .C(_0259_),
    .A(_0244_),
    .Y(_0260_));
 sg13g2_nand2_2 _2417_ (.Y(_0261_),
    .A(_0258_),
    .B(_0260_));
 sg13g2_nand2_1 _2418_ (.Y(_0262_),
    .A(_0143_),
    .B(_1386_));
 sg13g2_nor2_1 _2419_ (.A(_1308_),
    .B(_0262_),
    .Y(_0263_));
 sg13g2_a21oi_1 _2420_ (.A1(_0157_),
    .A2(_1411_),
    .Y(_0264_),
    .B1(_0172_));
 sg13g2_nor2b_1 _2421_ (.A(_0263_),
    .B_N(_0264_),
    .Y(_0265_));
 sg13g2_nor2_1 _2422_ (.A(_1274_),
    .B(_1113_),
    .Y(_0266_));
 sg13g2_nor2_1 _2423_ (.A(_1391_),
    .B(_0159_),
    .Y(_0267_));
 sg13g2_nand3_1 _2424_ (.B(_0267_),
    .C(_1033_),
    .A(_0266_),
    .Y(_0268_));
 sg13g2_nand2_1 _2425_ (.Y(_0269_),
    .A(_0265_),
    .B(_0268_));
 sg13g2_xnor2_1 _2426_ (.Y(_0270_),
    .A(_0261_),
    .B(_0269_));
 sg13g2_inv_1 _2427_ (.Y(_0271_),
    .A(_0270_));
 sg13g2_nand2_1 _2428_ (.Y(_0272_),
    .A(_0271_),
    .B(_0151_));
 sg13g2_nor2_1 _2429_ (.A(_0149_),
    .B(_1399_),
    .Y(_0273_));
 sg13g2_nand2_1 _2430_ (.Y(_0274_),
    .A(_0273_),
    .B(_0270_));
 sg13g2_nand3_1 _2431_ (.B(_0274_),
    .C(_1119_),
    .A(_0272_),
    .Y(_0275_));
 sg13g2_nor2_1 _2432_ (.A(_1401_),
    .B(_0161_),
    .Y(_0276_));
 sg13g2_nand2_1 _2433_ (.Y(_0277_),
    .A(_0276_),
    .B(_1402_));
 sg13g2_nand2_1 _2434_ (.Y(_0278_),
    .A(_1386_),
    .B(_1277_));
 sg13g2_nand2_1 _2435_ (.Y(_0279_),
    .A(_0155_),
    .B(_0278_));
 sg13g2_nand2_1 _2436_ (.Y(_0280_),
    .A(_0279_),
    .B(_0160_));
 sg13g2_inv_2 _2437_ (.Y(_0281_),
    .A(_0261_));
 sg13g2_nand2_1 _2438_ (.Y(_0282_),
    .A(_0142_),
    .B(_1423_));
 sg13g2_nand2_1 _2439_ (.Y(_0283_),
    .A(_0281_),
    .B(_0282_));
 sg13g2_nand2b_1 _2440_ (.Y(_0284_),
    .B(_0261_),
    .A_N(_0282_));
 sg13g2_nand2_1 _2441_ (.Y(_0285_),
    .A(_0283_),
    .B(_0284_));
 sg13g2_a21oi_1 _2442_ (.A1(_0277_),
    .A2(_0280_),
    .Y(_0286_),
    .B1(_0285_));
 sg13g2_nor2b_1 _2443_ (.A(_0286_),
    .B_N(_1152_),
    .Y(_0287_));
 sg13g2_nand3_1 _2444_ (.B(_0280_),
    .C(_0285_),
    .A(_0277_),
    .Y(_0288_));
 sg13g2_a221oi_1 _2445_ (.B2(_1127_),
    .C1(_1132_),
    .B1(_0254_),
    .A1(_1129_),
    .Y(_0289_),
    .A2(_0257_));
 sg13g2_nand2_1 _2446_ (.Y(_0290_),
    .A(_0281_),
    .B(_1136_));
 sg13g2_nand2_1 _2447_ (.Y(_0291_),
    .A(_0260_),
    .B(_1139_));
 sg13g2_nand3_1 _2448_ (.B(_1123_),
    .C(_0257_),
    .A(_0254_),
    .Y(_0292_));
 sg13g2_nand4_1 _2449_ (.B(_0290_),
    .C(_0291_),
    .A(_0289_),
    .Y(_0293_),
    .D(_0292_));
 sg13g2_a21oi_1 _2450_ (.A1(_0287_),
    .A2(_0288_),
    .Y(_0294_),
    .B1(_0293_));
 sg13g2_nand2_1 _2451_ (.Y(_0295_),
    .A(_0275_),
    .B(_0294_));
 sg13g2_nand2_1 _2452_ (.Y(_0296_),
    .A(_0271_),
    .B(net75));
 sg13g2_nand2_1 _2453_ (.Y(_0297_),
    .A(_0295_),
    .B(_0296_));
 sg13g2_nand2_1 _2454_ (.Y(_0298_),
    .A(_0297_),
    .B(_1162_));
 sg13g2_nand2b_1 _2455_ (.Y(_0299_),
    .B(_0298_),
    .A_N(_0183_));
 sg13g2_buf_1 _2456_ (.A(_0299_),
    .X(_0300_));
 sg13g2_nor2_1 _2457_ (.A(\DJ8.ACC[4] ),
    .B(net66),
    .Y(_0301_));
 sg13g2_a21oi_1 _2458_ (.A1(net29),
    .A2(net66),
    .Y(_0042_),
    .B1(_0301_));
 sg13g2_nand2_1 _2459_ (.Y(_0302_),
    .A(_1227_),
    .B(net31));
 sg13g2_nor2_1 _2460_ (.A(_0302_),
    .B(_1446_),
    .Y(_0303_));
 sg13g2_nand4_1 _2461_ (.B(_1365_),
    .C(_1045_),
    .A(_0884_),
    .Y(_0304_),
    .D(_1440_));
 sg13g2_nor2b_1 _2462_ (.A(_0303_),
    .B_N(_0304_),
    .Y(_0305_));
 sg13g2_nor3_1 _2463_ (.A(_1370_),
    .B(_1453_),
    .C(_1069_),
    .Y(_0306_));
 sg13g2_a21oi_1 _2464_ (.A1(_0854_),
    .A2(_0306_),
    .Y(_0307_),
    .B1(net32));
 sg13g2_o21ai_1 _2465_ (.B1(_0307_),
    .Y(_0308_),
    .A1(net43),
    .A2(_0305_));
 sg13g2_nand2b_1 _2466_ (.Y(_0309_),
    .B(_0951_),
    .A_N(_0189_));
 sg13g2_nand4_1 _2467_ (.B(net48),
    .C(_1078_),
    .A(_0309_),
    .Y(_0310_),
    .D(_1190_));
 sg13g2_a21oi_1 _2468_ (.A1(net37),
    .A2(_0894_),
    .Y(_0311_),
    .B1(net48));
 sg13g2_a21oi_1 _2469_ (.A1(_1424_),
    .A2(_0311_),
    .Y(_0312_),
    .B1(net47));
 sg13g2_a21oi_1 _2470_ (.A1(_0310_),
    .A2(_0312_),
    .Y(_0313_),
    .B1(_1062_));
 sg13g2_a21oi_1 _2471_ (.A1(_0308_),
    .A2(_0313_),
    .Y(_0314_),
    .B1(net41));
 sg13g2_o21ai_1 _2472_ (.B1(_0230_),
    .Y(_0315_),
    .A1(_0900_),
    .A2(_0919_));
 sg13g2_nand3_1 _2473_ (.B(_0899_),
    .C(_0836_),
    .A(net33),
    .Y(_0316_));
 sg13g2_nand3_1 _2474_ (.B(_1194_),
    .C(_0316_),
    .A(_0315_),
    .Y(_0317_));
 sg13g2_nand2_1 _2475_ (.Y(_0318_),
    .A(_0317_),
    .B(net32));
 sg13g2_nand3_1 _2476_ (.B(_1365_),
    .C(_0926_),
    .A(_1325_),
    .Y(_0319_));
 sg13g2_o21ai_1 _2477_ (.B1(net31),
    .Y(_0320_),
    .A1(_1445_),
    .A2(_0910_));
 sg13g2_nand3_1 _2478_ (.B(net47),
    .C(_0320_),
    .A(_0319_),
    .Y(_0321_));
 sg13g2_nand3_1 _2479_ (.B(_0321_),
    .C(net48),
    .A(_0318_),
    .Y(_0322_));
 sg13g2_o21ai_1 _2480_ (.B1(net30),
    .Y(_0323_),
    .A1(_1459_),
    .A2(_1324_));
 sg13g2_nand2_1 _2481_ (.Y(_0324_),
    .A(_0908_),
    .B(_0889_));
 sg13g2_a21oi_1 _2482_ (.A1(_0323_),
    .A2(_0324_),
    .Y(_0325_),
    .B1(_1439_));
 sg13g2_a21oi_1 _2483_ (.A1(_0883_),
    .A2(net33),
    .Y(_0326_),
    .B1(_0190_));
 sg13g2_nor2b_1 _2484_ (.A(_0862_),
    .B_N(_1220_),
    .Y(_0327_));
 sg13g2_o21ai_1 _2485_ (.B1(_0327_),
    .Y(_0328_),
    .A1(net40),
    .A2(_0326_));
 sg13g2_o21ai_1 _2486_ (.B1(_0965_),
    .Y(_0329_),
    .A1(_0959_),
    .A2(_0215_));
 sg13g2_a21oi_1 _2487_ (.A1(_0328_),
    .A2(_1047_),
    .Y(_0330_),
    .B1(_0329_));
 sg13g2_nand2b_1 _2488_ (.Y(_0331_),
    .B(_0330_),
    .A_N(_0325_));
 sg13g2_nand2_1 _2489_ (.Y(_0332_),
    .A(_0322_),
    .B(_0331_));
 sg13g2_nand2_1 _2490_ (.Y(_0333_),
    .A(_0332_),
    .B(_1062_));
 sg13g2_nand2_1 _2491_ (.Y(_0334_),
    .A(_0314_),
    .B(_0333_));
 sg13g2_nand2_1 _2492_ (.Y(_0335_),
    .A(net41),
    .B(net8));
 sg13g2_nand3_1 _2493_ (.B(net79),
    .C(_0335_),
    .A(_0334_),
    .Y(_0336_));
 sg13g2_inv_1 _2494_ (.Y(_0337_),
    .A(\DJ8.GH[14] ));
 sg13g2_nand2_1 _2495_ (.Y(_0338_),
    .A(_1013_),
    .B(\DJ8.GH[6] ));
 sg13g2_o21ai_1 _2496_ (.B1(_0338_),
    .Y(_0339_),
    .A1(_0337_),
    .A2(_1010_));
 sg13g2_a221oi_1 _2497_ (.B2(_1004_),
    .C1(_0339_),
    .B1(\DJ8.EF[14] ),
    .A1(\DJ8.EF[6] ),
    .Y(_0340_),
    .A2(_1007_));
 sg13g2_nand2_1 _2498_ (.Y(_0341_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][6] ));
 sg13g2_a22oi_1 _2499_ (.Y(_0342_),
    .B1(\DJ8.REGS.regs[2][6] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][6] ));
 sg13g2_nand2_1 _2500_ (.Y(_0343_),
    .A(net69),
    .B(\DJ8.ACC[6] ));
 sg13g2_nand4_1 _2501_ (.B(_0341_),
    .C(_0342_),
    .A(_0340_),
    .Y(_0344_),
    .D(_0343_));
 sg13g2_nand2b_1 _2502_ (.Y(_0345_),
    .B(_1103_),
    .A_N(_0344_));
 sg13g2_nand2_1 _2503_ (.Y(_0346_),
    .A(_0336_),
    .B(_0345_));
 sg13g2_nor2_1 _2504_ (.A(net83),
    .B(_0024_),
    .Y(_0347_));
 sg13g2_nand2b_1 _2505_ (.Y(_0348_),
    .B(net83),
    .A_N(_0023_));
 sg13g2_nand2b_1 _2506_ (.Y(_0349_),
    .B(_0348_),
    .A_N(_0347_));
 sg13g2_inv_1 _2507_ (.Y(_0350_),
    .A(_0349_));
 sg13g2_nand2_1 _2508_ (.Y(_0351_),
    .A(_0346_),
    .B(_0350_));
 sg13g2_nand3_1 _2509_ (.B(_0345_),
    .C(_0349_),
    .A(_0336_),
    .Y(_0352_));
 sg13g2_nand2_2 _2510_ (.Y(_0353_),
    .A(_0351_),
    .B(_0352_));
 sg13g2_nor2_1 _2511_ (.A(_0261_),
    .B(_0159_),
    .Y(_0354_));
 sg13g2_inv_1 _2512_ (.Y(_0355_),
    .A(_0260_));
 sg13g2_o21ai_1 _2513_ (.B1(_0258_),
    .Y(_0356_),
    .A1(_0158_),
    .A2(_0355_));
 sg13g2_a21oi_1 _2514_ (.A1(_0354_),
    .A2(_0145_),
    .Y(_0357_),
    .B1(_0356_));
 sg13g2_nand3_1 _2515_ (.B(_0146_),
    .C(_1292_),
    .A(_0354_),
    .Y(_0358_));
 sg13g2_nand2_1 _2516_ (.Y(_0359_),
    .A(_0357_),
    .B(_0358_));
 sg13g2_xnor2_1 _2517_ (.Y(_0360_),
    .A(_0353_),
    .B(_0359_));
 sg13g2_inv_1 _2518_ (.Y(_0361_),
    .A(_0360_));
 sg13g2_nand2_1 _2519_ (.Y(_0362_),
    .A(_0274_),
    .B(_0361_));
 sg13g2_nand3_1 _2520_ (.B(_0270_),
    .C(_0360_),
    .A(_0273_),
    .Y(_0363_));
 sg13g2_nand3_1 _2521_ (.B(_0363_),
    .C(_1119_),
    .A(_0362_),
    .Y(_0364_));
 sg13g2_nand2_1 _2522_ (.Y(_0365_),
    .A(_0283_),
    .B(_0155_));
 sg13g2_nor2_1 _2523_ (.A(_0365_),
    .B(_0165_),
    .Y(_0366_));
 sg13g2_nor2_1 _2524_ (.A(_0259_),
    .B(_0254_),
    .Y(_0367_));
 sg13g2_nor2_1 _2525_ (.A(_0367_),
    .B(_0353_),
    .Y(_0368_));
 sg13g2_nand2_1 _2526_ (.Y(_0369_),
    .A(_0353_),
    .B(_0367_));
 sg13g2_nand2b_1 _2527_ (.Y(_0370_),
    .B(_0369_),
    .A_N(_0368_));
 sg13g2_inv_1 _2528_ (.Y(_0371_),
    .A(_0370_));
 sg13g2_nand3b_1 _2529_ (.B(_0284_),
    .C(_0371_),
    .Y(_0372_),
    .A_N(_0366_));
 sg13g2_inv_1 _2530_ (.Y(_0373_),
    .A(_0284_));
 sg13g2_o21ai_1 _2531_ (.B1(_0370_),
    .Y(_0374_),
    .A1(_0373_),
    .A2(_0366_));
 sg13g2_nand3_1 _2532_ (.B(_0374_),
    .C(_1152_),
    .A(_0372_),
    .Y(_0375_));
 sg13g2_inv_1 _2533_ (.Y(_0376_),
    .A(_0353_));
 sg13g2_inv_1 _2534_ (.Y(_0377_),
    .A(_1123_));
 sg13g2_inv_1 _2535_ (.Y(_0378_),
    .A(_0346_));
 sg13g2_a221oi_1 _2536_ (.B2(_1127_),
    .C1(_1132_),
    .B1(_0378_),
    .A1(_1129_),
    .Y(_0379_),
    .A2(_0349_));
 sg13g2_o21ai_1 _2537_ (.B1(_0379_),
    .Y(_0380_),
    .A1(_0377_),
    .A2(_0352_));
 sg13g2_a221oi_1 _2538_ (.B2(_0351_),
    .C1(_0380_),
    .B1(_1139_),
    .A1(_1136_),
    .Y(_0381_),
    .A2(_0376_));
 sg13g2_nand3_1 _2539_ (.B(_0375_),
    .C(_0381_),
    .A(_0364_),
    .Y(_0382_));
 sg13g2_nand2_1 _2540_ (.Y(_0383_),
    .A(_0361_),
    .B(net75));
 sg13g2_nand2_1 _2541_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_nand2_1 _2542_ (.Y(_0385_),
    .A(_0384_),
    .B(_1162_));
 sg13g2_nand2_1 _2543_ (.Y(_0386_),
    .A(_0297_),
    .B(_1161_));
 sg13g2_nand2_1 _2544_ (.Y(_0387_),
    .A(_0385_),
    .B(_0386_));
 sg13g2_nor2_1 _2545_ (.A(\DJ8.ACC[5] ),
    .B(_0768_),
    .Y(_0388_));
 sg13g2_a21oi_1 _2546_ (.A1(net28),
    .A2(net66),
    .Y(_0043_),
    .B1(_0388_));
 sg13g2_nor2_1 _2547_ (.A(_0361_),
    .B(_0274_),
    .Y(_0389_));
 sg13g2_nor2_1 _2548_ (.A(net83),
    .B(\DJ8.ACC[7] ),
    .Y(_0390_));
 sg13g2_a21oi_1 _2549_ (.A1(net83),
    .A2(_0003_),
    .Y(_0391_),
    .B1(_0390_));
 sg13g2_inv_1 _2550_ (.Y(_0392_),
    .A(_0391_));
 sg13g2_nand2_1 _2551_ (.Y(_0393_),
    .A(_0821_),
    .B(net52));
 sg13g2_nor2b_1 _2552_ (.A(_0205_),
    .B_N(_0393_),
    .Y(_0394_));
 sg13g2_o21ai_1 _2553_ (.B1(_1328_),
    .Y(_0395_),
    .A1(_0931_),
    .A2(_1447_));
 sg13g2_o21ai_1 _2554_ (.B1(_0395_),
    .Y(_0396_),
    .A1(_1452_),
    .A2(_0394_));
 sg13g2_a21oi_1 _2555_ (.A1(net37),
    .A2(_0952_),
    .Y(_0397_),
    .B1(_0396_));
 sg13g2_nand2_1 _2556_ (.Y(_0398_),
    .A(_0397_),
    .B(net47));
 sg13g2_nand2_1 _2557_ (.Y(_0399_),
    .A(_0202_),
    .B(_1430_));
 sg13g2_a21oi_1 _2558_ (.A1(_0952_),
    .A2(net40),
    .Y(_0400_),
    .B1(_0399_));
 sg13g2_a21oi_1 _2559_ (.A1(_1237_),
    .A2(net35),
    .Y(_0401_),
    .B1(net31));
 sg13g2_a21oi_1 _2560_ (.A1(_0401_),
    .A2(_1044_),
    .Y(_0402_),
    .B1(net47));
 sg13g2_o21ai_1 _2561_ (.B1(_0402_),
    .Y(_0403_),
    .A1(net30),
    .A2(_0400_));
 sg13g2_nand3_1 _2562_ (.B(net48),
    .C(_0403_),
    .A(_0398_),
    .Y(_0404_));
 sg13g2_a22oi_1 _2563_ (.Y(_0405_),
    .B1(_0889_),
    .B2(_0949_),
    .A2(net39),
    .A1(_1182_));
 sg13g2_nand2b_1 _2564_ (.Y(_0406_),
    .B(_0393_),
    .A_N(_1240_));
 sg13g2_a21oi_1 _2565_ (.A1(_0406_),
    .A2(net37),
    .Y(_0407_),
    .B1(net32));
 sg13g2_nand3_1 _2566_ (.B(_0953_),
    .C(_0407_),
    .A(_0405_),
    .Y(_0408_));
 sg13g2_nor2_1 _2567_ (.A(_1316_),
    .B(_1363_),
    .Y(_0409_));
 sg13g2_o21ai_1 _2568_ (.B1(_0409_),
    .Y(_0410_),
    .A1(_0903_),
    .A2(_1190_));
 sg13g2_nand3_1 _2569_ (.B(net43),
    .C(_0410_),
    .A(_0408_),
    .Y(_0411_));
 sg13g2_nand3_1 _2570_ (.B(net49),
    .C(_0411_),
    .A(_0404_),
    .Y(_0412_));
 sg13g2_o21ai_1 _2571_ (.B1(net31),
    .Y(_0413_),
    .A1(_1350_),
    .A2(_1450_));
 sg13g2_a21oi_1 _2572_ (.A1(_0861_),
    .A2(_0865_),
    .Y(_0414_),
    .B1(_1441_));
 sg13g2_a221oi_1 _2573_ (.B2(net47),
    .C1(net43),
    .B1(_0414_),
    .A1(_0413_),
    .Y(_0415_),
    .A2(_1362_));
 sg13g2_nor2_1 _2574_ (.A(net49),
    .B(_0415_),
    .Y(_0416_));
 sg13g2_nor2_1 _2575_ (.A(net40),
    .B(_1081_),
    .Y(_0417_));
 sg13g2_o21ai_1 _2576_ (.B1(_0395_),
    .Y(_0418_),
    .A1(_1213_),
    .A2(_0417_));
 sg13g2_o21ai_1 _2577_ (.B1(_1227_),
    .Y(_0419_),
    .A1(net37),
    .A2(_1242_));
 sg13g2_nor2_1 _2578_ (.A(_1348_),
    .B(_1331_),
    .Y(_0420_));
 sg13g2_a21oi_1 _2579_ (.A1(_0419_),
    .A2(_0420_),
    .Y(_0421_),
    .B1(net48));
 sg13g2_o21ai_1 _2580_ (.B1(_0421_),
    .Y(_0422_),
    .A1(net47),
    .A2(_0418_));
 sg13g2_a21oi_1 _2581_ (.A1(_0416_),
    .A2(_0422_),
    .Y(_0423_),
    .B1(net41));
 sg13g2_nand2_1 _2582_ (.Y(_0424_),
    .A(_0412_),
    .B(_0423_));
 sg13g2_nand2_1 _2583_ (.Y(_0425_),
    .A(net41),
    .B(net9));
 sg13g2_nand2_1 _2584_ (.Y(_0426_),
    .A(_0424_),
    .B(_0425_));
 sg13g2_nand2_1 _2585_ (.Y(_0427_),
    .A(_1013_),
    .B(\DJ8.GH[7] ));
 sg13g2_o21ai_1 _2586_ (.B1(_0427_),
    .Y(_0428_),
    .A1(_0980_),
    .A2(_1010_));
 sg13g2_a221oi_1 _2587_ (.B2(_1007_),
    .C1(_0428_),
    .B1(\DJ8.EF[7] ),
    .A1(\DJ8.EF[15] ),
    .Y(_0429_),
    .A2(_1004_));
 sg13g2_nand2_1 _2588_ (.Y(_0430_),
    .A(_1018_),
    .B(\DJ8.REGS.regs[1][7] ));
 sg13g2_a22oi_1 _2589_ (.Y(_0431_),
    .B1(\DJ8.REGS.regs[2][7] ),
    .B2(_1022_),
    .A2(_1020_),
    .A1(\DJ8.REGS.regs[3][7] ));
 sg13g2_nand2_1 _2590_ (.Y(_0432_),
    .A(net69),
    .B(\DJ8.ACC[7] ));
 sg13g2_nand4_1 _2591_ (.B(_0430_),
    .C(_0431_),
    .A(_0429_),
    .Y(_0433_),
    .D(_0432_));
 sg13g2_nor2b_1 _2592_ (.A(net79),
    .B_N(_0433_),
    .Y(_0434_));
 sg13g2_a21oi_2 _2593_ (.B1(_0434_),
    .Y(_0435_),
    .A2(net79),
    .A1(_0426_));
 sg13g2_nor2_1 _2594_ (.A(_0392_),
    .B(_0435_),
    .Y(_0436_));
 sg13g2_nand2_1 _2595_ (.Y(_0437_),
    .A(_0435_),
    .B(_0392_));
 sg13g2_inv_1 _2596_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nor2_1 _2597_ (.A(_0436_),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_nor3_1 _2598_ (.A(_0261_),
    .B(_0353_),
    .C(_0262_),
    .Y(_0440_));
 sg13g2_nand2_1 _2599_ (.Y(_0441_),
    .A(_0440_),
    .B(_1309_));
 sg13g2_o21ai_1 _2600_ (.B1(_0352_),
    .Y(_0442_),
    .A1(_0258_),
    .A2(_0353_));
 sg13g2_nor3_1 _2601_ (.A(_0261_),
    .B(_0353_),
    .C(_0264_),
    .Y(_0443_));
 sg13g2_nor2_1 _2602_ (.A(_0442_),
    .B(_0443_),
    .Y(_0444_));
 sg13g2_nand2_1 _2603_ (.Y(_0445_),
    .A(_0441_),
    .B(_0444_));
 sg13g2_xnor2_1 _2604_ (.Y(_0446_),
    .A(_0439_),
    .B(_0445_));
 sg13g2_inv_1 _2605_ (.Y(_0447_),
    .A(_0446_));
 sg13g2_nand2_1 _2606_ (.Y(_0448_),
    .A(_0389_),
    .B(_0447_));
 sg13g2_nand2_1 _2607_ (.Y(_0449_),
    .A(_0363_),
    .B(_0446_));
 sg13g2_nand3_1 _2608_ (.B(_0449_),
    .C(_1119_),
    .A(_0448_),
    .Y(_0450_));
 sg13g2_inv_1 _2609_ (.Y(_0451_),
    .A(_0435_));
 sg13g2_a221oi_1 _2610_ (.B2(_1127_),
    .C1(_1163_),
    .B1(_0451_),
    .A1(_1129_),
    .Y(_0452_),
    .A2(_0391_));
 sg13g2_nand2_1 _2611_ (.Y(_0453_),
    .A(_0439_),
    .B(_1136_));
 sg13g2_nand2_1 _2612_ (.Y(_0454_),
    .A(_0437_),
    .B(_1139_));
 sg13g2_nand2_1 _2613_ (.Y(_0455_),
    .A(_0436_),
    .B(_1123_));
 sg13g2_nand4_1 _2614_ (.B(_0453_),
    .C(_0454_),
    .A(_0452_),
    .Y(_0456_),
    .D(_0455_));
 sg13g2_nor3_1 _2615_ (.A(_0285_),
    .B(_0370_),
    .C(_0280_),
    .Y(_0457_));
 sg13g2_inv_1 _2616_ (.Y(_0458_),
    .A(_0283_));
 sg13g2_o21ai_1 _2617_ (.B1(_0369_),
    .Y(_0459_),
    .A1(_0368_),
    .A2(_0458_));
 sg13g2_nor2b_1 _2618_ (.A(_0457_),
    .B_N(_0459_),
    .Y(_0460_));
 sg13g2_nor2_1 _2619_ (.A(_0285_),
    .B(_0370_),
    .Y(_0461_));
 sg13g2_nand3_1 _2620_ (.B(_1402_),
    .C(_0276_),
    .A(_0461_),
    .Y(_0462_));
 sg13g2_nor2_1 _2621_ (.A(_0350_),
    .B(_0378_),
    .Y(_0463_));
 sg13g2_o21ai_1 _2622_ (.B1(_0463_),
    .Y(_0464_),
    .A1(_0436_),
    .A2(_0438_));
 sg13g2_nand2b_1 _2623_ (.Y(_0465_),
    .B(_0439_),
    .A_N(_0463_));
 sg13g2_nand2_1 _2624_ (.Y(_0466_),
    .A(_0464_),
    .B(_0465_));
 sg13g2_a21oi_1 _2625_ (.A1(_0460_),
    .A2(_0462_),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_nand3_1 _2626_ (.B(_0466_),
    .C(_0462_),
    .A(_0460_),
    .Y(_0468_));
 sg13g2_nand2_1 _2627_ (.Y(_0469_),
    .A(_0468_),
    .B(_1152_));
 sg13g2_nor2_1 _2628_ (.A(_0467_),
    .B(_0469_),
    .Y(_0470_));
 sg13g2_nor2_1 _2629_ (.A(_0456_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nand2_1 _2630_ (.Y(_0472_),
    .A(_0450_),
    .B(_0471_));
 sg13g2_nand2_1 _2631_ (.Y(_0473_),
    .A(_0446_),
    .B(net75));
 sg13g2_nand2_1 _2632_ (.Y(_0474_),
    .A(_0472_),
    .B(_0473_));
 sg13g2_nand2_1 _2633_ (.Y(_0475_),
    .A(_0474_),
    .B(_1162_));
 sg13g2_nand2_1 _2634_ (.Y(_0476_),
    .A(_0384_),
    .B(_1161_));
 sg13g2_nand2_1 _2635_ (.Y(_0477_),
    .A(_0475_),
    .B(_0476_));
 sg13g2_nor2_1 _2636_ (.A(\DJ8.ACC[6] ),
    .B(_0768_),
    .Y(_0478_));
 sg13g2_a21oi_1 _2637_ (.A1(net26),
    .A2(net66),
    .Y(_0044_),
    .B1(_0478_));
 sg13g2_nor2_1 _2638_ (.A(_1158_),
    .B(_0474_),
    .Y(_0479_));
 sg13g2_nor2_1 _2639_ (.A(_0026_),
    .B(_0768_),
    .Y(_0480_));
 sg13g2_a21oi_1 _2640_ (.A1(net27),
    .A2(net66),
    .Y(_0045_),
    .B1(_0480_));
 sg13g2_nor3_2 _2641_ (.A(_0760_),
    .B(_0995_),
    .C(_0767_),
    .Y(_0481_));
 sg13g2_mux2_1 _2642_ (.A0(\DJ8.REGS.regs[1][0] ),
    .A1(_1178_),
    .S(_0481_),
    .X(_0046_));
 sg13g2_buf_1 _2643_ (.A(_0481_),
    .X(_0482_));
 sg13g2_nor2_1 _2644_ (.A(\DJ8.REGS.regs[1][1] ),
    .B(net62),
    .Y(_0483_));
 sg13g2_a21oi_1 _2645_ (.A1(_1305_),
    .A2(net62),
    .Y(_0047_),
    .B1(_0483_));
 sg13g2_mux2_1 _2646_ (.A0(\DJ8.REGS.regs[1][2] ),
    .A1(_1419_),
    .S(_0481_),
    .X(_0048_));
 sg13g2_nor2_1 _2647_ (.A(\DJ8.REGS.regs[1][3] ),
    .B(_0482_),
    .Y(_0484_));
 sg13g2_a21oi_1 _2648_ (.A1(_0181_),
    .A2(_0482_),
    .Y(_0049_),
    .B1(_0484_));
 sg13g2_nor2_1 _2649_ (.A(\DJ8.REGS.regs[1][4] ),
    .B(net62),
    .Y(_0485_));
 sg13g2_a21oi_1 _2650_ (.A1(net29),
    .A2(net62),
    .Y(_0050_),
    .B1(_0485_));
 sg13g2_nor2_1 _2651_ (.A(\DJ8.REGS.regs[1][5] ),
    .B(net62),
    .Y(_0486_));
 sg13g2_a21oi_1 _2652_ (.A1(net28),
    .A2(net62),
    .Y(_0051_),
    .B1(_0486_));
 sg13g2_nor2_1 _2653_ (.A(\DJ8.REGS.regs[1][6] ),
    .B(_0481_),
    .Y(_0487_));
 sg13g2_a21oi_1 _2654_ (.A1(_0477_),
    .A2(net62),
    .Y(_0052_),
    .B1(_0487_));
 sg13g2_nor2_1 _2655_ (.A(_0027_),
    .B(_0481_),
    .Y(_0488_));
 sg13g2_a21oi_1 _2656_ (.A1(net27),
    .A2(net62),
    .Y(_0053_),
    .B1(_0488_));
 sg13g2_inv_2 _2657_ (.Y(_0489_),
    .A(_0760_));
 sg13g2_nor3_2 _2658_ (.A(_0489_),
    .B(_0761_),
    .C(_0767_),
    .Y(_0490_));
 sg13g2_mux2_1 _2659_ (.A0(\DJ8.REGS.regs[2][0] ),
    .A1(_1178_),
    .S(_0490_),
    .X(_0054_));
 sg13g2_buf_1 _2660_ (.A(_0490_),
    .X(_0491_));
 sg13g2_nor2_1 _2661_ (.A(\DJ8.REGS.regs[2][1] ),
    .B(net61),
    .Y(_0492_));
 sg13g2_a21oi_1 _2662_ (.A1(_1305_),
    .A2(net61),
    .Y(_0055_),
    .B1(_0492_));
 sg13g2_mux2_1 _2663_ (.A0(\DJ8.REGS.regs[2][2] ),
    .A1(_1419_),
    .S(_0490_),
    .X(_0056_));
 sg13g2_nor2_1 _2664_ (.A(\DJ8.REGS.regs[2][3] ),
    .B(net61),
    .Y(_0493_));
 sg13g2_a21oi_1 _2665_ (.A1(_0181_),
    .A2(net61),
    .Y(_0057_),
    .B1(_0493_));
 sg13g2_nor2_1 _2666_ (.A(\DJ8.REGS.regs[2][4] ),
    .B(net61),
    .Y(_0494_));
 sg13g2_a21oi_1 _2667_ (.A1(net29),
    .A2(net61),
    .Y(_0058_),
    .B1(_0494_));
 sg13g2_nor2_1 _2668_ (.A(\DJ8.REGS.regs[2][5] ),
    .B(net61),
    .Y(_0495_));
 sg13g2_a21oi_1 _2669_ (.A1(net28),
    .A2(net61),
    .Y(_0059_),
    .B1(_0495_));
 sg13g2_nor2_1 _2670_ (.A(\DJ8.REGS.regs[2][6] ),
    .B(_0490_),
    .Y(_0496_));
 sg13g2_a21oi_1 _2671_ (.A1(net26),
    .A2(_0491_),
    .Y(_0060_),
    .B1(_0496_));
 sg13g2_nor2_1 _2672_ (.A(_0028_),
    .B(_0490_),
    .Y(_0497_));
 sg13g2_a21oi_1 _2673_ (.A1(net27),
    .A2(_0491_),
    .Y(_0061_),
    .B1(_0497_));
 sg13g2_nor3_2 _2674_ (.A(_0489_),
    .B(_0995_),
    .C(_0767_),
    .Y(_0498_));
 sg13g2_mux2_1 _2675_ (.A0(\DJ8.REGS.regs[3][0] ),
    .A1(_1178_),
    .S(_0498_),
    .X(_0062_));
 sg13g2_buf_1 _2676_ (.A(_0498_),
    .X(_0499_));
 sg13g2_nor2_1 _2677_ (.A(\DJ8.REGS.regs[3][1] ),
    .B(net60),
    .Y(_0500_));
 sg13g2_a21oi_1 _2678_ (.A1(_1305_),
    .A2(net60),
    .Y(_0063_),
    .B1(_0500_));
 sg13g2_mux2_1 _2679_ (.A0(\DJ8.REGS.regs[3][2] ),
    .A1(_1419_),
    .S(_0498_),
    .X(_0064_));
 sg13g2_nor2_1 _2680_ (.A(\DJ8.REGS.regs[3][3] ),
    .B(_0499_),
    .Y(_0501_));
 sg13g2_a21oi_1 _2681_ (.A1(_0181_),
    .A2(net60),
    .Y(_0065_),
    .B1(_0501_));
 sg13g2_nor2_1 _2682_ (.A(\DJ8.REGS.regs[3][4] ),
    .B(net60),
    .Y(_0502_));
 sg13g2_a21oi_1 _2683_ (.A1(net29),
    .A2(net60),
    .Y(_0066_),
    .B1(_0502_));
 sg13g2_nor2_1 _2684_ (.A(\DJ8.REGS.regs[3][5] ),
    .B(net60),
    .Y(_0503_));
 sg13g2_a21oi_1 _2685_ (.A1(net28),
    .A2(net60),
    .Y(_0067_),
    .B1(_0503_));
 sg13g2_nor2_1 _2686_ (.A(\DJ8.REGS.regs[3][6] ),
    .B(_0498_),
    .Y(_0504_));
 sg13g2_a21oi_1 _2687_ (.A1(net26),
    .A2(net60),
    .Y(_0068_),
    .B1(_0504_));
 sg13g2_nor2_1 _2688_ (.A(_0029_),
    .B(_0498_),
    .Y(_0505_));
 sg13g2_a21oi_1 _2689_ (.A1(net27),
    .A2(_0499_),
    .Y(_0069_),
    .B1(_0505_));
 sg13g2_nor2_1 _2690_ (.A(_0001_),
    .B(_0765_),
    .Y(_0506_));
 sg13g2_inv_2 _2691_ (.Y(_0507_),
    .A(_0506_));
 sg13g2_nor3_2 _2692_ (.A(_0760_),
    .B(_0761_),
    .C(_0507_),
    .Y(_0508_));
 sg13g2_mux2_1 _2693_ (.A0(\DJ8.EF[8] ),
    .A1(_1178_),
    .S(_0508_),
    .X(_0070_));
 sg13g2_buf_1 _2694_ (.A(_0508_),
    .X(_0509_));
 sg13g2_nor2_1 _2695_ (.A(\DJ8.EF[9] ),
    .B(net59),
    .Y(_0510_));
 sg13g2_a21oi_1 _2696_ (.A1(_1305_),
    .A2(net59),
    .Y(_0071_),
    .B1(_0510_));
 sg13g2_nand2_1 _2697_ (.Y(_0511_),
    .A(_1419_),
    .B(_0508_));
 sg13g2_o21ai_1 _2698_ (.B1(_0511_),
    .Y(_0072_),
    .A1(_1252_),
    .A2(net59));
 sg13g2_nor2_1 _2699_ (.A(\DJ8.EF[11] ),
    .B(_0509_),
    .Y(_0512_));
 sg13g2_a21oi_1 _2700_ (.A1(_0181_),
    .A2(_0509_),
    .Y(_0073_),
    .B1(_0512_));
 sg13g2_nor2_1 _2701_ (.A(\DJ8.EF[12] ),
    .B(net59),
    .Y(_0513_));
 sg13g2_a21oi_1 _2702_ (.A1(net29),
    .A2(net59),
    .Y(_0074_),
    .B1(_0513_));
 sg13g2_nor2_1 _2703_ (.A(\DJ8.EF[13] ),
    .B(_0508_),
    .Y(_0514_));
 sg13g2_a21oi_1 _2704_ (.A1(net28),
    .A2(net59),
    .Y(_0075_),
    .B1(_0514_));
 sg13g2_nor2_1 _2705_ (.A(\DJ8.EF[14] ),
    .B(_0508_),
    .Y(_0515_));
 sg13g2_a21oi_1 _2706_ (.A1(net26),
    .A2(net59),
    .Y(_0076_),
    .B1(_0515_));
 sg13g2_nor2_1 _2707_ (.A(_0030_),
    .B(_0508_),
    .Y(_0516_));
 sg13g2_a21oi_1 _2708_ (.A1(net27),
    .A2(net59),
    .Y(_0077_),
    .B1(_0516_));
 sg13g2_nor3_2 _2709_ (.A(_0760_),
    .B(_0995_),
    .C(_0507_),
    .Y(_0517_));
 sg13g2_inv_1 _2710_ (.Y(_0518_),
    .A(_0517_));
 sg13g2_nor2_1 _2711_ (.A(_0518_),
    .B(_1178_),
    .Y(_0519_));
 sg13g2_a21oi_1 _2712_ (.A1(_0812_),
    .A2(_0518_),
    .Y(_0078_),
    .B1(_0519_));
 sg13g2_buf_1 _2713_ (.A(_0517_),
    .X(_0520_));
 sg13g2_nor2_1 _2714_ (.A(\DJ8.EF[1] ),
    .B(net58),
    .Y(_0521_));
 sg13g2_a21oi_1 _2715_ (.A1(_1305_),
    .A2(net58),
    .Y(_0079_),
    .B1(_0521_));
 sg13g2_nor2_1 _2716_ (.A(_0518_),
    .B(_1419_),
    .Y(_0522_));
 sg13g2_a21oi_1 _2717_ (.A1(_1256_),
    .A2(_0518_),
    .Y(_0080_),
    .B1(_0522_));
 sg13g2_nor2_1 _2718_ (.A(\DJ8.EF[3] ),
    .B(net58),
    .Y(_0523_));
 sg13g2_a21oi_1 _2719_ (.A1(_0181_),
    .A2(net58),
    .Y(_0081_),
    .B1(_0523_));
 sg13g2_nor2_1 _2720_ (.A(\DJ8.EF[4] ),
    .B(net58),
    .Y(_0524_));
 sg13g2_a21oi_1 _2721_ (.A1(net29),
    .A2(net58),
    .Y(_0082_),
    .B1(_0524_));
 sg13g2_nor2_1 _2722_ (.A(\DJ8.EF[5] ),
    .B(net58),
    .Y(_0525_));
 sg13g2_a21oi_1 _2723_ (.A1(net28),
    .A2(net58),
    .Y(_0083_),
    .B1(_0525_));
 sg13g2_nor2_1 _2724_ (.A(\DJ8.EF[6] ),
    .B(_0517_),
    .Y(_0526_));
 sg13g2_a21oi_1 _2725_ (.A1(net26),
    .A2(_0520_),
    .Y(_0084_),
    .B1(_0526_));
 sg13g2_nor2_1 _2726_ (.A(_0031_),
    .B(_0517_),
    .Y(_0527_));
 sg13g2_a21oi_1 _2727_ (.A1(net27),
    .A2(_0520_),
    .Y(_0085_),
    .B1(_0527_));
 sg13g2_nor3_2 _2728_ (.A(_0489_),
    .B(_0761_),
    .C(_0507_),
    .Y(_0528_));
 sg13g2_inv_1 _2729_ (.Y(_0529_),
    .A(_0528_));
 sg13g2_nor2_1 _2730_ (.A(_0529_),
    .B(_1178_),
    .Y(_0530_));
 sg13g2_a21oi_1 _2731_ (.A1(_1008_),
    .A2(_0529_),
    .Y(_0086_),
    .B1(_0530_));
 sg13g2_buf_1 _2732_ (.A(_0528_),
    .X(_0531_));
 sg13g2_nor2_1 _2733_ (.A(\DJ8.GH[9] ),
    .B(net57),
    .Y(_0532_));
 sg13g2_a21oi_1 _2734_ (.A1(_1305_),
    .A2(net57),
    .Y(_0087_),
    .B1(_0532_));
 sg13g2_nor2_1 _2735_ (.A(_0529_),
    .B(_1419_),
    .Y(_0533_));
 sg13g2_a21oi_1 _2736_ (.A1(_1254_),
    .A2(_0529_),
    .Y(_0088_),
    .B1(_0533_));
 sg13g2_nor2_1 _2737_ (.A(\DJ8.GH[11] ),
    .B(net57),
    .Y(_0534_));
 sg13g2_a21oi_1 _2738_ (.A1(_0181_),
    .A2(net57),
    .Y(_0089_),
    .B1(_0534_));
 sg13g2_nor2_1 _2739_ (.A(\DJ8.GH[12] ),
    .B(net57),
    .Y(_0535_));
 sg13g2_a21oi_1 _2740_ (.A1(net29),
    .A2(net57),
    .Y(_0090_),
    .B1(_0535_));
 sg13g2_nor2_1 _2741_ (.A(\DJ8.GH[13] ),
    .B(_0531_),
    .Y(_0536_));
 sg13g2_a21oi_1 _2742_ (.A1(net28),
    .A2(_0531_),
    .Y(_0091_),
    .B1(_0536_));
 sg13g2_nor2_1 _2743_ (.A(\DJ8.GH[14] ),
    .B(_0528_),
    .Y(_0537_));
 sg13g2_a21oi_1 _2744_ (.A1(net26),
    .A2(net57),
    .Y(_0092_),
    .B1(_0537_));
 sg13g2_nor2_1 _2745_ (.A(_0032_),
    .B(_0528_),
    .Y(_0538_));
 sg13g2_a21oi_1 _2746_ (.A1(net27),
    .A2(net57),
    .Y(_0093_),
    .B1(_0538_));
 sg13g2_nor3_2 _2747_ (.A(_0489_),
    .B(_0995_),
    .C(_0507_),
    .Y(_0539_));
 sg13g2_inv_1 _2748_ (.Y(_0540_),
    .A(_0539_));
 sg13g2_nor2_1 _2749_ (.A(_0540_),
    .B(_1178_),
    .Y(_0541_));
 sg13g2_a21oi_1 _2750_ (.A1(_0810_),
    .A2(_0540_),
    .Y(_0094_),
    .B1(_0541_));
 sg13g2_buf_1 _2751_ (.A(_0539_),
    .X(_0542_));
 sg13g2_nor2_1 _2752_ (.A(\DJ8.GH[1] ),
    .B(net56),
    .Y(_0543_));
 sg13g2_a21oi_1 _2753_ (.A1(_1305_),
    .A2(net56),
    .Y(_0095_),
    .B1(_0543_));
 sg13g2_nor2_1 _2754_ (.A(_0540_),
    .B(_1419_),
    .Y(_0544_));
 sg13g2_a21oi_1 _2755_ (.A1(_1258_),
    .A2(_0540_),
    .Y(_0096_),
    .B1(_0544_));
 sg13g2_nor2_1 _2756_ (.A(\DJ8.GH[3] ),
    .B(net56),
    .Y(_0545_));
 sg13g2_a21oi_1 _2757_ (.A1(_0181_),
    .A2(net56),
    .Y(_0097_),
    .B1(_0545_));
 sg13g2_nor2_1 _2758_ (.A(\DJ8.GH[4] ),
    .B(_0542_),
    .Y(_0546_));
 sg13g2_a21oi_1 _2759_ (.A1(net29),
    .A2(_0542_),
    .Y(_0098_),
    .B1(_0546_));
 sg13g2_nor2_1 _2760_ (.A(\DJ8.GH[5] ),
    .B(net56),
    .Y(_0547_));
 sg13g2_a21oi_1 _2761_ (.A1(net28),
    .A2(net56),
    .Y(_0099_),
    .B1(_0547_));
 sg13g2_nor2_1 _2762_ (.A(\DJ8.GH[6] ),
    .B(_0539_),
    .Y(_0548_));
 sg13g2_a21oi_1 _2763_ (.A1(net26),
    .A2(net56),
    .Y(_0100_),
    .B1(_0548_));
 sg13g2_nor2_1 _2764_ (.A(_0033_),
    .B(_0539_),
    .Y(_0549_));
 sg13g2_a21oi_1 _2765_ (.A1(net27),
    .A2(net56),
    .Y(_0101_),
    .B1(_0549_));
 sg13g2_inv_1 _2766_ (.Y(_0550_),
    .A(_0763_));
 sg13g2_nand3b_1 _2767_ (.B(_0372_),
    .C(_0465_),
    .Y(_0551_),
    .A_N(_0368_));
 sg13g2_nand2_1 _2768_ (.Y(_0552_),
    .A(_0435_),
    .B(_0391_));
 sg13g2_nand3_1 _2769_ (.B(_0464_),
    .C(_0552_),
    .A(_0551_),
    .Y(_0553_));
 sg13g2_nand2_1 _2770_ (.Y(_0554_),
    .A(_0553_),
    .B(_1152_));
 sg13g2_nand2_1 _2771_ (.Y(_0555_),
    .A(_0359_),
    .B(_0376_));
 sg13g2_nor2b_1 _2772_ (.A(_0436_),
    .B_N(_0352_),
    .Y(_0556_));
 sg13g2_a21oi_1 _2773_ (.A1(_0555_),
    .A2(_0556_),
    .Y(_0557_),
    .B1(_0438_));
 sg13g2_inv_1 _2774_ (.Y(_0558_),
    .A(_0448_));
 sg13g2_o21ai_1 _2775_ (.B1(_1119_),
    .Y(_0559_),
    .A1(_0557_),
    .A2(_0558_));
 sg13g2_nand2_1 _2776_ (.Y(_0560_),
    .A(_0557_),
    .B(net75));
 sg13g2_nand3_1 _2777_ (.B(_0559_),
    .C(_0560_),
    .A(_0554_),
    .Y(_0561_));
 sg13g2_nand2_1 _2778_ (.Y(_0562_),
    .A(_0561_),
    .B(_0550_));
 sg13g2_o21ai_1 _2779_ (.B1(_0562_),
    .Y(_0102_),
    .A1(_1143_),
    .A2(_0550_));
 sg13g2_nand3_1 _2780_ (.B(_1177_),
    .C(_0550_),
    .A(_1165_),
    .Y(_0563_));
 sg13g2_nor2_1 _2781_ (.A(_0563_),
    .B(_1304_),
    .Y(_0564_));
 sg13g2_nand3_1 _2782_ (.B(_1417_),
    .C(_1418_),
    .A(_0564_),
    .Y(_0565_));
 sg13g2_nor2_1 _2783_ (.A(_0180_),
    .B(_0565_),
    .Y(_0566_));
 sg13g2_nand2_1 _2784_ (.Y(_0567_),
    .A(_0300_),
    .B(_0566_));
 sg13g2_nor2_1 _2785_ (.A(_0479_),
    .B(_0567_),
    .Y(_0568_));
 sg13g2_nand3_1 _2786_ (.B(_0387_),
    .C(net26),
    .A(_0568_),
    .Y(_0569_));
 sg13g2_nand2_1 _2787_ (.Y(_0570_),
    .A(_0763_),
    .B(\DJ8.flag_Z ));
 sg13g2_nand2_1 _2788_ (.Y(_0103_),
    .A(_0569_),
    .B(_0570_));
 sg13g2_and2_1 _2789_ (.A(_0985_),
    .B(_0990_),
    .X(_0571_));
 sg13g2_nor2_1 _2790_ (.A(_0752_),
    .B(net88),
    .Y(_0572_));
 sg13g2_a21oi_1 _2791_ (.A1(_0571_),
    .A2(net88),
    .Y(_0104_),
    .B1(_0572_));
 sg13g2_inv_1 _2792_ (.Y(_0573_),
    .A(\DJ8.REGS.write_addr[2] ));
 sg13g2_buf_1 _2793_ (.A(_0795_),
    .X(_0574_));
 sg13g2_nand2_1 _2794_ (.Y(_0575_),
    .A(_1249_),
    .B(_1250_));
 sg13g2_nor2_1 _2795_ (.A(net82),
    .B(_0575_),
    .Y(_0576_));
 sg13g2_a21oi_1 _2796_ (.A1(_0573_),
    .A2(net82),
    .Y(_0105_),
    .B1(_0576_));
 sg13g2_nor2_1 _2797_ (.A(_0574_),
    .B(_1404_),
    .Y(_0577_));
 sg13g2_a21oi_1 _2798_ (.A1(_0574_),
    .A2(_1117_),
    .Y(_0106_),
    .B1(_0577_));
 sg13g2_a22oi_1 _2799_ (.Y(_0578_),
    .B1(_1478_),
    .B2(_1458_),
    .A2(_1373_),
    .A1(net6));
 sg13g2_nor2_1 _2800_ (.A(_1115_),
    .B(net86),
    .Y(_0579_));
 sg13g2_a21oi_1 _2801_ (.A1(_0578_),
    .A2(net86),
    .Y(_0107_),
    .B1(_0579_));
 sg13g2_nand2_1 _2802_ (.Y(_0580_),
    .A(_0242_),
    .B(_0243_));
 sg13g2_nor2_1 _2803_ (.A(\DJ8.ALU.opalu[2] ),
    .B(net86),
    .Y(_0581_));
 sg13g2_a21oi_1 _2804_ (.A1(_0580_),
    .A2(net86),
    .Y(_0108_),
    .B1(_0581_));
 sg13g2_nand2_1 _2805_ (.Y(_0582_),
    .A(_0334_),
    .B(_0335_));
 sg13g2_nor2_1 _2806_ (.A(net82),
    .B(_0582_),
    .Y(_0583_));
 sg13g2_a21oi_1 _2807_ (.A1(_0755_),
    .A2(net82),
    .Y(_0109_),
    .B1(_0583_));
 sg13g2_nor2_1 _2808_ (.A(net82),
    .B(_0426_),
    .Y(_0584_));
 sg13g2_a21oi_1 _2809_ (.A1(_0787_),
    .A2(net82),
    .Y(_0110_),
    .B1(_0584_));
 sg13g2_inv_2 _2810_ (.Y(_0585_),
    .A(net88));
 sg13g2_nand2_1 _2811_ (.Y(_0586_),
    .A(_1091_),
    .B(_1093_));
 sg13g2_nor2_1 _2812_ (.A(_0585_),
    .B(_0586_),
    .Y(_0587_));
 sg13g2_a21oi_1 _2813_ (.A1(_0987_),
    .A2(_0585_),
    .Y(_0111_),
    .B1(_0587_));
 sg13g2_nor2_1 _2814_ (.A(_0585_),
    .B(_0575_),
    .Y(_0588_));
 sg13g2_a21oi_1 _2815_ (.A1(_0585_),
    .A2(_1157_),
    .Y(_0112_),
    .B1(_0588_));
 sg13g2_nor2_1 _2816_ (.A(_0585_),
    .B(_1404_),
    .Y(_0589_));
 sg13g2_a21oi_1 _2817_ (.A1(_0585_),
    .A2(_1159_),
    .Y(_0113_),
    .B1(_0589_));
 sg13g2_buf_1 _2818_ (.A(net84),
    .X(_0590_));
 sg13g2_nor2_1 _2819_ (.A(net78),
    .B(net88),
    .Y(_0591_));
 sg13g2_a21oi_1 _2820_ (.A1(_0578_),
    .A2(net88),
    .Y(_0114_),
    .B1(_0591_));
 sg13g2_nor2_1 _2821_ (.A(\DJ8.ir[5] ),
    .B(net88),
    .Y(_0592_));
 sg13g2_a21oi_1 _2822_ (.A1(_0580_),
    .A2(_0772_),
    .Y(_0115_),
    .B1(_0592_));
 sg13g2_nor2_1 _2823_ (.A(_0585_),
    .B(_0582_),
    .Y(_0593_));
 sg13g2_a21oi_1 _2824_ (.A1(_0992_),
    .A2(_0585_),
    .Y(_0116_),
    .B1(_0593_));
 sg13g2_mux2_1 _2825_ (.A0(\DJ8.ir[7] ),
    .A1(_0426_),
    .S(net88),
    .X(_0117_));
 sg13g2_nor2_1 _2826_ (.A(_0761_),
    .B(_0798_),
    .Y(_0594_));
 sg13g2_a21oi_1 _2827_ (.A1(_0571_),
    .A2(_0798_),
    .Y(_0118_),
    .B1(_0594_));
 sg13g2_nor2_1 _2828_ (.A(net82),
    .B(_0586_),
    .Y(_0595_));
 sg13g2_a21oi_1 _2829_ (.A1(_0489_),
    .A2(net82),
    .Y(_0119_),
    .B1(_0595_));
 sg13g2_inv_1 _2830_ (.Y(_0596_),
    .A(_0762_));
 sg13g2_buf_1 _2831_ (.A(_0596_),
    .X(_0597_));
 sg13g2_inv_1 _2832_ (.Y(_0598_),
    .A(\DJ8.pc[0] ));
 sg13g2_nor2_1 _2833_ (.A(\DJ8.ALU.opalu[2] ),
    .B(\DJ8.flag_Z ),
    .Y(_0599_));
 sg13g2_nand2_1 _2834_ (.Y(_0600_),
    .A(_1122_),
    .B(\DJ8.flag_Z ));
 sg13g2_nand3_1 _2835_ (.B(_0787_),
    .C(_0755_),
    .A(_0600_),
    .Y(_0601_));
 sg13g2_nor2_1 _2836_ (.A(_0599_),
    .B(_0601_),
    .Y(_0602_));
 sg13g2_buf_1 _2837_ (.A(_0602_),
    .X(_0603_));
 sg13g2_buf_1 _2838_ (.A(net73),
    .X(_0604_));
 sg13g2_nand2_1 _2839_ (.Y(_0605_),
    .A(net68),
    .B(_0752_));
 sg13g2_inv_1 _2840_ (.Y(_0606_),
    .A(_0602_));
 sg13g2_nor2_2 _2841_ (.A(\DJ8.ir[15] ),
    .B(_0755_),
    .Y(_0607_));
 sg13g2_inv_2 _2842_ (.Y(_0608_),
    .A(_0607_));
 sg13g2_nand2_1 _2843_ (.Y(_0609_),
    .A(_0608_),
    .B(_0006_));
 sg13g2_buf_1 _2844_ (.A(_0607_),
    .X(_0610_));
 sg13g2_nand2_1 _2845_ (.Y(_0611_),
    .A(_0610_),
    .B(\DJ8.GH[1] ));
 sg13g2_nand2_1 _2846_ (.Y(_0612_),
    .A(_0609_),
    .B(_0611_));
 sg13g2_a21oi_1 _2847_ (.A1(_0606_),
    .A2(_0612_),
    .Y(_0613_),
    .B1(net81));
 sg13g2_a22oi_1 _2848_ (.Y(_0120_),
    .B1(_0605_),
    .B2(_0613_),
    .A2(_0598_),
    .A1(net81));
 sg13g2_inv_1 _2849_ (.Y(_0614_),
    .A(\DJ8.pc[10] ));
 sg13g2_inv_1 _2850_ (.Y(_0615_),
    .A(\DJ8.pc[8] ));
 sg13g2_inv_1 _2851_ (.Y(_0616_),
    .A(\DJ8.pc[9] ));
 sg13g2_inv_1 _2852_ (.Y(_0617_),
    .A(\DJ8.pc[7] ));
 sg13g2_inv_1 _2853_ (.Y(_0618_),
    .A(\DJ8.pc[6] ));
 sg13g2_inv_1 _2854_ (.Y(_0619_),
    .A(\DJ8.pc[4] ));
 sg13g2_inv_1 _2855_ (.Y(_0620_),
    .A(\DJ8.pc[3] ));
 sg13g2_inv_1 _2856_ (.Y(_0621_),
    .A(\DJ8.pc[2] ));
 sg13g2_nand2_1 _2857_ (.Y(_0622_),
    .A(\DJ8.pc[1] ),
    .B(\DJ8.pc[0] ));
 sg13g2_nor2_1 _2858_ (.A(_0621_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_inv_1 _2859_ (.Y(_0624_),
    .A(_0623_));
 sg13g2_nor2_1 _2860_ (.A(_0620_),
    .B(_0624_),
    .Y(_0625_));
 sg13g2_inv_1 _2861_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_nor2_1 _2862_ (.A(_0619_),
    .B(_0626_),
    .Y(_0627_));
 sg13g2_nand2_1 _2863_ (.Y(_0628_),
    .A(_0627_),
    .B(\DJ8.pc[5] ));
 sg13g2_nor2_1 _2864_ (.A(_0618_),
    .B(_0628_),
    .Y(_0629_));
 sg13g2_inv_1 _2865_ (.Y(_0630_),
    .A(_0629_));
 sg13g2_nor2_1 _2866_ (.A(_0617_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_inv_1 _2867_ (.Y(_0632_),
    .A(_0631_));
 sg13g2_nor3_1 _2868_ (.A(_0615_),
    .B(_0616_),
    .C(_0632_),
    .Y(_0633_));
 sg13g2_inv_1 _2869_ (.Y(_0634_),
    .A(_0633_));
 sg13g2_a21oi_1 _2870_ (.A1(_0634_),
    .A2(_0614_),
    .Y(_0635_),
    .B1(_0607_));
 sg13g2_nor2_1 _2871_ (.A(_0614_),
    .B(_0634_),
    .Y(_0636_));
 sg13g2_inv_1 _2872_ (.Y(_0637_),
    .A(_0636_));
 sg13g2_nand2_1 _2873_ (.Y(_0638_),
    .A(_0635_),
    .B(_0637_));
 sg13g2_nand2_1 _2874_ (.Y(_0639_),
    .A(net77),
    .B(\DJ8.GH[11] ));
 sg13g2_nand3_1 _2875_ (.B(_0606_),
    .C(_0639_),
    .A(_0638_),
    .Y(_0640_));
 sg13g2_buf_1 _2876_ (.A(_0596_),
    .X(_0641_));
 sg13g2_a21oi_1 _2877_ (.A1(net73),
    .A2(_0573_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_nand2_1 _2878_ (.Y(_0643_),
    .A(_0640_),
    .B(_0642_));
 sg13g2_o21ai_1 _2879_ (.B1(_0643_),
    .Y(_0121_),
    .A1(_0762_),
    .A2(_0614_));
 sg13g2_inv_1 _2880_ (.Y(_0644_),
    .A(\DJ8.pc[11] ));
 sg13g2_a21oi_1 _2881_ (.A1(_0637_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(_0607_));
 sg13g2_nor2_1 _2882_ (.A(_0644_),
    .B(_0637_),
    .Y(_0646_));
 sg13g2_inv_1 _2883_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_nand2_1 _2884_ (.Y(_0648_),
    .A(_0645_),
    .B(_0647_));
 sg13g2_nand2_1 _2885_ (.Y(_0649_),
    .A(net77),
    .B(\DJ8.GH[12] ));
 sg13g2_nand3_1 _2886_ (.B(_0606_),
    .C(_0649_),
    .A(_0648_),
    .Y(_0650_));
 sg13g2_a21oi_1 _2887_ (.A1(_0603_),
    .A2(_1117_),
    .Y(_0651_),
    .B1(_0641_));
 sg13g2_nand2_1 _2888_ (.Y(_0652_),
    .A(_0650_),
    .B(_0651_));
 sg13g2_o21ai_1 _2889_ (.B1(_0652_),
    .Y(_0122_),
    .A1(_0762_),
    .A2(_0644_));
 sg13g2_inv_1 _2890_ (.Y(_0653_),
    .A(\DJ8.pc[12] ));
 sg13g2_nor2_1 _2891_ (.A(_0596_),
    .B(_0602_),
    .Y(_0654_));
 sg13g2_inv_1 _2892_ (.Y(_0655_),
    .A(_0654_));
 sg13g2_buf_1 _2893_ (.A(_0607_),
    .X(_0656_));
 sg13g2_a21oi_1 _2894_ (.A1(\DJ8.GH[13] ),
    .A2(net76),
    .Y(_0657_),
    .B1(_0655_));
 sg13g2_nor2_1 _2895_ (.A(_0653_),
    .B(_0647_),
    .Y(_0658_));
 sg13g2_inv_1 _2896_ (.Y(_0659_),
    .A(_0658_));
 sg13g2_nand2_1 _2897_ (.Y(_0660_),
    .A(_0647_),
    .B(_0653_));
 sg13g2_nand3_1 _2898_ (.B(_0608_),
    .C(_0660_),
    .A(_0659_),
    .Y(_0661_));
 sg13g2_a22oi_1 _2899_ (.Y(_0123_),
    .B1(_0657_),
    .B2(_0661_),
    .A2(_0655_),
    .A1(_0653_));
 sg13g2_inv_1 _2900_ (.Y(_0662_),
    .A(_0034_));
 sg13g2_inv_1 _2901_ (.Y(_0663_),
    .A(\DJ8.pc[13] ));
 sg13g2_nand2_1 _2902_ (.Y(_0664_),
    .A(_0659_),
    .B(_0663_));
 sg13g2_nand2_1 _2903_ (.Y(_0665_),
    .A(_0658_),
    .B(\DJ8.pc[13] ));
 sg13g2_nand3_1 _2904_ (.B(_0608_),
    .C(_0665_),
    .A(_0664_),
    .Y(_0666_));
 sg13g2_nand2_1 _2905_ (.Y(_0667_),
    .A(net76),
    .B(\DJ8.GH[14] ));
 sg13g2_nand3_1 _2906_ (.B(_0654_),
    .C(_0667_),
    .A(_0666_),
    .Y(_0668_));
 sg13g2_o21ai_1 _2907_ (.B1(_0668_),
    .Y(_0124_),
    .A1(_0662_),
    .A2(_0654_));
 sg13g2_inv_1 _2908_ (.Y(_0669_),
    .A(\DJ8.pc[14] ));
 sg13g2_a21oi_1 _2909_ (.A1(\DJ8.GH[15] ),
    .A2(net76),
    .Y(_0670_),
    .B1(_0655_));
 sg13g2_xnor2_1 _2910_ (.Y(_0671_),
    .A(\DJ8.pc[14] ),
    .B(_0665_));
 sg13g2_nand2_1 _2911_ (.Y(_0672_),
    .A(_0671_),
    .B(_0608_));
 sg13g2_a22oi_1 _2912_ (.Y(_0125_),
    .B1(_0670_),
    .B2(_0672_),
    .A2(_0655_),
    .A1(_0669_));
 sg13g2_inv_1 _2913_ (.Y(_0673_),
    .A(\DJ8.pc[1] ));
 sg13g2_a21oi_1 _2914_ (.A1(_0604_),
    .A2(\DJ8.ir[1] ),
    .Y(_0674_),
    .B1(net80));
 sg13g2_nand2_1 _2915_ (.Y(_0675_),
    .A(_0673_),
    .B(_0598_));
 sg13g2_a21oi_1 _2916_ (.A1(_0675_),
    .A2(_0622_),
    .Y(_0676_),
    .B1(net77));
 sg13g2_nor2_1 _2917_ (.A(_0676_),
    .B(net73),
    .Y(_0677_));
 sg13g2_o21ai_1 _2918_ (.B1(_0677_),
    .Y(_0678_),
    .A1(\DJ8.GH[2] ),
    .A2(_0608_));
 sg13g2_a22oi_1 _2919_ (.Y(_0126_),
    .B1(_0674_),
    .B2(_0678_),
    .A2(_0673_),
    .A1(net81));
 sg13g2_a21oi_1 _2920_ (.A1(net68),
    .A2(\DJ8.ir[2] ),
    .Y(_0679_),
    .B1(net80));
 sg13g2_nand2_1 _2921_ (.Y(_0680_),
    .A(_0622_),
    .B(_0621_));
 sg13g2_nand3_1 _2922_ (.B(_0608_),
    .C(_0680_),
    .A(_0624_),
    .Y(_0681_));
 sg13g2_nand2_1 _2923_ (.Y(_0682_),
    .A(net77),
    .B(\DJ8.GH[3] ));
 sg13g2_a21o_1 _2924_ (.A2(_0682_),
    .A1(_0681_),
    .B1(net68),
    .X(_0683_));
 sg13g2_a22oi_1 _2925_ (.Y(_0127_),
    .B1(_0679_),
    .B2(_0683_),
    .A2(_0621_),
    .A1(_0597_));
 sg13g2_a21oi_1 _2926_ (.A1(net68),
    .A2(\DJ8.ir[3] ),
    .Y(_0684_),
    .B1(net80));
 sg13g2_nand2_1 _2927_ (.Y(_0685_),
    .A(_0624_),
    .B(_0620_));
 sg13g2_a21oi_1 _2928_ (.A1(_0626_),
    .A2(_0685_),
    .Y(_0686_),
    .B1(net77));
 sg13g2_o21ai_1 _2929_ (.B1(_0606_),
    .Y(_0687_),
    .A1(\DJ8.GH[4] ),
    .A2(_0608_));
 sg13g2_or2_1 _2930_ (.X(_0688_),
    .B(_0687_),
    .A(_0686_));
 sg13g2_a22oi_1 _2931_ (.Y(_0128_),
    .B1(_0684_),
    .B2(_0688_),
    .A2(_0620_),
    .A1(net81));
 sg13g2_a21oi_1 _2932_ (.A1(net68),
    .A2(net78),
    .Y(_0689_),
    .B1(net80));
 sg13g2_xnor2_1 _2933_ (.Y(_0690_),
    .A(_0619_),
    .B(_0625_));
 sg13g2_a21oi_1 _2934_ (.A1(_0838_),
    .A2(net76),
    .Y(_0691_),
    .B1(net73));
 sg13g2_o21ai_1 _2935_ (.B1(_0691_),
    .Y(_0692_),
    .A1(net76),
    .A2(_0690_));
 sg13g2_a22oi_1 _2936_ (.Y(_0129_),
    .B1(_0689_),
    .B2(_0692_),
    .A2(_0619_),
    .A1(net81));
 sg13g2_inv_1 _2937_ (.Y(_0693_),
    .A(\DJ8.pc[5] ));
 sg13g2_a21oi_1 _2938_ (.A1(net68),
    .A2(\DJ8.ir[5] ),
    .Y(_0694_),
    .B1(net80));
 sg13g2_xnor2_1 _2939_ (.Y(_0695_),
    .A(_0693_),
    .B(_0627_));
 sg13g2_a21oi_1 _2940_ (.A1(_0873_),
    .A2(net76),
    .Y(_0696_),
    .B1(net73));
 sg13g2_o21ai_1 _2941_ (.B1(_0696_),
    .Y(_0697_),
    .A1(net76),
    .A2(_0695_));
 sg13g2_a22oi_1 _2942_ (.Y(_0130_),
    .B1(_0694_),
    .B2(_0697_),
    .A2(_0693_),
    .A1(net81));
 sg13g2_a21oi_1 _2943_ (.A1(net68),
    .A2(\DJ8.ir[6] ),
    .Y(_0698_),
    .B1(net80));
 sg13g2_xnor2_1 _2944_ (.Y(_0699_),
    .A(\DJ8.pc[6] ),
    .B(_0628_));
 sg13g2_a21oi_1 _2945_ (.A1(_0780_),
    .A2(net77),
    .Y(_0700_),
    .B1(net73));
 sg13g2_o21ai_1 _2946_ (.B1(_0700_),
    .Y(_0701_),
    .A1(net76),
    .A2(_0699_));
 sg13g2_a22oi_1 _2947_ (.Y(_0131_),
    .B1(_0698_),
    .B2(_0701_),
    .A2(_0618_),
    .A1(net81));
 sg13g2_a21oi_1 _2948_ (.A1(net68),
    .A2(\DJ8.ir[7] ),
    .Y(_0702_),
    .B1(net80));
 sg13g2_nand2_1 _2949_ (.Y(_0703_),
    .A(_0630_),
    .B(_0617_));
 sg13g2_nor2b_1 _2950_ (.A(_0631_),
    .B_N(_0703_),
    .Y(_0704_));
 sg13g2_a21oi_1 _2951_ (.A1(_1008_),
    .A2(_0610_),
    .Y(_0705_),
    .B1(_0603_));
 sg13g2_o21ai_1 _2952_ (.B1(_0705_),
    .Y(_0706_),
    .A1(_0656_),
    .A2(_0704_));
 sg13g2_a22oi_1 _2953_ (.Y(_0132_),
    .B1(_0702_),
    .B2(_0706_),
    .A2(_0617_),
    .A1(_0597_));
 sg13g2_a21oi_1 _2954_ (.A1(_0604_),
    .A2(_0761_),
    .Y(_0707_),
    .B1(net80));
 sg13g2_xnor2_1 _2955_ (.Y(_0708_),
    .A(_0615_),
    .B(_0631_));
 sg13g2_a21oi_1 _2956_ (.A1(_1097_),
    .A2(net77),
    .Y(_0709_),
    .B1(net73));
 sg13g2_o21ai_1 _2957_ (.B1(_0709_),
    .Y(_0710_),
    .A1(_0656_),
    .A2(_0708_));
 sg13g2_a22oi_1 _2958_ (.Y(_0133_),
    .B1(_0707_),
    .B2(_0710_),
    .A2(_0615_),
    .A1(net81));
 sg13g2_o21ai_1 _2959_ (.B1(_0616_),
    .Y(_0711_),
    .A1(_0615_),
    .A2(_0632_));
 sg13g2_nand3_1 _2960_ (.B(_0634_),
    .C(_0608_),
    .A(_0711_),
    .Y(_0712_));
 sg13g2_nand2_1 _2961_ (.Y(_0713_),
    .A(net77),
    .B(\DJ8.GH[10] ));
 sg13g2_nand3_1 _2962_ (.B(_0606_),
    .C(_0713_),
    .A(_0712_),
    .Y(_0714_));
 sg13g2_a21oi_1 _2963_ (.A1(net73),
    .A2(_0489_),
    .Y(_0715_),
    .B1(_0596_));
 sg13g2_nand2_1 _2964_ (.Y(_0716_),
    .A(_0714_),
    .B(_0715_));
 sg13g2_o21ai_1 _2965_ (.B1(_0716_),
    .Y(_0134_),
    .A1(_0762_),
    .A2(_0616_));
 sg13g2_nor2_1 _2966_ (.A(_0596_),
    .B(_0758_),
    .Y(_0717_));
 sg13g2_a21oi_1 _2967_ (.A1(_0596_),
    .A2(\DJ8.state[3] ),
    .Y(_0718_),
    .B1(_0717_));
 sg13g2_mux2_1 _2968_ (.A0(_0025_),
    .A1(_0035_),
    .S(_0718_),
    .X(_0135_));
 sg13g2_a21oi_1 _2969_ (.A1(_0758_),
    .A2(_0762_),
    .Y(_0036_),
    .B1(\DJ8.state[3] ));
 sg13g2_nand2_1 _2970_ (.Y(_0719_),
    .A(_0757_),
    .B(_0774_));
 sg13g2_buf_1 _2971_ (.A(_0719_),
    .X(_0720_));
 sg13g2_nor2_1 _2972_ (.A(net72),
    .B(_1027_),
    .Y(_0721_));
 sg13g2_a21oi_1 _2973_ (.A1(net65),
    .A2(_0720_),
    .Y(net10),
    .B1(_0721_));
 sg13g2_inv_1 _2974_ (.Y(_0722_),
    .A(_0719_));
 sg13g2_nor2_1 _2975_ (.A(_0722_),
    .B(_0198_),
    .Y(_0723_));
 sg13g2_a21oi_1 _2976_ (.A1(_1102_),
    .A2(_0722_),
    .Y(net11),
    .B1(_0723_));
 sg13g2_nor2_1 _2977_ (.A(net72),
    .B(_1265_),
    .Y(_0724_));
 sg13g2_a21oi_1 _2978_ (.A1(net52),
    .A2(net72),
    .Y(net12),
    .B1(_0724_));
 sg13g2_nor2_1 _2979_ (.A(net72),
    .B(_1383_),
    .Y(_0725_));
 sg13g2_a21oi_1 _2980_ (.A1(net35),
    .A2(_0720_),
    .Y(net13),
    .B1(_0725_));
 sg13g2_nor2_1 _2981_ (.A(net72),
    .B(_0139_),
    .Y(_0726_));
 sg13g2_a21oi_1 _2982_ (.A1(net30),
    .A2(net72),
    .Y(net14),
    .B1(_0726_));
 sg13g2_nor2_1 _2983_ (.A(_0722_),
    .B(net32),
    .Y(_0727_));
 sg13g2_a21oi_1 _2984_ (.A1(_0252_),
    .A2(_0722_),
    .Y(net15),
    .B1(_0727_));
 sg13g2_nor2_1 _2985_ (.A(_0719_),
    .B(_0344_),
    .Y(_0728_));
 sg13g2_a21oi_1 _2986_ (.A1(_1370_),
    .A2(net72),
    .Y(net16),
    .B1(_0728_));
 sg13g2_nor2_1 _2987_ (.A(_0719_),
    .B(_0433_),
    .Y(_0729_));
 sg13g2_a21oi_1 _2988_ (.A1(net49),
    .A2(net72),
    .Y(net17),
    .B1(_0729_));
 sg13g2_buf_1 _2989_ (.A(net74),
    .X(_0730_));
 sg13g2_nand2_1 _2990_ (.Y(_0731_),
    .A(\DJ8.EF[8] ),
    .B(_0779_));
 sg13g2_o21ai_1 _2991_ (.B1(_0731_),
    .Y(_0732_),
    .A1(_0590_),
    .A2(_1008_));
 sg13g2_nor2_1 _2992_ (.A(_0732_),
    .B(net67),
    .Y(_0733_));
 sg13g2_a21oi_1 _2993_ (.A1(_0617_),
    .A2(_0730_),
    .Y(net18),
    .B1(_0733_));
 sg13g2_nand2_1 _2994_ (.Y(_0734_),
    .A(net78),
    .B(\DJ8.EF[9] ));
 sg13g2_o21ai_1 _2995_ (.B1(_0734_),
    .Y(_0735_),
    .A1(net78),
    .A2(_1097_));
 sg13g2_nor2_1 _2996_ (.A(_0735_),
    .B(net67),
    .Y(_0736_));
 sg13g2_a21oi_1 _2997_ (.A1(_0615_),
    .A2(net67),
    .Y(net19),
    .B1(_0736_));
 sg13g2_nand2_1 _2998_ (.Y(_0737_),
    .A(_0779_),
    .B(\DJ8.EF[10] ));
 sg13g2_o21ai_1 _2999_ (.B1(_0737_),
    .Y(_0738_),
    .A1(_0590_),
    .A2(_1254_));
 sg13g2_nor2_1 _3000_ (.A(_0738_),
    .B(net67),
    .Y(_0739_));
 sg13g2_a21oi_1 _3001_ (.A1(_0616_),
    .A2(_0730_),
    .Y(net20),
    .B1(_0739_));
 sg13g2_nand2_1 _3002_ (.Y(_0740_),
    .A(net84),
    .B(\DJ8.EF[11] ));
 sg13g2_o21ai_1 _3003_ (.B1(_0740_),
    .Y(_0741_),
    .A1(net78),
    .A2(_1376_));
 sg13g2_nor2_1 _3004_ (.A(_0741_),
    .B(net74),
    .Y(_0742_));
 sg13g2_a21oi_1 _3005_ (.A1(_0614_),
    .A2(net67),
    .Y(net21),
    .B1(_0742_));
 sg13g2_nand2_1 _3006_ (.Y(_0743_),
    .A(net84),
    .B(\DJ8.EF[12] ));
 sg13g2_o21ai_1 _3007_ (.B1(_0743_),
    .Y(_0744_),
    .A1(net78),
    .A2(_1484_));
 sg13g2_nor2_1 _3008_ (.A(_0744_),
    .B(net74),
    .Y(_0745_));
 sg13g2_a21oi_1 _3009_ (.A1(_0644_),
    .A2(net67),
    .Y(net22),
    .B1(_0745_));
 sg13g2_nand2_1 _3010_ (.Y(_0746_),
    .A(net84),
    .B(\DJ8.EF[13] ));
 sg13g2_o21ai_1 _3011_ (.B1(_0746_),
    .Y(_0747_),
    .A1(net78),
    .A2(_0247_));
 sg13g2_nor2_1 _3012_ (.A(_0747_),
    .B(_0776_),
    .Y(_0748_));
 sg13g2_a21oi_1 _3013_ (.A1(_0653_),
    .A2(net67),
    .Y(net23),
    .B1(_0748_));
 sg13g2_nand2_1 _3014_ (.Y(_0749_),
    .A(net84),
    .B(\DJ8.EF[14] ));
 sg13g2_o21ai_1 _3015_ (.B1(_0749_),
    .Y(_0750_),
    .A1(net78),
    .A2(_0337_));
 sg13g2_nor2_1 _3016_ (.A(_0750_),
    .B(_0776_),
    .Y(_0751_));
 sg13g2_a21oi_1 _3017_ (.A1(_0663_),
    .A2(net67),
    .Y(net24),
    .B1(_0751_));
 sg13g2_inv_1 _1561__1 (.Y(net115),
    .A(clknet_4_7_0_clk));
 sg13g2_buf_1 _3019_ (.A(net107),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3020_ (.A(net108),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3021_ (.A(net109),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3022_ (.A(net110),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3023_ (.A(net111),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3024_ (.A(net112),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3025_ (.A(net113),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3026_ (.A(net114),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3027_ (.A(\DJ8.we ),
    .X(net25));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout26 (.A(_0477_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0479_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0387_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0300_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_1365_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_1328_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_1348_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_1210_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1067_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1051_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0914_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0892_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0853_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0836_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1445_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1373_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1042_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_0965_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_0911_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0864_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0847_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1439_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1370_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1062_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_0930_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0929_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0905_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_0871_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_0844_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_0785_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_0542_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_0531_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_0520_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0509_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0499_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_0491_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0482_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_1058_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_0878_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0869_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_0769_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_0730_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_0604_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1025_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0863_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0809_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0720_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0603_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_0776_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_1163_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_0656_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0610_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0590_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_1092_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0641_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_0597_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_0574_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1156_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_0779_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_0986_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0798_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0778_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_0772_),
    .X(net88));
 sg13g2_buf_4 fanout89 (.X(net89),
    .A(net90));
 sg13g2_buf_4 fanout90 (.X(net90),
    .A(net93));
 sg13g2_buf_4 fanout91 (.X(net91),
    .A(net92));
 sg13g2_buf_2 fanout92 (.A(net93),
    .X(net92));
 sg13g2_buf_1 fanout93 (.A(net106),
    .X(net93));
 sg13g2_buf_4 fanout94 (.X(net94),
    .A(net97));
 sg13g2_buf_2 fanout95 (.A(net97),
    .X(net95));
 sg13g2_buf_4 fanout96 (.X(net96),
    .A(net97));
 sg13g2_buf_1 fanout97 (.A(net106),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(net102));
 sg13g2_buf_4 fanout99 (.X(net99),
    .A(net102));
 sg13g2_buf_4 fanout100 (.X(net100),
    .A(net102));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(net102));
 sg13g2_buf_2 fanout102 (.A(net106),
    .X(net102));
 sg13g2_buf_4 fanout103 (.X(net103),
    .A(net105));
 sg13g2_buf_2 fanout104 (.A(net105),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(net1),
    .X(net106));
 sg13g2_tiehi _3019__107 (.L_HI(net107));
 sg13g2_tiehi _3020__108 (.L_HI(net108));
 sg13g2_tiehi _3021__109 (.L_HI(net109));
 sg13g2_tiehi _3022__110 (.L_HI(net110));
 sg13g2_tiehi _3023__111 (.L_HI(net111));
 sg13g2_tiehi _3024__112 (.L_HI(net112));
 sg13g2_tiehi _3025__113 (.L_HI(net113));
 sg13g2_tiehi _3026__114 (.L_HI(net114));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_6_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_4_14_0_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_fill_2 FILLER_1_315 ();
 sg13g2_fill_1 FILLER_1_317 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_327 ();
 sg13g2_decap_8 FILLER_1_334 ();
 sg13g2_decap_8 FILLER_1_341 ();
 sg13g2_decap_4 FILLER_1_348 ();
 sg13g2_decap_8 FILLER_1_360 ();
 sg13g2_decap_8 FILLER_1_367 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_409 ();
 sg13g2_decap_8 FILLER_1_416 ();
 sg13g2_decap_8 FILLER_1_423 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_4 FILLER_2_21 ();
 sg13g2_fill_2 FILLER_2_25 ();
 sg13g2_decap_4 FILLER_2_53 ();
 sg13g2_fill_2 FILLER_2_57 ();
 sg13g2_fill_1 FILLER_2_85 ();
 sg13g2_decap_4 FILLER_2_112 ();
 sg13g2_fill_1 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_121 ();
 sg13g2_decap_8 FILLER_2_128 ();
 sg13g2_decap_8 FILLER_2_135 ();
 sg13g2_decap_4 FILLER_2_168 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_4 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_226 ();
 sg13g2_decap_8 FILLER_2_233 ();
 sg13g2_decap_8 FILLER_2_240 ();
 sg13g2_decap_4 FILLER_2_247 ();
 sg13g2_fill_2 FILLER_2_251 ();
 sg13g2_fill_1 FILLER_2_265 ();
 sg13g2_fill_1 FILLER_2_270 ();
 sg13g2_decap_4 FILLER_2_285 ();
 sg13g2_decap_4 FILLER_2_293 ();
 sg13g2_fill_1 FILLER_2_313 ();
 sg13g2_fill_2 FILLER_2_318 ();
 sg13g2_fill_1 FILLER_2_323 ();
 sg13g2_decap_4 FILLER_2_333 ();
 sg13g2_fill_1 FILLER_2_362 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_4 FILLER_2_388 ();
 sg13g2_fill_1 FILLER_2_392 ();
 sg13g2_decap_4 FILLER_2_398 ();
 sg13g2_fill_1 FILLER_2_402 ();
 sg13g2_fill_2 FILLER_2_413 ();
 sg13g2_fill_1 FILLER_2_415 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_fill_1 FILLER_3_31 ();
 sg13g2_decap_4 FILLER_3_36 ();
 sg13g2_fill_2 FILLER_3_40 ();
 sg13g2_decap_8 FILLER_3_51 ();
 sg13g2_decap_4 FILLER_3_64 ();
 sg13g2_fill_2 FILLER_3_68 ();
 sg13g2_decap_4 FILLER_3_84 ();
 sg13g2_fill_1 FILLER_3_88 ();
 sg13g2_fill_1 FILLER_3_94 ();
 sg13g2_fill_2 FILLER_3_101 ();
 sg13g2_fill_1 FILLER_3_107 ();
 sg13g2_fill_1 FILLER_3_113 ();
 sg13g2_fill_2 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_155 ();
 sg13g2_decap_8 FILLER_3_198 ();
 sg13g2_decap_8 FILLER_3_205 ();
 sg13g2_decap_8 FILLER_3_212 ();
 sg13g2_decap_8 FILLER_3_219 ();
 sg13g2_decap_8 FILLER_3_226 ();
 sg13g2_decap_4 FILLER_3_233 ();
 sg13g2_fill_2 FILLER_3_237 ();
 sg13g2_decap_4 FILLER_3_243 ();
 sg13g2_fill_2 FILLER_3_255 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_decap_4 FILLER_3_271 ();
 sg13g2_decap_8 FILLER_3_284 ();
 sg13g2_decap_4 FILLER_3_295 ();
 sg13g2_fill_1 FILLER_3_303 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_4 FILLER_3_333 ();
 sg13g2_fill_1 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_346 ();
 sg13g2_fill_1 FILLER_3_348 ();
 sg13g2_fill_2 FILLER_3_384 ();
 sg13g2_fill_2 FILLER_3_391 ();
 sg13g2_fill_2 FILLER_3_398 ();
 sg13g2_fill_1 FILLER_3_400 ();
 sg13g2_fill_1 FILLER_3_418 ();
 sg13g2_decap_8 FILLER_3_423 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_4 FILLER_4_28 ();
 sg13g2_fill_1 FILLER_4_62 ();
 sg13g2_decap_4 FILLER_4_73 ();
 sg13g2_fill_2 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_83 ();
 sg13g2_decap_8 FILLER_4_90 ();
 sg13g2_decap_4 FILLER_4_97 ();
 sg13g2_fill_1 FILLER_4_101 ();
 sg13g2_fill_2 FILLER_4_107 ();
 sg13g2_fill_1 FILLER_4_109 ();
 sg13g2_fill_1 FILLER_4_115 ();
 sg13g2_decap_4 FILLER_4_125 ();
 sg13g2_fill_1 FILLER_4_129 ();
 sg13g2_fill_2 FILLER_4_140 ();
 sg13g2_fill_2 FILLER_4_146 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_4 FILLER_4_168 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_decap_8 FILLER_4_179 ();
 sg13g2_decap_4 FILLER_4_212 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_decap_4 FILLER_4_226 ();
 sg13g2_decap_4 FILLER_4_234 ();
 sg13g2_fill_2 FILLER_4_238 ();
 sg13g2_decap_4 FILLER_4_244 ();
 sg13g2_fill_1 FILLER_4_254 ();
 sg13g2_decap_8 FILLER_4_260 ();
 sg13g2_decap_4 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_271 ();
 sg13g2_fill_1 FILLER_4_278 ();
 sg13g2_decap_8 FILLER_4_284 ();
 sg13g2_decap_8 FILLER_4_291 ();
 sg13g2_decap_4 FILLER_4_298 ();
 sg13g2_decap_8 FILLER_4_311 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_335 ();
 sg13g2_decap_4 FILLER_4_342 ();
 sg13g2_fill_1 FILLER_4_346 ();
 sg13g2_fill_1 FILLER_4_354 ();
 sg13g2_fill_2 FILLER_4_358 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_385 ();
 sg13g2_fill_1 FILLER_4_396 ();
 sg13g2_fill_1 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_410 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_4 FILLER_5_21 ();
 sg13g2_fill_1 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_57 ();
 sg13g2_fill_2 FILLER_5_64 ();
 sg13g2_fill_1 FILLER_5_92 ();
 sg13g2_fill_2 FILLER_5_145 ();
 sg13g2_fill_1 FILLER_5_147 ();
 sg13g2_fill_2 FILLER_5_184 ();
 sg13g2_fill_2 FILLER_5_191 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_223 ();
 sg13g2_decap_4 FILLER_5_230 ();
 sg13g2_fill_2 FILLER_5_234 ();
 sg13g2_decap_4 FILLER_5_240 ();
 sg13g2_fill_2 FILLER_5_244 ();
 sg13g2_fill_1 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_271 ();
 sg13g2_fill_2 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_fill_1 FILLER_5_324 ();
 sg13g2_decap_4 FILLER_5_329 ();
 sg13g2_fill_1 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_fill_2 FILLER_5_345 ();
 sg13g2_fill_1 FILLER_5_366 ();
 sg13g2_decap_4 FILLER_5_390 ();
 sg13g2_fill_1 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_2 FILLER_6_11 ();
 sg13g2_fill_1 FILLER_6_43 ();
 sg13g2_decap_4 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_89 ();
 sg13g2_fill_2 FILLER_6_96 ();
 sg13g2_decap_8 FILLER_6_103 ();
 sg13g2_decap_8 FILLER_6_110 ();
 sg13g2_decap_4 FILLER_6_117 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_fill_1 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_181 ();
 sg13g2_fill_2 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_190 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_decap_8 FILLER_6_206 ();
 sg13g2_decap_4 FILLER_6_213 ();
 sg13g2_decap_8 FILLER_6_246 ();
 sg13g2_decap_8 FILLER_6_262 ();
 sg13g2_decap_8 FILLER_6_269 ();
 sg13g2_decap_8 FILLER_6_276 ();
 sg13g2_fill_2 FILLER_6_283 ();
 sg13g2_decap_4 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_297 ();
 sg13g2_fill_2 FILLER_6_304 ();
 sg13g2_fill_1 FILLER_6_306 ();
 sg13g2_fill_1 FILLER_6_311 ();
 sg13g2_fill_1 FILLER_6_325 ();
 sg13g2_decap_8 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_356 ();
 sg13g2_decap_8 FILLER_6_363 ();
 sg13g2_decap_4 FILLER_6_370 ();
 sg13g2_fill_1 FILLER_6_374 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_fill_1 FILLER_6_398 ();
 sg13g2_fill_1 FILLER_6_404 ();
 sg13g2_fill_2 FILLER_6_410 ();
 sg13g2_fill_1 FILLER_6_412 ();
 sg13g2_fill_1 FILLER_6_417 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_4 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_29 ();
 sg13g2_decap_4 FILLER_7_36 ();
 sg13g2_decap_8 FILLER_7_45 ();
 sg13g2_fill_1 FILLER_7_52 ();
 sg13g2_fill_2 FILLER_7_79 ();
 sg13g2_fill_1 FILLER_7_81 ();
 sg13g2_decap_4 FILLER_7_111 ();
 sg13g2_decap_8 FILLER_7_145 ();
 sg13g2_decap_8 FILLER_7_152 ();
 sg13g2_decap_8 FILLER_7_159 ();
 sg13g2_decap_4 FILLER_7_166 ();
 sg13g2_fill_2 FILLER_7_170 ();
 sg13g2_fill_1 FILLER_7_202 ();
 sg13g2_fill_1 FILLER_7_216 ();
 sg13g2_decap_8 FILLER_7_226 ();
 sg13g2_decap_8 FILLER_7_233 ();
 sg13g2_decap_8 FILLER_7_240 ();
 sg13g2_fill_2 FILLER_7_247 ();
 sg13g2_fill_1 FILLER_7_249 ();
 sg13g2_decap_4 FILLER_7_276 ();
 sg13g2_fill_1 FILLER_7_284 ();
 sg13g2_fill_2 FILLER_7_307 ();
 sg13g2_fill_1 FILLER_7_309 ();
 sg13g2_fill_2 FILLER_7_317 ();
 sg13g2_decap_4 FILLER_7_324 ();
 sg13g2_fill_2 FILLER_7_332 ();
 sg13g2_fill_1 FILLER_7_334 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_fill_2 FILLER_7_363 ();
 sg13g2_fill_2 FILLER_7_378 ();
 sg13g2_decap_4 FILLER_7_385 ();
 sg13g2_fill_1 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_394 ();
 sg13g2_decap_8 FILLER_7_401 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_fill_1 FILLER_8_31 ();
 sg13g2_decap_8 FILLER_8_62 ();
 sg13g2_decap_4 FILLER_8_69 ();
 sg13g2_fill_2 FILLER_8_73 ();
 sg13g2_decap_8 FILLER_8_80 ();
 sg13g2_fill_2 FILLER_8_87 ();
 sg13g2_fill_2 FILLER_8_94 ();
 sg13g2_fill_1 FILLER_8_100 ();
 sg13g2_fill_1 FILLER_8_105 ();
 sg13g2_decap_4 FILLER_8_111 ();
 sg13g2_fill_2 FILLER_8_115 ();
 sg13g2_decap_8 FILLER_8_122 ();
 sg13g2_decap_8 FILLER_8_129 ();
 sg13g2_decap_4 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_4 FILLER_8_168 ();
 sg13g2_fill_2 FILLER_8_172 ();
 sg13g2_decap_4 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_188 ();
 sg13g2_decap_4 FILLER_8_193 ();
 sg13g2_fill_1 FILLER_8_206 ();
 sg13g2_fill_1 FILLER_8_233 ();
 sg13g2_decap_8 FILLER_8_243 ();
 sg13g2_decap_8 FILLER_8_250 ();
 sg13g2_decap_8 FILLER_8_257 ();
 sg13g2_decap_8 FILLER_8_264 ();
 sg13g2_fill_2 FILLER_8_271 ();
 sg13g2_fill_1 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_295 ();
 sg13g2_decap_8 FILLER_8_302 ();
 sg13g2_decap_8 FILLER_8_309 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_decap_4 FILLER_8_324 ();
 sg13g2_fill_2 FILLER_8_328 ();
 sg13g2_fill_2 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_360 ();
 sg13g2_fill_1 FILLER_8_362 ();
 sg13g2_fill_2 FILLER_8_368 ();
 sg13g2_fill_1 FILLER_8_370 ();
 sg13g2_decap_8 FILLER_8_384 ();
 sg13g2_fill_2 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_8_397 ();
 sg13g2_fill_1 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_fill_2 FILLER_8_427 ();
 sg13g2_fill_1 FILLER_8_429 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_4 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_29 ();
 sg13g2_decap_8 FILLER_9_36 ();
 sg13g2_decap_8 FILLER_9_51 ();
 sg13g2_fill_2 FILLER_9_58 ();
 sg13g2_fill_1 FILLER_9_60 ();
 sg13g2_fill_1 FILLER_9_65 ();
 sg13g2_fill_2 FILLER_9_97 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_fill_1 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_212 ();
 sg13g2_fill_2 FILLER_9_219 ();
 sg13g2_decap_4 FILLER_9_226 ();
 sg13g2_decap_4 FILLER_9_265 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_fill_1 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_decap_8 FILLER_9_310 ();
 sg13g2_decap_4 FILLER_9_317 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_4 FILLER_9_342 ();
 sg13g2_fill_2 FILLER_9_346 ();
 sg13g2_fill_1 FILLER_9_372 ();
 sg13g2_fill_2 FILLER_9_410 ();
 sg13g2_fill_1 FILLER_9_417 ();
 sg13g2_decap_8 FILLER_9_423 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_75 ();
 sg13g2_fill_1 FILLER_10_83 ();
 sg13g2_decap_8 FILLER_10_89 ();
 sg13g2_decap_8 FILLER_10_96 ();
 sg13g2_fill_2 FILLER_10_103 ();
 sg13g2_fill_1 FILLER_10_105 ();
 sg13g2_decap_8 FILLER_10_114 ();
 sg13g2_decap_8 FILLER_10_121 ();
 sg13g2_decap_8 FILLER_10_128 ();
 sg13g2_fill_2 FILLER_10_135 ();
 sg13g2_fill_1 FILLER_10_137 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_decap_4 FILLER_10_151 ();
 sg13g2_fill_2 FILLER_10_155 ();
 sg13g2_decap_4 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_164 ();
 sg13g2_fill_2 FILLER_10_169 ();
 sg13g2_fill_1 FILLER_10_171 ();
 sg13g2_decap_4 FILLER_10_186 ();
 sg13g2_fill_1 FILLER_10_190 ();
 sg13g2_decap_4 FILLER_10_199 ();
 sg13g2_fill_2 FILLER_10_203 ();
 sg13g2_fill_1 FILLER_10_215 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_fill_2 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_312 ();
 sg13g2_decap_4 FILLER_10_317 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_fill_2 FILLER_10_346 ();
 sg13g2_fill_1 FILLER_10_362 ();
 sg13g2_fill_1 FILLER_10_368 ();
 sg13g2_fill_1 FILLER_10_377 ();
 sg13g2_fill_2 FILLER_10_384 ();
 sg13g2_fill_2 FILLER_10_405 ();
 sg13g2_decap_4 FILLER_10_413 ();
 sg13g2_fill_2 FILLER_10_417 ();
 sg13g2_fill_2 FILLER_10_427 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_fill_1 FILLER_11_21 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_55 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_2 FILLER_11_69 ();
 sg13g2_fill_1 FILLER_11_71 ();
 sg13g2_decap_8 FILLER_11_76 ();
 sg13g2_fill_1 FILLER_11_83 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_decap_8 FILLER_11_124 ();
 sg13g2_decap_4 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_145 ();
 sg13g2_fill_2 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_158 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_4 FILLER_11_188 ();
 sg13g2_decap_4 FILLER_11_197 ();
 sg13g2_decap_8 FILLER_11_206 ();
 sg13g2_decap_8 FILLER_11_218 ();
 sg13g2_fill_2 FILLER_11_225 ();
 sg13g2_decap_4 FILLER_11_274 ();
 sg13g2_fill_2 FILLER_11_278 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_295 ();
 sg13g2_decap_8 FILLER_11_306 ();
 sg13g2_decap_8 FILLER_11_313 ();
 sg13g2_decap_4 FILLER_11_320 ();
 sg13g2_fill_2 FILLER_11_324 ();
 sg13g2_decap_8 FILLER_11_334 ();
 sg13g2_decap_8 FILLER_11_341 ();
 sg13g2_fill_1 FILLER_11_348 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_fill_1 FILLER_11_383 ();
 sg13g2_fill_2 FILLER_11_392 ();
 sg13g2_fill_1 FILLER_11_402 ();
 sg13g2_decap_8 FILLER_11_411 ();
 sg13g2_decap_8 FILLER_11_418 ();
 sg13g2_decap_4 FILLER_11_425 ();
 sg13g2_fill_1 FILLER_11_429 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_78 ();
 sg13g2_decap_8 FILLER_12_85 ();
 sg13g2_decap_8 FILLER_12_92 ();
 sg13g2_fill_1 FILLER_12_99 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_153 ();
 sg13g2_decap_4 FILLER_12_160 ();
 sg13g2_fill_2 FILLER_12_169 ();
 sg13g2_fill_1 FILLER_12_171 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_229 ();
 sg13g2_fill_1 FILLER_12_236 ();
 sg13g2_fill_1 FILLER_12_241 ();
 sg13g2_fill_1 FILLER_12_246 ();
 sg13g2_decap_8 FILLER_12_266 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_288 ();
 sg13g2_decap_8 FILLER_12_314 ();
 sg13g2_decap_4 FILLER_12_321 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_4 FILLER_12_358 ();
 sg13g2_fill_2 FILLER_12_362 ();
 sg13g2_decap_8 FILLER_12_372 ();
 sg13g2_decap_4 FILLER_12_388 ();
 sg13g2_decap_4 FILLER_12_403 ();
 sg13g2_fill_2 FILLER_12_407 ();
 sg13g2_fill_2 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_fill_1 FILLER_13_28 ();
 sg13g2_decap_4 FILLER_13_34 ();
 sg13g2_fill_1 FILLER_13_38 ();
 sg13g2_fill_2 FILLER_13_48 ();
 sg13g2_fill_2 FILLER_13_125 ();
 sg13g2_fill_1 FILLER_13_127 ();
 sg13g2_decap_4 FILLER_13_136 ();
 sg13g2_fill_2 FILLER_13_140 ();
 sg13g2_fill_2 FILLER_13_167 ();
 sg13g2_fill_1 FILLER_13_169 ();
 sg13g2_decap_4 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_183 ();
 sg13g2_decap_8 FILLER_13_194 ();
 sg13g2_decap_8 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_208 ();
 sg13g2_decap_4 FILLER_13_218 ();
 sg13g2_fill_2 FILLER_13_222 ();
 sg13g2_decap_4 FILLER_13_232 ();
 sg13g2_fill_1 FILLER_13_236 ();
 sg13g2_fill_2 FILLER_13_242 ();
 sg13g2_fill_2 FILLER_13_249 ();
 sg13g2_fill_1 FILLER_13_251 ();
 sg13g2_fill_2 FILLER_13_257 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_297 ();
 sg13g2_fill_2 FILLER_13_311 ();
 sg13g2_fill_1 FILLER_13_313 ();
 sg13g2_fill_1 FILLER_13_319 ();
 sg13g2_fill_1 FILLER_13_325 ();
 sg13g2_fill_1 FILLER_13_331 ();
 sg13g2_fill_1 FILLER_13_336 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_2 FILLER_13_349 ();
 sg13g2_fill_1 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_372 ();
 sg13g2_decap_8 FILLER_13_379 ();
 sg13g2_decap_4 FILLER_13_386 ();
 sg13g2_fill_2 FILLER_13_390 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_4 FILLER_14_21 ();
 sg13g2_fill_1 FILLER_14_25 ();
 sg13g2_decap_8 FILLER_14_30 ();
 sg13g2_decap_8 FILLER_14_37 ();
 sg13g2_fill_2 FILLER_14_44 ();
 sg13g2_decap_8 FILLER_14_81 ();
 sg13g2_decap_8 FILLER_14_88 ();
 sg13g2_decap_4 FILLER_14_95 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_decap_4 FILLER_14_147 ();
 sg13g2_fill_2 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_178 ();
 sg13g2_fill_1 FILLER_14_180 ();
 sg13g2_decap_4 FILLER_14_185 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_fill_2 FILLER_14_207 ();
 sg13g2_decap_8 FILLER_14_227 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_243 ();
 sg13g2_fill_2 FILLER_14_262 ();
 sg13g2_decap_8 FILLER_14_267 ();
 sg13g2_decap_8 FILLER_14_274 ();
 sg13g2_decap_4 FILLER_14_281 ();
 sg13g2_decap_8 FILLER_14_303 ();
 sg13g2_fill_1 FILLER_14_310 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_fill_2 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_4 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_4 FILLER_14_383 ();
 sg13g2_fill_2 FILLER_14_387 ();
 sg13g2_fill_1 FILLER_14_403 ();
 sg13g2_decap_4 FILLER_14_407 ();
 sg13g2_fill_1 FILLER_14_411 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_4 FILLER_14_424 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_32 ();
 sg13g2_fill_1 FILLER_15_43 ();
 sg13g2_decap_8 FILLER_15_52 ();
 sg13g2_fill_2 FILLER_15_59 ();
 sg13g2_fill_1 FILLER_15_61 ();
 sg13g2_fill_1 FILLER_15_79 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_fill_1 FILLER_15_91 ();
 sg13g2_decap_8 FILLER_15_100 ();
 sg13g2_decap_8 FILLER_15_107 ();
 sg13g2_decap_4 FILLER_15_123 ();
 sg13g2_decap_4 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_134 ();
 sg13g2_fill_1 FILLER_15_139 ();
 sg13g2_fill_1 FILLER_15_149 ();
 sg13g2_fill_2 FILLER_15_169 ();
 sg13g2_decap_4 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_184 ();
 sg13g2_fill_2 FILLER_15_214 ();
 sg13g2_fill_1 FILLER_15_216 ();
 sg13g2_decap_4 FILLER_15_222 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_1 FILLER_15_254 ();
 sg13g2_fill_1 FILLER_15_293 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_fill_2 FILLER_15_310 ();
 sg13g2_fill_1 FILLER_15_312 ();
 sg13g2_fill_1 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_370 ();
 sg13g2_fill_2 FILLER_15_405 ();
 sg13g2_fill_2 FILLER_15_410 ();
 sg13g2_fill_1 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_4 FILLER_16_14 ();
 sg13g2_fill_2 FILLER_16_18 ();
 sg13g2_fill_2 FILLER_16_46 ();
 sg13g2_fill_1 FILLER_16_48 ();
 sg13g2_fill_2 FILLER_16_75 ();
 sg13g2_decap_4 FILLER_16_82 ();
 sg13g2_fill_2 FILLER_16_91 ();
 sg13g2_decap_4 FILLER_16_97 ();
 sg13g2_decap_8 FILLER_16_107 ();
 sg13g2_decap_8 FILLER_16_114 ();
 sg13g2_decap_4 FILLER_16_121 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_decap_4 FILLER_16_154 ();
 sg13g2_fill_2 FILLER_16_158 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_4 FILLER_16_177 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_2 FILLER_16_185 ();
 sg13g2_fill_1 FILLER_16_187 ();
 sg13g2_fill_2 FILLER_16_197 ();
 sg13g2_decap_4 FILLER_16_204 ();
 sg13g2_decap_8 FILLER_16_216 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_8 FILLER_16_230 ();
 sg13g2_fill_1 FILLER_16_237 ();
 sg13g2_fill_1 FILLER_16_243 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_255 ();
 sg13g2_decap_8 FILLER_16_261 ();
 sg13g2_decap_8 FILLER_16_268 ();
 sg13g2_fill_2 FILLER_16_275 ();
 sg13g2_fill_1 FILLER_16_282 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_4 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_2 FILLER_16_328 ();
 sg13g2_fill_1 FILLER_16_330 ();
 sg13g2_fill_1 FILLER_16_343 ();
 sg13g2_fill_2 FILLER_16_353 ();
 sg13g2_fill_1 FILLER_16_355 ();
 sg13g2_fill_2 FILLER_16_364 ();
 sg13g2_fill_1 FILLER_16_366 ();
 sg13g2_fill_1 FILLER_16_375 ();
 sg13g2_fill_2 FILLER_16_381 ();
 sg13g2_fill_1 FILLER_16_383 ();
 sg13g2_decap_4 FILLER_16_387 ();
 sg13g2_fill_2 FILLER_16_399 ();
 sg13g2_fill_1 FILLER_16_401 ();
 sg13g2_decap_8 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_16_414 ();
 sg13g2_decap_8 FILLER_16_421 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_decap_8 FILLER_17_26 ();
 sg13g2_decap_8 FILLER_17_33 ();
 sg13g2_fill_2 FILLER_17_40 ();
 sg13g2_fill_1 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_51 ();
 sg13g2_decap_8 FILLER_17_65 ();
 sg13g2_decap_8 FILLER_17_72 ();
 sg13g2_decap_4 FILLER_17_79 ();
 sg13g2_fill_1 FILLER_17_83 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_8 FILLER_17_117 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_decap_4 FILLER_17_161 ();
 sg13g2_fill_2 FILLER_17_165 ();
 sg13g2_fill_1 FILLER_17_182 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_fill_1 FILLER_17_193 ();
 sg13g2_fill_1 FILLER_17_227 ();
 sg13g2_decap_8 FILLER_17_258 ();
 sg13g2_fill_1 FILLER_17_265 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_308 ();
 sg13g2_fill_2 FILLER_17_315 ();
 sg13g2_fill_2 FILLER_17_343 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_fill_1 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_364 ();
 sg13g2_decap_4 FILLER_17_371 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_fill_2 FILLER_17_393 ();
 sg13g2_fill_1 FILLER_17_395 ();
 sg13g2_decap_8 FILLER_17_422 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_2 FILLER_18_76 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_4 FILLER_18_91 ();
 sg13g2_fill_1 FILLER_18_95 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_4 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_156 ();
 sg13g2_fill_2 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_decap_4 FILLER_18_199 ();
 sg13g2_fill_2 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_209 ();
 sg13g2_decap_4 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_2 FILLER_18_229 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_250 ();
 sg13g2_fill_1 FILLER_18_255 ();
 sg13g2_fill_2 FILLER_18_261 ();
 sg13g2_decap_8 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_303 ();
 sg13g2_decap_4 FILLER_18_310 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_335 ();
 sg13g2_decap_8 FILLER_18_342 ();
 sg13g2_decap_4 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_353 ();
 sg13g2_decap_8 FILLER_18_363 ();
 sg13g2_decap_8 FILLER_18_379 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_decap_4 FILLER_18_392 ();
 sg13g2_fill_2 FILLER_18_427 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_1 FILLER_19_30 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_decap_8 FILLER_19_40 ();
 sg13g2_fill_1 FILLER_19_56 ();
 sg13g2_fill_2 FILLER_19_60 ();
 sg13g2_fill_2 FILLER_19_66 ();
 sg13g2_fill_1 FILLER_19_68 ();
 sg13g2_fill_2 FILLER_19_137 ();
 sg13g2_fill_1 FILLER_19_139 ();
 sg13g2_fill_2 FILLER_19_144 ();
 sg13g2_fill_2 FILLER_19_149 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_176 ();
 sg13g2_fill_1 FILLER_19_204 ();
 sg13g2_decap_8 FILLER_19_209 ();
 sg13g2_decap_8 FILLER_19_216 ();
 sg13g2_decap_4 FILLER_19_223 ();
 sg13g2_fill_1 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_4 FILLER_19_259 ();
 sg13g2_decap_4 FILLER_19_270 ();
 sg13g2_fill_1 FILLER_19_274 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_fill_2 FILLER_19_287 ();
 sg13g2_fill_1 FILLER_19_289 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_fill_2 FILLER_19_302 ();
 sg13g2_decap_8 FILLER_19_318 ();
 sg13g2_fill_2 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_335 ();
 sg13g2_decap_4 FILLER_19_342 ();
 sg13g2_fill_2 FILLER_19_346 ();
 sg13g2_fill_2 FILLER_19_366 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_fill_2 FILLER_19_379 ();
 sg13g2_decap_4 FILLER_19_386 ();
 sg13g2_decap_8 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_411 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_4 FILLER_20_66 ();
 sg13g2_fill_1 FILLER_20_75 ();
 sg13g2_decap_4 FILLER_20_117 ();
 sg13g2_fill_2 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_166 ();
 sg13g2_decap_8 FILLER_20_173 ();
 sg13g2_decap_8 FILLER_20_180 ();
 sg13g2_decap_8 FILLER_20_187 ();
 sg13g2_decap_4 FILLER_20_194 ();
 sg13g2_fill_2 FILLER_20_198 ();
 sg13g2_fill_2 FILLER_20_209 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_fill_2 FILLER_20_238 ();
 sg13g2_fill_1 FILLER_20_240 ();
 sg13g2_decap_8 FILLER_20_250 ();
 sg13g2_decap_8 FILLER_20_257 ();
 sg13g2_decap_8 FILLER_20_264 ();
 sg13g2_decap_8 FILLER_20_271 ();
 sg13g2_decap_8 FILLER_20_278 ();
 sg13g2_decap_4 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_289 ();
 sg13g2_fill_1 FILLER_20_295 ();
 sg13g2_fill_1 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_306 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_355 ();
 sg13g2_decap_8 FILLER_20_362 ();
 sg13g2_decap_4 FILLER_20_369 ();
 sg13g2_fill_1 FILLER_20_373 ();
 sg13g2_fill_2 FILLER_20_382 ();
 sg13g2_fill_1 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_404 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_4 FILLER_20_424 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_21_26 ();
 sg13g2_decap_8 FILLER_21_33 ();
 sg13g2_decap_8 FILLER_21_40 ();
 sg13g2_decap_4 FILLER_21_47 ();
 sg13g2_fill_2 FILLER_21_51 ();
 sg13g2_fill_2 FILLER_21_56 ();
 sg13g2_fill_1 FILLER_21_58 ();
 sg13g2_decap_8 FILLER_21_68 ();
 sg13g2_fill_2 FILLER_21_75 ();
 sg13g2_decap_4 FILLER_21_82 ();
 sg13g2_fill_1 FILLER_21_99 ();
 sg13g2_fill_1 FILLER_21_105 ();
 sg13g2_fill_2 FILLER_21_115 ();
 sg13g2_decap_4 FILLER_21_125 ();
 sg13g2_fill_2 FILLER_21_129 ();
 sg13g2_decap_4 FILLER_21_140 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_fill_1 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_166 ();
 sg13g2_decap_8 FILLER_21_208 ();
 sg13g2_decap_8 FILLER_21_284 ();
 sg13g2_decap_8 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_fill_1 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_321 ();
 sg13g2_decap_8 FILLER_21_328 ();
 sg13g2_decap_4 FILLER_21_339 ();
 sg13g2_decap_4 FILLER_21_347 ();
 sg13g2_fill_2 FILLER_21_351 ();
 sg13g2_fill_2 FILLER_21_358 ();
 sg13g2_decap_4 FILLER_21_364 ();
 sg13g2_fill_1 FILLER_21_368 ();
 sg13g2_fill_1 FILLER_21_373 ();
 sg13g2_decap_4 FILLER_21_383 ();
 sg13g2_fill_2 FILLER_21_387 ();
 sg13g2_fill_1 FILLER_21_397 ();
 sg13g2_fill_1 FILLER_21_402 ();
 sg13g2_decap_8 FILLER_21_407 ();
 sg13g2_decap_4 FILLER_21_414 ();
 sg13g2_fill_2 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_424 ();
 sg13g2_fill_2 FILLER_21_428 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_fill_1 FILLER_22_39 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_49 ();
 sg13g2_decap_8 FILLER_22_69 ();
 sg13g2_fill_2 FILLER_22_76 ();
 sg13g2_fill_1 FILLER_22_78 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_decap_4 FILLER_22_98 ();
 sg13g2_fill_1 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_129 ();
 sg13g2_decap_4 FILLER_22_136 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_decap_4 FILLER_22_146 ();
 sg13g2_fill_1 FILLER_22_150 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_fill_1 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_decap_8 FILLER_22_225 ();
 sg13g2_decap_8 FILLER_22_232 ();
 sg13g2_decap_8 FILLER_22_239 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_264 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_292 ();
 sg13g2_fill_2 FILLER_22_301 ();
 sg13g2_decap_4 FILLER_22_307 ();
 sg13g2_decap_8 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_329 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_fill_2 FILLER_22_361 ();
 sg13g2_fill_2 FILLER_22_367 ();
 sg13g2_fill_2 FILLER_22_374 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_390 ();
 sg13g2_decap_4 FILLER_22_416 ();
 sg13g2_decap_4 FILLER_22_424 ();
 sg13g2_fill_2 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_fill_2 FILLER_23_14 ();
 sg13g2_decap_4 FILLER_23_25 ();
 sg13g2_fill_1 FILLER_23_55 ();
 sg13g2_fill_1 FILLER_23_59 ();
 sg13g2_decap_8 FILLER_23_86 ();
 sg13g2_fill_1 FILLER_23_93 ();
 sg13g2_decap_8 FILLER_23_107 ();
 sg13g2_fill_1 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_124 ();
 sg13g2_decap_8 FILLER_23_131 ();
 sg13g2_decap_4 FILLER_23_138 ();
 sg13g2_fill_2 FILLER_23_142 ();
 sg13g2_fill_1 FILLER_23_148 ();
 sg13g2_decap_8 FILLER_23_153 ();
 sg13g2_decap_4 FILLER_23_160 ();
 sg13g2_decap_8 FILLER_23_202 ();
 sg13g2_decap_8 FILLER_23_209 ();
 sg13g2_decap_4 FILLER_23_216 ();
 sg13g2_fill_1 FILLER_23_220 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_fill_2 FILLER_23_252 ();
 sg13g2_fill_2 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_278 ();
 sg13g2_decap_8 FILLER_23_283 ();
 sg13g2_fill_1 FILLER_23_290 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_2 FILLER_23_322 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_329 ();
 sg13g2_fill_1 FILLER_23_331 ();
 sg13g2_decap_4 FILLER_23_345 ();
 sg13g2_fill_1 FILLER_23_349 ();
 sg13g2_fill_1 FILLER_23_355 ();
 sg13g2_decap_4 FILLER_23_361 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_2 FILLER_23_385 ();
 sg13g2_fill_1 FILLER_23_387 ();
 sg13g2_fill_2 FILLER_23_401 ();
 sg13g2_decap_4 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_23_411 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_26 ();
 sg13g2_decap_8 FILLER_24_33 ();
 sg13g2_decap_8 FILLER_24_40 ();
 sg13g2_decap_8 FILLER_24_47 ();
 sg13g2_fill_2 FILLER_24_54 ();
 sg13g2_fill_1 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_92 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_decap_8 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_161 ();
 sg13g2_decap_4 FILLER_24_181 ();
 sg13g2_decap_8 FILLER_24_201 ();
 sg13g2_decap_4 FILLER_24_208 ();
 sg13g2_fill_2 FILLER_24_212 ();
 sg13g2_fill_2 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_226 ();
 sg13g2_decap_8 FILLER_24_233 ();
 sg13g2_decap_4 FILLER_24_240 ();
 sg13g2_fill_1 FILLER_24_244 ();
 sg13g2_fill_2 FILLER_24_266 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_273 ();
 sg13g2_fill_1 FILLER_24_286 ();
 sg13g2_fill_2 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_294 ();
 sg13g2_decap_4 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_1 FILLER_24_320 ();
 sg13g2_fill_2 FILLER_24_326 ();
 sg13g2_fill_1 FILLER_24_328 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_2 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_351 ();
 sg13g2_fill_1 FILLER_24_353 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_1 FILLER_24_375 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_fill_2 FILLER_24_390 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_4 FILLER_24_403 ();
 sg13g2_fill_1 FILLER_24_407 ();
 sg13g2_fill_2 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_422 ();
 sg13g2_fill_1 FILLER_24_429 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_14 ();
 sg13g2_fill_1 FILLER_25_16 ();
 sg13g2_decap_4 FILLER_25_26 ();
 sg13g2_decap_8 FILLER_25_39 ();
 sg13g2_decap_8 FILLER_25_46 ();
 sg13g2_fill_2 FILLER_25_53 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_2 FILLER_25_70 ();
 sg13g2_decap_4 FILLER_25_75 ();
 sg13g2_fill_1 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_4 FILLER_25_91 ();
 sg13g2_fill_1 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_106 ();
 sg13g2_decap_4 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_117 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_decap_4 FILLER_25_141 ();
 sg13g2_fill_2 FILLER_25_156 ();
 sg13g2_fill_1 FILLER_25_158 ();
 sg13g2_fill_2 FILLER_25_166 ();
 sg13g2_fill_1 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_173 ();
 sg13g2_decap_8 FILLER_25_180 ();
 sg13g2_fill_2 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_197 ();
 sg13g2_fill_2 FILLER_25_204 ();
 sg13g2_fill_1 FILLER_25_206 ();
 sg13g2_decap_8 FILLER_25_225 ();
 sg13g2_decap_8 FILLER_25_232 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_decap_4 FILLER_25_261 ();
 sg13g2_fill_1 FILLER_25_265 ();
 sg13g2_decap_4 FILLER_25_283 ();
 sg13g2_fill_1 FILLER_25_301 ();
 sg13g2_decap_4 FILLER_25_319 ();
 sg13g2_decap_4 FILLER_25_333 ();
 sg13g2_fill_2 FILLER_25_337 ();
 sg13g2_fill_2 FILLER_25_344 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_fill_1 FILLER_25_356 ();
 sg13g2_decap_4 FILLER_25_362 ();
 sg13g2_fill_2 FILLER_25_393 ();
 sg13g2_fill_1 FILLER_25_395 ();
 sg13g2_decap_4 FILLER_25_404 ();
 sg13g2_decap_4 FILLER_25_416 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_fill_1 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_58 ();
 sg13g2_fill_1 FILLER_26_65 ();
 sg13g2_fill_2 FILLER_26_70 ();
 sg13g2_fill_2 FILLER_26_76 ();
 sg13g2_decap_8 FILLER_26_83 ();
 sg13g2_fill_1 FILLER_26_90 ();
 sg13g2_decap_8 FILLER_26_99 ();
 sg13g2_fill_1 FILLER_26_106 ();
 sg13g2_fill_1 FILLER_26_112 ();
 sg13g2_fill_1 FILLER_26_123 ();
 sg13g2_fill_1 FILLER_26_128 ();
 sg13g2_fill_2 FILLER_26_139 ();
 sg13g2_decap_8 FILLER_26_180 ();
 sg13g2_fill_2 FILLER_26_187 ();
 sg13g2_decap_4 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_208 ();
 sg13g2_fill_2 FILLER_26_215 ();
 sg13g2_decap_8 FILLER_26_221 ();
 sg13g2_decap_8 FILLER_26_228 ();
 sg13g2_decap_4 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_fill_2 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_279 ();
 sg13g2_fill_2 FILLER_26_284 ();
 sg13g2_fill_2 FILLER_26_295 ();
 sg13g2_fill_2 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_308 ();
 sg13g2_decap_4 FILLER_26_322 ();
 sg13g2_fill_1 FILLER_26_342 ();
 sg13g2_decap_4 FILLER_26_351 ();
 sg13g2_decap_4 FILLER_26_365 ();
 sg13g2_decap_8 FILLER_26_380 ();
 sg13g2_decap_8 FILLER_26_387 ();
 sg13g2_decap_8 FILLER_26_394 ();
 sg13g2_decap_4 FILLER_26_401 ();
 sg13g2_decap_8 FILLER_26_419 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_1 FILLER_27_30 ();
 sg13g2_decap_4 FILLER_27_42 ();
 sg13g2_fill_2 FILLER_27_46 ();
 sg13g2_decap_4 FILLER_27_58 ();
 sg13g2_decap_4 FILLER_27_70 ();
 sg13g2_fill_2 FILLER_27_78 ();
 sg13g2_decap_4 FILLER_27_84 ();
 sg13g2_fill_1 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_94 ();
 sg13g2_decap_8 FILLER_27_101 ();
 sg13g2_decap_4 FILLER_27_123 ();
 sg13g2_fill_1 FILLER_27_127 ();
 sg13g2_decap_8 FILLER_27_156 ();
 sg13g2_decap_8 FILLER_27_163 ();
 sg13g2_fill_1 FILLER_27_170 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_4 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_190 ();
 sg13g2_decap_8 FILLER_27_208 ();
 sg13g2_fill_2 FILLER_27_215 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_4 FILLER_27_235 ();
 sg13g2_fill_2 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_decap_4 FILLER_27_261 ();
 sg13g2_fill_1 FILLER_27_265 ();
 sg13g2_fill_1 FILLER_27_270 ();
 sg13g2_fill_2 FILLER_27_275 ();
 sg13g2_fill_2 FILLER_27_287 ();
 sg13g2_fill_1 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_300 ();
 sg13g2_fill_2 FILLER_27_309 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_fill_2 FILLER_27_322 ();
 sg13g2_fill_1 FILLER_27_337 ();
 sg13g2_fill_1 FILLER_27_347 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_359 ();
 sg13g2_fill_2 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_fill_2 FILLER_28_35 ();
 sg13g2_fill_2 FILLER_28_48 ();
 sg13g2_fill_1 FILLER_28_50 ();
 sg13g2_fill_1 FILLER_28_59 ();
 sg13g2_fill_2 FILLER_28_64 ();
 sg13g2_fill_1 FILLER_28_66 ();
 sg13g2_decap_8 FILLER_28_72 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_85 ();
 sg13g2_decap_8 FILLER_28_102 ();
 sg13g2_decap_8 FILLER_28_109 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_decap_4 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_212 ();
 sg13g2_decap_4 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_1 FILLER_28_238 ();
 sg13g2_fill_1 FILLER_28_248 ();
 sg13g2_fill_1 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_263 ();
 sg13g2_fill_2 FILLER_28_272 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_307 ();
 sg13g2_decap_8 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_319 ();
 sg13g2_fill_2 FILLER_28_326 ();
 sg13g2_fill_1 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_353 ();
 sg13g2_fill_2 FILLER_28_364 ();
 sg13g2_fill_1 FILLER_28_366 ();
 sg13g2_fill_2 FILLER_28_372 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_fill_1 FILLER_28_379 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_391 ();
 sg13g2_fill_1 FILLER_28_393 ();
 sg13g2_fill_2 FILLER_28_399 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_decap_8 FILLER_28_414 ();
 sg13g2_decap_8 FILLER_28_421 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_4 FILLER_29_28 ();
 sg13g2_fill_1 FILLER_29_32 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_4 FILLER_29_81 ();
 sg13g2_fill_1 FILLER_29_85 ();
 sg13g2_decap_8 FILLER_29_90 ();
 sg13g2_fill_2 FILLER_29_97 ();
 sg13g2_fill_1 FILLER_29_99 ();
 sg13g2_fill_2 FILLER_29_114 ();
 sg13g2_fill_2 FILLER_29_135 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_fill_1 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_147 ();
 sg13g2_fill_1 FILLER_29_149 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_fill_1 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_4 FILLER_29_186 ();
 sg13g2_fill_1 FILLER_29_195 ();
 sg13g2_decap_4 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_208 ();
 sg13g2_decap_4 FILLER_29_214 ();
 sg13g2_fill_1 FILLER_29_228 ();
 sg13g2_decap_4 FILLER_29_244 ();
 sg13g2_fill_1 FILLER_29_248 ();
 sg13g2_decap_4 FILLER_29_254 ();
 sg13g2_fill_2 FILLER_29_262 ();
 sg13g2_fill_1 FILLER_29_272 ();
 sg13g2_fill_1 FILLER_29_301 ();
 sg13g2_fill_1 FILLER_29_311 ();
 sg13g2_decap_4 FILLER_29_316 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_326 ();
 sg13g2_fill_1 FILLER_29_340 ();
 sg13g2_fill_1 FILLER_29_346 ();
 sg13g2_fill_1 FILLER_29_370 ();
 sg13g2_fill_1 FILLER_29_376 ();
 sg13g2_fill_1 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_1 FILLER_29_402 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_29_409 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_27 ();
 sg13g2_fill_1 FILLER_30_29 ();
 sg13g2_fill_2 FILLER_30_49 ();
 sg13g2_fill_1 FILLER_30_51 ();
 sg13g2_fill_2 FILLER_30_69 ();
 sg13g2_fill_1 FILLER_30_71 ();
 sg13g2_fill_2 FILLER_30_77 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_121 ();
 sg13g2_decap_8 FILLER_30_128 ();
 sg13g2_decap_8 FILLER_30_135 ();
 sg13g2_fill_2 FILLER_30_142 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_fill_1 FILLER_30_194 ();
 sg13g2_decap_8 FILLER_30_205 ();
 sg13g2_decap_8 FILLER_30_212 ();
 sg13g2_decap_4 FILLER_30_219 ();
 sg13g2_fill_1 FILLER_30_223 ();
 sg13g2_fill_1 FILLER_30_232 ();
 sg13g2_fill_1 FILLER_30_238 ();
 sg13g2_fill_2 FILLER_30_243 ();
 sg13g2_decap_4 FILLER_30_258 ();
 sg13g2_fill_2 FILLER_30_266 ();
 sg13g2_fill_1 FILLER_30_277 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_287 ();
 sg13g2_fill_2 FILLER_30_296 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_337 ();
 sg13g2_fill_2 FILLER_30_343 ();
 sg13g2_fill_1 FILLER_30_345 ();
 sg13g2_fill_1 FILLER_30_356 ();
 sg13g2_fill_1 FILLER_30_370 ();
 sg13g2_fill_2 FILLER_30_374 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_4 FILLER_30_410 ();
 sg13g2_decap_8 FILLER_30_419 ();
 sg13g2_decap_4 FILLER_30_426 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_4 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_18 ();
 sg13g2_fill_1 FILLER_31_24 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_fill_2 FILLER_31_73 ();
 sg13g2_fill_1 FILLER_31_75 ();
 sg13g2_decap_8 FILLER_31_79 ();
 sg13g2_decap_4 FILLER_31_86 ();
 sg13g2_fill_2 FILLER_31_90 ();
 sg13g2_decap_4 FILLER_31_96 ();
 sg13g2_fill_2 FILLER_31_100 ();
 sg13g2_decap_4 FILLER_31_110 ();
 sg13g2_fill_1 FILLER_31_119 ();
 sg13g2_fill_1 FILLER_31_151 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_decap_4 FILLER_31_163 ();
 sg13g2_decap_8 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_decap_8 FILLER_31_205 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_decap_8 FILLER_31_219 ();
 sg13g2_decap_8 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_fill_1 FILLER_31_240 ();
 sg13g2_fill_1 FILLER_31_260 ();
 sg13g2_decap_8 FILLER_31_269 ();
 sg13g2_fill_2 FILLER_31_280 ();
 sg13g2_fill_2 FILLER_31_303 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_311 ();
 sg13g2_fill_2 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_318 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_338 ();
 sg13g2_fill_1 FILLER_31_355 ();
 sg13g2_fill_1 FILLER_31_360 ();
 sg13g2_fill_1 FILLER_31_366 ();
 sg13g2_fill_2 FILLER_31_377 ();
 sg13g2_fill_1 FILLER_31_379 ();
 sg13g2_decap_4 FILLER_31_388 ();
 sg13g2_fill_2 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_411 ();
 sg13g2_decap_8 FILLER_31_418 ();
 sg13g2_decap_4 FILLER_31_425 ();
 sg13g2_fill_1 FILLER_31_429 ();
 sg13g2_fill_1 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_27 ();
 sg13g2_fill_2 FILLER_32_33 ();
 sg13g2_fill_2 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_73 ();
 sg13g2_fill_1 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_85 ();
 sg13g2_fill_1 FILLER_32_90 ();
 sg13g2_fill_1 FILLER_32_101 ();
 sg13g2_decap_8 FILLER_32_108 ();
 sg13g2_decap_4 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_124 ();
 sg13g2_fill_2 FILLER_32_129 ();
 sg13g2_fill_1 FILLER_32_131 ();
 sg13g2_decap_4 FILLER_32_151 ();
 sg13g2_fill_2 FILLER_32_155 ();
 sg13g2_fill_2 FILLER_32_166 ();
 sg13g2_fill_1 FILLER_32_177 ();
 sg13g2_decap_8 FILLER_32_199 ();
 sg13g2_decap_8 FILLER_32_206 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_fill_2 FILLER_32_235 ();
 sg13g2_fill_1 FILLER_32_237 ();
 sg13g2_fill_1 FILLER_32_247 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_4 FILLER_32_277 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_decap_4 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_300 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_311 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_decap_4 FILLER_32_335 ();
 sg13g2_fill_1 FILLER_32_339 ();
 sg13g2_fill_2 FILLER_32_345 ();
 sg13g2_fill_1 FILLER_32_347 ();
 sg13g2_fill_1 FILLER_32_357 ();
 sg13g2_fill_1 FILLER_32_362 ();
 sg13g2_decap_4 FILLER_32_373 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_383 ();
 sg13g2_fill_2 FILLER_32_388 ();
 sg13g2_fill_2 FILLER_32_404 ();
 sg13g2_decap_8 FILLER_32_415 ();
 sg13g2_decap_8 FILLER_32_422 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_fill_1 FILLER_33_14 ();
 sg13g2_fill_2 FILLER_33_24 ();
 sg13g2_decap_4 FILLER_33_34 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_2 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_92 ();
 sg13g2_decap_4 FILLER_33_99 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_131 ();
 sg13g2_fill_1 FILLER_33_136 ();
 sg13g2_decap_4 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_151 ();
 sg13g2_fill_1 FILLER_33_158 ();
 sg13g2_decap_4 FILLER_33_164 ();
 sg13g2_fill_1 FILLER_33_168 ();
 sg13g2_decap_4 FILLER_33_174 ();
 sg13g2_fill_1 FILLER_33_178 ();
 sg13g2_fill_1 FILLER_33_183 ();
 sg13g2_fill_2 FILLER_33_189 ();
 sg13g2_decap_4 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_199 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_fill_2 FILLER_33_217 ();
 sg13g2_fill_1 FILLER_33_219 ();
 sg13g2_fill_2 FILLER_33_233 ();
 sg13g2_fill_2 FILLER_33_252 ();
 sg13g2_fill_1 FILLER_33_258 ();
 sg13g2_fill_1 FILLER_33_264 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_fill_1 FILLER_33_287 ();
 sg13g2_fill_2 FILLER_33_292 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_decap_4 FILLER_33_312 ();
 sg13g2_fill_1 FILLER_33_316 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_339 ();
 sg13g2_fill_1 FILLER_33_341 ();
 sg13g2_decap_4 FILLER_33_352 ();
 sg13g2_fill_2 FILLER_33_356 ();
 sg13g2_fill_2 FILLER_33_363 ();
 sg13g2_fill_1 FILLER_33_370 ();
 sg13g2_fill_2 FILLER_33_380 ();
 sg13g2_fill_2 FILLER_33_386 ();
 sg13g2_fill_2 FILLER_33_391 ();
 sg13g2_fill_1 FILLER_33_403 ();
 sg13g2_fill_1 FILLER_33_414 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_decap_8 FILLER_34_42 ();
 sg13g2_decap_8 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_56 ();
 sg13g2_fill_2 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_77 ();
 sg13g2_decap_4 FILLER_34_83 ();
 sg13g2_fill_1 FILLER_34_87 ();
 sg13g2_fill_1 FILLER_34_103 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_143 ();
 sg13g2_decap_8 FILLER_34_150 ();
 sg13g2_decap_8 FILLER_34_157 ();
 sg13g2_decap_8 FILLER_34_164 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_204 ();
 sg13g2_decap_8 FILLER_34_212 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_1 FILLER_34_238 ();
 sg13g2_decap_4 FILLER_34_245 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_fill_1 FILLER_34_261 ();
 sg13g2_fill_1 FILLER_34_266 ();
 sg13g2_fill_2 FILLER_34_280 ();
 sg13g2_fill_1 FILLER_34_282 ();
 sg13g2_fill_1 FILLER_34_288 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_331 ();
 sg13g2_decap_4 FILLER_34_338 ();
 sg13g2_fill_2 FILLER_34_346 ();
 sg13g2_fill_1 FILLER_34_353 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_fill_2 FILLER_34_381 ();
 sg13g2_fill_2 FILLER_34_393 ();
 sg13g2_fill_2 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_402 ();
 sg13g2_fill_2 FILLER_34_408 ();
 sg13g2_fill_1 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_fill_1 FILLER_35_32 ();
 sg13g2_decap_8 FILLER_35_51 ();
 sg13g2_fill_2 FILLER_35_62 ();
 sg13g2_fill_2 FILLER_35_68 ();
 sg13g2_fill_1 FILLER_35_79 ();
 sg13g2_fill_2 FILLER_35_89 ();
 sg13g2_decap_8 FILLER_35_104 ();
 sg13g2_decap_4 FILLER_35_111 ();
 sg13g2_decap_8 FILLER_35_123 ();
 sg13g2_fill_2 FILLER_35_160 ();
 sg13g2_decap_8 FILLER_35_165 ();
 sg13g2_decap_8 FILLER_35_172 ();
 sg13g2_decap_8 FILLER_35_179 ();
 sg13g2_decap_8 FILLER_35_186 ();
 sg13g2_decap_8 FILLER_35_193 ();
 sg13g2_decap_4 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_204 ();
 sg13g2_fill_2 FILLER_35_219 ();
 sg13g2_fill_1 FILLER_35_221 ();
 sg13g2_decap_4 FILLER_35_227 ();
 sg13g2_decap_4 FILLER_35_245 ();
 sg13g2_decap_4 FILLER_35_262 ();
 sg13g2_decap_4 FILLER_35_270 ();
 sg13g2_fill_2 FILLER_35_286 ();
 sg13g2_fill_1 FILLER_35_288 ();
 sg13g2_fill_2 FILLER_35_297 ();
 sg13g2_decap_4 FILLER_35_312 ();
 sg13g2_fill_2 FILLER_35_316 ();
 sg13g2_fill_2 FILLER_35_327 ();
 sg13g2_fill_1 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_339 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_365 ();
 sg13g2_decap_4 FILLER_35_381 ();
 sg13g2_decap_4 FILLER_35_389 ();
 sg13g2_fill_2 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_399 ();
 sg13g2_fill_2 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_decap_4 FILLER_35_426 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_2 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_33 ();
 sg13g2_fill_1 FILLER_36_39 ();
 sg13g2_decap_8 FILLER_36_43 ();
 sg13g2_fill_2 FILLER_36_50 ();
 sg13g2_fill_1 FILLER_36_52 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_63 ();
 sg13g2_fill_1 FILLER_36_67 ();
 sg13g2_fill_2 FILLER_36_78 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_1 FILLER_36_116 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_4 FILLER_36_140 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_decap_8 FILLER_36_188 ();
 sg13g2_decap_8 FILLER_36_199 ();
 sg13g2_decap_8 FILLER_36_206 ();
 sg13g2_decap_8 FILLER_36_213 ();
 sg13g2_fill_1 FILLER_36_220 ();
 sg13g2_decap_8 FILLER_36_226 ();
 sg13g2_decap_8 FILLER_36_233 ();
 sg13g2_fill_2 FILLER_36_240 ();
 sg13g2_fill_1 FILLER_36_242 ();
 sg13g2_fill_1 FILLER_36_256 ();
 sg13g2_fill_1 FILLER_36_262 ();
 sg13g2_fill_1 FILLER_36_272 ();
 sg13g2_fill_1 FILLER_36_291 ();
 sg13g2_decap_4 FILLER_36_300 ();
 sg13g2_fill_1 FILLER_36_304 ();
 sg13g2_fill_1 FILLER_36_310 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_fill_2 FILLER_36_322 ();
 sg13g2_decap_4 FILLER_36_337 ();
 sg13g2_fill_1 FILLER_36_341 ();
 sg13g2_decap_4 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_380 ();
 sg13g2_fill_1 FILLER_36_382 ();
 sg13g2_decap_4 FILLER_36_387 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_decap_4 FILLER_36_396 ();
 sg13g2_fill_1 FILLER_36_400 ();
 sg13g2_decap_8 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_36_414 ();
 sg13g2_decap_8 FILLER_36_421 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_75 ();
 sg13g2_decap_4 FILLER_37_82 ();
 sg13g2_fill_2 FILLER_37_86 ();
 sg13g2_decap_4 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_128 ();
 sg13g2_fill_2 FILLER_37_166 ();
 sg13g2_fill_2 FILLER_37_185 ();
 sg13g2_fill_1 FILLER_37_187 ();
 sg13g2_decap_8 FILLER_37_192 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_decap_4 FILLER_37_204 ();
 sg13g2_fill_1 FILLER_37_208 ();
 sg13g2_decap_8 FILLER_37_213 ();
 sg13g2_decap_8 FILLER_37_220 ();
 sg13g2_decap_8 FILLER_37_227 ();
 sg13g2_fill_2 FILLER_37_234 ();
 sg13g2_fill_1 FILLER_37_236 ();
 sg13g2_fill_1 FILLER_37_250 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_decap_4 FILLER_37_260 ();
 sg13g2_fill_2 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_278 ();
 sg13g2_fill_1 FILLER_37_284 ();
 sg13g2_decap_4 FILLER_37_298 ();
 sg13g2_fill_2 FILLER_37_306 ();
 sg13g2_fill_1 FILLER_37_308 ();
 sg13g2_decap_8 FILLER_37_322 ();
 sg13g2_fill_2 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_393 ();
 sg13g2_decap_8 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_405 ();
 sg13g2_fill_1 FILLER_37_407 ();
 sg13g2_decap_8 FILLER_37_421 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_fill_2 FILLER_38_21 ();
 sg13g2_fill_1 FILLER_38_23 ();
 sg13g2_fill_1 FILLER_38_27 ();
 sg13g2_decap_4 FILLER_38_67 ();
 sg13g2_fill_1 FILLER_38_103 ();
 sg13g2_fill_2 FILLER_38_132 ();
 sg13g2_decap_4 FILLER_38_138 ();
 sg13g2_decap_4 FILLER_38_146 ();
 sg13g2_fill_2 FILLER_38_154 ();
 sg13g2_fill_1 FILLER_38_156 ();
 sg13g2_fill_1 FILLER_38_171 ();
 sg13g2_fill_2 FILLER_38_209 ();
 sg13g2_fill_1 FILLER_38_211 ();
 sg13g2_decap_4 FILLER_38_216 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_fill_1 FILLER_38_231 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_2 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_252 ();
 sg13g2_fill_1 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_272 ();
 sg13g2_decap_8 FILLER_38_279 ();
 sg13g2_decap_8 FILLER_38_286 ();
 sg13g2_decap_8 FILLER_38_293 ();
 sg13g2_decap_8 FILLER_38_300 ();
 sg13g2_decap_8 FILLER_38_307 ();
 sg13g2_decap_8 FILLER_38_314 ();
 sg13g2_decap_8 FILLER_38_321 ();
 sg13g2_decap_4 FILLER_38_328 ();
 sg13g2_fill_1 FILLER_38_332 ();
 sg13g2_fill_2 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_348 ();
 sg13g2_fill_1 FILLER_38_350 ();
 sg13g2_fill_2 FILLER_38_355 ();
 sg13g2_fill_1 FILLER_38_357 ();
 sg13g2_decap_4 FILLER_38_362 ();
 sg13g2_decap_4 FILLER_38_370 ();
 sg13g2_fill_2 FILLER_38_386 ();
 sg13g2_fill_1 FILLER_38_388 ();
 sg13g2_decap_4 FILLER_38_393 ();
 sg13g2_decap_8 FILLER_38_401 ();
 sg13g2_decap_8 FILLER_38_408 ();
 sg13g2_decap_8 FILLER_38_415 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_429 ();
endmodule
