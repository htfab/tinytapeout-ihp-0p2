module tt_um_froith_goldcrest (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire clknet_leaf_0_clk;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire _09004_;
 wire _09005_;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire net2007;
 wire _13703_;
 wire _13704_;
 wire \top_ihp.gpio_o_1 ;
 wire \top_ihp.gpio_o_2 ;
 wire \top_ihp.gpio_o_3 ;
 wire \top_ihp.gpio_o_4 ;
 wire \top_ihp.oisc.decoder.decoded[0] ;
 wire \top_ihp.oisc.decoder.decoded[10] ;
 wire \top_ihp.oisc.decoder.decoded[11] ;
 wire \top_ihp.oisc.decoder.decoded[12] ;
 wire \top_ihp.oisc.decoder.decoded[13] ;
 wire \top_ihp.oisc.decoder.decoded[14] ;
 wire \top_ihp.oisc.decoder.decoded[15] ;
 wire \top_ihp.oisc.decoder.decoded[1] ;
 wire \top_ihp.oisc.decoder.decoded[2] ;
 wire \top_ihp.oisc.decoder.decoded[3] ;
 wire \top_ihp.oisc.decoder.decoded[4] ;
 wire \top_ihp.oisc.decoder.decoded[5] ;
 wire \top_ihp.oisc.decoder.decoded[6] ;
 wire \top_ihp.oisc.decoder.decoded[7] ;
 wire \top_ihp.oisc.decoder.instruction[10] ;
 wire \top_ihp.oisc.decoder.instruction[11] ;
 wire \top_ihp.oisc.decoder.instruction[12] ;
 wire \top_ihp.oisc.decoder.instruction[13] ;
 wire \top_ihp.oisc.decoder.instruction[14] ;
 wire \top_ihp.oisc.decoder.instruction[15] ;
 wire \top_ihp.oisc.decoder.instruction[16] ;
 wire \top_ihp.oisc.decoder.instruction[17] ;
 wire \top_ihp.oisc.decoder.instruction[18] ;
 wire \top_ihp.oisc.decoder.instruction[19] ;
 wire \top_ihp.oisc.decoder.instruction[20] ;
 wire \top_ihp.oisc.decoder.instruction[21] ;
 wire \top_ihp.oisc.decoder.instruction[22] ;
 wire \top_ihp.oisc.decoder.instruction[23] ;
 wire \top_ihp.oisc.decoder.instruction[24] ;
 wire \top_ihp.oisc.decoder.instruction[25] ;
 wire \top_ihp.oisc.decoder.instruction[26] ;
 wire \top_ihp.oisc.decoder.instruction[27] ;
 wire \top_ihp.oisc.decoder.instruction[28] ;
 wire \top_ihp.oisc.decoder.instruction[29] ;
 wire \top_ihp.oisc.decoder.instruction[30] ;
 wire \top_ihp.oisc.decoder.instruction[31] ;
 wire \top_ihp.oisc.decoder.instruction[7] ;
 wire \top_ihp.oisc.decoder.instruction[8] ;
 wire \top_ihp.oisc.decoder.instruction[9] ;
 wire \top_ihp.oisc.mem_addr_lowbits[0] ;
 wire \top_ihp.oisc.mem_addr_lowbits[1] ;
 wire \top_ihp.oisc.micro_op[0] ;
 wire \top_ihp.oisc.micro_op[10] ;
 wire \top_ihp.oisc.micro_op[11] ;
 wire \top_ihp.oisc.micro_op[12] ;
 wire \top_ihp.oisc.micro_op[13] ;
 wire \top_ihp.oisc.micro_op[14] ;
 wire \top_ihp.oisc.micro_op[15] ;
 wire \top_ihp.oisc.micro_op[1] ;
 wire \top_ihp.oisc.micro_op[2] ;
 wire \top_ihp.oisc.micro_op[3] ;
 wire \top_ihp.oisc.micro_op[4] ;
 wire \top_ihp.oisc.micro_op[5] ;
 wire \top_ihp.oisc.micro_op[8] ;
 wire \top_ihp.oisc.micro_op[9] ;
 wire \top_ihp.oisc.micro_pc[0] ;
 wire \top_ihp.oisc.micro_pc[1] ;
 wire \top_ihp.oisc.micro_pc[2] ;
 wire \top_ihp.oisc.micro_pc[3] ;
 wire \top_ihp.oisc.micro_pc[4] ;
 wire \top_ihp.oisc.micro_pc[5] ;
 wire \top_ihp.oisc.micro_pc[6] ;
 wire \top_ihp.oisc.micro_pc[7] ;
 wire \top_ihp.oisc.micro_res_addr[0] ;
 wire \top_ihp.oisc.micro_res_addr[1] ;
 wire \top_ihp.oisc.micro_res_addr[2] ;
 wire \top_ihp.oisc.micro_res_addr[3] ;
 wire \top_ihp.oisc.micro_state[0] ;
 wire \top_ihp.oisc.micro_state[1] ;
 wire \top_ihp.oisc.micro_state[2] ;
 wire \top_ihp.oisc.op_a[0] ;
 wire \top_ihp.oisc.op_a[10] ;
 wire \top_ihp.oisc.op_a[11] ;
 wire \top_ihp.oisc.op_a[12] ;
 wire \top_ihp.oisc.op_a[13] ;
 wire \top_ihp.oisc.op_a[14] ;
 wire \top_ihp.oisc.op_a[15] ;
 wire \top_ihp.oisc.op_a[16] ;
 wire \top_ihp.oisc.op_a[17] ;
 wire \top_ihp.oisc.op_a[18] ;
 wire \top_ihp.oisc.op_a[19] ;
 wire \top_ihp.oisc.op_a[1] ;
 wire \top_ihp.oisc.op_a[20] ;
 wire \top_ihp.oisc.op_a[21] ;
 wire \top_ihp.oisc.op_a[22] ;
 wire \top_ihp.oisc.op_a[23] ;
 wire \top_ihp.oisc.op_a[24] ;
 wire \top_ihp.oisc.op_a[25] ;
 wire \top_ihp.oisc.op_a[26] ;
 wire \top_ihp.oisc.op_a[27] ;
 wire \top_ihp.oisc.op_a[28] ;
 wire \top_ihp.oisc.op_a[29] ;
 wire \top_ihp.oisc.op_a[2] ;
 wire \top_ihp.oisc.op_a[30] ;
 wire \top_ihp.oisc.op_a[31] ;
 wire \top_ihp.oisc.op_a[3] ;
 wire \top_ihp.oisc.op_a[4] ;
 wire \top_ihp.oisc.op_a[5] ;
 wire \top_ihp.oisc.op_a[6] ;
 wire \top_ihp.oisc.op_a[7] ;
 wire \top_ihp.oisc.op_a[8] ;
 wire \top_ihp.oisc.op_a[9] ;
 wire \top_ihp.oisc.op_b[0] ;
 wire \top_ihp.oisc.op_b[10] ;
 wire \top_ihp.oisc.op_b[11] ;
 wire \top_ihp.oisc.op_b[12] ;
 wire \top_ihp.oisc.op_b[13] ;
 wire \top_ihp.oisc.op_b[14] ;
 wire \top_ihp.oisc.op_b[15] ;
 wire \top_ihp.oisc.op_b[16] ;
 wire \top_ihp.oisc.op_b[17] ;
 wire \top_ihp.oisc.op_b[18] ;
 wire \top_ihp.oisc.op_b[19] ;
 wire \top_ihp.oisc.op_b[1] ;
 wire \top_ihp.oisc.op_b[20] ;
 wire \top_ihp.oisc.op_b[21] ;
 wire \top_ihp.oisc.op_b[22] ;
 wire \top_ihp.oisc.op_b[23] ;
 wire \top_ihp.oisc.op_b[24] ;
 wire \top_ihp.oisc.op_b[25] ;
 wire \top_ihp.oisc.op_b[26] ;
 wire \top_ihp.oisc.op_b[27] ;
 wire \top_ihp.oisc.op_b[28] ;
 wire \top_ihp.oisc.op_b[29] ;
 wire \top_ihp.oisc.op_b[2] ;
 wire \top_ihp.oisc.op_b[30] ;
 wire \top_ihp.oisc.op_b[31] ;
 wire \top_ihp.oisc.op_b[3] ;
 wire \top_ihp.oisc.op_b[4] ;
 wire \top_ihp.oisc.op_b[5] ;
 wire \top_ihp.oisc.op_b[6] ;
 wire \top_ihp.oisc.op_b[7] ;
 wire \top_ihp.oisc.op_b[8] ;
 wire \top_ihp.oisc.op_b[9] ;
 wire \top_ihp.oisc.reg_rb[0] ;
 wire \top_ihp.oisc.reg_rb[1] ;
 wire \top_ihp.oisc.reg_rb[2] ;
 wire \top_ihp.oisc.reg_rb[3] ;
 wire \top_ihp.oisc.regs[0][0] ;
 wire \top_ihp.oisc.regs[0][10] ;
 wire \top_ihp.oisc.regs[0][11] ;
 wire \top_ihp.oisc.regs[0][12] ;
 wire \top_ihp.oisc.regs[0][13] ;
 wire \top_ihp.oisc.regs[0][14] ;
 wire \top_ihp.oisc.regs[0][15] ;
 wire \top_ihp.oisc.regs[0][16] ;
 wire \top_ihp.oisc.regs[0][17] ;
 wire \top_ihp.oisc.regs[0][18] ;
 wire \top_ihp.oisc.regs[0][19] ;
 wire \top_ihp.oisc.regs[0][1] ;
 wire \top_ihp.oisc.regs[0][20] ;
 wire \top_ihp.oisc.regs[0][21] ;
 wire \top_ihp.oisc.regs[0][22] ;
 wire \top_ihp.oisc.regs[0][23] ;
 wire \top_ihp.oisc.regs[0][24] ;
 wire \top_ihp.oisc.regs[0][25] ;
 wire \top_ihp.oisc.regs[0][26] ;
 wire \top_ihp.oisc.regs[0][27] ;
 wire \top_ihp.oisc.regs[0][28] ;
 wire \top_ihp.oisc.regs[0][29] ;
 wire \top_ihp.oisc.regs[0][2] ;
 wire \top_ihp.oisc.regs[0][30] ;
 wire \top_ihp.oisc.regs[0][31] ;
 wire \top_ihp.oisc.regs[0][3] ;
 wire \top_ihp.oisc.regs[0][4] ;
 wire \top_ihp.oisc.regs[0][5] ;
 wire \top_ihp.oisc.regs[0][6] ;
 wire \top_ihp.oisc.regs[0][7] ;
 wire \top_ihp.oisc.regs[0][8] ;
 wire \top_ihp.oisc.regs[0][9] ;
 wire \top_ihp.oisc.regs[10][0] ;
 wire \top_ihp.oisc.regs[10][10] ;
 wire \top_ihp.oisc.regs[10][11] ;
 wire \top_ihp.oisc.regs[10][12] ;
 wire \top_ihp.oisc.regs[10][13] ;
 wire \top_ihp.oisc.regs[10][14] ;
 wire \top_ihp.oisc.regs[10][15] ;
 wire \top_ihp.oisc.regs[10][16] ;
 wire \top_ihp.oisc.regs[10][17] ;
 wire \top_ihp.oisc.regs[10][18] ;
 wire \top_ihp.oisc.regs[10][19] ;
 wire \top_ihp.oisc.regs[10][1] ;
 wire \top_ihp.oisc.regs[10][20] ;
 wire \top_ihp.oisc.regs[10][21] ;
 wire \top_ihp.oisc.regs[10][22] ;
 wire \top_ihp.oisc.regs[10][23] ;
 wire \top_ihp.oisc.regs[10][24] ;
 wire \top_ihp.oisc.regs[10][25] ;
 wire \top_ihp.oisc.regs[10][26] ;
 wire \top_ihp.oisc.regs[10][27] ;
 wire \top_ihp.oisc.regs[10][28] ;
 wire \top_ihp.oisc.regs[10][29] ;
 wire \top_ihp.oisc.regs[10][2] ;
 wire \top_ihp.oisc.regs[10][30] ;
 wire \top_ihp.oisc.regs[10][31] ;
 wire \top_ihp.oisc.regs[10][3] ;
 wire \top_ihp.oisc.regs[10][4] ;
 wire \top_ihp.oisc.regs[10][5] ;
 wire \top_ihp.oisc.regs[10][6] ;
 wire \top_ihp.oisc.regs[10][7] ;
 wire \top_ihp.oisc.regs[10][8] ;
 wire \top_ihp.oisc.regs[10][9] ;
 wire \top_ihp.oisc.regs[11][0] ;
 wire \top_ihp.oisc.regs[11][10] ;
 wire \top_ihp.oisc.regs[11][11] ;
 wire \top_ihp.oisc.regs[11][12] ;
 wire \top_ihp.oisc.regs[11][13] ;
 wire \top_ihp.oisc.regs[11][14] ;
 wire \top_ihp.oisc.regs[11][15] ;
 wire \top_ihp.oisc.regs[11][16] ;
 wire \top_ihp.oisc.regs[11][17] ;
 wire \top_ihp.oisc.regs[11][18] ;
 wire \top_ihp.oisc.regs[11][19] ;
 wire \top_ihp.oisc.regs[11][1] ;
 wire \top_ihp.oisc.regs[11][20] ;
 wire \top_ihp.oisc.regs[11][21] ;
 wire \top_ihp.oisc.regs[11][22] ;
 wire \top_ihp.oisc.regs[11][23] ;
 wire \top_ihp.oisc.regs[11][24] ;
 wire \top_ihp.oisc.regs[11][25] ;
 wire \top_ihp.oisc.regs[11][26] ;
 wire \top_ihp.oisc.regs[11][27] ;
 wire \top_ihp.oisc.regs[11][28] ;
 wire \top_ihp.oisc.regs[11][29] ;
 wire \top_ihp.oisc.regs[11][2] ;
 wire \top_ihp.oisc.regs[11][30] ;
 wire \top_ihp.oisc.regs[11][31] ;
 wire \top_ihp.oisc.regs[11][3] ;
 wire \top_ihp.oisc.regs[11][4] ;
 wire \top_ihp.oisc.regs[11][5] ;
 wire \top_ihp.oisc.regs[11][6] ;
 wire \top_ihp.oisc.regs[11][7] ;
 wire \top_ihp.oisc.regs[11][8] ;
 wire \top_ihp.oisc.regs[11][9] ;
 wire \top_ihp.oisc.regs[12][0] ;
 wire \top_ihp.oisc.regs[12][10] ;
 wire \top_ihp.oisc.regs[12][11] ;
 wire \top_ihp.oisc.regs[12][12] ;
 wire \top_ihp.oisc.regs[12][13] ;
 wire \top_ihp.oisc.regs[12][14] ;
 wire \top_ihp.oisc.regs[12][15] ;
 wire \top_ihp.oisc.regs[12][16] ;
 wire \top_ihp.oisc.regs[12][17] ;
 wire \top_ihp.oisc.regs[12][18] ;
 wire \top_ihp.oisc.regs[12][19] ;
 wire \top_ihp.oisc.regs[12][1] ;
 wire \top_ihp.oisc.regs[12][20] ;
 wire \top_ihp.oisc.regs[12][21] ;
 wire \top_ihp.oisc.regs[12][22] ;
 wire \top_ihp.oisc.regs[12][23] ;
 wire \top_ihp.oisc.regs[12][24] ;
 wire \top_ihp.oisc.regs[12][25] ;
 wire \top_ihp.oisc.regs[12][26] ;
 wire \top_ihp.oisc.regs[12][27] ;
 wire \top_ihp.oisc.regs[12][28] ;
 wire \top_ihp.oisc.regs[12][29] ;
 wire \top_ihp.oisc.regs[12][2] ;
 wire \top_ihp.oisc.regs[12][30] ;
 wire \top_ihp.oisc.regs[12][31] ;
 wire \top_ihp.oisc.regs[12][3] ;
 wire \top_ihp.oisc.regs[12][4] ;
 wire \top_ihp.oisc.regs[12][5] ;
 wire \top_ihp.oisc.regs[12][6] ;
 wire \top_ihp.oisc.regs[12][7] ;
 wire \top_ihp.oisc.regs[12][8] ;
 wire \top_ihp.oisc.regs[12][9] ;
 wire \top_ihp.oisc.regs[13][0] ;
 wire \top_ihp.oisc.regs[13][10] ;
 wire \top_ihp.oisc.regs[13][11] ;
 wire \top_ihp.oisc.regs[13][12] ;
 wire \top_ihp.oisc.regs[13][13] ;
 wire \top_ihp.oisc.regs[13][14] ;
 wire \top_ihp.oisc.regs[13][15] ;
 wire \top_ihp.oisc.regs[13][16] ;
 wire \top_ihp.oisc.regs[13][17] ;
 wire \top_ihp.oisc.regs[13][18] ;
 wire \top_ihp.oisc.regs[13][19] ;
 wire \top_ihp.oisc.regs[13][1] ;
 wire \top_ihp.oisc.regs[13][20] ;
 wire \top_ihp.oisc.regs[13][21] ;
 wire \top_ihp.oisc.regs[13][22] ;
 wire \top_ihp.oisc.regs[13][23] ;
 wire \top_ihp.oisc.regs[13][24] ;
 wire \top_ihp.oisc.regs[13][25] ;
 wire \top_ihp.oisc.regs[13][26] ;
 wire \top_ihp.oisc.regs[13][27] ;
 wire \top_ihp.oisc.regs[13][28] ;
 wire \top_ihp.oisc.regs[13][29] ;
 wire \top_ihp.oisc.regs[13][2] ;
 wire \top_ihp.oisc.regs[13][30] ;
 wire \top_ihp.oisc.regs[13][31] ;
 wire \top_ihp.oisc.regs[13][3] ;
 wire \top_ihp.oisc.regs[13][4] ;
 wire \top_ihp.oisc.regs[13][5] ;
 wire \top_ihp.oisc.regs[13][6] ;
 wire \top_ihp.oisc.regs[13][7] ;
 wire \top_ihp.oisc.regs[13][8] ;
 wire \top_ihp.oisc.regs[13][9] ;
 wire \top_ihp.oisc.regs[14][0] ;
 wire \top_ihp.oisc.regs[14][10] ;
 wire \top_ihp.oisc.regs[14][11] ;
 wire \top_ihp.oisc.regs[14][12] ;
 wire \top_ihp.oisc.regs[14][13] ;
 wire \top_ihp.oisc.regs[14][14] ;
 wire \top_ihp.oisc.regs[14][15] ;
 wire \top_ihp.oisc.regs[14][16] ;
 wire \top_ihp.oisc.regs[14][17] ;
 wire \top_ihp.oisc.regs[14][18] ;
 wire \top_ihp.oisc.regs[14][19] ;
 wire \top_ihp.oisc.regs[14][1] ;
 wire \top_ihp.oisc.regs[14][20] ;
 wire \top_ihp.oisc.regs[14][21] ;
 wire \top_ihp.oisc.regs[14][22] ;
 wire \top_ihp.oisc.regs[14][23] ;
 wire \top_ihp.oisc.regs[14][24] ;
 wire \top_ihp.oisc.regs[14][25] ;
 wire \top_ihp.oisc.regs[14][26] ;
 wire \top_ihp.oisc.regs[14][27] ;
 wire \top_ihp.oisc.regs[14][28] ;
 wire \top_ihp.oisc.regs[14][29] ;
 wire \top_ihp.oisc.regs[14][2] ;
 wire \top_ihp.oisc.regs[14][30] ;
 wire \top_ihp.oisc.regs[14][31] ;
 wire \top_ihp.oisc.regs[14][3] ;
 wire \top_ihp.oisc.regs[14][4] ;
 wire \top_ihp.oisc.regs[14][5] ;
 wire \top_ihp.oisc.regs[14][6] ;
 wire \top_ihp.oisc.regs[14][7] ;
 wire \top_ihp.oisc.regs[14][8] ;
 wire \top_ihp.oisc.regs[14][9] ;
 wire \top_ihp.oisc.regs[15][0] ;
 wire \top_ihp.oisc.regs[15][10] ;
 wire \top_ihp.oisc.regs[15][11] ;
 wire \top_ihp.oisc.regs[15][12] ;
 wire \top_ihp.oisc.regs[15][13] ;
 wire \top_ihp.oisc.regs[15][14] ;
 wire \top_ihp.oisc.regs[15][15] ;
 wire \top_ihp.oisc.regs[15][16] ;
 wire \top_ihp.oisc.regs[15][17] ;
 wire \top_ihp.oisc.regs[15][18] ;
 wire \top_ihp.oisc.regs[15][19] ;
 wire \top_ihp.oisc.regs[15][1] ;
 wire \top_ihp.oisc.regs[15][20] ;
 wire \top_ihp.oisc.regs[15][21] ;
 wire \top_ihp.oisc.regs[15][22] ;
 wire \top_ihp.oisc.regs[15][23] ;
 wire \top_ihp.oisc.regs[15][24] ;
 wire \top_ihp.oisc.regs[15][25] ;
 wire \top_ihp.oisc.regs[15][26] ;
 wire \top_ihp.oisc.regs[15][27] ;
 wire \top_ihp.oisc.regs[15][28] ;
 wire \top_ihp.oisc.regs[15][29] ;
 wire \top_ihp.oisc.regs[15][2] ;
 wire \top_ihp.oisc.regs[15][30] ;
 wire \top_ihp.oisc.regs[15][31] ;
 wire \top_ihp.oisc.regs[15][3] ;
 wire \top_ihp.oisc.regs[15][4] ;
 wire \top_ihp.oisc.regs[15][5] ;
 wire \top_ihp.oisc.regs[15][6] ;
 wire \top_ihp.oisc.regs[15][7] ;
 wire \top_ihp.oisc.regs[15][8] ;
 wire \top_ihp.oisc.regs[15][9] ;
 wire \top_ihp.oisc.regs[16][0] ;
 wire \top_ihp.oisc.regs[16][10] ;
 wire \top_ihp.oisc.regs[16][11] ;
 wire \top_ihp.oisc.regs[16][12] ;
 wire \top_ihp.oisc.regs[16][13] ;
 wire \top_ihp.oisc.regs[16][14] ;
 wire \top_ihp.oisc.regs[16][15] ;
 wire \top_ihp.oisc.regs[16][16] ;
 wire \top_ihp.oisc.regs[16][17] ;
 wire \top_ihp.oisc.regs[16][18] ;
 wire \top_ihp.oisc.regs[16][19] ;
 wire \top_ihp.oisc.regs[16][1] ;
 wire \top_ihp.oisc.regs[16][20] ;
 wire \top_ihp.oisc.regs[16][21] ;
 wire \top_ihp.oisc.regs[16][22] ;
 wire \top_ihp.oisc.regs[16][23] ;
 wire \top_ihp.oisc.regs[16][24] ;
 wire \top_ihp.oisc.regs[16][25] ;
 wire \top_ihp.oisc.regs[16][26] ;
 wire \top_ihp.oisc.regs[16][27] ;
 wire \top_ihp.oisc.regs[16][28] ;
 wire \top_ihp.oisc.regs[16][29] ;
 wire \top_ihp.oisc.regs[16][2] ;
 wire \top_ihp.oisc.regs[16][30] ;
 wire \top_ihp.oisc.regs[16][31] ;
 wire \top_ihp.oisc.regs[16][3] ;
 wire \top_ihp.oisc.regs[16][4] ;
 wire \top_ihp.oisc.regs[16][5] ;
 wire \top_ihp.oisc.regs[16][6] ;
 wire \top_ihp.oisc.regs[16][7] ;
 wire \top_ihp.oisc.regs[16][8] ;
 wire \top_ihp.oisc.regs[16][9] ;
 wire \top_ihp.oisc.regs[17][0] ;
 wire \top_ihp.oisc.regs[17][10] ;
 wire \top_ihp.oisc.regs[17][11] ;
 wire \top_ihp.oisc.regs[17][12] ;
 wire \top_ihp.oisc.regs[17][13] ;
 wire \top_ihp.oisc.regs[17][14] ;
 wire \top_ihp.oisc.regs[17][15] ;
 wire \top_ihp.oisc.regs[17][16] ;
 wire \top_ihp.oisc.regs[17][17] ;
 wire \top_ihp.oisc.regs[17][18] ;
 wire \top_ihp.oisc.regs[17][19] ;
 wire \top_ihp.oisc.regs[17][1] ;
 wire \top_ihp.oisc.regs[17][20] ;
 wire \top_ihp.oisc.regs[17][21] ;
 wire \top_ihp.oisc.regs[17][22] ;
 wire \top_ihp.oisc.regs[17][23] ;
 wire \top_ihp.oisc.regs[17][24] ;
 wire \top_ihp.oisc.regs[17][25] ;
 wire \top_ihp.oisc.regs[17][26] ;
 wire \top_ihp.oisc.regs[17][27] ;
 wire \top_ihp.oisc.regs[17][28] ;
 wire \top_ihp.oisc.regs[17][29] ;
 wire \top_ihp.oisc.regs[17][2] ;
 wire \top_ihp.oisc.regs[17][30] ;
 wire \top_ihp.oisc.regs[17][31] ;
 wire \top_ihp.oisc.regs[17][3] ;
 wire \top_ihp.oisc.regs[17][4] ;
 wire \top_ihp.oisc.regs[17][5] ;
 wire \top_ihp.oisc.regs[17][6] ;
 wire \top_ihp.oisc.regs[17][7] ;
 wire \top_ihp.oisc.regs[17][8] ;
 wire \top_ihp.oisc.regs[17][9] ;
 wire \top_ihp.oisc.regs[18][0] ;
 wire \top_ihp.oisc.regs[18][10] ;
 wire \top_ihp.oisc.regs[18][11] ;
 wire \top_ihp.oisc.regs[18][12] ;
 wire \top_ihp.oisc.regs[18][13] ;
 wire \top_ihp.oisc.regs[18][14] ;
 wire \top_ihp.oisc.regs[18][15] ;
 wire \top_ihp.oisc.regs[18][16] ;
 wire \top_ihp.oisc.regs[18][17] ;
 wire \top_ihp.oisc.regs[18][18] ;
 wire \top_ihp.oisc.regs[18][19] ;
 wire \top_ihp.oisc.regs[18][1] ;
 wire \top_ihp.oisc.regs[18][20] ;
 wire \top_ihp.oisc.regs[18][21] ;
 wire \top_ihp.oisc.regs[18][22] ;
 wire \top_ihp.oisc.regs[18][23] ;
 wire \top_ihp.oisc.regs[18][24] ;
 wire \top_ihp.oisc.regs[18][25] ;
 wire \top_ihp.oisc.regs[18][26] ;
 wire \top_ihp.oisc.regs[18][27] ;
 wire \top_ihp.oisc.regs[18][28] ;
 wire \top_ihp.oisc.regs[18][29] ;
 wire \top_ihp.oisc.regs[18][2] ;
 wire \top_ihp.oisc.regs[18][30] ;
 wire \top_ihp.oisc.regs[18][31] ;
 wire \top_ihp.oisc.regs[18][3] ;
 wire \top_ihp.oisc.regs[18][4] ;
 wire \top_ihp.oisc.regs[18][5] ;
 wire \top_ihp.oisc.regs[18][6] ;
 wire \top_ihp.oisc.regs[18][7] ;
 wire \top_ihp.oisc.regs[18][8] ;
 wire \top_ihp.oisc.regs[18][9] ;
 wire \top_ihp.oisc.regs[19][0] ;
 wire \top_ihp.oisc.regs[19][10] ;
 wire \top_ihp.oisc.regs[19][11] ;
 wire \top_ihp.oisc.regs[19][12] ;
 wire \top_ihp.oisc.regs[19][13] ;
 wire \top_ihp.oisc.regs[19][14] ;
 wire \top_ihp.oisc.regs[19][15] ;
 wire \top_ihp.oisc.regs[19][16] ;
 wire \top_ihp.oisc.regs[19][17] ;
 wire \top_ihp.oisc.regs[19][18] ;
 wire \top_ihp.oisc.regs[19][19] ;
 wire \top_ihp.oisc.regs[19][1] ;
 wire \top_ihp.oisc.regs[19][20] ;
 wire \top_ihp.oisc.regs[19][21] ;
 wire \top_ihp.oisc.regs[19][22] ;
 wire \top_ihp.oisc.regs[19][23] ;
 wire \top_ihp.oisc.regs[19][24] ;
 wire \top_ihp.oisc.regs[19][25] ;
 wire \top_ihp.oisc.regs[19][26] ;
 wire \top_ihp.oisc.regs[19][27] ;
 wire \top_ihp.oisc.regs[19][28] ;
 wire \top_ihp.oisc.regs[19][29] ;
 wire \top_ihp.oisc.regs[19][2] ;
 wire \top_ihp.oisc.regs[19][30] ;
 wire \top_ihp.oisc.regs[19][31] ;
 wire \top_ihp.oisc.regs[19][3] ;
 wire \top_ihp.oisc.regs[19][4] ;
 wire \top_ihp.oisc.regs[19][5] ;
 wire \top_ihp.oisc.regs[19][6] ;
 wire \top_ihp.oisc.regs[19][7] ;
 wire \top_ihp.oisc.regs[19][8] ;
 wire \top_ihp.oisc.regs[19][9] ;
 wire \top_ihp.oisc.regs[1][0] ;
 wire \top_ihp.oisc.regs[1][10] ;
 wire \top_ihp.oisc.regs[1][11] ;
 wire \top_ihp.oisc.regs[1][12] ;
 wire \top_ihp.oisc.regs[1][13] ;
 wire \top_ihp.oisc.regs[1][14] ;
 wire \top_ihp.oisc.regs[1][15] ;
 wire \top_ihp.oisc.regs[1][16] ;
 wire \top_ihp.oisc.regs[1][17] ;
 wire \top_ihp.oisc.regs[1][18] ;
 wire \top_ihp.oisc.regs[1][19] ;
 wire \top_ihp.oisc.regs[1][1] ;
 wire \top_ihp.oisc.regs[1][20] ;
 wire \top_ihp.oisc.regs[1][21] ;
 wire \top_ihp.oisc.regs[1][22] ;
 wire \top_ihp.oisc.regs[1][23] ;
 wire \top_ihp.oisc.regs[1][24] ;
 wire \top_ihp.oisc.regs[1][25] ;
 wire \top_ihp.oisc.regs[1][26] ;
 wire \top_ihp.oisc.regs[1][27] ;
 wire \top_ihp.oisc.regs[1][28] ;
 wire \top_ihp.oisc.regs[1][29] ;
 wire \top_ihp.oisc.regs[1][2] ;
 wire \top_ihp.oisc.regs[1][30] ;
 wire \top_ihp.oisc.regs[1][31] ;
 wire \top_ihp.oisc.regs[1][3] ;
 wire \top_ihp.oisc.regs[1][4] ;
 wire \top_ihp.oisc.regs[1][5] ;
 wire \top_ihp.oisc.regs[1][6] ;
 wire \top_ihp.oisc.regs[1][7] ;
 wire \top_ihp.oisc.regs[1][8] ;
 wire \top_ihp.oisc.regs[1][9] ;
 wire \top_ihp.oisc.regs[20][0] ;
 wire \top_ihp.oisc.regs[20][10] ;
 wire \top_ihp.oisc.regs[20][11] ;
 wire \top_ihp.oisc.regs[20][12] ;
 wire \top_ihp.oisc.regs[20][13] ;
 wire \top_ihp.oisc.regs[20][14] ;
 wire \top_ihp.oisc.regs[20][15] ;
 wire \top_ihp.oisc.regs[20][16] ;
 wire \top_ihp.oisc.regs[20][17] ;
 wire \top_ihp.oisc.regs[20][18] ;
 wire \top_ihp.oisc.regs[20][19] ;
 wire \top_ihp.oisc.regs[20][1] ;
 wire \top_ihp.oisc.regs[20][20] ;
 wire \top_ihp.oisc.regs[20][21] ;
 wire \top_ihp.oisc.regs[20][22] ;
 wire \top_ihp.oisc.regs[20][23] ;
 wire \top_ihp.oisc.regs[20][24] ;
 wire \top_ihp.oisc.regs[20][25] ;
 wire \top_ihp.oisc.regs[20][26] ;
 wire \top_ihp.oisc.regs[20][27] ;
 wire \top_ihp.oisc.regs[20][28] ;
 wire \top_ihp.oisc.regs[20][29] ;
 wire \top_ihp.oisc.regs[20][2] ;
 wire \top_ihp.oisc.regs[20][30] ;
 wire \top_ihp.oisc.regs[20][31] ;
 wire \top_ihp.oisc.regs[20][3] ;
 wire \top_ihp.oisc.regs[20][4] ;
 wire \top_ihp.oisc.regs[20][5] ;
 wire \top_ihp.oisc.regs[20][6] ;
 wire \top_ihp.oisc.regs[20][7] ;
 wire \top_ihp.oisc.regs[20][8] ;
 wire \top_ihp.oisc.regs[20][9] ;
 wire \top_ihp.oisc.regs[21][0] ;
 wire \top_ihp.oisc.regs[21][10] ;
 wire \top_ihp.oisc.regs[21][11] ;
 wire \top_ihp.oisc.regs[21][12] ;
 wire \top_ihp.oisc.regs[21][13] ;
 wire \top_ihp.oisc.regs[21][14] ;
 wire \top_ihp.oisc.regs[21][15] ;
 wire \top_ihp.oisc.regs[21][16] ;
 wire \top_ihp.oisc.regs[21][17] ;
 wire \top_ihp.oisc.regs[21][18] ;
 wire \top_ihp.oisc.regs[21][19] ;
 wire \top_ihp.oisc.regs[21][1] ;
 wire \top_ihp.oisc.regs[21][20] ;
 wire \top_ihp.oisc.regs[21][21] ;
 wire \top_ihp.oisc.regs[21][22] ;
 wire \top_ihp.oisc.regs[21][23] ;
 wire \top_ihp.oisc.regs[21][24] ;
 wire \top_ihp.oisc.regs[21][25] ;
 wire \top_ihp.oisc.regs[21][26] ;
 wire \top_ihp.oisc.regs[21][27] ;
 wire \top_ihp.oisc.regs[21][28] ;
 wire \top_ihp.oisc.regs[21][29] ;
 wire \top_ihp.oisc.regs[21][2] ;
 wire \top_ihp.oisc.regs[21][30] ;
 wire \top_ihp.oisc.regs[21][31] ;
 wire \top_ihp.oisc.regs[21][3] ;
 wire \top_ihp.oisc.regs[21][4] ;
 wire \top_ihp.oisc.regs[21][5] ;
 wire \top_ihp.oisc.regs[21][6] ;
 wire \top_ihp.oisc.regs[21][7] ;
 wire \top_ihp.oisc.regs[21][8] ;
 wire \top_ihp.oisc.regs[21][9] ;
 wire \top_ihp.oisc.regs[22][0] ;
 wire \top_ihp.oisc.regs[22][10] ;
 wire \top_ihp.oisc.regs[22][11] ;
 wire \top_ihp.oisc.regs[22][12] ;
 wire \top_ihp.oisc.regs[22][13] ;
 wire \top_ihp.oisc.regs[22][14] ;
 wire \top_ihp.oisc.regs[22][15] ;
 wire \top_ihp.oisc.regs[22][16] ;
 wire \top_ihp.oisc.regs[22][17] ;
 wire \top_ihp.oisc.regs[22][18] ;
 wire \top_ihp.oisc.regs[22][19] ;
 wire \top_ihp.oisc.regs[22][1] ;
 wire \top_ihp.oisc.regs[22][20] ;
 wire \top_ihp.oisc.regs[22][21] ;
 wire \top_ihp.oisc.regs[22][22] ;
 wire \top_ihp.oisc.regs[22][23] ;
 wire \top_ihp.oisc.regs[22][24] ;
 wire \top_ihp.oisc.regs[22][25] ;
 wire \top_ihp.oisc.regs[22][26] ;
 wire \top_ihp.oisc.regs[22][27] ;
 wire \top_ihp.oisc.regs[22][28] ;
 wire \top_ihp.oisc.regs[22][29] ;
 wire \top_ihp.oisc.regs[22][2] ;
 wire \top_ihp.oisc.regs[22][30] ;
 wire \top_ihp.oisc.regs[22][31] ;
 wire \top_ihp.oisc.regs[22][3] ;
 wire \top_ihp.oisc.regs[22][4] ;
 wire \top_ihp.oisc.regs[22][5] ;
 wire \top_ihp.oisc.regs[22][6] ;
 wire \top_ihp.oisc.regs[22][7] ;
 wire \top_ihp.oisc.regs[22][8] ;
 wire \top_ihp.oisc.regs[22][9] ;
 wire \top_ihp.oisc.regs[23][0] ;
 wire \top_ihp.oisc.regs[23][10] ;
 wire \top_ihp.oisc.regs[23][11] ;
 wire \top_ihp.oisc.regs[23][12] ;
 wire \top_ihp.oisc.regs[23][13] ;
 wire \top_ihp.oisc.regs[23][14] ;
 wire \top_ihp.oisc.regs[23][15] ;
 wire \top_ihp.oisc.regs[23][16] ;
 wire \top_ihp.oisc.regs[23][17] ;
 wire \top_ihp.oisc.regs[23][18] ;
 wire \top_ihp.oisc.regs[23][19] ;
 wire \top_ihp.oisc.regs[23][1] ;
 wire \top_ihp.oisc.regs[23][20] ;
 wire \top_ihp.oisc.regs[23][21] ;
 wire \top_ihp.oisc.regs[23][22] ;
 wire \top_ihp.oisc.regs[23][23] ;
 wire \top_ihp.oisc.regs[23][24] ;
 wire \top_ihp.oisc.regs[23][25] ;
 wire \top_ihp.oisc.regs[23][26] ;
 wire \top_ihp.oisc.regs[23][27] ;
 wire \top_ihp.oisc.regs[23][28] ;
 wire \top_ihp.oisc.regs[23][29] ;
 wire \top_ihp.oisc.regs[23][2] ;
 wire \top_ihp.oisc.regs[23][30] ;
 wire \top_ihp.oisc.regs[23][31] ;
 wire \top_ihp.oisc.regs[23][3] ;
 wire \top_ihp.oisc.regs[23][4] ;
 wire \top_ihp.oisc.regs[23][5] ;
 wire \top_ihp.oisc.regs[23][6] ;
 wire \top_ihp.oisc.regs[23][7] ;
 wire \top_ihp.oisc.regs[23][8] ;
 wire \top_ihp.oisc.regs[23][9] ;
 wire \top_ihp.oisc.regs[24][0] ;
 wire \top_ihp.oisc.regs[24][10] ;
 wire \top_ihp.oisc.regs[24][11] ;
 wire \top_ihp.oisc.regs[24][12] ;
 wire \top_ihp.oisc.regs[24][13] ;
 wire \top_ihp.oisc.regs[24][14] ;
 wire \top_ihp.oisc.regs[24][15] ;
 wire \top_ihp.oisc.regs[24][16] ;
 wire \top_ihp.oisc.regs[24][17] ;
 wire \top_ihp.oisc.regs[24][18] ;
 wire \top_ihp.oisc.regs[24][19] ;
 wire \top_ihp.oisc.regs[24][1] ;
 wire \top_ihp.oisc.regs[24][20] ;
 wire \top_ihp.oisc.regs[24][21] ;
 wire \top_ihp.oisc.regs[24][22] ;
 wire \top_ihp.oisc.regs[24][23] ;
 wire \top_ihp.oisc.regs[24][24] ;
 wire \top_ihp.oisc.regs[24][25] ;
 wire \top_ihp.oisc.regs[24][26] ;
 wire \top_ihp.oisc.regs[24][27] ;
 wire \top_ihp.oisc.regs[24][28] ;
 wire \top_ihp.oisc.regs[24][29] ;
 wire \top_ihp.oisc.regs[24][2] ;
 wire \top_ihp.oisc.regs[24][30] ;
 wire \top_ihp.oisc.regs[24][31] ;
 wire \top_ihp.oisc.regs[24][3] ;
 wire \top_ihp.oisc.regs[24][4] ;
 wire \top_ihp.oisc.regs[24][5] ;
 wire \top_ihp.oisc.regs[24][6] ;
 wire \top_ihp.oisc.regs[24][7] ;
 wire \top_ihp.oisc.regs[24][8] ;
 wire \top_ihp.oisc.regs[24][9] ;
 wire \top_ihp.oisc.regs[25][0] ;
 wire \top_ihp.oisc.regs[25][10] ;
 wire \top_ihp.oisc.regs[25][11] ;
 wire \top_ihp.oisc.regs[25][12] ;
 wire \top_ihp.oisc.regs[25][13] ;
 wire \top_ihp.oisc.regs[25][14] ;
 wire \top_ihp.oisc.regs[25][15] ;
 wire \top_ihp.oisc.regs[25][16] ;
 wire \top_ihp.oisc.regs[25][17] ;
 wire \top_ihp.oisc.regs[25][18] ;
 wire \top_ihp.oisc.regs[25][19] ;
 wire \top_ihp.oisc.regs[25][1] ;
 wire \top_ihp.oisc.regs[25][20] ;
 wire \top_ihp.oisc.regs[25][21] ;
 wire \top_ihp.oisc.regs[25][22] ;
 wire \top_ihp.oisc.regs[25][23] ;
 wire \top_ihp.oisc.regs[25][24] ;
 wire \top_ihp.oisc.regs[25][25] ;
 wire \top_ihp.oisc.regs[25][26] ;
 wire \top_ihp.oisc.regs[25][27] ;
 wire \top_ihp.oisc.regs[25][28] ;
 wire \top_ihp.oisc.regs[25][29] ;
 wire \top_ihp.oisc.regs[25][2] ;
 wire \top_ihp.oisc.regs[25][30] ;
 wire \top_ihp.oisc.regs[25][31] ;
 wire \top_ihp.oisc.regs[25][3] ;
 wire \top_ihp.oisc.regs[25][4] ;
 wire \top_ihp.oisc.regs[25][5] ;
 wire \top_ihp.oisc.regs[25][6] ;
 wire \top_ihp.oisc.regs[25][7] ;
 wire \top_ihp.oisc.regs[25][8] ;
 wire \top_ihp.oisc.regs[25][9] ;
 wire \top_ihp.oisc.regs[26][0] ;
 wire \top_ihp.oisc.regs[26][10] ;
 wire \top_ihp.oisc.regs[26][11] ;
 wire \top_ihp.oisc.regs[26][12] ;
 wire \top_ihp.oisc.regs[26][13] ;
 wire \top_ihp.oisc.regs[26][14] ;
 wire \top_ihp.oisc.regs[26][15] ;
 wire \top_ihp.oisc.regs[26][16] ;
 wire \top_ihp.oisc.regs[26][17] ;
 wire \top_ihp.oisc.regs[26][18] ;
 wire \top_ihp.oisc.regs[26][19] ;
 wire \top_ihp.oisc.regs[26][1] ;
 wire \top_ihp.oisc.regs[26][20] ;
 wire \top_ihp.oisc.regs[26][21] ;
 wire \top_ihp.oisc.regs[26][22] ;
 wire \top_ihp.oisc.regs[26][23] ;
 wire \top_ihp.oisc.regs[26][24] ;
 wire \top_ihp.oisc.regs[26][25] ;
 wire \top_ihp.oisc.regs[26][26] ;
 wire \top_ihp.oisc.regs[26][27] ;
 wire \top_ihp.oisc.regs[26][28] ;
 wire \top_ihp.oisc.regs[26][29] ;
 wire \top_ihp.oisc.regs[26][2] ;
 wire \top_ihp.oisc.regs[26][30] ;
 wire \top_ihp.oisc.regs[26][31] ;
 wire \top_ihp.oisc.regs[26][3] ;
 wire \top_ihp.oisc.regs[26][4] ;
 wire \top_ihp.oisc.regs[26][5] ;
 wire \top_ihp.oisc.regs[26][6] ;
 wire \top_ihp.oisc.regs[26][7] ;
 wire \top_ihp.oisc.regs[26][8] ;
 wire \top_ihp.oisc.regs[26][9] ;
 wire \top_ihp.oisc.regs[27][0] ;
 wire \top_ihp.oisc.regs[27][10] ;
 wire \top_ihp.oisc.regs[27][11] ;
 wire \top_ihp.oisc.regs[27][12] ;
 wire \top_ihp.oisc.regs[27][13] ;
 wire \top_ihp.oisc.regs[27][14] ;
 wire \top_ihp.oisc.regs[27][15] ;
 wire \top_ihp.oisc.regs[27][16] ;
 wire \top_ihp.oisc.regs[27][17] ;
 wire \top_ihp.oisc.regs[27][18] ;
 wire \top_ihp.oisc.regs[27][19] ;
 wire \top_ihp.oisc.regs[27][1] ;
 wire \top_ihp.oisc.regs[27][20] ;
 wire \top_ihp.oisc.regs[27][21] ;
 wire \top_ihp.oisc.regs[27][22] ;
 wire \top_ihp.oisc.regs[27][23] ;
 wire \top_ihp.oisc.regs[27][24] ;
 wire \top_ihp.oisc.regs[27][25] ;
 wire \top_ihp.oisc.regs[27][26] ;
 wire \top_ihp.oisc.regs[27][27] ;
 wire \top_ihp.oisc.regs[27][28] ;
 wire \top_ihp.oisc.regs[27][29] ;
 wire \top_ihp.oisc.regs[27][2] ;
 wire \top_ihp.oisc.regs[27][30] ;
 wire \top_ihp.oisc.regs[27][31] ;
 wire \top_ihp.oisc.regs[27][3] ;
 wire \top_ihp.oisc.regs[27][4] ;
 wire \top_ihp.oisc.regs[27][5] ;
 wire \top_ihp.oisc.regs[27][6] ;
 wire \top_ihp.oisc.regs[27][7] ;
 wire \top_ihp.oisc.regs[27][8] ;
 wire \top_ihp.oisc.regs[27][9] ;
 wire \top_ihp.oisc.regs[28][0] ;
 wire \top_ihp.oisc.regs[28][10] ;
 wire \top_ihp.oisc.regs[28][11] ;
 wire \top_ihp.oisc.regs[28][12] ;
 wire \top_ihp.oisc.regs[28][13] ;
 wire \top_ihp.oisc.regs[28][14] ;
 wire \top_ihp.oisc.regs[28][15] ;
 wire \top_ihp.oisc.regs[28][16] ;
 wire \top_ihp.oisc.regs[28][17] ;
 wire \top_ihp.oisc.regs[28][18] ;
 wire \top_ihp.oisc.regs[28][19] ;
 wire \top_ihp.oisc.regs[28][1] ;
 wire \top_ihp.oisc.regs[28][20] ;
 wire \top_ihp.oisc.regs[28][21] ;
 wire \top_ihp.oisc.regs[28][22] ;
 wire \top_ihp.oisc.regs[28][23] ;
 wire \top_ihp.oisc.regs[28][24] ;
 wire \top_ihp.oisc.regs[28][25] ;
 wire \top_ihp.oisc.regs[28][26] ;
 wire \top_ihp.oisc.regs[28][27] ;
 wire \top_ihp.oisc.regs[28][28] ;
 wire \top_ihp.oisc.regs[28][29] ;
 wire \top_ihp.oisc.regs[28][2] ;
 wire \top_ihp.oisc.regs[28][30] ;
 wire \top_ihp.oisc.regs[28][31] ;
 wire \top_ihp.oisc.regs[28][3] ;
 wire \top_ihp.oisc.regs[28][4] ;
 wire \top_ihp.oisc.regs[28][5] ;
 wire \top_ihp.oisc.regs[28][6] ;
 wire \top_ihp.oisc.regs[28][7] ;
 wire \top_ihp.oisc.regs[28][8] ;
 wire \top_ihp.oisc.regs[28][9] ;
 wire \top_ihp.oisc.regs[29][0] ;
 wire \top_ihp.oisc.regs[29][10] ;
 wire \top_ihp.oisc.regs[29][11] ;
 wire \top_ihp.oisc.regs[29][12] ;
 wire \top_ihp.oisc.regs[29][13] ;
 wire \top_ihp.oisc.regs[29][14] ;
 wire \top_ihp.oisc.regs[29][15] ;
 wire \top_ihp.oisc.regs[29][16] ;
 wire \top_ihp.oisc.regs[29][17] ;
 wire \top_ihp.oisc.regs[29][18] ;
 wire \top_ihp.oisc.regs[29][19] ;
 wire \top_ihp.oisc.regs[29][1] ;
 wire \top_ihp.oisc.regs[29][20] ;
 wire \top_ihp.oisc.regs[29][21] ;
 wire \top_ihp.oisc.regs[29][22] ;
 wire \top_ihp.oisc.regs[29][23] ;
 wire \top_ihp.oisc.regs[29][24] ;
 wire \top_ihp.oisc.regs[29][25] ;
 wire \top_ihp.oisc.regs[29][26] ;
 wire \top_ihp.oisc.regs[29][27] ;
 wire \top_ihp.oisc.regs[29][28] ;
 wire \top_ihp.oisc.regs[29][29] ;
 wire \top_ihp.oisc.regs[29][2] ;
 wire \top_ihp.oisc.regs[29][30] ;
 wire \top_ihp.oisc.regs[29][31] ;
 wire \top_ihp.oisc.regs[29][3] ;
 wire \top_ihp.oisc.regs[29][4] ;
 wire \top_ihp.oisc.regs[29][5] ;
 wire \top_ihp.oisc.regs[29][6] ;
 wire \top_ihp.oisc.regs[29][7] ;
 wire \top_ihp.oisc.regs[29][8] ;
 wire \top_ihp.oisc.regs[29][9] ;
 wire \top_ihp.oisc.regs[2][0] ;
 wire \top_ihp.oisc.regs[2][10] ;
 wire \top_ihp.oisc.regs[2][11] ;
 wire \top_ihp.oisc.regs[2][12] ;
 wire \top_ihp.oisc.regs[2][13] ;
 wire \top_ihp.oisc.regs[2][14] ;
 wire \top_ihp.oisc.regs[2][15] ;
 wire \top_ihp.oisc.regs[2][16] ;
 wire \top_ihp.oisc.regs[2][17] ;
 wire \top_ihp.oisc.regs[2][18] ;
 wire \top_ihp.oisc.regs[2][19] ;
 wire \top_ihp.oisc.regs[2][1] ;
 wire \top_ihp.oisc.regs[2][20] ;
 wire \top_ihp.oisc.regs[2][21] ;
 wire \top_ihp.oisc.regs[2][22] ;
 wire \top_ihp.oisc.regs[2][23] ;
 wire \top_ihp.oisc.regs[2][24] ;
 wire \top_ihp.oisc.regs[2][25] ;
 wire \top_ihp.oisc.regs[2][26] ;
 wire \top_ihp.oisc.regs[2][27] ;
 wire \top_ihp.oisc.regs[2][28] ;
 wire \top_ihp.oisc.regs[2][29] ;
 wire \top_ihp.oisc.regs[2][2] ;
 wire \top_ihp.oisc.regs[2][30] ;
 wire \top_ihp.oisc.regs[2][31] ;
 wire \top_ihp.oisc.regs[2][3] ;
 wire \top_ihp.oisc.regs[2][4] ;
 wire \top_ihp.oisc.regs[2][5] ;
 wire \top_ihp.oisc.regs[2][6] ;
 wire \top_ihp.oisc.regs[2][7] ;
 wire \top_ihp.oisc.regs[2][8] ;
 wire \top_ihp.oisc.regs[2][9] ;
 wire \top_ihp.oisc.regs[30][0] ;
 wire \top_ihp.oisc.regs[30][10] ;
 wire \top_ihp.oisc.regs[30][11] ;
 wire \top_ihp.oisc.regs[30][12] ;
 wire \top_ihp.oisc.regs[30][13] ;
 wire \top_ihp.oisc.regs[30][14] ;
 wire \top_ihp.oisc.regs[30][15] ;
 wire \top_ihp.oisc.regs[30][16] ;
 wire \top_ihp.oisc.regs[30][17] ;
 wire \top_ihp.oisc.regs[30][18] ;
 wire \top_ihp.oisc.regs[30][19] ;
 wire \top_ihp.oisc.regs[30][1] ;
 wire \top_ihp.oisc.regs[30][20] ;
 wire \top_ihp.oisc.regs[30][21] ;
 wire \top_ihp.oisc.regs[30][22] ;
 wire \top_ihp.oisc.regs[30][23] ;
 wire \top_ihp.oisc.regs[30][24] ;
 wire \top_ihp.oisc.regs[30][25] ;
 wire \top_ihp.oisc.regs[30][26] ;
 wire \top_ihp.oisc.regs[30][27] ;
 wire \top_ihp.oisc.regs[30][28] ;
 wire \top_ihp.oisc.regs[30][29] ;
 wire \top_ihp.oisc.regs[30][2] ;
 wire \top_ihp.oisc.regs[30][30] ;
 wire \top_ihp.oisc.regs[30][31] ;
 wire \top_ihp.oisc.regs[30][3] ;
 wire \top_ihp.oisc.regs[30][4] ;
 wire \top_ihp.oisc.regs[30][5] ;
 wire \top_ihp.oisc.regs[30][6] ;
 wire \top_ihp.oisc.regs[30][7] ;
 wire \top_ihp.oisc.regs[30][8] ;
 wire \top_ihp.oisc.regs[30][9] ;
 wire \top_ihp.oisc.regs[31][0] ;
 wire \top_ihp.oisc.regs[31][10] ;
 wire \top_ihp.oisc.regs[31][11] ;
 wire \top_ihp.oisc.regs[31][12] ;
 wire \top_ihp.oisc.regs[31][13] ;
 wire \top_ihp.oisc.regs[31][14] ;
 wire \top_ihp.oisc.regs[31][15] ;
 wire \top_ihp.oisc.regs[31][16] ;
 wire \top_ihp.oisc.regs[31][17] ;
 wire \top_ihp.oisc.regs[31][18] ;
 wire \top_ihp.oisc.regs[31][19] ;
 wire \top_ihp.oisc.regs[31][1] ;
 wire \top_ihp.oisc.regs[31][20] ;
 wire \top_ihp.oisc.regs[31][21] ;
 wire \top_ihp.oisc.regs[31][22] ;
 wire \top_ihp.oisc.regs[31][23] ;
 wire \top_ihp.oisc.regs[31][24] ;
 wire \top_ihp.oisc.regs[31][25] ;
 wire \top_ihp.oisc.regs[31][26] ;
 wire \top_ihp.oisc.regs[31][27] ;
 wire \top_ihp.oisc.regs[31][28] ;
 wire \top_ihp.oisc.regs[31][29] ;
 wire \top_ihp.oisc.regs[31][2] ;
 wire \top_ihp.oisc.regs[31][30] ;
 wire \top_ihp.oisc.regs[31][31] ;
 wire \top_ihp.oisc.regs[31][3] ;
 wire \top_ihp.oisc.regs[31][4] ;
 wire \top_ihp.oisc.regs[31][5] ;
 wire \top_ihp.oisc.regs[31][6] ;
 wire \top_ihp.oisc.regs[31][7] ;
 wire \top_ihp.oisc.regs[31][8] ;
 wire \top_ihp.oisc.regs[31][9] ;
 wire \top_ihp.oisc.regs[32][0] ;
 wire \top_ihp.oisc.regs[32][10] ;
 wire \top_ihp.oisc.regs[32][11] ;
 wire \top_ihp.oisc.regs[32][12] ;
 wire \top_ihp.oisc.regs[32][13] ;
 wire \top_ihp.oisc.regs[32][14] ;
 wire \top_ihp.oisc.regs[32][15] ;
 wire \top_ihp.oisc.regs[32][16] ;
 wire \top_ihp.oisc.regs[32][17] ;
 wire \top_ihp.oisc.regs[32][18] ;
 wire \top_ihp.oisc.regs[32][19] ;
 wire \top_ihp.oisc.regs[32][1] ;
 wire \top_ihp.oisc.regs[32][20] ;
 wire \top_ihp.oisc.regs[32][21] ;
 wire \top_ihp.oisc.regs[32][22] ;
 wire \top_ihp.oisc.regs[32][23] ;
 wire \top_ihp.oisc.regs[32][24] ;
 wire \top_ihp.oisc.regs[32][25] ;
 wire \top_ihp.oisc.regs[32][26] ;
 wire \top_ihp.oisc.regs[32][27] ;
 wire \top_ihp.oisc.regs[32][28] ;
 wire \top_ihp.oisc.regs[32][29] ;
 wire \top_ihp.oisc.regs[32][2] ;
 wire \top_ihp.oisc.regs[32][30] ;
 wire \top_ihp.oisc.regs[32][31] ;
 wire \top_ihp.oisc.regs[32][3] ;
 wire \top_ihp.oisc.regs[32][4] ;
 wire \top_ihp.oisc.regs[32][5] ;
 wire \top_ihp.oisc.regs[32][6] ;
 wire \top_ihp.oisc.regs[32][7] ;
 wire \top_ihp.oisc.regs[32][8] ;
 wire \top_ihp.oisc.regs[32][9] ;
 wire \top_ihp.oisc.regs[33][0] ;
 wire \top_ihp.oisc.regs[33][10] ;
 wire \top_ihp.oisc.regs[33][11] ;
 wire \top_ihp.oisc.regs[33][12] ;
 wire \top_ihp.oisc.regs[33][13] ;
 wire \top_ihp.oisc.regs[33][14] ;
 wire \top_ihp.oisc.regs[33][15] ;
 wire \top_ihp.oisc.regs[33][16] ;
 wire \top_ihp.oisc.regs[33][17] ;
 wire \top_ihp.oisc.regs[33][18] ;
 wire \top_ihp.oisc.regs[33][19] ;
 wire \top_ihp.oisc.regs[33][1] ;
 wire \top_ihp.oisc.regs[33][20] ;
 wire \top_ihp.oisc.regs[33][21] ;
 wire \top_ihp.oisc.regs[33][22] ;
 wire \top_ihp.oisc.regs[33][23] ;
 wire \top_ihp.oisc.regs[33][24] ;
 wire \top_ihp.oisc.regs[33][25] ;
 wire \top_ihp.oisc.regs[33][26] ;
 wire \top_ihp.oisc.regs[33][27] ;
 wire \top_ihp.oisc.regs[33][28] ;
 wire \top_ihp.oisc.regs[33][29] ;
 wire \top_ihp.oisc.regs[33][2] ;
 wire \top_ihp.oisc.regs[33][30] ;
 wire \top_ihp.oisc.regs[33][31] ;
 wire \top_ihp.oisc.regs[33][3] ;
 wire \top_ihp.oisc.regs[33][4] ;
 wire \top_ihp.oisc.regs[33][5] ;
 wire \top_ihp.oisc.regs[33][6] ;
 wire \top_ihp.oisc.regs[33][7] ;
 wire \top_ihp.oisc.regs[33][8] ;
 wire \top_ihp.oisc.regs[33][9] ;
 wire \top_ihp.oisc.regs[34][0] ;
 wire \top_ihp.oisc.regs[34][10] ;
 wire \top_ihp.oisc.regs[34][11] ;
 wire \top_ihp.oisc.regs[34][12] ;
 wire \top_ihp.oisc.regs[34][13] ;
 wire \top_ihp.oisc.regs[34][14] ;
 wire \top_ihp.oisc.regs[34][15] ;
 wire \top_ihp.oisc.regs[34][16] ;
 wire \top_ihp.oisc.regs[34][17] ;
 wire \top_ihp.oisc.regs[34][18] ;
 wire \top_ihp.oisc.regs[34][19] ;
 wire \top_ihp.oisc.regs[34][1] ;
 wire \top_ihp.oisc.regs[34][20] ;
 wire \top_ihp.oisc.regs[34][21] ;
 wire \top_ihp.oisc.regs[34][22] ;
 wire \top_ihp.oisc.regs[34][23] ;
 wire \top_ihp.oisc.regs[34][24] ;
 wire \top_ihp.oisc.regs[34][25] ;
 wire \top_ihp.oisc.regs[34][26] ;
 wire \top_ihp.oisc.regs[34][27] ;
 wire \top_ihp.oisc.regs[34][28] ;
 wire \top_ihp.oisc.regs[34][29] ;
 wire \top_ihp.oisc.regs[34][2] ;
 wire \top_ihp.oisc.regs[34][30] ;
 wire \top_ihp.oisc.regs[34][31] ;
 wire \top_ihp.oisc.regs[34][3] ;
 wire \top_ihp.oisc.regs[34][4] ;
 wire \top_ihp.oisc.regs[34][5] ;
 wire \top_ihp.oisc.regs[34][6] ;
 wire \top_ihp.oisc.regs[34][7] ;
 wire \top_ihp.oisc.regs[34][8] ;
 wire \top_ihp.oisc.regs[34][9] ;
 wire \top_ihp.oisc.regs[35][0] ;
 wire \top_ihp.oisc.regs[35][10] ;
 wire \top_ihp.oisc.regs[35][11] ;
 wire \top_ihp.oisc.regs[35][12] ;
 wire \top_ihp.oisc.regs[35][13] ;
 wire \top_ihp.oisc.regs[35][14] ;
 wire \top_ihp.oisc.regs[35][15] ;
 wire \top_ihp.oisc.regs[35][16] ;
 wire \top_ihp.oisc.regs[35][17] ;
 wire \top_ihp.oisc.regs[35][18] ;
 wire \top_ihp.oisc.regs[35][19] ;
 wire \top_ihp.oisc.regs[35][1] ;
 wire \top_ihp.oisc.regs[35][20] ;
 wire \top_ihp.oisc.regs[35][21] ;
 wire \top_ihp.oisc.regs[35][22] ;
 wire \top_ihp.oisc.regs[35][23] ;
 wire \top_ihp.oisc.regs[35][24] ;
 wire \top_ihp.oisc.regs[35][25] ;
 wire \top_ihp.oisc.regs[35][26] ;
 wire \top_ihp.oisc.regs[35][27] ;
 wire \top_ihp.oisc.regs[35][28] ;
 wire \top_ihp.oisc.regs[35][29] ;
 wire \top_ihp.oisc.regs[35][2] ;
 wire \top_ihp.oisc.regs[35][30] ;
 wire \top_ihp.oisc.regs[35][31] ;
 wire \top_ihp.oisc.regs[35][3] ;
 wire \top_ihp.oisc.regs[35][4] ;
 wire \top_ihp.oisc.regs[35][5] ;
 wire \top_ihp.oisc.regs[35][6] ;
 wire \top_ihp.oisc.regs[35][7] ;
 wire \top_ihp.oisc.regs[35][8] ;
 wire \top_ihp.oisc.regs[35][9] ;
 wire \top_ihp.oisc.regs[36][0] ;
 wire \top_ihp.oisc.regs[36][10] ;
 wire \top_ihp.oisc.regs[36][11] ;
 wire \top_ihp.oisc.regs[36][12] ;
 wire \top_ihp.oisc.regs[36][13] ;
 wire \top_ihp.oisc.regs[36][14] ;
 wire \top_ihp.oisc.regs[36][15] ;
 wire \top_ihp.oisc.regs[36][16] ;
 wire \top_ihp.oisc.regs[36][17] ;
 wire \top_ihp.oisc.regs[36][18] ;
 wire \top_ihp.oisc.regs[36][19] ;
 wire \top_ihp.oisc.regs[36][1] ;
 wire \top_ihp.oisc.regs[36][20] ;
 wire \top_ihp.oisc.regs[36][21] ;
 wire \top_ihp.oisc.regs[36][22] ;
 wire \top_ihp.oisc.regs[36][23] ;
 wire \top_ihp.oisc.regs[36][24] ;
 wire \top_ihp.oisc.regs[36][25] ;
 wire \top_ihp.oisc.regs[36][26] ;
 wire \top_ihp.oisc.regs[36][27] ;
 wire \top_ihp.oisc.regs[36][28] ;
 wire \top_ihp.oisc.regs[36][29] ;
 wire \top_ihp.oisc.regs[36][2] ;
 wire \top_ihp.oisc.regs[36][30] ;
 wire \top_ihp.oisc.regs[36][31] ;
 wire \top_ihp.oisc.regs[36][3] ;
 wire \top_ihp.oisc.regs[36][4] ;
 wire \top_ihp.oisc.regs[36][5] ;
 wire \top_ihp.oisc.regs[36][6] ;
 wire \top_ihp.oisc.regs[36][7] ;
 wire \top_ihp.oisc.regs[36][8] ;
 wire \top_ihp.oisc.regs[36][9] ;
 wire \top_ihp.oisc.regs[37][0] ;
 wire \top_ihp.oisc.regs[37][10] ;
 wire \top_ihp.oisc.regs[37][11] ;
 wire \top_ihp.oisc.regs[37][12] ;
 wire \top_ihp.oisc.regs[37][13] ;
 wire \top_ihp.oisc.regs[37][14] ;
 wire \top_ihp.oisc.regs[37][15] ;
 wire \top_ihp.oisc.regs[37][16] ;
 wire \top_ihp.oisc.regs[37][17] ;
 wire \top_ihp.oisc.regs[37][18] ;
 wire \top_ihp.oisc.regs[37][19] ;
 wire \top_ihp.oisc.regs[37][1] ;
 wire \top_ihp.oisc.regs[37][20] ;
 wire \top_ihp.oisc.regs[37][21] ;
 wire \top_ihp.oisc.regs[37][22] ;
 wire \top_ihp.oisc.regs[37][23] ;
 wire \top_ihp.oisc.regs[37][24] ;
 wire \top_ihp.oisc.regs[37][25] ;
 wire \top_ihp.oisc.regs[37][26] ;
 wire \top_ihp.oisc.regs[37][27] ;
 wire \top_ihp.oisc.regs[37][28] ;
 wire \top_ihp.oisc.regs[37][29] ;
 wire \top_ihp.oisc.regs[37][2] ;
 wire \top_ihp.oisc.regs[37][30] ;
 wire \top_ihp.oisc.regs[37][31] ;
 wire \top_ihp.oisc.regs[37][3] ;
 wire \top_ihp.oisc.regs[37][4] ;
 wire \top_ihp.oisc.regs[37][5] ;
 wire \top_ihp.oisc.regs[37][6] ;
 wire \top_ihp.oisc.regs[37][7] ;
 wire \top_ihp.oisc.regs[37][8] ;
 wire \top_ihp.oisc.regs[37][9] ;
 wire \top_ihp.oisc.regs[38][0] ;
 wire \top_ihp.oisc.regs[38][10] ;
 wire \top_ihp.oisc.regs[38][11] ;
 wire \top_ihp.oisc.regs[38][12] ;
 wire \top_ihp.oisc.regs[38][13] ;
 wire \top_ihp.oisc.regs[38][14] ;
 wire \top_ihp.oisc.regs[38][15] ;
 wire \top_ihp.oisc.regs[38][16] ;
 wire \top_ihp.oisc.regs[38][17] ;
 wire \top_ihp.oisc.regs[38][18] ;
 wire \top_ihp.oisc.regs[38][19] ;
 wire \top_ihp.oisc.regs[38][1] ;
 wire \top_ihp.oisc.regs[38][20] ;
 wire \top_ihp.oisc.regs[38][21] ;
 wire \top_ihp.oisc.regs[38][22] ;
 wire \top_ihp.oisc.regs[38][23] ;
 wire \top_ihp.oisc.regs[38][24] ;
 wire \top_ihp.oisc.regs[38][25] ;
 wire \top_ihp.oisc.regs[38][26] ;
 wire \top_ihp.oisc.regs[38][27] ;
 wire \top_ihp.oisc.regs[38][28] ;
 wire \top_ihp.oisc.regs[38][29] ;
 wire \top_ihp.oisc.regs[38][2] ;
 wire \top_ihp.oisc.regs[38][30] ;
 wire \top_ihp.oisc.regs[38][31] ;
 wire \top_ihp.oisc.regs[38][3] ;
 wire \top_ihp.oisc.regs[38][4] ;
 wire \top_ihp.oisc.regs[38][5] ;
 wire \top_ihp.oisc.regs[38][6] ;
 wire \top_ihp.oisc.regs[38][7] ;
 wire \top_ihp.oisc.regs[38][8] ;
 wire \top_ihp.oisc.regs[38][9] ;
 wire \top_ihp.oisc.regs[39][0] ;
 wire \top_ihp.oisc.regs[39][10] ;
 wire \top_ihp.oisc.regs[39][11] ;
 wire \top_ihp.oisc.regs[39][12] ;
 wire \top_ihp.oisc.regs[39][13] ;
 wire \top_ihp.oisc.regs[39][14] ;
 wire \top_ihp.oisc.regs[39][15] ;
 wire \top_ihp.oisc.regs[39][16] ;
 wire \top_ihp.oisc.regs[39][17] ;
 wire \top_ihp.oisc.regs[39][18] ;
 wire \top_ihp.oisc.regs[39][19] ;
 wire \top_ihp.oisc.regs[39][1] ;
 wire \top_ihp.oisc.regs[39][20] ;
 wire \top_ihp.oisc.regs[39][21] ;
 wire \top_ihp.oisc.regs[39][22] ;
 wire \top_ihp.oisc.regs[39][23] ;
 wire \top_ihp.oisc.regs[39][24] ;
 wire \top_ihp.oisc.regs[39][25] ;
 wire \top_ihp.oisc.regs[39][26] ;
 wire \top_ihp.oisc.regs[39][27] ;
 wire \top_ihp.oisc.regs[39][28] ;
 wire \top_ihp.oisc.regs[39][29] ;
 wire \top_ihp.oisc.regs[39][2] ;
 wire \top_ihp.oisc.regs[39][30] ;
 wire \top_ihp.oisc.regs[39][31] ;
 wire \top_ihp.oisc.regs[39][3] ;
 wire \top_ihp.oisc.regs[39][4] ;
 wire \top_ihp.oisc.regs[39][5] ;
 wire \top_ihp.oisc.regs[39][6] ;
 wire \top_ihp.oisc.regs[39][7] ;
 wire \top_ihp.oisc.regs[39][8] ;
 wire \top_ihp.oisc.regs[39][9] ;
 wire \top_ihp.oisc.regs[3][0] ;
 wire \top_ihp.oisc.regs[3][10] ;
 wire \top_ihp.oisc.regs[3][11] ;
 wire \top_ihp.oisc.regs[3][12] ;
 wire \top_ihp.oisc.regs[3][13] ;
 wire \top_ihp.oisc.regs[3][14] ;
 wire \top_ihp.oisc.regs[3][15] ;
 wire \top_ihp.oisc.regs[3][16] ;
 wire \top_ihp.oisc.regs[3][17] ;
 wire \top_ihp.oisc.regs[3][18] ;
 wire \top_ihp.oisc.regs[3][19] ;
 wire \top_ihp.oisc.regs[3][1] ;
 wire \top_ihp.oisc.regs[3][20] ;
 wire \top_ihp.oisc.regs[3][21] ;
 wire \top_ihp.oisc.regs[3][22] ;
 wire \top_ihp.oisc.regs[3][23] ;
 wire \top_ihp.oisc.regs[3][24] ;
 wire \top_ihp.oisc.regs[3][25] ;
 wire \top_ihp.oisc.regs[3][26] ;
 wire \top_ihp.oisc.regs[3][27] ;
 wire \top_ihp.oisc.regs[3][28] ;
 wire \top_ihp.oisc.regs[3][29] ;
 wire \top_ihp.oisc.regs[3][2] ;
 wire \top_ihp.oisc.regs[3][30] ;
 wire \top_ihp.oisc.regs[3][31] ;
 wire \top_ihp.oisc.regs[3][3] ;
 wire \top_ihp.oisc.regs[3][4] ;
 wire \top_ihp.oisc.regs[3][5] ;
 wire \top_ihp.oisc.regs[3][6] ;
 wire \top_ihp.oisc.regs[3][7] ;
 wire \top_ihp.oisc.regs[3][8] ;
 wire \top_ihp.oisc.regs[3][9] ;
 wire \top_ihp.oisc.regs[40][0] ;
 wire \top_ihp.oisc.regs[40][10] ;
 wire \top_ihp.oisc.regs[40][11] ;
 wire \top_ihp.oisc.regs[40][12] ;
 wire \top_ihp.oisc.regs[40][13] ;
 wire \top_ihp.oisc.regs[40][14] ;
 wire \top_ihp.oisc.regs[40][15] ;
 wire \top_ihp.oisc.regs[40][16] ;
 wire \top_ihp.oisc.regs[40][17] ;
 wire \top_ihp.oisc.regs[40][18] ;
 wire \top_ihp.oisc.regs[40][19] ;
 wire \top_ihp.oisc.regs[40][1] ;
 wire \top_ihp.oisc.regs[40][20] ;
 wire \top_ihp.oisc.regs[40][21] ;
 wire \top_ihp.oisc.regs[40][22] ;
 wire \top_ihp.oisc.regs[40][23] ;
 wire \top_ihp.oisc.regs[40][24] ;
 wire \top_ihp.oisc.regs[40][25] ;
 wire \top_ihp.oisc.regs[40][26] ;
 wire \top_ihp.oisc.regs[40][27] ;
 wire \top_ihp.oisc.regs[40][28] ;
 wire \top_ihp.oisc.regs[40][29] ;
 wire \top_ihp.oisc.regs[40][2] ;
 wire \top_ihp.oisc.regs[40][30] ;
 wire \top_ihp.oisc.regs[40][31] ;
 wire \top_ihp.oisc.regs[40][3] ;
 wire \top_ihp.oisc.regs[40][4] ;
 wire \top_ihp.oisc.regs[40][5] ;
 wire \top_ihp.oisc.regs[40][6] ;
 wire \top_ihp.oisc.regs[40][7] ;
 wire \top_ihp.oisc.regs[40][8] ;
 wire \top_ihp.oisc.regs[40][9] ;
 wire \top_ihp.oisc.regs[41][0] ;
 wire \top_ihp.oisc.regs[41][10] ;
 wire \top_ihp.oisc.regs[41][11] ;
 wire \top_ihp.oisc.regs[41][12] ;
 wire \top_ihp.oisc.regs[41][13] ;
 wire \top_ihp.oisc.regs[41][14] ;
 wire \top_ihp.oisc.regs[41][15] ;
 wire \top_ihp.oisc.regs[41][16] ;
 wire \top_ihp.oisc.regs[41][17] ;
 wire \top_ihp.oisc.regs[41][18] ;
 wire \top_ihp.oisc.regs[41][19] ;
 wire \top_ihp.oisc.regs[41][1] ;
 wire \top_ihp.oisc.regs[41][20] ;
 wire \top_ihp.oisc.regs[41][21] ;
 wire \top_ihp.oisc.regs[41][22] ;
 wire \top_ihp.oisc.regs[41][23] ;
 wire \top_ihp.oisc.regs[41][24] ;
 wire \top_ihp.oisc.regs[41][25] ;
 wire \top_ihp.oisc.regs[41][26] ;
 wire \top_ihp.oisc.regs[41][27] ;
 wire \top_ihp.oisc.regs[41][28] ;
 wire \top_ihp.oisc.regs[41][29] ;
 wire \top_ihp.oisc.regs[41][2] ;
 wire \top_ihp.oisc.regs[41][30] ;
 wire \top_ihp.oisc.regs[41][31] ;
 wire \top_ihp.oisc.regs[41][3] ;
 wire \top_ihp.oisc.regs[41][4] ;
 wire \top_ihp.oisc.regs[41][5] ;
 wire \top_ihp.oisc.regs[41][6] ;
 wire \top_ihp.oisc.regs[41][7] ;
 wire \top_ihp.oisc.regs[41][8] ;
 wire \top_ihp.oisc.regs[41][9] ;
 wire \top_ihp.oisc.regs[42][0] ;
 wire \top_ihp.oisc.regs[42][10] ;
 wire \top_ihp.oisc.regs[42][11] ;
 wire \top_ihp.oisc.regs[42][12] ;
 wire \top_ihp.oisc.regs[42][13] ;
 wire \top_ihp.oisc.regs[42][14] ;
 wire \top_ihp.oisc.regs[42][15] ;
 wire \top_ihp.oisc.regs[42][16] ;
 wire \top_ihp.oisc.regs[42][17] ;
 wire \top_ihp.oisc.regs[42][18] ;
 wire \top_ihp.oisc.regs[42][19] ;
 wire \top_ihp.oisc.regs[42][1] ;
 wire \top_ihp.oisc.regs[42][20] ;
 wire \top_ihp.oisc.regs[42][21] ;
 wire \top_ihp.oisc.regs[42][22] ;
 wire \top_ihp.oisc.regs[42][23] ;
 wire \top_ihp.oisc.regs[42][24] ;
 wire \top_ihp.oisc.regs[42][25] ;
 wire \top_ihp.oisc.regs[42][26] ;
 wire \top_ihp.oisc.regs[42][27] ;
 wire \top_ihp.oisc.regs[42][28] ;
 wire \top_ihp.oisc.regs[42][29] ;
 wire \top_ihp.oisc.regs[42][2] ;
 wire \top_ihp.oisc.regs[42][30] ;
 wire \top_ihp.oisc.regs[42][31] ;
 wire \top_ihp.oisc.regs[42][3] ;
 wire \top_ihp.oisc.regs[42][4] ;
 wire \top_ihp.oisc.regs[42][5] ;
 wire \top_ihp.oisc.regs[42][6] ;
 wire \top_ihp.oisc.regs[42][7] ;
 wire \top_ihp.oisc.regs[42][8] ;
 wire \top_ihp.oisc.regs[42][9] ;
 wire \top_ihp.oisc.regs[43][0] ;
 wire \top_ihp.oisc.regs[43][10] ;
 wire \top_ihp.oisc.regs[43][11] ;
 wire \top_ihp.oisc.regs[43][12] ;
 wire \top_ihp.oisc.regs[43][13] ;
 wire \top_ihp.oisc.regs[43][14] ;
 wire \top_ihp.oisc.regs[43][15] ;
 wire \top_ihp.oisc.regs[43][16] ;
 wire \top_ihp.oisc.regs[43][17] ;
 wire \top_ihp.oisc.regs[43][18] ;
 wire \top_ihp.oisc.regs[43][19] ;
 wire \top_ihp.oisc.regs[43][1] ;
 wire \top_ihp.oisc.regs[43][20] ;
 wire \top_ihp.oisc.regs[43][21] ;
 wire \top_ihp.oisc.regs[43][22] ;
 wire \top_ihp.oisc.regs[43][23] ;
 wire \top_ihp.oisc.regs[43][24] ;
 wire \top_ihp.oisc.regs[43][25] ;
 wire \top_ihp.oisc.regs[43][26] ;
 wire \top_ihp.oisc.regs[43][27] ;
 wire \top_ihp.oisc.regs[43][28] ;
 wire \top_ihp.oisc.regs[43][29] ;
 wire \top_ihp.oisc.regs[43][2] ;
 wire \top_ihp.oisc.regs[43][30] ;
 wire \top_ihp.oisc.regs[43][31] ;
 wire \top_ihp.oisc.regs[43][3] ;
 wire \top_ihp.oisc.regs[43][4] ;
 wire \top_ihp.oisc.regs[43][5] ;
 wire \top_ihp.oisc.regs[43][6] ;
 wire \top_ihp.oisc.regs[43][7] ;
 wire \top_ihp.oisc.regs[43][8] ;
 wire \top_ihp.oisc.regs[43][9] ;
 wire \top_ihp.oisc.regs[44][0] ;
 wire \top_ihp.oisc.regs[44][10] ;
 wire \top_ihp.oisc.regs[44][11] ;
 wire \top_ihp.oisc.regs[44][12] ;
 wire \top_ihp.oisc.regs[44][13] ;
 wire \top_ihp.oisc.regs[44][14] ;
 wire \top_ihp.oisc.regs[44][15] ;
 wire \top_ihp.oisc.regs[44][16] ;
 wire \top_ihp.oisc.regs[44][17] ;
 wire \top_ihp.oisc.regs[44][18] ;
 wire \top_ihp.oisc.regs[44][19] ;
 wire \top_ihp.oisc.regs[44][1] ;
 wire \top_ihp.oisc.regs[44][20] ;
 wire \top_ihp.oisc.regs[44][21] ;
 wire \top_ihp.oisc.regs[44][22] ;
 wire \top_ihp.oisc.regs[44][23] ;
 wire \top_ihp.oisc.regs[44][24] ;
 wire \top_ihp.oisc.regs[44][25] ;
 wire \top_ihp.oisc.regs[44][26] ;
 wire \top_ihp.oisc.regs[44][27] ;
 wire \top_ihp.oisc.regs[44][28] ;
 wire \top_ihp.oisc.regs[44][29] ;
 wire \top_ihp.oisc.regs[44][2] ;
 wire \top_ihp.oisc.regs[44][30] ;
 wire \top_ihp.oisc.regs[44][31] ;
 wire \top_ihp.oisc.regs[44][3] ;
 wire \top_ihp.oisc.regs[44][4] ;
 wire \top_ihp.oisc.regs[44][5] ;
 wire \top_ihp.oisc.regs[44][6] ;
 wire \top_ihp.oisc.regs[44][7] ;
 wire \top_ihp.oisc.regs[44][8] ;
 wire \top_ihp.oisc.regs[44][9] ;
 wire \top_ihp.oisc.regs[45][0] ;
 wire \top_ihp.oisc.regs[45][10] ;
 wire \top_ihp.oisc.regs[45][11] ;
 wire \top_ihp.oisc.regs[45][12] ;
 wire \top_ihp.oisc.regs[45][13] ;
 wire \top_ihp.oisc.regs[45][14] ;
 wire \top_ihp.oisc.regs[45][15] ;
 wire \top_ihp.oisc.regs[45][16] ;
 wire \top_ihp.oisc.regs[45][17] ;
 wire \top_ihp.oisc.regs[45][18] ;
 wire \top_ihp.oisc.regs[45][19] ;
 wire \top_ihp.oisc.regs[45][1] ;
 wire \top_ihp.oisc.regs[45][20] ;
 wire \top_ihp.oisc.regs[45][21] ;
 wire \top_ihp.oisc.regs[45][22] ;
 wire \top_ihp.oisc.regs[45][23] ;
 wire \top_ihp.oisc.regs[45][24] ;
 wire \top_ihp.oisc.regs[45][25] ;
 wire \top_ihp.oisc.regs[45][26] ;
 wire \top_ihp.oisc.regs[45][27] ;
 wire \top_ihp.oisc.regs[45][28] ;
 wire \top_ihp.oisc.regs[45][29] ;
 wire \top_ihp.oisc.regs[45][2] ;
 wire \top_ihp.oisc.regs[45][30] ;
 wire \top_ihp.oisc.regs[45][31] ;
 wire \top_ihp.oisc.regs[45][3] ;
 wire \top_ihp.oisc.regs[45][4] ;
 wire \top_ihp.oisc.regs[45][5] ;
 wire \top_ihp.oisc.regs[45][6] ;
 wire \top_ihp.oisc.regs[45][7] ;
 wire \top_ihp.oisc.regs[45][8] ;
 wire \top_ihp.oisc.regs[45][9] ;
 wire \top_ihp.oisc.regs[46][0] ;
 wire \top_ihp.oisc.regs[46][10] ;
 wire \top_ihp.oisc.regs[46][11] ;
 wire \top_ihp.oisc.regs[46][12] ;
 wire \top_ihp.oisc.regs[46][13] ;
 wire \top_ihp.oisc.regs[46][14] ;
 wire \top_ihp.oisc.regs[46][15] ;
 wire \top_ihp.oisc.regs[46][16] ;
 wire \top_ihp.oisc.regs[46][17] ;
 wire \top_ihp.oisc.regs[46][18] ;
 wire \top_ihp.oisc.regs[46][19] ;
 wire \top_ihp.oisc.regs[46][1] ;
 wire \top_ihp.oisc.regs[46][20] ;
 wire \top_ihp.oisc.regs[46][21] ;
 wire \top_ihp.oisc.regs[46][22] ;
 wire \top_ihp.oisc.regs[46][23] ;
 wire \top_ihp.oisc.regs[46][24] ;
 wire \top_ihp.oisc.regs[46][25] ;
 wire \top_ihp.oisc.regs[46][26] ;
 wire \top_ihp.oisc.regs[46][27] ;
 wire \top_ihp.oisc.regs[46][28] ;
 wire \top_ihp.oisc.regs[46][29] ;
 wire \top_ihp.oisc.regs[46][2] ;
 wire \top_ihp.oisc.regs[46][30] ;
 wire \top_ihp.oisc.regs[46][31] ;
 wire \top_ihp.oisc.regs[46][3] ;
 wire \top_ihp.oisc.regs[46][4] ;
 wire \top_ihp.oisc.regs[46][5] ;
 wire \top_ihp.oisc.regs[46][6] ;
 wire \top_ihp.oisc.regs[46][7] ;
 wire \top_ihp.oisc.regs[46][8] ;
 wire \top_ihp.oisc.regs[46][9] ;
 wire \top_ihp.oisc.regs[47][0] ;
 wire \top_ihp.oisc.regs[47][10] ;
 wire \top_ihp.oisc.regs[47][11] ;
 wire \top_ihp.oisc.regs[47][12] ;
 wire \top_ihp.oisc.regs[47][13] ;
 wire \top_ihp.oisc.regs[47][14] ;
 wire \top_ihp.oisc.regs[47][15] ;
 wire \top_ihp.oisc.regs[47][16] ;
 wire \top_ihp.oisc.regs[47][17] ;
 wire \top_ihp.oisc.regs[47][18] ;
 wire \top_ihp.oisc.regs[47][19] ;
 wire \top_ihp.oisc.regs[47][1] ;
 wire \top_ihp.oisc.regs[47][20] ;
 wire \top_ihp.oisc.regs[47][21] ;
 wire \top_ihp.oisc.regs[47][22] ;
 wire \top_ihp.oisc.regs[47][23] ;
 wire \top_ihp.oisc.regs[47][24] ;
 wire \top_ihp.oisc.regs[47][25] ;
 wire \top_ihp.oisc.regs[47][26] ;
 wire \top_ihp.oisc.regs[47][27] ;
 wire \top_ihp.oisc.regs[47][28] ;
 wire \top_ihp.oisc.regs[47][29] ;
 wire \top_ihp.oisc.regs[47][2] ;
 wire \top_ihp.oisc.regs[47][30] ;
 wire \top_ihp.oisc.regs[47][31] ;
 wire \top_ihp.oisc.regs[47][3] ;
 wire \top_ihp.oisc.regs[47][4] ;
 wire \top_ihp.oisc.regs[47][5] ;
 wire \top_ihp.oisc.regs[47][6] ;
 wire \top_ihp.oisc.regs[47][7] ;
 wire \top_ihp.oisc.regs[47][8] ;
 wire \top_ihp.oisc.regs[47][9] ;
 wire \top_ihp.oisc.regs[48][0] ;
 wire \top_ihp.oisc.regs[48][10] ;
 wire \top_ihp.oisc.regs[48][11] ;
 wire \top_ihp.oisc.regs[48][12] ;
 wire \top_ihp.oisc.regs[48][13] ;
 wire \top_ihp.oisc.regs[48][14] ;
 wire \top_ihp.oisc.regs[48][15] ;
 wire \top_ihp.oisc.regs[48][16] ;
 wire \top_ihp.oisc.regs[48][17] ;
 wire \top_ihp.oisc.regs[48][18] ;
 wire \top_ihp.oisc.regs[48][19] ;
 wire \top_ihp.oisc.regs[48][1] ;
 wire \top_ihp.oisc.regs[48][20] ;
 wire \top_ihp.oisc.regs[48][21] ;
 wire \top_ihp.oisc.regs[48][22] ;
 wire \top_ihp.oisc.regs[48][23] ;
 wire \top_ihp.oisc.regs[48][24] ;
 wire \top_ihp.oisc.regs[48][25] ;
 wire \top_ihp.oisc.regs[48][26] ;
 wire \top_ihp.oisc.regs[48][27] ;
 wire \top_ihp.oisc.regs[48][28] ;
 wire \top_ihp.oisc.regs[48][29] ;
 wire \top_ihp.oisc.regs[48][2] ;
 wire \top_ihp.oisc.regs[48][30] ;
 wire \top_ihp.oisc.regs[48][31] ;
 wire \top_ihp.oisc.regs[48][3] ;
 wire \top_ihp.oisc.regs[48][4] ;
 wire \top_ihp.oisc.regs[48][5] ;
 wire \top_ihp.oisc.regs[48][6] ;
 wire \top_ihp.oisc.regs[48][7] ;
 wire \top_ihp.oisc.regs[48][8] ;
 wire \top_ihp.oisc.regs[48][9] ;
 wire \top_ihp.oisc.regs[49][0] ;
 wire \top_ihp.oisc.regs[49][10] ;
 wire \top_ihp.oisc.regs[49][11] ;
 wire \top_ihp.oisc.regs[49][12] ;
 wire \top_ihp.oisc.regs[49][13] ;
 wire \top_ihp.oisc.regs[49][14] ;
 wire \top_ihp.oisc.regs[49][15] ;
 wire \top_ihp.oisc.regs[49][16] ;
 wire \top_ihp.oisc.regs[49][17] ;
 wire \top_ihp.oisc.regs[49][18] ;
 wire \top_ihp.oisc.regs[49][19] ;
 wire \top_ihp.oisc.regs[49][1] ;
 wire \top_ihp.oisc.regs[49][20] ;
 wire \top_ihp.oisc.regs[49][21] ;
 wire \top_ihp.oisc.regs[49][22] ;
 wire \top_ihp.oisc.regs[49][23] ;
 wire \top_ihp.oisc.regs[49][24] ;
 wire \top_ihp.oisc.regs[49][25] ;
 wire \top_ihp.oisc.regs[49][26] ;
 wire \top_ihp.oisc.regs[49][27] ;
 wire \top_ihp.oisc.regs[49][28] ;
 wire \top_ihp.oisc.regs[49][29] ;
 wire \top_ihp.oisc.regs[49][2] ;
 wire \top_ihp.oisc.regs[49][30] ;
 wire \top_ihp.oisc.regs[49][31] ;
 wire \top_ihp.oisc.regs[49][3] ;
 wire \top_ihp.oisc.regs[49][4] ;
 wire \top_ihp.oisc.regs[49][5] ;
 wire \top_ihp.oisc.regs[49][6] ;
 wire \top_ihp.oisc.regs[49][7] ;
 wire \top_ihp.oisc.regs[49][8] ;
 wire \top_ihp.oisc.regs[49][9] ;
 wire \top_ihp.oisc.regs[4][0] ;
 wire \top_ihp.oisc.regs[4][10] ;
 wire \top_ihp.oisc.regs[4][11] ;
 wire \top_ihp.oisc.regs[4][12] ;
 wire \top_ihp.oisc.regs[4][13] ;
 wire \top_ihp.oisc.regs[4][14] ;
 wire \top_ihp.oisc.regs[4][15] ;
 wire \top_ihp.oisc.regs[4][16] ;
 wire \top_ihp.oisc.regs[4][17] ;
 wire \top_ihp.oisc.regs[4][18] ;
 wire \top_ihp.oisc.regs[4][19] ;
 wire \top_ihp.oisc.regs[4][1] ;
 wire \top_ihp.oisc.regs[4][20] ;
 wire \top_ihp.oisc.regs[4][21] ;
 wire \top_ihp.oisc.regs[4][22] ;
 wire \top_ihp.oisc.regs[4][23] ;
 wire \top_ihp.oisc.regs[4][24] ;
 wire \top_ihp.oisc.regs[4][25] ;
 wire \top_ihp.oisc.regs[4][26] ;
 wire \top_ihp.oisc.regs[4][27] ;
 wire \top_ihp.oisc.regs[4][28] ;
 wire \top_ihp.oisc.regs[4][29] ;
 wire \top_ihp.oisc.regs[4][2] ;
 wire \top_ihp.oisc.regs[4][30] ;
 wire \top_ihp.oisc.regs[4][31] ;
 wire \top_ihp.oisc.regs[4][3] ;
 wire \top_ihp.oisc.regs[4][4] ;
 wire \top_ihp.oisc.regs[4][5] ;
 wire \top_ihp.oisc.regs[4][6] ;
 wire \top_ihp.oisc.regs[4][7] ;
 wire \top_ihp.oisc.regs[4][8] ;
 wire \top_ihp.oisc.regs[4][9] ;
 wire \top_ihp.oisc.regs[50][0] ;
 wire \top_ihp.oisc.regs[50][10] ;
 wire \top_ihp.oisc.regs[50][11] ;
 wire \top_ihp.oisc.regs[50][12] ;
 wire \top_ihp.oisc.regs[50][13] ;
 wire \top_ihp.oisc.regs[50][14] ;
 wire \top_ihp.oisc.regs[50][15] ;
 wire \top_ihp.oisc.regs[50][16] ;
 wire \top_ihp.oisc.regs[50][17] ;
 wire \top_ihp.oisc.regs[50][18] ;
 wire \top_ihp.oisc.regs[50][19] ;
 wire \top_ihp.oisc.regs[50][1] ;
 wire \top_ihp.oisc.regs[50][20] ;
 wire \top_ihp.oisc.regs[50][21] ;
 wire \top_ihp.oisc.regs[50][22] ;
 wire \top_ihp.oisc.regs[50][23] ;
 wire \top_ihp.oisc.regs[50][24] ;
 wire \top_ihp.oisc.regs[50][25] ;
 wire \top_ihp.oisc.regs[50][26] ;
 wire \top_ihp.oisc.regs[50][27] ;
 wire \top_ihp.oisc.regs[50][28] ;
 wire \top_ihp.oisc.regs[50][29] ;
 wire \top_ihp.oisc.regs[50][2] ;
 wire \top_ihp.oisc.regs[50][30] ;
 wire \top_ihp.oisc.regs[50][31] ;
 wire \top_ihp.oisc.regs[50][3] ;
 wire \top_ihp.oisc.regs[50][4] ;
 wire \top_ihp.oisc.regs[50][5] ;
 wire \top_ihp.oisc.regs[50][6] ;
 wire \top_ihp.oisc.regs[50][7] ;
 wire \top_ihp.oisc.regs[50][8] ;
 wire \top_ihp.oisc.regs[50][9] ;
 wire \top_ihp.oisc.regs[51][0] ;
 wire \top_ihp.oisc.regs[51][10] ;
 wire \top_ihp.oisc.regs[51][11] ;
 wire \top_ihp.oisc.regs[51][12] ;
 wire \top_ihp.oisc.regs[51][13] ;
 wire \top_ihp.oisc.regs[51][14] ;
 wire \top_ihp.oisc.regs[51][15] ;
 wire \top_ihp.oisc.regs[51][16] ;
 wire \top_ihp.oisc.regs[51][17] ;
 wire \top_ihp.oisc.regs[51][18] ;
 wire \top_ihp.oisc.regs[51][19] ;
 wire \top_ihp.oisc.regs[51][1] ;
 wire \top_ihp.oisc.regs[51][20] ;
 wire \top_ihp.oisc.regs[51][21] ;
 wire \top_ihp.oisc.regs[51][22] ;
 wire \top_ihp.oisc.regs[51][23] ;
 wire \top_ihp.oisc.regs[51][24] ;
 wire \top_ihp.oisc.regs[51][25] ;
 wire \top_ihp.oisc.regs[51][26] ;
 wire \top_ihp.oisc.regs[51][27] ;
 wire \top_ihp.oisc.regs[51][28] ;
 wire \top_ihp.oisc.regs[51][29] ;
 wire \top_ihp.oisc.regs[51][2] ;
 wire \top_ihp.oisc.regs[51][30] ;
 wire \top_ihp.oisc.regs[51][31] ;
 wire \top_ihp.oisc.regs[51][3] ;
 wire \top_ihp.oisc.regs[51][4] ;
 wire \top_ihp.oisc.regs[51][5] ;
 wire \top_ihp.oisc.regs[51][6] ;
 wire \top_ihp.oisc.regs[51][7] ;
 wire \top_ihp.oisc.regs[51][8] ;
 wire \top_ihp.oisc.regs[51][9] ;
 wire \top_ihp.oisc.regs[52][0] ;
 wire \top_ihp.oisc.regs[52][10] ;
 wire \top_ihp.oisc.regs[52][11] ;
 wire \top_ihp.oisc.regs[52][12] ;
 wire \top_ihp.oisc.regs[52][13] ;
 wire \top_ihp.oisc.regs[52][14] ;
 wire \top_ihp.oisc.regs[52][15] ;
 wire \top_ihp.oisc.regs[52][16] ;
 wire \top_ihp.oisc.regs[52][17] ;
 wire \top_ihp.oisc.regs[52][18] ;
 wire \top_ihp.oisc.regs[52][19] ;
 wire \top_ihp.oisc.regs[52][1] ;
 wire \top_ihp.oisc.regs[52][20] ;
 wire \top_ihp.oisc.regs[52][21] ;
 wire \top_ihp.oisc.regs[52][22] ;
 wire \top_ihp.oisc.regs[52][23] ;
 wire \top_ihp.oisc.regs[52][24] ;
 wire \top_ihp.oisc.regs[52][25] ;
 wire \top_ihp.oisc.regs[52][26] ;
 wire \top_ihp.oisc.regs[52][27] ;
 wire \top_ihp.oisc.regs[52][28] ;
 wire \top_ihp.oisc.regs[52][29] ;
 wire \top_ihp.oisc.regs[52][2] ;
 wire \top_ihp.oisc.regs[52][30] ;
 wire \top_ihp.oisc.regs[52][31] ;
 wire \top_ihp.oisc.regs[52][3] ;
 wire \top_ihp.oisc.regs[52][4] ;
 wire \top_ihp.oisc.regs[52][5] ;
 wire \top_ihp.oisc.regs[52][6] ;
 wire \top_ihp.oisc.regs[52][7] ;
 wire \top_ihp.oisc.regs[52][8] ;
 wire \top_ihp.oisc.regs[52][9] ;
 wire \top_ihp.oisc.regs[53][0] ;
 wire \top_ihp.oisc.regs[53][10] ;
 wire \top_ihp.oisc.regs[53][11] ;
 wire \top_ihp.oisc.regs[53][12] ;
 wire \top_ihp.oisc.regs[53][13] ;
 wire \top_ihp.oisc.regs[53][14] ;
 wire \top_ihp.oisc.regs[53][15] ;
 wire \top_ihp.oisc.regs[53][16] ;
 wire \top_ihp.oisc.regs[53][17] ;
 wire \top_ihp.oisc.regs[53][18] ;
 wire \top_ihp.oisc.regs[53][19] ;
 wire \top_ihp.oisc.regs[53][1] ;
 wire \top_ihp.oisc.regs[53][20] ;
 wire \top_ihp.oisc.regs[53][21] ;
 wire \top_ihp.oisc.regs[53][22] ;
 wire \top_ihp.oisc.regs[53][23] ;
 wire \top_ihp.oisc.regs[53][24] ;
 wire \top_ihp.oisc.regs[53][25] ;
 wire \top_ihp.oisc.regs[53][26] ;
 wire \top_ihp.oisc.regs[53][27] ;
 wire \top_ihp.oisc.regs[53][28] ;
 wire \top_ihp.oisc.regs[53][29] ;
 wire \top_ihp.oisc.regs[53][2] ;
 wire \top_ihp.oisc.regs[53][30] ;
 wire \top_ihp.oisc.regs[53][31] ;
 wire \top_ihp.oisc.regs[53][3] ;
 wire \top_ihp.oisc.regs[53][4] ;
 wire \top_ihp.oisc.regs[53][5] ;
 wire \top_ihp.oisc.regs[53][6] ;
 wire \top_ihp.oisc.regs[53][7] ;
 wire \top_ihp.oisc.regs[53][8] ;
 wire \top_ihp.oisc.regs[53][9] ;
 wire \top_ihp.oisc.regs[54][0] ;
 wire \top_ihp.oisc.regs[54][10] ;
 wire \top_ihp.oisc.regs[54][11] ;
 wire \top_ihp.oisc.regs[54][12] ;
 wire \top_ihp.oisc.regs[54][13] ;
 wire \top_ihp.oisc.regs[54][14] ;
 wire \top_ihp.oisc.regs[54][15] ;
 wire \top_ihp.oisc.regs[54][16] ;
 wire \top_ihp.oisc.regs[54][17] ;
 wire \top_ihp.oisc.regs[54][18] ;
 wire \top_ihp.oisc.regs[54][19] ;
 wire \top_ihp.oisc.regs[54][1] ;
 wire \top_ihp.oisc.regs[54][20] ;
 wire \top_ihp.oisc.regs[54][21] ;
 wire \top_ihp.oisc.regs[54][22] ;
 wire \top_ihp.oisc.regs[54][23] ;
 wire \top_ihp.oisc.regs[54][24] ;
 wire \top_ihp.oisc.regs[54][25] ;
 wire \top_ihp.oisc.regs[54][26] ;
 wire \top_ihp.oisc.regs[54][27] ;
 wire \top_ihp.oisc.regs[54][28] ;
 wire \top_ihp.oisc.regs[54][29] ;
 wire \top_ihp.oisc.regs[54][2] ;
 wire \top_ihp.oisc.regs[54][30] ;
 wire \top_ihp.oisc.regs[54][31] ;
 wire \top_ihp.oisc.regs[54][3] ;
 wire \top_ihp.oisc.regs[54][4] ;
 wire \top_ihp.oisc.regs[54][5] ;
 wire \top_ihp.oisc.regs[54][6] ;
 wire \top_ihp.oisc.regs[54][7] ;
 wire \top_ihp.oisc.regs[54][8] ;
 wire \top_ihp.oisc.regs[54][9] ;
 wire \top_ihp.oisc.regs[55][0] ;
 wire \top_ihp.oisc.regs[55][10] ;
 wire \top_ihp.oisc.regs[55][11] ;
 wire \top_ihp.oisc.regs[55][12] ;
 wire \top_ihp.oisc.regs[55][13] ;
 wire \top_ihp.oisc.regs[55][14] ;
 wire \top_ihp.oisc.regs[55][15] ;
 wire \top_ihp.oisc.regs[55][16] ;
 wire \top_ihp.oisc.regs[55][17] ;
 wire \top_ihp.oisc.regs[55][18] ;
 wire \top_ihp.oisc.regs[55][19] ;
 wire \top_ihp.oisc.regs[55][1] ;
 wire \top_ihp.oisc.regs[55][20] ;
 wire \top_ihp.oisc.regs[55][21] ;
 wire \top_ihp.oisc.regs[55][22] ;
 wire \top_ihp.oisc.regs[55][23] ;
 wire \top_ihp.oisc.regs[55][24] ;
 wire \top_ihp.oisc.regs[55][25] ;
 wire \top_ihp.oisc.regs[55][26] ;
 wire \top_ihp.oisc.regs[55][27] ;
 wire \top_ihp.oisc.regs[55][28] ;
 wire \top_ihp.oisc.regs[55][29] ;
 wire \top_ihp.oisc.regs[55][2] ;
 wire \top_ihp.oisc.regs[55][30] ;
 wire \top_ihp.oisc.regs[55][31] ;
 wire \top_ihp.oisc.regs[55][3] ;
 wire \top_ihp.oisc.regs[55][4] ;
 wire \top_ihp.oisc.regs[55][5] ;
 wire \top_ihp.oisc.regs[55][6] ;
 wire \top_ihp.oisc.regs[55][7] ;
 wire \top_ihp.oisc.regs[55][8] ;
 wire \top_ihp.oisc.regs[55][9] ;
 wire \top_ihp.oisc.regs[56][0] ;
 wire \top_ihp.oisc.regs[56][10] ;
 wire \top_ihp.oisc.regs[56][11] ;
 wire \top_ihp.oisc.regs[56][12] ;
 wire \top_ihp.oisc.regs[56][13] ;
 wire \top_ihp.oisc.regs[56][14] ;
 wire \top_ihp.oisc.regs[56][15] ;
 wire \top_ihp.oisc.regs[56][16] ;
 wire \top_ihp.oisc.regs[56][17] ;
 wire \top_ihp.oisc.regs[56][18] ;
 wire \top_ihp.oisc.regs[56][19] ;
 wire \top_ihp.oisc.regs[56][1] ;
 wire \top_ihp.oisc.regs[56][20] ;
 wire \top_ihp.oisc.regs[56][21] ;
 wire \top_ihp.oisc.regs[56][22] ;
 wire \top_ihp.oisc.regs[56][23] ;
 wire \top_ihp.oisc.regs[56][24] ;
 wire \top_ihp.oisc.regs[56][25] ;
 wire \top_ihp.oisc.regs[56][26] ;
 wire \top_ihp.oisc.regs[56][27] ;
 wire \top_ihp.oisc.regs[56][28] ;
 wire \top_ihp.oisc.regs[56][29] ;
 wire \top_ihp.oisc.regs[56][2] ;
 wire \top_ihp.oisc.regs[56][30] ;
 wire \top_ihp.oisc.regs[56][31] ;
 wire \top_ihp.oisc.regs[56][3] ;
 wire \top_ihp.oisc.regs[56][4] ;
 wire \top_ihp.oisc.regs[56][5] ;
 wire \top_ihp.oisc.regs[56][6] ;
 wire \top_ihp.oisc.regs[56][7] ;
 wire \top_ihp.oisc.regs[56][8] ;
 wire \top_ihp.oisc.regs[56][9] ;
 wire \top_ihp.oisc.regs[57][0] ;
 wire \top_ihp.oisc.regs[57][10] ;
 wire \top_ihp.oisc.regs[57][11] ;
 wire \top_ihp.oisc.regs[57][12] ;
 wire \top_ihp.oisc.regs[57][13] ;
 wire \top_ihp.oisc.regs[57][14] ;
 wire \top_ihp.oisc.regs[57][15] ;
 wire \top_ihp.oisc.regs[57][16] ;
 wire \top_ihp.oisc.regs[57][17] ;
 wire \top_ihp.oisc.regs[57][18] ;
 wire \top_ihp.oisc.regs[57][19] ;
 wire \top_ihp.oisc.regs[57][1] ;
 wire \top_ihp.oisc.regs[57][20] ;
 wire \top_ihp.oisc.regs[57][21] ;
 wire \top_ihp.oisc.regs[57][22] ;
 wire \top_ihp.oisc.regs[57][23] ;
 wire \top_ihp.oisc.regs[57][24] ;
 wire \top_ihp.oisc.regs[57][25] ;
 wire \top_ihp.oisc.regs[57][26] ;
 wire \top_ihp.oisc.regs[57][27] ;
 wire \top_ihp.oisc.regs[57][28] ;
 wire \top_ihp.oisc.regs[57][29] ;
 wire \top_ihp.oisc.regs[57][2] ;
 wire \top_ihp.oisc.regs[57][30] ;
 wire \top_ihp.oisc.regs[57][31] ;
 wire \top_ihp.oisc.regs[57][3] ;
 wire \top_ihp.oisc.regs[57][4] ;
 wire \top_ihp.oisc.regs[57][5] ;
 wire \top_ihp.oisc.regs[57][6] ;
 wire \top_ihp.oisc.regs[57][7] ;
 wire \top_ihp.oisc.regs[57][8] ;
 wire \top_ihp.oisc.regs[57][9] ;
 wire \top_ihp.oisc.regs[58][0] ;
 wire \top_ihp.oisc.regs[58][10] ;
 wire \top_ihp.oisc.regs[58][11] ;
 wire \top_ihp.oisc.regs[58][12] ;
 wire \top_ihp.oisc.regs[58][13] ;
 wire \top_ihp.oisc.regs[58][14] ;
 wire \top_ihp.oisc.regs[58][15] ;
 wire \top_ihp.oisc.regs[58][16] ;
 wire \top_ihp.oisc.regs[58][17] ;
 wire \top_ihp.oisc.regs[58][18] ;
 wire \top_ihp.oisc.regs[58][19] ;
 wire \top_ihp.oisc.regs[58][1] ;
 wire \top_ihp.oisc.regs[58][20] ;
 wire \top_ihp.oisc.regs[58][21] ;
 wire \top_ihp.oisc.regs[58][22] ;
 wire \top_ihp.oisc.regs[58][23] ;
 wire \top_ihp.oisc.regs[58][24] ;
 wire \top_ihp.oisc.regs[58][25] ;
 wire \top_ihp.oisc.regs[58][26] ;
 wire \top_ihp.oisc.regs[58][27] ;
 wire \top_ihp.oisc.regs[58][28] ;
 wire \top_ihp.oisc.regs[58][29] ;
 wire \top_ihp.oisc.regs[58][2] ;
 wire \top_ihp.oisc.regs[58][30] ;
 wire \top_ihp.oisc.regs[58][31] ;
 wire \top_ihp.oisc.regs[58][3] ;
 wire \top_ihp.oisc.regs[58][4] ;
 wire \top_ihp.oisc.regs[58][5] ;
 wire \top_ihp.oisc.regs[58][6] ;
 wire \top_ihp.oisc.regs[58][7] ;
 wire \top_ihp.oisc.regs[58][8] ;
 wire \top_ihp.oisc.regs[58][9] ;
 wire \top_ihp.oisc.regs[59][0] ;
 wire \top_ihp.oisc.regs[59][10] ;
 wire \top_ihp.oisc.regs[59][11] ;
 wire \top_ihp.oisc.regs[59][12] ;
 wire \top_ihp.oisc.regs[59][13] ;
 wire \top_ihp.oisc.regs[59][14] ;
 wire \top_ihp.oisc.regs[59][15] ;
 wire \top_ihp.oisc.regs[59][16] ;
 wire \top_ihp.oisc.regs[59][17] ;
 wire \top_ihp.oisc.regs[59][18] ;
 wire \top_ihp.oisc.regs[59][19] ;
 wire \top_ihp.oisc.regs[59][1] ;
 wire \top_ihp.oisc.regs[59][20] ;
 wire \top_ihp.oisc.regs[59][21] ;
 wire \top_ihp.oisc.regs[59][22] ;
 wire \top_ihp.oisc.regs[59][23] ;
 wire \top_ihp.oisc.regs[59][24] ;
 wire \top_ihp.oisc.regs[59][25] ;
 wire \top_ihp.oisc.regs[59][26] ;
 wire \top_ihp.oisc.regs[59][27] ;
 wire \top_ihp.oisc.regs[59][28] ;
 wire \top_ihp.oisc.regs[59][29] ;
 wire \top_ihp.oisc.regs[59][2] ;
 wire \top_ihp.oisc.regs[59][30] ;
 wire \top_ihp.oisc.regs[59][31] ;
 wire \top_ihp.oisc.regs[59][3] ;
 wire \top_ihp.oisc.regs[59][4] ;
 wire \top_ihp.oisc.regs[59][5] ;
 wire \top_ihp.oisc.regs[59][6] ;
 wire \top_ihp.oisc.regs[59][7] ;
 wire \top_ihp.oisc.regs[59][8] ;
 wire \top_ihp.oisc.regs[59][9] ;
 wire \top_ihp.oisc.regs[5][0] ;
 wire \top_ihp.oisc.regs[5][10] ;
 wire \top_ihp.oisc.regs[5][11] ;
 wire \top_ihp.oisc.regs[5][12] ;
 wire \top_ihp.oisc.regs[5][13] ;
 wire \top_ihp.oisc.regs[5][14] ;
 wire \top_ihp.oisc.regs[5][15] ;
 wire \top_ihp.oisc.regs[5][16] ;
 wire \top_ihp.oisc.regs[5][17] ;
 wire \top_ihp.oisc.regs[5][18] ;
 wire \top_ihp.oisc.regs[5][19] ;
 wire \top_ihp.oisc.regs[5][1] ;
 wire \top_ihp.oisc.regs[5][20] ;
 wire \top_ihp.oisc.regs[5][21] ;
 wire \top_ihp.oisc.regs[5][22] ;
 wire \top_ihp.oisc.regs[5][23] ;
 wire \top_ihp.oisc.regs[5][24] ;
 wire \top_ihp.oisc.regs[5][25] ;
 wire \top_ihp.oisc.regs[5][26] ;
 wire \top_ihp.oisc.regs[5][27] ;
 wire \top_ihp.oisc.regs[5][28] ;
 wire \top_ihp.oisc.regs[5][29] ;
 wire \top_ihp.oisc.regs[5][2] ;
 wire \top_ihp.oisc.regs[5][30] ;
 wire \top_ihp.oisc.regs[5][31] ;
 wire \top_ihp.oisc.regs[5][3] ;
 wire \top_ihp.oisc.regs[5][4] ;
 wire \top_ihp.oisc.regs[5][5] ;
 wire \top_ihp.oisc.regs[5][6] ;
 wire \top_ihp.oisc.regs[5][7] ;
 wire \top_ihp.oisc.regs[5][8] ;
 wire \top_ihp.oisc.regs[5][9] ;
 wire \top_ihp.oisc.regs[60][0] ;
 wire \top_ihp.oisc.regs[60][10] ;
 wire \top_ihp.oisc.regs[60][11] ;
 wire \top_ihp.oisc.regs[60][12] ;
 wire \top_ihp.oisc.regs[60][13] ;
 wire \top_ihp.oisc.regs[60][14] ;
 wire \top_ihp.oisc.regs[60][15] ;
 wire \top_ihp.oisc.regs[60][16] ;
 wire \top_ihp.oisc.regs[60][17] ;
 wire \top_ihp.oisc.regs[60][18] ;
 wire \top_ihp.oisc.regs[60][19] ;
 wire \top_ihp.oisc.regs[60][1] ;
 wire \top_ihp.oisc.regs[60][20] ;
 wire \top_ihp.oisc.regs[60][21] ;
 wire \top_ihp.oisc.regs[60][22] ;
 wire \top_ihp.oisc.regs[60][23] ;
 wire \top_ihp.oisc.regs[60][24] ;
 wire \top_ihp.oisc.regs[60][25] ;
 wire \top_ihp.oisc.regs[60][26] ;
 wire \top_ihp.oisc.regs[60][27] ;
 wire \top_ihp.oisc.regs[60][28] ;
 wire \top_ihp.oisc.regs[60][29] ;
 wire \top_ihp.oisc.regs[60][2] ;
 wire \top_ihp.oisc.regs[60][30] ;
 wire \top_ihp.oisc.regs[60][31] ;
 wire \top_ihp.oisc.regs[60][3] ;
 wire \top_ihp.oisc.regs[60][4] ;
 wire \top_ihp.oisc.regs[60][5] ;
 wire \top_ihp.oisc.regs[60][6] ;
 wire \top_ihp.oisc.regs[60][7] ;
 wire \top_ihp.oisc.regs[60][8] ;
 wire \top_ihp.oisc.regs[60][9] ;
 wire \top_ihp.oisc.regs[61][0] ;
 wire \top_ihp.oisc.regs[61][10] ;
 wire \top_ihp.oisc.regs[61][11] ;
 wire \top_ihp.oisc.regs[61][12] ;
 wire \top_ihp.oisc.regs[61][13] ;
 wire \top_ihp.oisc.regs[61][14] ;
 wire \top_ihp.oisc.regs[61][15] ;
 wire \top_ihp.oisc.regs[61][16] ;
 wire \top_ihp.oisc.regs[61][17] ;
 wire \top_ihp.oisc.regs[61][18] ;
 wire \top_ihp.oisc.regs[61][19] ;
 wire \top_ihp.oisc.regs[61][1] ;
 wire \top_ihp.oisc.regs[61][20] ;
 wire \top_ihp.oisc.regs[61][21] ;
 wire \top_ihp.oisc.regs[61][22] ;
 wire \top_ihp.oisc.regs[61][23] ;
 wire \top_ihp.oisc.regs[61][24] ;
 wire \top_ihp.oisc.regs[61][25] ;
 wire \top_ihp.oisc.regs[61][26] ;
 wire \top_ihp.oisc.regs[61][27] ;
 wire \top_ihp.oisc.regs[61][28] ;
 wire \top_ihp.oisc.regs[61][29] ;
 wire \top_ihp.oisc.regs[61][2] ;
 wire \top_ihp.oisc.regs[61][30] ;
 wire \top_ihp.oisc.regs[61][31] ;
 wire \top_ihp.oisc.regs[61][3] ;
 wire \top_ihp.oisc.regs[61][4] ;
 wire \top_ihp.oisc.regs[61][5] ;
 wire \top_ihp.oisc.regs[61][6] ;
 wire \top_ihp.oisc.regs[61][7] ;
 wire \top_ihp.oisc.regs[61][8] ;
 wire \top_ihp.oisc.regs[61][9] ;
 wire \top_ihp.oisc.regs[62][0] ;
 wire \top_ihp.oisc.regs[62][10] ;
 wire \top_ihp.oisc.regs[62][11] ;
 wire \top_ihp.oisc.regs[62][12] ;
 wire \top_ihp.oisc.regs[62][13] ;
 wire \top_ihp.oisc.regs[62][14] ;
 wire \top_ihp.oisc.regs[62][15] ;
 wire \top_ihp.oisc.regs[62][16] ;
 wire \top_ihp.oisc.regs[62][17] ;
 wire \top_ihp.oisc.regs[62][18] ;
 wire \top_ihp.oisc.regs[62][19] ;
 wire \top_ihp.oisc.regs[62][1] ;
 wire \top_ihp.oisc.regs[62][20] ;
 wire \top_ihp.oisc.regs[62][21] ;
 wire \top_ihp.oisc.regs[62][22] ;
 wire \top_ihp.oisc.regs[62][23] ;
 wire \top_ihp.oisc.regs[62][24] ;
 wire \top_ihp.oisc.regs[62][25] ;
 wire \top_ihp.oisc.regs[62][26] ;
 wire \top_ihp.oisc.regs[62][27] ;
 wire \top_ihp.oisc.regs[62][28] ;
 wire \top_ihp.oisc.regs[62][29] ;
 wire \top_ihp.oisc.regs[62][2] ;
 wire \top_ihp.oisc.regs[62][30] ;
 wire \top_ihp.oisc.regs[62][31] ;
 wire \top_ihp.oisc.regs[62][3] ;
 wire \top_ihp.oisc.regs[62][4] ;
 wire \top_ihp.oisc.regs[62][5] ;
 wire \top_ihp.oisc.regs[62][6] ;
 wire \top_ihp.oisc.regs[62][7] ;
 wire \top_ihp.oisc.regs[62][8] ;
 wire \top_ihp.oisc.regs[62][9] ;
 wire \top_ihp.oisc.regs[63][0] ;
 wire \top_ihp.oisc.regs[63][10] ;
 wire \top_ihp.oisc.regs[63][11] ;
 wire \top_ihp.oisc.regs[63][12] ;
 wire \top_ihp.oisc.regs[63][13] ;
 wire \top_ihp.oisc.regs[63][14] ;
 wire \top_ihp.oisc.regs[63][15] ;
 wire \top_ihp.oisc.regs[63][16] ;
 wire \top_ihp.oisc.regs[63][17] ;
 wire \top_ihp.oisc.regs[63][18] ;
 wire \top_ihp.oisc.regs[63][19] ;
 wire \top_ihp.oisc.regs[63][1] ;
 wire \top_ihp.oisc.regs[63][20] ;
 wire \top_ihp.oisc.regs[63][21] ;
 wire \top_ihp.oisc.regs[63][22] ;
 wire \top_ihp.oisc.regs[63][23] ;
 wire \top_ihp.oisc.regs[63][24] ;
 wire \top_ihp.oisc.regs[63][25] ;
 wire \top_ihp.oisc.regs[63][26] ;
 wire \top_ihp.oisc.regs[63][27] ;
 wire \top_ihp.oisc.regs[63][28] ;
 wire \top_ihp.oisc.regs[63][29] ;
 wire \top_ihp.oisc.regs[63][2] ;
 wire \top_ihp.oisc.regs[63][30] ;
 wire \top_ihp.oisc.regs[63][31] ;
 wire \top_ihp.oisc.regs[63][3] ;
 wire \top_ihp.oisc.regs[63][4] ;
 wire \top_ihp.oisc.regs[63][5] ;
 wire \top_ihp.oisc.regs[63][6] ;
 wire \top_ihp.oisc.regs[63][7] ;
 wire \top_ihp.oisc.regs[63][8] ;
 wire \top_ihp.oisc.regs[63][9] ;
 wire \top_ihp.oisc.regs[6][0] ;
 wire \top_ihp.oisc.regs[6][10] ;
 wire \top_ihp.oisc.regs[6][11] ;
 wire \top_ihp.oisc.regs[6][12] ;
 wire \top_ihp.oisc.regs[6][13] ;
 wire \top_ihp.oisc.regs[6][14] ;
 wire \top_ihp.oisc.regs[6][15] ;
 wire \top_ihp.oisc.regs[6][16] ;
 wire \top_ihp.oisc.regs[6][17] ;
 wire \top_ihp.oisc.regs[6][18] ;
 wire \top_ihp.oisc.regs[6][19] ;
 wire \top_ihp.oisc.regs[6][1] ;
 wire \top_ihp.oisc.regs[6][20] ;
 wire \top_ihp.oisc.regs[6][21] ;
 wire \top_ihp.oisc.regs[6][22] ;
 wire \top_ihp.oisc.regs[6][23] ;
 wire \top_ihp.oisc.regs[6][24] ;
 wire \top_ihp.oisc.regs[6][25] ;
 wire \top_ihp.oisc.regs[6][26] ;
 wire \top_ihp.oisc.regs[6][27] ;
 wire \top_ihp.oisc.regs[6][28] ;
 wire \top_ihp.oisc.regs[6][29] ;
 wire \top_ihp.oisc.regs[6][2] ;
 wire \top_ihp.oisc.regs[6][30] ;
 wire \top_ihp.oisc.regs[6][31] ;
 wire \top_ihp.oisc.regs[6][3] ;
 wire \top_ihp.oisc.regs[6][4] ;
 wire \top_ihp.oisc.regs[6][5] ;
 wire \top_ihp.oisc.regs[6][6] ;
 wire \top_ihp.oisc.regs[6][7] ;
 wire \top_ihp.oisc.regs[6][8] ;
 wire \top_ihp.oisc.regs[6][9] ;
 wire \top_ihp.oisc.regs[7][0] ;
 wire \top_ihp.oisc.regs[7][10] ;
 wire \top_ihp.oisc.regs[7][11] ;
 wire \top_ihp.oisc.regs[7][12] ;
 wire \top_ihp.oisc.regs[7][13] ;
 wire \top_ihp.oisc.regs[7][14] ;
 wire \top_ihp.oisc.regs[7][15] ;
 wire \top_ihp.oisc.regs[7][16] ;
 wire \top_ihp.oisc.regs[7][17] ;
 wire \top_ihp.oisc.regs[7][18] ;
 wire \top_ihp.oisc.regs[7][19] ;
 wire \top_ihp.oisc.regs[7][1] ;
 wire \top_ihp.oisc.regs[7][20] ;
 wire \top_ihp.oisc.regs[7][21] ;
 wire \top_ihp.oisc.regs[7][22] ;
 wire \top_ihp.oisc.regs[7][23] ;
 wire \top_ihp.oisc.regs[7][24] ;
 wire \top_ihp.oisc.regs[7][25] ;
 wire \top_ihp.oisc.regs[7][26] ;
 wire \top_ihp.oisc.regs[7][27] ;
 wire \top_ihp.oisc.regs[7][28] ;
 wire \top_ihp.oisc.regs[7][29] ;
 wire \top_ihp.oisc.regs[7][2] ;
 wire \top_ihp.oisc.regs[7][30] ;
 wire \top_ihp.oisc.regs[7][31] ;
 wire \top_ihp.oisc.regs[7][3] ;
 wire \top_ihp.oisc.regs[7][4] ;
 wire \top_ihp.oisc.regs[7][5] ;
 wire \top_ihp.oisc.regs[7][6] ;
 wire \top_ihp.oisc.regs[7][7] ;
 wire \top_ihp.oisc.regs[7][8] ;
 wire \top_ihp.oisc.regs[7][9] ;
 wire \top_ihp.oisc.regs[8][0] ;
 wire \top_ihp.oisc.regs[8][10] ;
 wire \top_ihp.oisc.regs[8][11] ;
 wire \top_ihp.oisc.regs[8][12] ;
 wire \top_ihp.oisc.regs[8][13] ;
 wire \top_ihp.oisc.regs[8][14] ;
 wire \top_ihp.oisc.regs[8][15] ;
 wire \top_ihp.oisc.regs[8][16] ;
 wire \top_ihp.oisc.regs[8][17] ;
 wire \top_ihp.oisc.regs[8][18] ;
 wire \top_ihp.oisc.regs[8][19] ;
 wire \top_ihp.oisc.regs[8][1] ;
 wire \top_ihp.oisc.regs[8][20] ;
 wire \top_ihp.oisc.regs[8][21] ;
 wire \top_ihp.oisc.regs[8][22] ;
 wire \top_ihp.oisc.regs[8][23] ;
 wire \top_ihp.oisc.regs[8][24] ;
 wire \top_ihp.oisc.regs[8][25] ;
 wire \top_ihp.oisc.regs[8][26] ;
 wire \top_ihp.oisc.regs[8][27] ;
 wire \top_ihp.oisc.regs[8][28] ;
 wire \top_ihp.oisc.regs[8][29] ;
 wire \top_ihp.oisc.regs[8][2] ;
 wire \top_ihp.oisc.regs[8][30] ;
 wire \top_ihp.oisc.regs[8][31] ;
 wire \top_ihp.oisc.regs[8][3] ;
 wire \top_ihp.oisc.regs[8][4] ;
 wire \top_ihp.oisc.regs[8][5] ;
 wire \top_ihp.oisc.regs[8][6] ;
 wire \top_ihp.oisc.regs[8][7] ;
 wire \top_ihp.oisc.regs[8][8] ;
 wire \top_ihp.oisc.regs[8][9] ;
 wire \top_ihp.oisc.regs[9][0] ;
 wire \top_ihp.oisc.regs[9][10] ;
 wire \top_ihp.oisc.regs[9][11] ;
 wire \top_ihp.oisc.regs[9][12] ;
 wire \top_ihp.oisc.regs[9][13] ;
 wire \top_ihp.oisc.regs[9][14] ;
 wire \top_ihp.oisc.regs[9][15] ;
 wire \top_ihp.oisc.regs[9][16] ;
 wire \top_ihp.oisc.regs[9][17] ;
 wire \top_ihp.oisc.regs[9][18] ;
 wire \top_ihp.oisc.regs[9][19] ;
 wire \top_ihp.oisc.regs[9][1] ;
 wire \top_ihp.oisc.regs[9][20] ;
 wire \top_ihp.oisc.regs[9][21] ;
 wire \top_ihp.oisc.regs[9][22] ;
 wire \top_ihp.oisc.regs[9][23] ;
 wire \top_ihp.oisc.regs[9][24] ;
 wire \top_ihp.oisc.regs[9][25] ;
 wire \top_ihp.oisc.regs[9][26] ;
 wire \top_ihp.oisc.regs[9][27] ;
 wire \top_ihp.oisc.regs[9][28] ;
 wire \top_ihp.oisc.regs[9][29] ;
 wire \top_ihp.oisc.regs[9][2] ;
 wire \top_ihp.oisc.regs[9][30] ;
 wire \top_ihp.oisc.regs[9][31] ;
 wire \top_ihp.oisc.regs[9][3] ;
 wire \top_ihp.oisc.regs[9][4] ;
 wire \top_ihp.oisc.regs[9][5] ;
 wire \top_ihp.oisc.regs[9][6] ;
 wire \top_ihp.oisc.regs[9][7] ;
 wire \top_ihp.oisc.regs[9][8] ;
 wire \top_ihp.oisc.regs[9][9] ;
 wire \top_ihp.oisc.state[0] ;
 wire \top_ihp.oisc.state[1] ;
 wire \top_ihp.oisc.state[2] ;
 wire \top_ihp.oisc.state[3] ;
 wire \top_ihp.oisc.state[4] ;
 wire \top_ihp.oisc.state[5] ;
 wire \top_ihp.oisc.state[6] ;
 wire \top_ihp.oisc.wb_adr_o[0] ;
 wire \top_ihp.oisc.wb_adr_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[0] ;
 wire \top_ihp.oisc.wb_dat_o[10] ;
 wire \top_ihp.oisc.wb_dat_o[11] ;
 wire \top_ihp.oisc.wb_dat_o[12] ;
 wire \top_ihp.oisc.wb_dat_o[13] ;
 wire \top_ihp.oisc.wb_dat_o[14] ;
 wire \top_ihp.oisc.wb_dat_o[15] ;
 wire \top_ihp.oisc.wb_dat_o[16] ;
 wire \top_ihp.oisc.wb_dat_o[17] ;
 wire \top_ihp.oisc.wb_dat_o[18] ;
 wire \top_ihp.oisc.wb_dat_o[19] ;
 wire \top_ihp.oisc.wb_dat_o[1] ;
 wire \top_ihp.oisc.wb_dat_o[20] ;
 wire \top_ihp.oisc.wb_dat_o[21] ;
 wire \top_ihp.oisc.wb_dat_o[22] ;
 wire \top_ihp.oisc.wb_dat_o[23] ;
 wire \top_ihp.oisc.wb_dat_o[24] ;
 wire \top_ihp.oisc.wb_dat_o[25] ;
 wire \top_ihp.oisc.wb_dat_o[26] ;
 wire \top_ihp.oisc.wb_dat_o[27] ;
 wire \top_ihp.oisc.wb_dat_o[28] ;
 wire \top_ihp.oisc.wb_dat_o[29] ;
 wire \top_ihp.oisc.wb_dat_o[2] ;
 wire \top_ihp.oisc.wb_dat_o[30] ;
 wire \top_ihp.oisc.wb_dat_o[31] ;
 wire \top_ihp.oisc.wb_dat_o[3] ;
 wire \top_ihp.oisc.wb_dat_o[4] ;
 wire \top_ihp.oisc.wb_dat_o[5] ;
 wire \top_ihp.oisc.wb_dat_o[6] ;
 wire \top_ihp.oisc.wb_dat_o[7] ;
 wire \top_ihp.oisc.wb_dat_o[8] ;
 wire \top_ihp.oisc.wb_dat_o[9] ;
 wire \top_ihp.ram_clk_o ;
 wire \top_ihp.ram_cs_o ;
 wire \top_ihp.ram_data_o ;
 wire \top_ihp.rom_clk_o ;
 wire \top_ihp.rom_cs_o ;
 wire \top_ihp.rom_data_o ;
 wire \top_ihp.spi_clk_o ;
 wire \top_ihp.spi_cs_o_1 ;
 wire \top_ihp.spi_cs_o_2 ;
 wire \top_ihp.spi_cs_o_3 ;
 wire \top_ihp.spi_data_o ;
 wire \top_ihp.tx ;
 wire \top_ihp.wb_ack_coproc ;
 wire \top_ihp.wb_ack_gpio ;
 wire \top_ihp.wb_ack_spi ;
 wire \top_ihp.wb_ack_uart ;
 wire \top_ihp.wb_coproc.dat_o[0] ;
 wire \top_ihp.wb_coproc.dat_o[10] ;
 wire \top_ihp.wb_coproc.dat_o[11] ;
 wire \top_ihp.wb_coproc.dat_o[12] ;
 wire \top_ihp.wb_coproc.dat_o[13] ;
 wire \top_ihp.wb_coproc.dat_o[14] ;
 wire \top_ihp.wb_coproc.dat_o[15] ;
 wire \top_ihp.wb_coproc.dat_o[16] ;
 wire \top_ihp.wb_coproc.dat_o[17] ;
 wire \top_ihp.wb_coproc.dat_o[18] ;
 wire \top_ihp.wb_coproc.dat_o[19] ;
 wire \top_ihp.wb_coproc.dat_o[1] ;
 wire \top_ihp.wb_coproc.dat_o[20] ;
 wire \top_ihp.wb_coproc.dat_o[21] ;
 wire \top_ihp.wb_coproc.dat_o[22] ;
 wire \top_ihp.wb_coproc.dat_o[23] ;
 wire \top_ihp.wb_coproc.dat_o[24] ;
 wire \top_ihp.wb_coproc.dat_o[25] ;
 wire \top_ihp.wb_coproc.dat_o[26] ;
 wire \top_ihp.wb_coproc.dat_o[27] ;
 wire \top_ihp.wb_coproc.dat_o[28] ;
 wire \top_ihp.wb_coproc.dat_o[29] ;
 wire \top_ihp.wb_coproc.dat_o[2] ;
 wire \top_ihp.wb_coproc.dat_o[30] ;
 wire \top_ihp.wb_coproc.dat_o[31] ;
 wire \top_ihp.wb_coproc.dat_o[3] ;
 wire \top_ihp.wb_coproc.dat_o[4] ;
 wire \top_ihp.wb_coproc.dat_o[5] ;
 wire \top_ihp.wb_coproc.dat_o[6] ;
 wire \top_ihp.wb_coproc.dat_o[7] ;
 wire \top_ihp.wb_coproc.dat_o[8] ;
 wire \top_ihp.wb_coproc.dat_o[9] ;
 wire \top_ihp.wb_coproc.opa[0] ;
 wire \top_ihp.wb_coproc.opa[10] ;
 wire \top_ihp.wb_coproc.opa[11] ;
 wire \top_ihp.wb_coproc.opa[12] ;
 wire \top_ihp.wb_coproc.opa[13] ;
 wire \top_ihp.wb_coproc.opa[14] ;
 wire \top_ihp.wb_coproc.opa[15] ;
 wire \top_ihp.wb_coproc.opa[16] ;
 wire \top_ihp.wb_coproc.opa[17] ;
 wire \top_ihp.wb_coproc.opa[18] ;
 wire \top_ihp.wb_coproc.opa[19] ;
 wire \top_ihp.wb_coproc.opa[1] ;
 wire \top_ihp.wb_coproc.opa[20] ;
 wire \top_ihp.wb_coproc.opa[21] ;
 wire \top_ihp.wb_coproc.opa[22] ;
 wire \top_ihp.wb_coproc.opa[23] ;
 wire \top_ihp.wb_coproc.opa[24] ;
 wire \top_ihp.wb_coproc.opa[25] ;
 wire \top_ihp.wb_coproc.opa[26] ;
 wire \top_ihp.wb_coproc.opa[27] ;
 wire \top_ihp.wb_coproc.opa[28] ;
 wire \top_ihp.wb_coproc.opa[29] ;
 wire \top_ihp.wb_coproc.opa[2] ;
 wire \top_ihp.wb_coproc.opa[30] ;
 wire \top_ihp.wb_coproc.opa[31] ;
 wire \top_ihp.wb_coproc.opa[3] ;
 wire \top_ihp.wb_coproc.opa[4] ;
 wire \top_ihp.wb_coproc.opa[5] ;
 wire \top_ihp.wb_coproc.opa[6] ;
 wire \top_ihp.wb_coproc.opa[7] ;
 wire \top_ihp.wb_coproc.opa[8] ;
 wire \top_ihp.wb_coproc.opa[9] ;
 wire \top_ihp.wb_coproc.opb[0] ;
 wire \top_ihp.wb_coproc.opb[10] ;
 wire \top_ihp.wb_coproc.opb[11] ;
 wire \top_ihp.wb_coproc.opb[12] ;
 wire \top_ihp.wb_coproc.opb[13] ;
 wire \top_ihp.wb_coproc.opb[14] ;
 wire \top_ihp.wb_coproc.opb[15] ;
 wire \top_ihp.wb_coproc.opb[16] ;
 wire \top_ihp.wb_coproc.opb[17] ;
 wire \top_ihp.wb_coproc.opb[18] ;
 wire \top_ihp.wb_coproc.opb[19] ;
 wire \top_ihp.wb_coproc.opb[1] ;
 wire \top_ihp.wb_coproc.opb[20] ;
 wire \top_ihp.wb_coproc.opb[21] ;
 wire \top_ihp.wb_coproc.opb[22] ;
 wire \top_ihp.wb_coproc.opb[23] ;
 wire \top_ihp.wb_coproc.opb[24] ;
 wire \top_ihp.wb_coproc.opb[25] ;
 wire \top_ihp.wb_coproc.opb[26] ;
 wire \top_ihp.wb_coproc.opb[27] ;
 wire \top_ihp.wb_coproc.opb[28] ;
 wire \top_ihp.wb_coproc.opb[29] ;
 wire \top_ihp.wb_coproc.opb[2] ;
 wire \top_ihp.wb_coproc.opb[30] ;
 wire \top_ihp.wb_coproc.opb[31] ;
 wire \top_ihp.wb_coproc.opb[3] ;
 wire \top_ihp.wb_coproc.opb[4] ;
 wire \top_ihp.wb_coproc.opb[5] ;
 wire \top_ihp.wb_coproc.opb[6] ;
 wire \top_ihp.wb_coproc.opb[7] ;
 wire \top_ihp.wb_coproc.opb[8] ;
 wire \top_ihp.wb_coproc.opb[9] ;
 wire \top_ihp.wb_dati_gpio[0] ;
 wire \top_ihp.wb_dati_ram[0] ;
 wire \top_ihp.wb_dati_ram[10] ;
 wire \top_ihp.wb_dati_ram[11] ;
 wire \top_ihp.wb_dati_ram[12] ;
 wire \top_ihp.wb_dati_ram[13] ;
 wire \top_ihp.wb_dati_ram[14] ;
 wire \top_ihp.wb_dati_ram[15] ;
 wire \top_ihp.wb_dati_ram[16] ;
 wire \top_ihp.wb_dati_ram[17] ;
 wire \top_ihp.wb_dati_ram[18] ;
 wire \top_ihp.wb_dati_ram[19] ;
 wire \top_ihp.wb_dati_ram[1] ;
 wire \top_ihp.wb_dati_ram[20] ;
 wire \top_ihp.wb_dati_ram[21] ;
 wire \top_ihp.wb_dati_ram[22] ;
 wire \top_ihp.wb_dati_ram[23] ;
 wire \top_ihp.wb_dati_ram[24] ;
 wire \top_ihp.wb_dati_ram[25] ;
 wire \top_ihp.wb_dati_ram[26] ;
 wire \top_ihp.wb_dati_ram[27] ;
 wire \top_ihp.wb_dati_ram[28] ;
 wire \top_ihp.wb_dati_ram[29] ;
 wire \top_ihp.wb_dati_ram[2] ;
 wire \top_ihp.wb_dati_ram[30] ;
 wire \top_ihp.wb_dati_ram[31] ;
 wire \top_ihp.wb_dati_ram[3] ;
 wire \top_ihp.wb_dati_ram[4] ;
 wire \top_ihp.wb_dati_ram[5] ;
 wire \top_ihp.wb_dati_ram[6] ;
 wire \top_ihp.wb_dati_ram[7] ;
 wire \top_ihp.wb_dati_ram[8] ;
 wire \top_ihp.wb_dati_ram[9] ;
 wire \top_ihp.wb_dati_rom[0] ;
 wire \top_ihp.wb_dati_rom[10] ;
 wire \top_ihp.wb_dati_rom[11] ;
 wire \top_ihp.wb_dati_rom[12] ;
 wire \top_ihp.wb_dati_rom[13] ;
 wire \top_ihp.wb_dati_rom[14] ;
 wire \top_ihp.wb_dati_rom[15] ;
 wire \top_ihp.wb_dati_rom[16] ;
 wire \top_ihp.wb_dati_rom[17] ;
 wire \top_ihp.wb_dati_rom[18] ;
 wire \top_ihp.wb_dati_rom[19] ;
 wire \top_ihp.wb_dati_rom[1] ;
 wire \top_ihp.wb_dati_rom[20] ;
 wire \top_ihp.wb_dati_rom[21] ;
 wire \top_ihp.wb_dati_rom[22] ;
 wire \top_ihp.wb_dati_rom[23] ;
 wire \top_ihp.wb_dati_rom[24] ;
 wire \top_ihp.wb_dati_rom[25] ;
 wire \top_ihp.wb_dati_rom[26] ;
 wire \top_ihp.wb_dati_rom[27] ;
 wire \top_ihp.wb_dati_rom[28] ;
 wire \top_ihp.wb_dati_rom[29] ;
 wire \top_ihp.wb_dati_rom[2] ;
 wire \top_ihp.wb_dati_rom[30] ;
 wire \top_ihp.wb_dati_rom[31] ;
 wire \top_ihp.wb_dati_rom[3] ;
 wire \top_ihp.wb_dati_rom[4] ;
 wire \top_ihp.wb_dati_rom[5] ;
 wire \top_ihp.wb_dati_rom[6] ;
 wire \top_ihp.wb_dati_rom[7] ;
 wire \top_ihp.wb_dati_rom[8] ;
 wire \top_ihp.wb_dati_rom[9] ;
 wire \top_ihp.wb_dati_spi[0] ;
 wire \top_ihp.wb_dati_spi[10] ;
 wire \top_ihp.wb_dati_spi[11] ;
 wire \top_ihp.wb_dati_spi[12] ;
 wire \top_ihp.wb_dati_spi[13] ;
 wire \top_ihp.wb_dati_spi[14] ;
 wire \top_ihp.wb_dati_spi[15] ;
 wire \top_ihp.wb_dati_spi[16] ;
 wire \top_ihp.wb_dati_spi[17] ;
 wire \top_ihp.wb_dati_spi[18] ;
 wire \top_ihp.wb_dati_spi[19] ;
 wire \top_ihp.wb_dati_spi[1] ;
 wire \top_ihp.wb_dati_spi[20] ;
 wire \top_ihp.wb_dati_spi[21] ;
 wire \top_ihp.wb_dati_spi[22] ;
 wire \top_ihp.wb_dati_spi[23] ;
 wire \top_ihp.wb_dati_spi[24] ;
 wire \top_ihp.wb_dati_spi[25] ;
 wire \top_ihp.wb_dati_spi[26] ;
 wire \top_ihp.wb_dati_spi[27] ;
 wire \top_ihp.wb_dati_spi[28] ;
 wire \top_ihp.wb_dati_spi[29] ;
 wire \top_ihp.wb_dati_spi[2] ;
 wire \top_ihp.wb_dati_spi[30] ;
 wire \top_ihp.wb_dati_spi[31] ;
 wire \top_ihp.wb_dati_spi[3] ;
 wire \top_ihp.wb_dati_spi[4] ;
 wire \top_ihp.wb_dati_spi[5] ;
 wire \top_ihp.wb_dati_spi[6] ;
 wire \top_ihp.wb_dati_spi[7] ;
 wire \top_ihp.wb_dati_spi[8] ;
 wire \top_ihp.wb_dati_spi[9] ;
 wire \top_ihp.wb_dati_uart[0] ;
 wire \top_ihp.wb_dati_uart[1] ;
 wire \top_ihp.wb_dati_uart[2] ;
 wire \top_ihp.wb_dati_uart[3] ;
 wire \top_ihp.wb_dati_uart[4] ;
 wire \top_ihp.wb_dati_uart[5] ;
 wire \top_ihp.wb_dati_uart[6] ;
 wire \top_ihp.wb_dati_uart[7] ;
 wire \top_ihp.wb_emem.bit_counter[0] ;
 wire \top_ihp.wb_emem.bit_counter[1] ;
 wire \top_ihp.wb_emem.bit_counter[2] ;
 wire \top_ihp.wb_emem.bit_counter[3] ;
 wire \top_ihp.wb_emem.bit_counter[4] ;
 wire \top_ihp.wb_emem.bit_counter[5] ;
 wire \top_ihp.wb_emem.bit_counter[6] ;
 wire \top_ihp.wb_emem.bit_counter[7] ;
 wire \top_ihp.wb_emem.cmd[32] ;
 wire \top_ihp.wb_emem.cmd[33] ;
 wire \top_ihp.wb_emem.cmd[34] ;
 wire \top_ihp.wb_emem.cmd[35] ;
 wire \top_ihp.wb_emem.cmd[36] ;
 wire \top_ihp.wb_emem.cmd[37] ;
 wire \top_ihp.wb_emem.cmd[38] ;
 wire \top_ihp.wb_emem.cmd[39] ;
 wire \top_ihp.wb_emem.cmd[40] ;
 wire \top_ihp.wb_emem.cmd[41] ;
 wire \top_ihp.wb_emem.cmd[42] ;
 wire \top_ihp.wb_emem.cmd[43] ;
 wire \top_ihp.wb_emem.cmd[44] ;
 wire \top_ihp.wb_emem.cmd[45] ;
 wire \top_ihp.wb_emem.cmd[46] ;
 wire \top_ihp.wb_emem.cmd[47] ;
 wire \top_ihp.wb_emem.cmd[48] ;
 wire \top_ihp.wb_emem.cmd[49] ;
 wire \top_ihp.wb_emem.cmd[50] ;
 wire \top_ihp.wb_emem.cmd[51] ;
 wire \top_ihp.wb_emem.cmd[52] ;
 wire \top_ihp.wb_emem.cmd[53] ;
 wire \top_ihp.wb_emem.cmd[54] ;
 wire \top_ihp.wb_emem.cmd[55] ;
 wire \top_ihp.wb_emem.cmd[56] ;
 wire \top_ihp.wb_emem.cmd[57] ;
 wire \top_ihp.wb_emem.cmd[58] ;
 wire \top_ihp.wb_emem.cmd[59] ;
 wire \top_ihp.wb_emem.cmd[60] ;
 wire \top_ihp.wb_emem.cmd[61] ;
 wire \top_ihp.wb_emem.cmd[62] ;
 wire \top_ihp.wb_emem.cmd[63] ;
 wire \top_ihp.wb_emem.last_bit ;
 wire \top_ihp.wb_emem.last_wait ;
 wire \top_ihp.wb_emem.nbits[3] ;
 wire \top_ihp.wb_emem.nbits[4] ;
 wire \top_ihp.wb_emem.nbits[5] ;
 wire \top_ihp.wb_emem.nbits[6] ;
 wire \top_ihp.wb_emem.state[0] ;
 wire \top_ihp.wb_emem.state[1] ;
 wire \top_ihp.wb_emem.state[2] ;
 wire \top_ihp.wb_emem.state[3] ;
 wire \top_ihp.wb_emem.wait_counter[0] ;
 wire \top_ihp.wb_emem.wait_counter[1] ;
 wire \top_ihp.wb_emem.wait_counter[2] ;
 wire \top_ihp.wb_emem.wait_counter[3] ;
 wire \top_ihp.wb_emem.wait_counter[4] ;
 wire \top_ihp.wb_emem.wait_counter[5] ;
 wire \top_ihp.wb_emem.wait_counter[6] ;
 wire \top_ihp.wb_emem.wait_counter[7] ;
 wire \top_ihp.wb_imem.bits_left[0] ;
 wire \top_ihp.wb_imem.bits_left[1] ;
 wire \top_ihp.wb_imem.bits_left[2] ;
 wire \top_ihp.wb_imem.bits_left[3] ;
 wire \top_ihp.wb_imem.bits_left[4] ;
 wire \top_ihp.wb_imem.bits_left[5] ;
 wire \top_ihp.wb_imem.state[0] ;
 wire \top_ihp.wb_imem.state[1] ;
 wire \top_ihp.wb_imem.state[2] ;
 wire \top_ihp.wb_spi.bits_left[0] ;
 wire \top_ihp.wb_spi.bits_left[1] ;
 wire \top_ihp.wb_spi.bits_left[2] ;
 wire \top_ihp.wb_spi.bits_left[3] ;
 wire \top_ihp.wb_spi.bits_left[4] ;
 wire \top_ihp.wb_spi.bits_left[5] ;
 wire \top_ihp.wb_spi.spi_clk_cnt[0] ;
 wire \top_ihp.wb_spi.state ;
 wire \top_ihp.wb_uart.rx_ready ;
 wire \top_ihp.wb_uart.state[0] ;
 wire \top_ihp.wb_uart.state[1] ;
 wire \top_ihp.wb_uart.tx_ready ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_rx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_rx.next_state[2] ;
 wire \top_ihp.wb_uart.uart_rx.state[0] ;
 wire \top_ihp.wb_uart.uart_rx.state[1] ;
 wire \top_ihp.wb_uart.uart_rx.state[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.bit_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[0] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[10] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[11] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[12] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[13] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[14] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[15] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[16] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[17] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[18] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[19] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[1] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[20] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[21] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[22] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[23] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[24] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[25] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[26] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[27] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[28] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[29] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[2] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[30] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[31] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[3] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[4] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[5] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[6] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[7] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[8] ;
 wire \top_ihp.wb_uart.uart_tx.cycle_cnt[9] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[0] ;
 wire \top_ihp.wb_uart.uart_tx.next_state[1] ;
 wire \top_ihp.wb_uart.uart_tx.state[0] ;
 wire \top_ihp.wb_uart.uart_tx.state[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[0] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[1] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[2] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[3] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[4] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[5] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[6] ;
 wire \top_ihp.wb_uart.uart_tx.tx_data_latch[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_252_clk;
 wire clknet_leaf_253_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_leaf_303_clk;
 wire clknet_leaf_304_clk;
 wire clknet_leaf_305_clk;
 wire clknet_leaf_306_clk;
 wire clknet_leaf_307_clk;
 wire clknet_leaf_308_clk;
 wire clknet_leaf_309_clk;
 wire clknet_leaf_310_clk;
 wire clknet_leaf_311_clk;
 wire clknet_leaf_312_clk;
 wire clknet_leaf_313_clk;
 wire clknet_leaf_314_clk;
 wire clknet_leaf_315_clk;
 wire clknet_leaf_316_clk;
 wire clknet_leaf_317_clk;
 wire clknet_leaf_318_clk;
 wire clknet_leaf_319_clk;
 wire clknet_leaf_320_clk;
 wire clknet_leaf_321_clk;
 wire clknet_leaf_322_clk;
 wire clknet_leaf_323_clk;
 wire clknet_leaf_324_clk;
 wire clknet_leaf_325_clk;
 wire clknet_leaf_326_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire clknet_6_0__leaf_clk;
 wire clknet_6_1__leaf_clk;
 wire clknet_6_2__leaf_clk;
 wire clknet_6_3__leaf_clk;
 wire clknet_6_4__leaf_clk;
 wire clknet_6_5__leaf_clk;
 wire clknet_6_6__leaf_clk;
 wire clknet_6_7__leaf_clk;
 wire clknet_6_8__leaf_clk;
 wire clknet_6_9__leaf_clk;
 wire clknet_6_10__leaf_clk;
 wire clknet_6_11__leaf_clk;
 wire clknet_6_12__leaf_clk;
 wire clknet_6_13__leaf_clk;
 wire clknet_6_14__leaf_clk;
 wire clknet_6_15__leaf_clk;
 wire clknet_6_16__leaf_clk;
 wire clknet_6_17__leaf_clk;
 wire clknet_6_18__leaf_clk;
 wire clknet_6_19__leaf_clk;
 wire clknet_6_20__leaf_clk;
 wire clknet_6_21__leaf_clk;
 wire clknet_6_22__leaf_clk;
 wire clknet_6_23__leaf_clk;
 wire clknet_6_24__leaf_clk;
 wire clknet_6_25__leaf_clk;
 wire clknet_6_26__leaf_clk;
 wire clknet_6_27__leaf_clk;
 wire clknet_6_28__leaf_clk;
 wire clknet_6_29__leaf_clk;
 wire clknet_6_30__leaf_clk;
 wire clknet_6_31__leaf_clk;
 wire clknet_6_32__leaf_clk;
 wire clknet_6_33__leaf_clk;
 wire clknet_6_34__leaf_clk;
 wire clknet_6_35__leaf_clk;
 wire clknet_6_36__leaf_clk;
 wire clknet_6_37__leaf_clk;
 wire clknet_6_38__leaf_clk;
 wire clknet_6_39__leaf_clk;
 wire clknet_6_40__leaf_clk;
 wire clknet_6_41__leaf_clk;
 wire clknet_6_42__leaf_clk;
 wire clknet_6_43__leaf_clk;
 wire clknet_6_44__leaf_clk;
 wire clknet_6_45__leaf_clk;
 wire clknet_6_46__leaf_clk;
 wire clknet_6_47__leaf_clk;
 wire clknet_6_48__leaf_clk;
 wire clknet_6_49__leaf_clk;
 wire clknet_6_50__leaf_clk;
 wire clknet_6_51__leaf_clk;
 wire clknet_6_52__leaf_clk;
 wire clknet_6_53__leaf_clk;
 wire clknet_6_54__leaf_clk;
 wire clknet_6_55__leaf_clk;
 wire clknet_6_56__leaf_clk;
 wire clknet_6_57__leaf_clk;
 wire clknet_6_58__leaf_clk;
 wire clknet_6_59__leaf_clk;
 wire clknet_6_60__leaf_clk;
 wire clknet_6_61__leaf_clk;
 wire clknet_6_62__leaf_clk;
 wire clknet_6_63__leaf_clk;

 sg13g2_buf_2 _13705_ (.A(\top_ihp.oisc.state[5] ),
    .X(_08199_));
 sg13g2_buf_1 _13706_ (.A(_08199_),
    .X(_08200_));
 sg13g2_buf_2 _13707_ (.A(\top_ihp.oisc.decoder.decoded[10] ),
    .X(_08201_));
 sg13g2_buf_1 _13708_ (.A(\top_ihp.oisc.micro_op[1] ),
    .X(_08202_));
 sg13g2_buf_1 _13709_ (.A(\top_ihp.oisc.micro_op[0] ),
    .X(_08203_));
 sg13g2_buf_1 _13710_ (.A(\top_ihp.oisc.micro_op[3] ),
    .X(_08204_));
 sg13g2_buf_2 _13711_ (.A(\top_ihp.oisc.micro_op[2] ),
    .X(_08205_));
 sg13g2_buf_2 _13712_ (.A(\top_ihp.oisc.micro_op[4] ),
    .X(_08206_));
 sg13g2_buf_2 _13713_ (.A(\top_ihp.oisc.micro_op[5] ),
    .X(_08207_));
 sg13g2_and4_1 _13714_ (.A(_08205_),
    .B(_08206_),
    .C(_08207_),
    .D(\top_ihp.oisc.micro_state[2] ),
    .X(_08208_));
 sg13g2_and4_1 _13715_ (.A(_08202_),
    .B(_08203_),
    .C(_08204_),
    .D(_08208_),
    .X(_08209_));
 sg13g2_buf_2 _13716_ (.A(_08209_),
    .X(_08210_));
 sg13g2_buf_8 _13717_ (.A(_08210_),
    .X(_08211_));
 sg13g2_nand3_1 _13718_ (.B(_08201_),
    .C(net892),
    .A(net1032),
    .Y(_08212_));
 sg13g2_buf_2 _13719_ (.A(_08212_),
    .X(_08213_));
 sg13g2_buf_2 _13720_ (.A(\top_ihp.wb_spi.state ),
    .X(_08214_));
 sg13g2_inv_1 _13721_ (.Y(_08215_),
    .A(_08214_));
 sg13g2_buf_1 _13722_ (.A(\top_ihp.oisc.op_a[26] ),
    .X(_08216_));
 sg13g2_buf_1 _13723_ (.A(_08216_),
    .X(_08217_));
 sg13g2_inv_1 _13724_ (.Y(_08218_),
    .A(\top_ihp.oisc.op_b[26] ));
 sg13g2_buf_2 _13725_ (.A(\top_ihp.oisc.op_b[19] ),
    .X(_08219_));
 sg13g2_buf_2 _13726_ (.A(\top_ihp.oisc.op_b[18] ),
    .X(_08220_));
 sg13g2_buf_2 _13727_ (.A(\top_ihp.oisc.op_a[18] ),
    .X(_08221_));
 sg13g2_nand2b_1 _13728_ (.Y(_08222_),
    .B(net1059),
    .A_N(_08220_));
 sg13g2_buf_2 _13729_ (.A(\top_ihp.oisc.op_a[19] ),
    .X(_08223_));
 sg13g2_inv_1 _13730_ (.Y(_08224_),
    .A(net1058));
 sg13g2_o21ai_1 _13731_ (.B1(_08224_),
    .Y(_08225_),
    .A1(_08219_),
    .A2(_08222_));
 sg13g2_nand2_1 _13732_ (.Y(_08226_),
    .A(_08219_),
    .B(_08222_));
 sg13g2_buf_1 _13733_ (.A(\top_ihp.oisc.op_b[20] ),
    .X(_08227_));
 sg13g2_buf_2 _13734_ (.A(\top_ihp.oisc.op_a[20] ),
    .X(_08228_));
 sg13g2_nor2b_1 _13735_ (.A(net1057),
    .B_N(net1056),
    .Y(_08229_));
 sg13g2_a21oi_1 _13736_ (.A1(_08225_),
    .A2(_08226_),
    .Y(_08230_),
    .B1(_08229_));
 sg13g2_buf_2 _13737_ (.A(\top_ihp.oisc.op_b[21] ),
    .X(_08231_));
 sg13g2_nor2b_1 _13738_ (.A(\top_ihp.oisc.op_a[20] ),
    .B_N(net1057),
    .Y(_08232_));
 sg13g2_buf_1 _13739_ (.A(_08232_),
    .X(_08233_));
 sg13g2_or2_1 _13740_ (.X(_08234_),
    .B(_08233_),
    .A(_08231_));
 sg13g2_buf_8 _13741_ (.A(\top_ihp.oisc.op_a[21] ),
    .X(_08235_));
 sg13g2_inv_1 _13742_ (.Y(_08236_),
    .A(_08235_));
 sg13g2_o21ai_1 _13743_ (.B1(_08236_),
    .Y(_08237_),
    .A1(_08230_),
    .A2(_08234_));
 sg13g2_o21ai_1 _13744_ (.B1(_08231_),
    .Y(_08238_),
    .A1(_08230_),
    .A2(_08233_));
 sg13g2_nand2_1 _13745_ (.Y(_08239_),
    .A(_08237_),
    .B(_08238_));
 sg13g2_nand2b_1 _13746_ (.Y(_08240_),
    .B(_08231_),
    .A_N(_08235_));
 sg13g2_buf_1 _13747_ (.A(_08240_),
    .X(_08241_));
 sg13g2_nand3b_1 _13748_ (.B(_08220_),
    .C(_08219_),
    .Y(_08242_),
    .A_N(net1059));
 sg13g2_nand3b_1 _13749_ (.B(_08241_),
    .C(_08242_),
    .Y(_08243_),
    .A_N(net1057));
 sg13g2_nand3_1 _13750_ (.B(_08241_),
    .C(_08242_),
    .A(net1056),
    .Y(_08244_));
 sg13g2_inv_1 _13751_ (.Y(_08245_),
    .A(_08219_));
 sg13g2_nand2b_1 _13752_ (.Y(_08246_),
    .B(_08220_),
    .A_N(net1059));
 sg13g2_a21oi_1 _13753_ (.A1(_08245_),
    .A2(_08246_),
    .Y(_08247_),
    .B1(\top_ihp.oisc.op_a[19] ));
 sg13g2_a21o_1 _13754_ (.A2(_08244_),
    .A1(_08243_),
    .B1(_08247_),
    .X(_08248_));
 sg13g2_nor2_1 _13755_ (.A(_08236_),
    .B(_08231_),
    .Y(_08249_));
 sg13g2_a21oi_1 _13756_ (.A1(_08241_),
    .A2(_08229_),
    .Y(_08250_),
    .B1(_08249_));
 sg13g2_buf_2 _13757_ (.A(\top_ihp.oisc.op_b[13] ),
    .X(_08251_));
 sg13g2_buf_2 _13758_ (.A(\top_ihp.oisc.op_a[12] ),
    .X(_08252_));
 sg13g2_buf_2 _13759_ (.A(\top_ihp.oisc.op_b[12] ),
    .X(_08253_));
 sg13g2_nor2b_1 _13760_ (.A(_08252_),
    .B_N(_08253_),
    .Y(_08254_));
 sg13g2_or2_1 _13761_ (.X(_08255_),
    .B(_08254_),
    .A(_08251_));
 sg13g2_buf_2 _13762_ (.A(\top_ihp.oisc.op_a[13] ),
    .X(_08256_));
 sg13g2_nand2_1 _13763_ (.Y(_08257_),
    .A(_08251_),
    .B(_08254_));
 sg13g2_nand2_1 _13764_ (.Y(_08258_),
    .A(net1055),
    .B(_08257_));
 sg13g2_buf_1 _13765_ (.A(\top_ihp.oisc.op_a[11] ),
    .X(_08259_));
 sg13g2_buf_2 _13766_ (.A(_08259_),
    .X(_08260_));
 sg13g2_buf_1 _13767_ (.A(\top_ihp.oisc.op_b[11] ),
    .X(_08261_));
 sg13g2_buf_1 _13768_ (.A(\top_ihp.oisc.op_a[10] ),
    .X(_08262_));
 sg13g2_buf_2 _13769_ (.A(\top_ihp.oisc.op_b[10] ),
    .X(_08263_));
 sg13g2_nor2b_1 _13770_ (.A(net1053),
    .B_N(_08263_),
    .Y(_08264_));
 sg13g2_nand2_1 _13771_ (.Y(_08265_),
    .A(net1054),
    .B(_08264_));
 sg13g2_nand2b_1 _13772_ (.Y(_08266_),
    .B(_08252_),
    .A_N(_08253_));
 sg13g2_nand2_1 _13773_ (.Y(_08267_),
    .A(_08251_),
    .B(_08266_));
 sg13g2_nand2b_1 _13774_ (.Y(_08268_),
    .B(_08266_),
    .A_N(net1055));
 sg13g2_nor2_1 _13775_ (.A(net1054),
    .B(_08264_),
    .Y(_08269_));
 sg13g2_a221oi_1 _13776_ (.B2(_08268_),
    .C1(_08269_),
    .B1(_08267_),
    .A1(net1030),
    .Y(_08270_),
    .A2(_08265_));
 sg13g2_a221oi_1 _13777_ (.B2(_08258_),
    .C1(_08270_),
    .B1(_08255_),
    .A1(_08248_),
    .Y(_08271_),
    .A2(_08250_));
 sg13g2_buf_2 _13778_ (.A(\top_ihp.oisc.op_b[16] ),
    .X(_08272_));
 sg13g2_inv_1 _13779_ (.Y(_08273_),
    .A(_08272_));
 sg13g2_buf_1 _13780_ (.A(\top_ihp.oisc.op_a[17] ),
    .X(_08274_));
 sg13g2_buf_2 _13781_ (.A(\top_ihp.oisc.op_b[17] ),
    .X(_08275_));
 sg13g2_nand2b_1 _13782_ (.Y(_08276_),
    .B(_08275_),
    .A_N(net1052));
 sg13g2_buf_2 _13783_ (.A(_08276_),
    .X(_08277_));
 sg13g2_buf_2 _13784_ (.A(\top_ihp.oisc.op_b[14] ),
    .X(_08278_));
 sg13g2_buf_2 _13785_ (.A(\top_ihp.oisc.op_b[15] ),
    .X(_08279_));
 sg13g2_nand3b_1 _13786_ (.B(_08278_),
    .C(_08279_),
    .Y(_08280_),
    .A_N(\top_ihp.oisc.op_a[14] ));
 sg13g2_nand3_1 _13787_ (.B(_08277_),
    .C(_08280_),
    .A(_08273_),
    .Y(_08281_));
 sg13g2_buf_2 _13788_ (.A(\top_ihp.oisc.op_a[16] ),
    .X(_08282_));
 sg13g2_nand3_1 _13789_ (.B(_08277_),
    .C(_08280_),
    .A(_08282_),
    .Y(_08283_));
 sg13g2_inv_1 _13790_ (.Y(_08284_),
    .A(_08279_));
 sg13g2_buf_2 _13791_ (.A(\top_ihp.oisc.op_a[14] ),
    .X(_08285_));
 sg13g2_nand2b_1 _13792_ (.Y(_08286_),
    .B(_08278_),
    .A_N(net1051));
 sg13g2_buf_4 _13793_ (.X(_08287_),
    .A(\top_ihp.oisc.op_a[15] ));
 sg13g2_a21oi_1 _13794_ (.A1(_08284_),
    .A2(_08286_),
    .Y(_08288_),
    .B1(_08287_));
 sg13g2_a21o_1 _13795_ (.A2(_08283_),
    .A1(_08281_),
    .B1(_08288_),
    .X(_08289_));
 sg13g2_buf_1 _13796_ (.A(_08289_),
    .X(_08290_));
 sg13g2_inv_1 _13797_ (.Y(_08291_),
    .A(_08282_));
 sg13g2_nor2_1 _13798_ (.A(_08291_),
    .B(_08272_),
    .Y(_08292_));
 sg13g2_nor2b_1 _13799_ (.A(_08275_),
    .B_N(net1052),
    .Y(_08293_));
 sg13g2_a21oi_2 _13800_ (.B1(_08293_),
    .Y(_08294_),
    .A2(_08292_),
    .A1(_08277_));
 sg13g2_xor2_1 _13801_ (.B(_08251_),
    .A(_08256_),
    .X(_08295_));
 sg13g2_xor2_1 _13802_ (.B(_08253_),
    .A(_08252_),
    .X(_08296_));
 sg13g2_nor2b_1 _13803_ (.A(_08259_),
    .B_N(net1054),
    .Y(_08297_));
 sg13g2_buf_1 _13804_ (.A(_08297_),
    .X(_08298_));
 sg13g2_nor2b_1 _13805_ (.A(net1054),
    .B_N(_08259_),
    .Y(_08299_));
 sg13g2_nor4_2 _13806_ (.A(_08295_),
    .B(_08296_),
    .C(_08298_),
    .Y(_08300_),
    .D(_08299_));
 sg13g2_xnor2_1 _13807_ (.Y(_08301_),
    .A(net1053),
    .B(_08263_));
 sg13g2_and2_1 _13808_ (.A(_08300_),
    .B(_08301_),
    .X(_08302_));
 sg13g2_a21oi_1 _13809_ (.A1(_08290_),
    .A2(_08294_),
    .Y(_08303_),
    .B1(_08302_));
 sg13g2_xor2_1 _13810_ (.B(_08279_),
    .A(_08287_),
    .X(_08304_));
 sg13g2_xnor2_1 _13811_ (.Y(_08305_),
    .A(net1051),
    .B(_08278_));
 sg13g2_nor2b_1 _13812_ (.A(_08304_),
    .B_N(_08305_),
    .Y(_08306_));
 sg13g2_xor2_1 _13813_ (.B(_08272_),
    .A(_08282_),
    .X(_08307_));
 sg13g2_xor2_1 _13814_ (.B(_08275_),
    .A(net1052),
    .X(_08308_));
 sg13g2_nor2_1 _13815_ (.A(_08307_),
    .B(_08308_),
    .Y(_08309_));
 sg13g2_and2_1 _13816_ (.A(_08306_),
    .B(_08309_),
    .X(_08310_));
 sg13g2_a221oi_1 _13817_ (.B2(_08250_),
    .C1(_08310_),
    .B1(_08248_),
    .A1(_08290_),
    .Y(_08311_),
    .A2(_08294_));
 sg13g2_a21oi_1 _13818_ (.A1(_08271_),
    .A2(_08303_),
    .Y(_08312_),
    .B1(_08311_));
 sg13g2_nand2_1 _13819_ (.Y(_08313_),
    .A(_08290_),
    .B(_08294_));
 sg13g2_buf_8 _13820_ (.A(\top_ihp.oisc.op_a[7] ),
    .X(_08314_));
 sg13g2_buf_2 _13821_ (.A(\top_ihp.oisc.op_b[7] ),
    .X(_08315_));
 sg13g2_nor2b_1 _13822_ (.A(_08314_),
    .B_N(_08315_),
    .Y(_08316_));
 sg13g2_buf_8 _13823_ (.A(\top_ihp.oisc.op_a[1] ),
    .X(_08317_));
 sg13g2_inv_1 _13824_ (.Y(_08318_),
    .A(_08317_));
 sg13g2_buf_2 _13825_ (.A(\top_ihp.oisc.op_b[1] ),
    .X(_08319_));
 sg13g2_buf_2 _13826_ (.A(\top_ihp.oisc.op_b[0] ),
    .X(_08320_));
 sg13g2_buf_2 _13827_ (.A(\top_ihp.oisc.op_a[0] ),
    .X(_08321_));
 sg13g2_nand2b_1 _13828_ (.Y(_08322_),
    .B(_08321_),
    .A_N(_08320_));
 sg13g2_buf_2 _13829_ (.A(_08322_),
    .X(_08323_));
 sg13g2_o21ai_1 _13830_ (.B1(_08323_),
    .Y(_08324_),
    .A1(_08318_),
    .A2(_08319_));
 sg13g2_buf_1 _13831_ (.A(_08324_),
    .X(_08325_));
 sg13g2_buf_2 _13832_ (.A(\top_ihp.oisc.op_a[3] ),
    .X(_08326_));
 sg13g2_inv_1 _13833_ (.Y(_08327_),
    .A(_08326_));
 sg13g2_buf_2 _13834_ (.A(\top_ihp.oisc.op_b[3] ),
    .X(_08328_));
 sg13g2_buf_8 _13835_ (.A(\top_ihp.oisc.op_a[2] ),
    .X(_08329_));
 sg13g2_buf_2 _13836_ (.A(\top_ihp.oisc.op_b[2] ),
    .X(_08330_));
 sg13g2_nor2b_1 _13837_ (.A(net1050),
    .B_N(_08330_),
    .Y(_08331_));
 sg13g2_a221oi_1 _13838_ (.B2(_08319_),
    .C1(_08331_),
    .B1(_08318_),
    .A1(_08327_),
    .Y(_08332_),
    .A2(_08328_));
 sg13g2_buf_1 _13839_ (.A(_08332_),
    .X(_08333_));
 sg13g2_nand2b_1 _13840_ (.Y(_08334_),
    .B(net1050),
    .A_N(_08330_));
 sg13g2_nand2_1 _13841_ (.Y(_08335_),
    .A(_08328_),
    .B(_08334_));
 sg13g2_o21ai_1 _13842_ (.B1(_08327_),
    .Y(_08336_),
    .A1(_08328_),
    .A2(_08334_));
 sg13g2_buf_1 _13843_ (.A(_08336_),
    .X(_08337_));
 sg13g2_buf_2 _13844_ (.A(\top_ihp.oisc.op_a[4] ),
    .X(_08338_));
 sg13g2_buf_2 _13845_ (.A(\top_ihp.oisc.op_b[4] ),
    .X(_08339_));
 sg13g2_xnor2_1 _13846_ (.Y(_08340_),
    .A(net1049),
    .B(_08339_));
 sg13g2_buf_2 _13847_ (.A(\top_ihp.oisc.op_a[5] ),
    .X(_08341_));
 sg13g2_buf_2 _13848_ (.A(\top_ihp.oisc.op_b[5] ),
    .X(_08342_));
 sg13g2_xnor2_1 _13849_ (.Y(_08343_),
    .A(_08341_),
    .B(_08342_));
 sg13g2_xnor2_1 _13850_ (.Y(_08344_),
    .A(_08314_),
    .B(_08315_));
 sg13g2_buf_4 _13851_ (.X(_08345_),
    .A(\top_ihp.oisc.op_a[6] ));
 sg13g2_buf_1 _13852_ (.A(\top_ihp.oisc.op_b[6] ),
    .X(_08346_));
 sg13g2_xnor2_1 _13853_ (.Y(_08347_),
    .A(_08345_),
    .B(_08346_));
 sg13g2_nand4_1 _13854_ (.B(_08343_),
    .C(_08344_),
    .A(_08340_),
    .Y(_08348_),
    .D(_08347_));
 sg13g2_a221oi_1 _13855_ (.B2(_08337_),
    .C1(_08348_),
    .B1(_08335_),
    .A1(_08325_),
    .Y(_08349_),
    .A2(_08333_));
 sg13g2_buf_2 _13856_ (.A(\top_ihp.oisc.op_a[8] ),
    .X(_08350_));
 sg13g2_buf_2 _13857_ (.A(\top_ihp.oisc.op_b[8] ),
    .X(_08351_));
 sg13g2_xnor2_1 _13858_ (.Y(_08352_),
    .A(_08350_),
    .B(_08351_));
 sg13g2_buf_2 _13859_ (.A(\top_ihp.oisc.op_a[9] ),
    .X(_08353_));
 sg13g2_buf_2 _13860_ (.A(\top_ihp.oisc.op_b[9] ),
    .X(_08354_));
 sg13g2_xnor2_1 _13861_ (.Y(_08355_),
    .A(_08353_),
    .B(_08354_));
 sg13g2_nand2_1 _13862_ (.Y(_08356_),
    .A(_08352_),
    .B(_08355_));
 sg13g2_inv_1 _13863_ (.Y(_08357_),
    .A(_08356_));
 sg13g2_o21ai_1 _13864_ (.B1(_08357_),
    .Y(_08358_),
    .A1(_08316_),
    .A2(_08349_));
 sg13g2_inv_1 _13865_ (.Y(_08359_),
    .A(_08351_));
 sg13g2_nor2_1 _13866_ (.A(_08350_),
    .B(_08359_),
    .Y(_08360_));
 sg13g2_nor2b_1 _13867_ (.A(net1049),
    .B_N(_08339_),
    .Y(_08361_));
 sg13g2_nor2_1 _13868_ (.A(_08342_),
    .B(_08361_),
    .Y(_08362_));
 sg13g2_inv_1 _13869_ (.Y(_08363_),
    .A(_08341_));
 sg13g2_a21oi_1 _13870_ (.A1(_08342_),
    .A2(_08361_),
    .Y(_08364_),
    .B1(_08363_));
 sg13g2_inv_1 _13871_ (.Y(_08365_),
    .A(_08345_));
 sg13g2_buf_2 _13872_ (.A(_08346_),
    .X(_08366_));
 sg13g2_nand2_1 _13873_ (.Y(_08367_),
    .A(_08365_),
    .B(net1029));
 sg13g2_o21ai_1 _13874_ (.B1(_08367_),
    .Y(_08368_),
    .A1(_08362_),
    .A2(_08364_));
 sg13g2_nand2b_1 _13875_ (.Y(_08369_),
    .B(_08314_),
    .A_N(_08315_));
 sg13g2_o21ai_1 _13876_ (.B1(_08369_),
    .Y(_08370_),
    .A1(_08365_),
    .A2(net1029));
 sg13g2_nor2_1 _13877_ (.A(_08356_),
    .B(_08370_),
    .Y(_08371_));
 sg13g2_inv_1 _13878_ (.Y(_08372_),
    .A(_08354_));
 sg13g2_nand2b_1 _13879_ (.Y(_08373_),
    .B(_08351_),
    .A_N(_08350_));
 sg13g2_a21oi_1 _13880_ (.A1(_08372_),
    .A2(_08373_),
    .Y(_08374_),
    .B1(_08353_));
 sg13g2_a221oi_1 _13881_ (.B2(_08371_),
    .C1(_08374_),
    .B1(_08368_),
    .A1(_08354_),
    .Y(_08375_),
    .A2(_08360_));
 sg13g2_nand4_1 _13882_ (.B(_08271_),
    .C(_08358_),
    .A(_08313_),
    .Y(_08376_),
    .D(_08375_));
 sg13g2_nand3_1 _13883_ (.B(_08312_),
    .C(_08376_),
    .A(_08239_),
    .Y(_08377_));
 sg13g2_buf_2 _13884_ (.A(_08377_),
    .X(_08378_));
 sg13g2_buf_2 _13885_ (.A(\top_ihp.oisc.op_b[24] ),
    .X(_08379_));
 sg13g2_buf_2 _13886_ (.A(\top_ihp.oisc.op_a[24] ),
    .X(_08380_));
 sg13g2_nand2b_1 _13887_ (.Y(_08381_),
    .B(net1048),
    .A_N(_08379_));
 sg13g2_nand2b_1 _13888_ (.Y(_08382_),
    .B(_08379_),
    .A_N(net1048));
 sg13g2_nand2_1 _13889_ (.Y(_08383_),
    .A(_08381_),
    .B(_08382_));
 sg13g2_buf_2 _13890_ (.A(\top_ihp.oisc.op_a[25] ),
    .X(_08384_));
 sg13g2_buf_1 _13891_ (.A(\top_ihp.oisc.op_b[25] ),
    .X(_08385_));
 sg13g2_nor2b_1 _13892_ (.A(_08384_),
    .B_N(_08385_),
    .Y(_08386_));
 sg13g2_buf_1 _13893_ (.A(_08386_),
    .X(_08387_));
 sg13g2_nand2b_1 _13894_ (.Y(_08388_),
    .B(_08384_),
    .A_N(_08385_));
 sg13g2_nand2b_1 _13895_ (.Y(_08389_),
    .B(_08388_),
    .A_N(_08387_));
 sg13g2_nor2_1 _13896_ (.A(_08383_),
    .B(_08389_),
    .Y(_08390_));
 sg13g2_buf_2 _13897_ (.A(\top_ihp.oisc.op_a[22] ),
    .X(_08391_));
 sg13g2_buf_2 _13898_ (.A(\top_ihp.oisc.op_b[22] ),
    .X(_08392_));
 sg13g2_xor2_1 _13899_ (.B(_08392_),
    .A(_08391_),
    .X(_08393_));
 sg13g2_buf_1 _13900_ (.A(\top_ihp.oisc.op_a[23] ),
    .X(_08394_));
 sg13g2_buf_2 _13901_ (.A(\top_ihp.oisc.op_b[23] ),
    .X(_08395_));
 sg13g2_xor2_1 _13902_ (.B(_08395_),
    .A(net1047),
    .X(_08396_));
 sg13g2_nor2_1 _13903_ (.A(_08393_),
    .B(_08396_),
    .Y(_08397_));
 sg13g2_nand2_1 _13904_ (.Y(_08398_),
    .A(_08390_),
    .B(_08397_));
 sg13g2_inv_1 _13905_ (.Y(_08399_),
    .A(_08395_));
 sg13g2_nand2b_1 _13906_ (.Y(_08400_),
    .B(_08392_),
    .A_N(_08391_));
 sg13g2_o21ai_1 _13907_ (.B1(net1047),
    .Y(_08401_),
    .A1(_08399_),
    .A2(_08400_));
 sg13g2_inv_1 _13908_ (.Y(_08402_),
    .A(_08379_));
 sg13g2_inv_1 _13909_ (.Y(_08403_),
    .A(_08385_));
 sg13g2_a221oi_1 _13910_ (.B2(_08400_),
    .C1(_08403_),
    .B1(_08399_),
    .A1(net1048),
    .Y(_08404_),
    .A2(_08402_));
 sg13g2_a21oi_1 _13911_ (.A1(_08384_),
    .A2(_08403_),
    .Y(_08405_),
    .B1(_08382_));
 sg13g2_a21oi_1 _13912_ (.A1(_08401_),
    .A2(_08404_),
    .Y(_08406_),
    .B1(_08405_));
 sg13g2_a221oi_1 _13913_ (.B2(_08400_),
    .C1(_08384_),
    .B1(_08399_),
    .A1(net1048),
    .Y(_08407_),
    .A2(_08402_));
 sg13g2_a21oi_1 _13914_ (.A1(_08401_),
    .A2(_08407_),
    .Y(_08408_),
    .B1(_08387_));
 sg13g2_and2_1 _13915_ (.A(_08406_),
    .B(_08408_),
    .X(_08409_));
 sg13g2_o21ai_1 _13916_ (.B1(_08409_),
    .Y(_08410_),
    .A1(_08378_),
    .A2(_08398_));
 sg13g2_xnor2_1 _13917_ (.Y(_08411_),
    .A(_08218_),
    .B(_08410_));
 sg13g2_buf_1 _13918_ (.A(\top_ihp.oisc.state[1] ),
    .X(_08412_));
 sg13g2_buf_1 _13919_ (.A(_08412_),
    .X(_08413_));
 sg13g2_nand2_2 _13920_ (.Y(_08414_),
    .A(_08200_),
    .B(net892));
 sg13g2_buf_1 _13921_ (.A(\top_ihp.oisc.decoder.decoded[11] ),
    .X(_08415_));
 sg13g2_nor2_2 _13922_ (.A(_08201_),
    .B(_08415_),
    .Y(_08416_));
 sg13g2_nor3_1 _13923_ (.A(net1028),
    .B(_08414_),
    .C(_08416_),
    .Y(_08417_));
 sg13g2_buf_1 _13924_ (.A(_08417_),
    .X(_08418_));
 sg13g2_buf_1 _13925_ (.A(net1028),
    .X(_08419_));
 sg13g2_buf_1 _13926_ (.A(net984),
    .X(_08420_));
 sg13g2_a21o_1 _13927_ (.A2(net832),
    .A1(_08411_),
    .B1(net934),
    .X(_08421_));
 sg13g2_or3_1 _13928_ (.A(net1028),
    .B(_08414_),
    .C(_08416_),
    .X(_08422_));
 sg13g2_buf_1 _13929_ (.A(_08422_),
    .X(_08423_));
 sg13g2_buf_1 _13930_ (.A(_08423_),
    .X(_08424_));
 sg13g2_nor3_1 _13931_ (.A(net1031),
    .B(_08411_),
    .C(_08424_),
    .Y(_08425_));
 sg13g2_a21o_1 _13932_ (.A2(_08421_),
    .A1(net1031),
    .B1(_08425_),
    .X(_08426_));
 sg13g2_nand2_1 _13933_ (.Y(_08427_),
    .A(_08215_),
    .B(_08426_));
 sg13g2_buf_2 _13934_ (.A(\top_ihp.wb_spi.bits_left[0] ),
    .X(_08428_));
 sg13g2_buf_1 _13935_ (.A(\top_ihp.wb_spi.bits_left[1] ),
    .X(_08429_));
 sg13g2_nor4_2 _13936_ (.A(_08429_),
    .B(\top_ihp.wb_spi.bits_left[3] ),
    .C(\top_ihp.wb_spi.bits_left[2] ),
    .Y(_08430_),
    .D(\top_ihp.wb_spi.bits_left[4] ));
 sg13g2_nor2b_1 _13937_ (.A(\top_ihp.wb_spi.bits_left[5] ),
    .B_N(_08430_),
    .Y(_08431_));
 sg13g2_nand2_1 _13938_ (.Y(_08432_),
    .A(_08428_),
    .B(_08431_));
 sg13g2_nand2b_1 _13939_ (.Y(_08433_),
    .B(\top_ihp.spi_clk_o ),
    .A_N(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_buf_1 _13940_ (.A(_08433_),
    .X(_08434_));
 sg13g2_buf_1 _13941_ (.A(_08214_),
    .X(_08435_));
 sg13g2_buf_1 _13942_ (.A(net1027),
    .X(_08436_));
 sg13g2_o21ai_1 _13943_ (.B1(net983),
    .Y(_08437_),
    .A1(_08432_),
    .A2(_08434_));
 sg13g2_o21ai_1 _13944_ (.B1(_08437_),
    .Y(_13704_),
    .A1(_08213_),
    .A2(_08427_));
 sg13g2_and3_1 _13945_ (.X(_08438_),
    .A(_08200_),
    .B(_08201_),
    .C(net892));
 sg13g2_buf_1 _13946_ (.A(_08438_),
    .X(_08439_));
 sg13g2_buf_1 _13947_ (.A(_08439_),
    .X(_08440_));
 sg13g2_buf_1 _13948_ (.A(net831),
    .X(_08441_));
 sg13g2_or3_1 _13949_ (.A(_08215_),
    .B(_08432_),
    .C(_08434_),
    .X(_08442_));
 sg13g2_o21ai_1 _13950_ (.B1(_08442_),
    .Y(_13703_),
    .A1(_08441_),
    .A2(_08427_));
 sg13g2_buf_2 _13951_ (.A(\top_ihp.oisc.op_a[28] ),
    .X(_08443_));
 sg13g2_buf_2 _13952_ (.A(\top_ihp.oisc.op_b[28] ),
    .X(_08444_));
 sg13g2_nand2b_1 _13953_ (.Y(_08445_),
    .B(_08444_),
    .A_N(_08443_));
 sg13g2_buf_1 _13954_ (.A(_08445_),
    .X(_08446_));
 sg13g2_inv_1 _13955_ (.Y(_08447_),
    .A(_08444_));
 sg13g2_nand2_1 _13956_ (.Y(_08448_),
    .A(_08443_),
    .B(_08447_));
 sg13g2_nand2_1 _13957_ (.Y(_08449_),
    .A(_08446_),
    .B(_08448_));
 sg13g2_buf_1 _13958_ (.A(\top_ihp.oisc.op_a[27] ),
    .X(_08450_));
 sg13g2_inv_1 _13959_ (.Y(_08451_),
    .A(\top_ihp.oisc.op_b[27] ));
 sg13g2_inv_1 _13960_ (.Y(_08452_),
    .A(_08278_));
 sg13g2_nor2b_1 _13961_ (.A(_08353_),
    .B_N(_08354_),
    .Y(_08453_));
 sg13g2_nor2_1 _13962_ (.A(_08263_),
    .B(_08453_),
    .Y(_08454_));
 sg13g2_nand2_1 _13963_ (.Y(_08455_),
    .A(_08263_),
    .B(_08453_));
 sg13g2_o21ai_1 _13964_ (.B1(_08455_),
    .Y(_08456_),
    .A1(net1053),
    .A2(_08454_));
 sg13g2_buf_1 _13965_ (.A(_08456_),
    .X(_08457_));
 sg13g2_nor2_1 _13966_ (.A(_08253_),
    .B(_08298_),
    .Y(_08458_));
 sg13g2_nand2_1 _13967_ (.Y(_08459_),
    .A(_08253_),
    .B(_08298_));
 sg13g2_o21ai_1 _13968_ (.B1(_08459_),
    .Y(_08460_),
    .A1(_08252_),
    .A2(_08458_));
 sg13g2_nand2b_1 _13969_ (.Y(_08461_),
    .B(net1055),
    .A_N(_08251_));
 sg13g2_nor2b_1 _13970_ (.A(net1055),
    .B_N(_08251_),
    .Y(_08462_));
 sg13g2_a221oi_1 _13971_ (.B2(_08461_),
    .C1(_08462_),
    .B1(_08460_),
    .A1(_08300_),
    .Y(_08463_),
    .A2(_08457_));
 sg13g2_o21ai_1 _13972_ (.B1(net1051),
    .Y(_08464_),
    .A1(_08452_),
    .A2(_08463_));
 sg13g2_nand2_1 _13973_ (.Y(_08465_),
    .A(_08452_),
    .B(_08463_));
 sg13g2_nor2b_1 _13974_ (.A(_08341_),
    .B_N(_08342_),
    .Y(_08466_));
 sg13g2_o21ai_1 _13975_ (.B1(_08365_),
    .Y(_08467_),
    .A1(net1029),
    .A2(_08466_));
 sg13g2_a21oi_1 _13976_ (.A1(net1029),
    .A2(_08466_),
    .Y(_08468_),
    .B1(_08361_));
 sg13g2_nand2_1 _13977_ (.Y(_08469_),
    .A(_08467_),
    .B(_08468_));
 sg13g2_nor2b_1 _13978_ (.A(_08339_),
    .B_N(net1049),
    .Y(_08470_));
 sg13g2_a221oi_1 _13979_ (.B2(_08337_),
    .C1(_08470_),
    .B1(_08335_),
    .A1(_08325_),
    .Y(_08471_),
    .A2(_08333_));
 sg13g2_nand2b_1 _13980_ (.Y(_08472_),
    .B(_08341_),
    .A_N(_08342_));
 sg13g2_o21ai_1 _13981_ (.B1(_08365_),
    .Y(_08473_),
    .A1(net1029),
    .A2(_08472_));
 sg13g2_nand2_1 _13982_ (.Y(_08474_),
    .A(net1029),
    .B(_08472_));
 sg13g2_nand2_1 _13983_ (.Y(_08475_),
    .A(_08352_),
    .B(_08344_));
 sg13g2_a21oi_1 _13984_ (.A1(_08473_),
    .A2(_08474_),
    .Y(_08476_),
    .B1(_08475_));
 sg13g2_o21ai_1 _13985_ (.B1(_08476_),
    .Y(_08477_),
    .A1(_08469_),
    .A2(_08471_));
 sg13g2_buf_1 _13986_ (.A(_08477_),
    .X(_08478_));
 sg13g2_nand2b_1 _13987_ (.Y(_08479_),
    .B(_08315_),
    .A_N(_08314_));
 sg13g2_o21ai_1 _13988_ (.B1(_08350_),
    .Y(_08480_),
    .A1(_08359_),
    .A2(_08479_));
 sg13g2_o21ai_1 _13989_ (.B1(_08480_),
    .Y(_08481_),
    .A1(_08351_),
    .A2(_08316_));
 sg13g2_buf_1 _13990_ (.A(_08481_),
    .X(_08482_));
 sg13g2_and3_1 _13991_ (.X(_08483_),
    .A(_08300_),
    .B(_08301_),
    .C(_08355_));
 sg13g2_nand2_1 _13992_ (.Y(_08484_),
    .A(_08305_),
    .B(_08483_));
 sg13g2_a21oi_1 _13993_ (.A1(_08478_),
    .A2(_08482_),
    .Y(_08485_),
    .B1(_08484_));
 sg13g2_a21o_1 _13994_ (.A2(_08465_),
    .A1(_08464_),
    .B1(_08485_),
    .X(_08486_));
 sg13g2_buf_2 _13995_ (.A(_08486_),
    .X(_08487_));
 sg13g2_nor2_1 _13996_ (.A(_08304_),
    .B(_08307_),
    .Y(_08488_));
 sg13g2_xor2_1 _13997_ (.B(_08219_),
    .A(net1058),
    .X(_08489_));
 sg13g2_or2_1 _13998_ (.X(_08490_),
    .B(_08233_),
    .A(_08229_));
 sg13g2_buf_1 _13999_ (.A(_08490_),
    .X(_08491_));
 sg13g2_xnor2_1 _14000_ (.Y(_08492_),
    .A(net1059),
    .B(_08220_));
 sg13g2_nand2b_1 _14001_ (.Y(_08493_),
    .B(_08492_),
    .A_N(_08308_));
 sg13g2_buf_1 _14002_ (.A(_08493_),
    .X(_08494_));
 sg13g2_or3_1 _14003_ (.A(_08489_),
    .B(_08491_),
    .C(_08494_),
    .X(_08495_));
 sg13g2_buf_1 _14004_ (.A(_08495_),
    .X(_08496_));
 sg13g2_nor2b_1 _14005_ (.A(_08235_),
    .B_N(_08231_),
    .Y(_08497_));
 sg13g2_or2_1 _14006_ (.X(_08498_),
    .B(_08249_),
    .A(_08497_));
 sg13g2_buf_1 _14007_ (.A(_08498_),
    .X(_08499_));
 sg13g2_or2_1 _14008_ (.X(_08500_),
    .B(_08499_),
    .A(_08393_));
 sg13g2_nor2_1 _14009_ (.A(_08496_),
    .B(_08500_),
    .Y(_08501_));
 sg13g2_nand2_1 _14010_ (.Y(_08502_),
    .A(_08218_),
    .B(_08216_));
 sg13g2_nand2b_1 _14011_ (.Y(_08503_),
    .B(\top_ihp.oisc.op_b[26] ),
    .A_N(_08216_));
 sg13g2_nand3_1 _14012_ (.B(_08502_),
    .C(_08503_),
    .A(_08390_),
    .Y(_08504_));
 sg13g2_buf_1 _14013_ (.A(_08504_),
    .X(_08505_));
 sg13g2_nor2_1 _14014_ (.A(_08396_),
    .B(_08505_),
    .Y(_08506_));
 sg13g2_and3_1 _14015_ (.X(_08507_),
    .A(_08488_),
    .B(_08501_),
    .C(_08506_));
 sg13g2_inv_1 _14016_ (.Y(_08508_),
    .A(_08391_));
 sg13g2_nand2b_1 _14017_ (.Y(_08509_),
    .B(_08279_),
    .A_N(_08287_));
 sg13g2_o21ai_1 _14018_ (.B1(_08282_),
    .Y(_08510_),
    .A1(_08273_),
    .A2(_08509_));
 sg13g2_nand2_1 _14019_ (.Y(_08511_),
    .A(_08273_),
    .B(_08509_));
 sg13g2_nand3b_1 _14020_ (.B(_08510_),
    .C(_08511_),
    .Y(_08512_),
    .A_N(_08494_));
 sg13g2_nor2_1 _14021_ (.A(net1058),
    .B(_08245_),
    .Y(_08513_));
 sg13g2_inv_1 _14022_ (.Y(_08514_),
    .A(_08220_));
 sg13g2_nor2_1 _14023_ (.A(_08514_),
    .B(_08277_),
    .Y(_08515_));
 sg13g2_a21oi_1 _14024_ (.A1(_08514_),
    .A2(_08277_),
    .Y(_08516_),
    .B1(net1059));
 sg13g2_nor4_1 _14025_ (.A(_08233_),
    .B(_08513_),
    .C(_08515_),
    .D(_08516_),
    .Y(_08517_));
 sg13g2_nand2_1 _14026_ (.Y(_08518_),
    .A(net1058),
    .B(_08245_));
 sg13g2_nand2_1 _14027_ (.Y(_08519_),
    .A(net1057),
    .B(_08518_));
 sg13g2_nor2_1 _14028_ (.A(net1057),
    .B(_08518_),
    .Y(_08520_));
 sg13g2_a221oi_1 _14029_ (.B2(net1056),
    .C1(_08520_),
    .B1(_08519_),
    .A1(_08512_),
    .Y(_08521_),
    .A2(_08517_));
 sg13g2_a221oi_1 _14030_ (.B2(_08231_),
    .C1(_08521_),
    .B1(_08236_),
    .A1(_08508_),
    .Y(_08522_),
    .A2(_08392_));
 sg13g2_inv_1 _14031_ (.Y(_08523_),
    .A(_08392_));
 sg13g2_o21ai_1 _14032_ (.B1(_08249_),
    .Y(_08524_),
    .A1(_08391_),
    .A2(_08523_));
 sg13g2_o21ai_1 _14033_ (.B1(_08524_),
    .Y(_08525_),
    .A1(_08508_),
    .A2(_08392_));
 sg13g2_nor2_1 _14034_ (.A(_08522_),
    .B(_08525_),
    .Y(_08526_));
 sg13g2_nor2b_1 _14035_ (.A(net1047),
    .B_N(_08395_),
    .Y(_08527_));
 sg13g2_buf_1 _14036_ (.A(_08527_),
    .X(_08528_));
 sg13g2_nor2_1 _14037_ (.A(_08379_),
    .B(_08528_),
    .Y(_08529_));
 sg13g2_nand2_1 _14038_ (.Y(_08530_),
    .A(_08379_),
    .B(_08528_));
 sg13g2_o21ai_1 _14039_ (.B1(_08530_),
    .Y(_08531_),
    .A1(net1048),
    .A2(_08529_));
 sg13g2_a21oi_1 _14040_ (.A1(_08388_),
    .A2(_08531_),
    .Y(_08532_),
    .B1(_08387_));
 sg13g2_a21o_1 _14041_ (.A2(_08532_),
    .A1(net1031),
    .B1(_08218_),
    .X(_08533_));
 sg13g2_o21ai_1 _14042_ (.B1(_08533_),
    .Y(_08534_),
    .A1(net1031),
    .A2(_08532_));
 sg13g2_a221oi_1 _14043_ (.B2(_08506_),
    .C1(_08534_),
    .B1(_08526_),
    .A1(_08487_),
    .Y(_08535_),
    .A2(_08507_));
 sg13g2_a21oi_1 _14044_ (.A1(net1046),
    .A2(_08451_),
    .Y(_08536_),
    .B1(_08535_));
 sg13g2_nor2_1 _14045_ (.A(net1046),
    .B(_08451_),
    .Y(_08537_));
 sg13g2_buf_1 _14046_ (.A(_08537_),
    .X(_08538_));
 sg13g2_nor2_1 _14047_ (.A(_08536_),
    .B(_08538_),
    .Y(_08539_));
 sg13g2_xor2_1 _14048_ (.B(_08539_),
    .A(_08449_),
    .X(_08540_));
 sg13g2_a22oi_1 _14049_ (.Y(_08541_),
    .B1(net832),
    .B2(_08540_),
    .A2(_08443_),
    .A1(net934));
 sg13g2_buf_1 _14050_ (.A(_08541_),
    .X(_08542_));
 sg13g2_buf_1 _14051_ (.A(_00094_),
    .X(_08543_));
 sg13g2_nor2b_1 _14052_ (.A(_08542_),
    .B_N(_08543_),
    .Y(_00004_));
 sg13g2_buf_1 _14053_ (.A(\top_ihp.wb_imem.state[0] ),
    .X(_08544_));
 sg13g2_buf_1 _14054_ (.A(\top_ihp.oisc.op_a[30] ),
    .X(_08545_));
 sg13g2_buf_2 _14055_ (.A(_08545_),
    .X(_08546_));
 sg13g2_nand2_1 _14056_ (.Y(_08547_),
    .A(net984),
    .B(net1026));
 sg13g2_buf_1 _14057_ (.A(_08418_),
    .X(_08548_));
 sg13g2_inv_1 _14058_ (.Y(_08549_),
    .A(\top_ihp.oisc.op_b[30] ));
 sg13g2_nand2_1 _14059_ (.Y(_08550_),
    .A(_08312_),
    .B(_08376_));
 sg13g2_or2_1 _14060_ (.X(_08551_),
    .B(_08396_),
    .A(_08393_));
 sg13g2_a21oi_1 _14061_ (.A1(_08237_),
    .A2(_08238_),
    .Y(_08552_),
    .B1(_08551_));
 sg13g2_nor2b_1 _14062_ (.A(\top_ihp.oisc.op_b[27] ),
    .B_N(net1046),
    .Y(_08553_));
 sg13g2_buf_1 _14063_ (.A(_08553_),
    .X(_08554_));
 sg13g2_nor2_1 _14064_ (.A(_08538_),
    .B(_08554_),
    .Y(_08555_));
 sg13g2_nand2b_1 _14065_ (.Y(_08556_),
    .B(_08555_),
    .A_N(_08449_));
 sg13g2_buf_1 _14066_ (.A(\top_ihp.oisc.op_a[29] ),
    .X(_08557_));
 sg13g2_buf_2 _14067_ (.A(\top_ihp.oisc.op_b[29] ),
    .X(_08558_));
 sg13g2_xor2_1 _14068_ (.B(_08558_),
    .A(net1045),
    .X(_08559_));
 sg13g2_buf_2 _14069_ (.A(_08559_),
    .X(_08560_));
 sg13g2_nor3_1 _14070_ (.A(_08505_),
    .B(_08556_),
    .C(_08560_),
    .Y(_08561_));
 sg13g2_nand2_1 _14071_ (.Y(_08562_),
    .A(_08552_),
    .B(_08561_));
 sg13g2_nand2b_1 _14072_ (.Y(_08563_),
    .B(_08558_),
    .A_N(net1045));
 sg13g2_nor2_1 _14073_ (.A(_08447_),
    .B(_08554_),
    .Y(_08564_));
 sg13g2_a21oi_1 _14074_ (.A1(_08447_),
    .A2(_08554_),
    .Y(_08565_),
    .B1(_08443_));
 sg13g2_nor2_1 _14075_ (.A(_08564_),
    .B(_08565_),
    .Y(_08566_));
 sg13g2_nor2b_1 _14076_ (.A(_08558_),
    .B_N(net1045),
    .Y(_08567_));
 sg13g2_a21oi_1 _14077_ (.A1(_08563_),
    .A2(_08566_),
    .Y(_08568_),
    .B1(_08567_));
 sg13g2_inv_1 _14078_ (.Y(_08569_),
    .A(_08558_));
 sg13g2_o21ai_1 _14079_ (.B1(net1045),
    .Y(_08570_),
    .A1(_08569_),
    .A2(_08446_));
 sg13g2_nand2_1 _14080_ (.Y(_08571_),
    .A(_08569_),
    .B(_08446_));
 sg13g2_a21oi_1 _14081_ (.A1(_08570_),
    .A2(_08571_),
    .Y(_08572_),
    .B1(_08538_));
 sg13g2_nand4_1 _14082_ (.B(_08406_),
    .C(_08408_),
    .A(_08216_),
    .Y(_08573_),
    .D(_08572_));
 sg13g2_nand4_1 _14083_ (.B(_08406_),
    .C(_08408_),
    .A(_08218_),
    .Y(_08574_),
    .D(_08572_));
 sg13g2_nand2b_1 _14084_ (.Y(_08575_),
    .B(_08572_),
    .A_N(_08502_));
 sg13g2_nand4_1 _14085_ (.B(_08573_),
    .C(_08574_),
    .A(_08568_),
    .Y(_08576_),
    .D(_08575_));
 sg13g2_o21ai_1 _14086_ (.B1(_08576_),
    .Y(_08577_),
    .A1(_08550_),
    .A2(_08562_));
 sg13g2_xnor2_1 _14087_ (.Y(_08578_),
    .A(_08549_),
    .B(_08577_));
 sg13g2_xnor2_1 _14088_ (.Y(_08579_),
    .A(net1026),
    .B(_08578_));
 sg13g2_nand2_1 _14089_ (.Y(_08580_),
    .A(net796),
    .B(_08579_));
 sg13g2_buf_1 _14090_ (.A(_08440_),
    .X(_08581_));
 sg13g2_a21oi_1 _14091_ (.A1(_08547_),
    .A2(_08580_),
    .Y(_08582_),
    .B1(net795));
 sg13g2_buf_2 _14092_ (.A(\top_ihp.wb_imem.bits_left[2] ),
    .X(_08583_));
 sg13g2_nor4_2 _14093_ (.A(_08583_),
    .B(\top_ihp.wb_imem.bits_left[3] ),
    .C(\top_ihp.wb_imem.bits_left[5] ),
    .Y(_08584_),
    .D(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_buf_1 _14094_ (.A(\top_ihp.wb_imem.bits_left[1] ),
    .X(_08585_));
 sg13g2_buf_2 _14095_ (.A(\top_ihp.wb_imem.bits_left[0] ),
    .X(_08586_));
 sg13g2_nor2b_1 _14096_ (.A(_08585_),
    .B_N(_08586_),
    .Y(_08587_));
 sg13g2_nand2_1 _14097_ (.Y(_08588_),
    .A(_08584_),
    .B(_08587_));
 sg13g2_buf_1 _14098_ (.A(\top_ihp.wb_imem.state[2] ),
    .X(_08589_));
 sg13g2_a22oi_1 _14099_ (.Y(_08590_),
    .B1(_08588_),
    .B2(_08589_),
    .A2(_08582_),
    .A1(_08544_));
 sg13g2_inv_1 _14100_ (.Y(_00001_),
    .A(_08590_));
 sg13g2_buf_1 _14101_ (.A(_00095_),
    .X(_08591_));
 sg13g2_nor2_1 _14102_ (.A(_08586_),
    .B(_08585_),
    .Y(_08592_));
 sg13g2_and2_1 _14103_ (.A(_08584_),
    .B(_08592_),
    .X(_08593_));
 sg13g2_buf_1 _14104_ (.A(_08593_),
    .X(_08594_));
 sg13g2_buf_1 _14105_ (.A(_08594_),
    .X(_08595_));
 sg13g2_and2_1 _14106_ (.A(_08584_),
    .B(_08587_),
    .X(_08596_));
 sg13g2_nand2_1 _14107_ (.Y(_08597_),
    .A(_08589_),
    .B(_08596_));
 sg13g2_o21ai_1 _14108_ (.B1(_08597_),
    .Y(_00000_),
    .A1(_08591_),
    .A2(net862));
 sg13g2_buf_2 _14109_ (.A(\top_ihp.wb_ack_coproc ),
    .X(_08598_));
 sg13g2_nand3_1 _14110_ (.B(_08488_),
    .C(_08501_),
    .A(_08487_),
    .Y(_08599_));
 sg13g2_nand2b_1 _14111_ (.Y(_08600_),
    .B(_08599_),
    .A_N(_08526_));
 sg13g2_a21oi_1 _14112_ (.A1(_08506_),
    .A2(_08600_),
    .Y(_08601_),
    .B1(_08534_));
 sg13g2_xor2_1 _14113_ (.B(_08601_),
    .A(_08555_),
    .X(_08602_));
 sg13g2_nand2_1 _14114_ (.Y(_08603_),
    .A(net934),
    .B(net1046));
 sg13g2_o21ai_1 _14115_ (.B1(_08603_),
    .Y(_08604_),
    .A1(net798),
    .A2(_08602_));
 sg13g2_nor2b_1 _14116_ (.A(_08598_),
    .B_N(_08604_),
    .Y(_00003_));
 sg13g2_xor2_1 _14117_ (.B(_08323_),
    .A(_08319_),
    .X(_08605_));
 sg13g2_a21o_1 _14118_ (.A2(_08605_),
    .A1(net832),
    .B1(net984),
    .X(_08606_));
 sg13g2_nor2_1 _14119_ (.A(_08317_),
    .B(_08605_),
    .Y(_08607_));
 sg13g2_nor3_1 _14120_ (.A(_08419_),
    .B(_08414_),
    .C(_08416_),
    .Y(_08608_));
 sg13g2_buf_2 _14121_ (.A(_08608_),
    .X(_08609_));
 sg13g2_a22oi_1 _14122_ (.Y(_08610_),
    .B1(_08607_),
    .B2(_08609_),
    .A2(_08606_),
    .A1(_08317_));
 sg13g2_buf_1 _14123_ (.A(_08610_),
    .X(_08611_));
 sg13g2_inv_1 _14124_ (.Y(\top_ihp.oisc.wb_adr_o[1] ),
    .A(_08611_));
 sg13g2_or3_1 _14125_ (.A(net1028),
    .B(_08414_),
    .C(_08416_),
    .X(_08612_));
 sg13g2_buf_1 _14126_ (.A(_08612_),
    .X(_08613_));
 sg13g2_nand2b_1 _14127_ (.Y(_08614_),
    .B(_08320_),
    .A_N(_08321_));
 sg13g2_inv_1 _14128_ (.Y(_08615_),
    .A(_08412_));
 sg13g2_o21ai_1 _14129_ (.B1(_08615_),
    .Y(_08616_),
    .A1(_08320_),
    .A2(net798));
 sg13g2_nand2_1 _14130_ (.Y(_08617_),
    .A(_08321_),
    .B(_08616_));
 sg13g2_o21ai_1 _14131_ (.B1(_08617_),
    .Y(_08618_),
    .A1(_08613_),
    .A2(_08614_));
 sg13g2_buf_2 _14132_ (.A(_08618_),
    .X(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_buf_1 _14133_ (.A(\top_ihp.wb_uart.uart_rx.state[0] ),
    .X(_08619_));
 sg13g2_buf_1 _14134_ (.A(_00098_),
    .X(_08620_));
 sg13g2_nor2b_1 _14135_ (.A(_08449_),
    .B_N(_08555_),
    .Y(_08621_));
 sg13g2_nand3b_1 _14136_ (.B(_08506_),
    .C(_08621_),
    .Y(_08622_),
    .A_N(_08500_));
 sg13g2_buf_1 _14137_ (.A(_08622_),
    .X(_08623_));
 sg13g2_or3_1 _14138_ (.A(_08496_),
    .B(_08560_),
    .C(_08623_),
    .X(_08624_));
 sg13g2_a21oi_1 _14139_ (.A1(_08392_),
    .A2(_08497_),
    .Y(_08625_),
    .B1(_08508_));
 sg13g2_a221oi_1 _14140_ (.B2(_08241_),
    .C1(_08625_),
    .B1(_08523_),
    .A1(net1047),
    .Y(_08626_),
    .A2(_08399_));
 sg13g2_buf_1 _14141_ (.A(_08626_),
    .X(_08627_));
 sg13g2_o21ai_1 _14142_ (.B1(_08379_),
    .Y(_08628_),
    .A1(_08528_),
    .A2(_08627_));
 sg13g2_nor3_1 _14143_ (.A(_08379_),
    .B(_08528_),
    .C(_08627_),
    .Y(_08629_));
 sg13g2_a21oi_1 _14144_ (.A1(net1048),
    .A2(_08628_),
    .Y(_08630_),
    .B1(_08629_));
 sg13g2_and3_1 _14145_ (.X(_08631_),
    .A(_08388_),
    .B(_08502_),
    .C(_08621_));
 sg13g2_o21ai_1 _14146_ (.B1(_08631_),
    .Y(_08632_),
    .A1(_08387_),
    .A2(_08630_));
 sg13g2_buf_1 _14147_ (.A(_08632_),
    .X(_08633_));
 sg13g2_nor2_1 _14148_ (.A(_08503_),
    .B(_08554_),
    .Y(_08634_));
 sg13g2_o21ai_1 _14149_ (.B1(_08448_),
    .Y(_08635_),
    .A1(_08538_),
    .A2(_08634_));
 sg13g2_and2_1 _14150_ (.A(_08446_),
    .B(_08635_),
    .X(_08636_));
 sg13g2_buf_1 _14151_ (.A(_08636_),
    .X(_08637_));
 sg13g2_nor2_1 _14152_ (.A(_08515_),
    .B(_08516_),
    .Y(_08638_));
 sg13g2_buf_2 _14153_ (.A(_08638_),
    .X(_08639_));
 sg13g2_a21o_1 _14154_ (.A2(_08639_),
    .A1(_08245_),
    .B1(net1058),
    .X(_08640_));
 sg13g2_o21ai_1 _14155_ (.B1(_08640_),
    .Y(_08641_),
    .A1(_08245_),
    .A2(_08639_));
 sg13g2_nand2b_1 _14156_ (.Y(_08642_),
    .B(net1056),
    .A_N(net1057));
 sg13g2_o21ai_1 _14157_ (.B1(_08642_),
    .Y(_08643_),
    .A1(_08233_),
    .A2(_08641_));
 sg13g2_buf_1 _14158_ (.A(_08643_),
    .X(_08644_));
 sg13g2_nand4_1 _14159_ (.B(_08633_),
    .C(_08637_),
    .A(_08560_),
    .Y(_08645_),
    .D(_08644_));
 sg13g2_a22oi_1 _14160_ (.Y(_08646_),
    .B1(_08510_),
    .B2(_08511_),
    .A2(_08488_),
    .A1(_08487_));
 sg13g2_buf_2 _14161_ (.A(_08646_),
    .X(_08647_));
 sg13g2_mux2_1 _14162_ (.A0(_08624_),
    .A1(_08645_),
    .S(_08647_),
    .X(_08648_));
 sg13g2_nand4_1 _14163_ (.B(_08633_),
    .C(_08637_),
    .A(_08560_),
    .Y(_08649_),
    .D(_08623_));
 sg13g2_a21o_1 _14164_ (.A2(_08637_),
    .A1(_08633_),
    .B1(_08560_),
    .X(_08650_));
 sg13g2_and2_1 _14165_ (.A(_08496_),
    .B(_08560_),
    .X(_08651_));
 sg13g2_nand4_1 _14166_ (.B(_08637_),
    .C(_08644_),
    .A(_08633_),
    .Y(_08652_),
    .D(_08651_));
 sg13g2_or3_1 _14167_ (.A(_08560_),
    .B(_08623_),
    .C(_08644_),
    .X(_08653_));
 sg13g2_and4_1 _14168_ (.A(_08649_),
    .B(_08650_),
    .C(_08652_),
    .D(_08653_),
    .X(_08654_));
 sg13g2_nand2_1 _14169_ (.Y(_08655_),
    .A(_08648_),
    .B(_08654_));
 sg13g2_buf_2 _14170_ (.A(\top_ihp.oisc.decoder.instruction[12] ),
    .X(_08656_));
 sg13g2_buf_1 _14171_ (.A(\top_ihp.oisc.decoder.instruction[13] ),
    .X(_08657_));
 sg13g2_buf_1 _14172_ (.A(_08657_),
    .X(_08658_));
 sg13g2_buf_1 _14173_ (.A(_00079_),
    .X(_08659_));
 sg13g2_inv_1 _14174_ (.Y(_08660_),
    .A(_08659_));
 sg13g2_a21oi_1 _14175_ (.A1(_08656_),
    .A2(net1025),
    .Y(_08661_),
    .B1(_08660_));
 sg13g2_buf_1 _14176_ (.A(_08661_),
    .X(_08662_));
 sg13g2_nand3_1 _14177_ (.B(_08609_),
    .C(_08662_),
    .A(_08213_),
    .Y(_08663_));
 sg13g2_and2_1 _14178_ (.A(net984),
    .B(net1045),
    .X(_08664_));
 sg13g2_buf_1 _14179_ (.A(_08664_),
    .X(_08665_));
 sg13g2_nand3_1 _14180_ (.B(_08662_),
    .C(_08665_),
    .A(_08213_),
    .Y(_08666_));
 sg13g2_o21ai_1 _14181_ (.B1(_08666_),
    .Y(_08667_),
    .A1(_08655_),
    .A2(_08663_));
 sg13g2_nand3b_1 _14182_ (.B(_08620_),
    .C(_08667_),
    .Y(_08668_),
    .A_N(_08619_));
 sg13g2_buf_1 _14183_ (.A(net2),
    .X(_08669_));
 sg13g2_buf_1 _14184_ (.A(\top_ihp.wb_uart.uart_rx.state[2] ),
    .X(_08670_));
 sg13g2_nor2b_1 _14185_ (.A(_08670_),
    .B_N(_08619_),
    .Y(_08671_));
 sg13g2_buf_2 _14186_ (.A(\top_ihp.wb_uart.uart_rx.state[1] ),
    .X(_08672_));
 sg13g2_a21oi_1 _14187_ (.A1(net1060),
    .A2(_08671_),
    .Y(_08673_),
    .B1(_08672_));
 sg13g2_buf_1 _14188_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ),
    .X(_08674_));
 sg13g2_buf_1 _14189_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ),
    .X(_08675_));
 sg13g2_nor4_1 _14190_ (.A(_08674_),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ),
    .C(_08675_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .Y(_08676_));
 sg13g2_buf_2 _14191_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ),
    .X(_08677_));
 sg13g2_buf_1 _14192_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ),
    .X(_08678_));
 sg13g2_buf_1 _14193_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ),
    .X(_08679_));
 sg13g2_nor4_1 _14194_ (.A(_08677_),
    .B(_08678_),
    .C(_08679_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ),
    .Y(_08680_));
 sg13g2_buf_1 _14195_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ),
    .X(_08681_));
 sg13g2_buf_1 _14196_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ),
    .X(_08682_));
 sg13g2_nor4_1 _14197_ (.A(_08681_),
    .B(_08682_),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ),
    .Y(_08683_));
 sg13g2_buf_2 _14198_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ),
    .X(_08684_));
 sg13g2_nor3_1 _14199_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ),
    .C(_08684_),
    .Y(_08685_));
 sg13g2_nand4_1 _14200_ (.B(_08680_),
    .C(_08683_),
    .A(_08676_),
    .Y(_08686_),
    .D(_08685_));
 sg13g2_buf_2 _14201_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ),
    .X(_08687_));
 sg13g2_nor4_1 _14202_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .B(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .C(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .D(_08687_),
    .Y(_08688_));
 sg13g2_buf_1 _14203_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ),
    .X(_08689_));
 sg13g2_buf_1 _14204_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ),
    .X(_08690_));
 sg13g2_nor4_1 _14205_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_08689_),
    .C(_08690_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .Y(_08691_));
 sg13g2_nand2_1 _14206_ (.Y(_08692_),
    .A(_08688_),
    .B(_08691_));
 sg13g2_inv_1 _14207_ (.Y(_08693_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ));
 sg13g2_buf_1 _14208_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ),
    .X(_08694_));
 sg13g2_buf_8 _14209_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ),
    .X(_08695_));
 sg13g2_buf_2 _14210_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ),
    .X(_08696_));
 sg13g2_inv_1 _14211_ (.Y(_08697_),
    .A(_08696_));
 sg13g2_buf_1 _14212_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ),
    .X(_08698_));
 sg13g2_inv_2 _14213_ (.Y(_08699_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ));
 sg13g2_nor4_1 _14214_ (.A(_08695_),
    .B(_08697_),
    .C(_08698_),
    .D(_08699_),
    .Y(_08700_));
 sg13g2_nand3_1 _14215_ (.B(_08694_),
    .C(_08700_),
    .A(_08693_),
    .Y(_08701_));
 sg13g2_buf_8 _14216_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ),
    .X(_08702_));
 sg13g2_buf_8 _14217_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ),
    .X(_08703_));
 sg13g2_buf_8 _14218_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ),
    .X(_08704_));
 sg13g2_nand3b_1 _14219_ (.B(_08703_),
    .C(_08704_),
    .Y(_08705_),
    .A_N(_08702_));
 sg13g2_nor4_2 _14220_ (.A(_08686_),
    .B(_08692_),
    .C(_08701_),
    .Y(_08706_),
    .D(_08705_));
 sg13g2_buf_2 _14221_ (.A(_08706_),
    .X(_08707_));
 sg13g2_buf_1 _14222_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ),
    .X(_08708_));
 sg13g2_buf_1 _14223_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ),
    .X(_08709_));
 sg13g2_buf_1 _14224_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ),
    .X(_08710_));
 sg13g2_nand3_1 _14225_ (.B(net1043),
    .C(net1042),
    .A(net1044),
    .Y(_08711_));
 sg13g2_buf_1 _14226_ (.A(_08711_),
    .X(_08712_));
 sg13g2_nor2_1 _14227_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .B(_08712_),
    .Y(_08713_));
 sg13g2_nand3_1 _14228_ (.B(_08707_),
    .C(_08713_),
    .A(_08619_),
    .Y(_08714_));
 sg13g2_and2_1 _14229_ (.A(_08620_),
    .B(_08714_),
    .X(_08715_));
 sg13g2_o21ai_1 _14230_ (.B1(_08715_),
    .Y(_08716_),
    .A1(_08619_),
    .A2(_08707_));
 sg13g2_a22oi_1 _14231_ (.Y(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .B1(_08716_),
    .B2(_08672_),
    .A2(_08673_),
    .A1(_08668_));
 sg13g2_nor2_1 _14232_ (.A(_08672_),
    .B(net1060),
    .Y(_08717_));
 sg13g2_a22oi_1 _14233_ (.Y(_08718_),
    .B1(_08717_),
    .B2(_08671_),
    .A2(_08715_),
    .A1(_08672_));
 sg13g2_inv_1 _14234_ (.Y(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .A(_08718_));
 sg13g2_nor2_1 _14235_ (.A(_08672_),
    .B(_08619_),
    .Y(_08719_));
 sg13g2_and2_1 _14236_ (.A(_08670_),
    .B(_08719_),
    .X(_08720_));
 sg13g2_nand3_1 _14237_ (.B(_08619_),
    .C(_08620_),
    .A(_08672_),
    .Y(_08721_));
 sg13g2_buf_2 _14238_ (.A(_08721_),
    .X(_08722_));
 sg13g2_nor3_1 _14239_ (.A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .B(_08712_),
    .C(_08722_),
    .Y(_08723_));
 sg13g2_mux2_1 _14240_ (.A0(_08720_),
    .A1(_08723_),
    .S(_08707_),
    .X(\top_ihp.wb_uart.uart_rx.next_state[2] ));
 sg13g2_nand3_1 _14241_ (.B(_08667_),
    .C(_08673_),
    .A(_08620_),
    .Y(_08724_));
 sg13g2_xnor2_1 _14242_ (.Y(_08725_),
    .A(_08670_),
    .B(\top_ihp.wb_uart.uart_rx.next_state[2] ));
 sg13g2_nand2_1 _14243_ (.Y(_08726_),
    .A(_08672_),
    .B(_08620_));
 sg13g2_nand2b_1 _14244_ (.Y(_08727_),
    .B(net2),
    .A_N(_08670_));
 sg13g2_a21o_1 _14245_ (.A2(_08727_),
    .A1(_08619_),
    .B1(_08672_),
    .X(_08728_));
 sg13g2_o21ai_1 _14246_ (.B1(_08728_),
    .Y(_08729_),
    .A1(_08707_),
    .A2(_08726_));
 sg13g2_nand3_1 _14247_ (.B(_08725_),
    .C(_08729_),
    .A(_08724_),
    .Y(_08730_));
 sg13g2_buf_2 _14248_ (.A(_08730_),
    .X(_08731_));
 sg13g2_buf_8 _14249_ (.A(_08731_),
    .X(_08732_));
 sg13g2_nor2_1 _14250_ (.A(_08695_),
    .B(net149),
    .Y(_00005_));
 sg13g2_xnor2_1 _14251_ (.Y(_08733_),
    .A(_08695_),
    .B(_08704_));
 sg13g2_nor2_1 _14252_ (.A(net149),
    .B(_08733_),
    .Y(_00016_));
 sg13g2_nand2_1 _14253_ (.Y(_08734_),
    .A(_08695_),
    .B(_08704_));
 sg13g2_xor2_1 _14254_ (.B(_08734_),
    .A(_08702_),
    .X(_08735_));
 sg13g2_nor2_1 _14255_ (.A(net149),
    .B(_08735_),
    .Y(_00027_));
 sg13g2_nand3_1 _14256_ (.B(_08704_),
    .C(_08702_),
    .A(_08695_),
    .Y(_08736_));
 sg13g2_xor2_1 _14257_ (.B(_08736_),
    .A(_08703_),
    .X(_08737_));
 sg13g2_nor2_1 _14258_ (.A(net149),
    .B(_08737_),
    .Y(_00030_));
 sg13g2_nand4_1 _14259_ (.B(_08704_),
    .C(_08703_),
    .A(_08695_),
    .Y(_08738_),
    .D(_08702_));
 sg13g2_buf_1 _14260_ (.A(_08738_),
    .X(_08739_));
 sg13g2_xnor2_1 _14261_ (.Y(_08740_),
    .A(_08699_),
    .B(_08739_));
 sg13g2_nor2_1 _14262_ (.A(net149),
    .B(_08740_),
    .Y(_00031_));
 sg13g2_nor2_1 _14263_ (.A(_08699_),
    .B(_08739_),
    .Y(_08741_));
 sg13g2_xnor2_1 _14264_ (.Y(_08742_),
    .A(_00097_),
    .B(_08741_));
 sg13g2_nor2b_1 _14265_ (.A(net149),
    .B_N(_08742_),
    .Y(_00032_));
 sg13g2_nor3_2 _14266_ (.A(_08699_),
    .B(_08693_),
    .C(_08739_),
    .Y(_08743_));
 sg13g2_xnor2_1 _14267_ (.Y(_08744_),
    .A(_08696_),
    .B(_08743_));
 sg13g2_nor2_1 _14268_ (.A(net149),
    .B(_08744_),
    .Y(_00033_));
 sg13g2_inv_1 _14269_ (.Y(_08745_),
    .A(_08698_));
 sg13g2_nand2_1 _14270_ (.Y(_08746_),
    .A(_08696_),
    .B(_08743_));
 sg13g2_xnor2_1 _14271_ (.Y(_08747_),
    .A(_08745_),
    .B(_08746_));
 sg13g2_nor2_1 _14272_ (.A(_08732_),
    .B(_08747_),
    .Y(_00034_));
 sg13g2_nand3_1 _14273_ (.B(_08698_),
    .C(_08743_),
    .A(_08696_),
    .Y(_08748_));
 sg13g2_xor2_1 _14274_ (.B(_08748_),
    .A(_08694_),
    .X(_08749_));
 sg13g2_nor2_1 _14275_ (.A(_08732_),
    .B(_08749_),
    .Y(_00035_));
 sg13g2_and4_1 _14276_ (.A(_08696_),
    .B(_08698_),
    .C(_08694_),
    .D(_08743_),
    .X(_08750_));
 sg13g2_buf_8 _14277_ (.A(_08750_),
    .X(_08751_));
 sg13g2_xnor2_1 _14278_ (.Y(_08752_),
    .A(_08690_),
    .B(_08751_));
 sg13g2_nor2_1 _14279_ (.A(net149),
    .B(_08752_),
    .Y(_00036_));
 sg13g2_buf_1 _14280_ (.A(_08731_),
    .X(_08753_));
 sg13g2_nand2_1 _14281_ (.Y(_08754_),
    .A(_08690_),
    .B(_08751_));
 sg13g2_xor2_1 _14282_ (.B(_08754_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .X(_08755_));
 sg13g2_nor2_1 _14283_ (.A(net148),
    .B(_08755_),
    .Y(_00006_));
 sg13g2_and3_1 _14284_ (.X(_08756_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ),
    .B(_08690_),
    .C(_08751_));
 sg13g2_buf_8 _14285_ (.A(_08756_),
    .X(_08757_));
 sg13g2_xnor2_1 _14286_ (.Y(_08758_),
    .A(_08689_),
    .B(_08757_));
 sg13g2_nor2_1 _14287_ (.A(net148),
    .B(_08758_),
    .Y(_00007_));
 sg13g2_nand2_1 _14288_ (.Y(_08759_),
    .A(_08689_),
    .B(_08757_));
 sg13g2_xor2_1 _14289_ (.B(_08759_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .X(_08760_));
 sg13g2_nor2_1 _14290_ (.A(net148),
    .B(_08760_),
    .Y(_00008_));
 sg13g2_and3_1 _14291_ (.X(_08761_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ),
    .B(_08689_),
    .C(_08757_));
 sg13g2_buf_8 _14292_ (.A(_08761_),
    .X(_08762_));
 sg13g2_xnor2_1 _14293_ (.Y(_08763_),
    .A(_08675_),
    .B(_08762_));
 sg13g2_nor2_1 _14294_ (.A(net148),
    .B(_08763_),
    .Y(_00009_));
 sg13g2_nand2_1 _14295_ (.Y(_08764_),
    .A(_08675_),
    .B(_08762_));
 sg13g2_xor2_1 _14296_ (.B(_08764_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ),
    .X(_08765_));
 sg13g2_nor2_1 _14297_ (.A(_08753_),
    .B(_08765_),
    .Y(_00010_));
 sg13g2_and2_1 _14298_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ),
    .B(_08675_),
    .X(_08766_));
 sg13g2_buf_1 _14299_ (.A(_08766_),
    .X(_08767_));
 sg13g2_nand2_1 _14300_ (.Y(_08768_),
    .A(_08762_),
    .B(_08767_));
 sg13g2_xor2_1 _14301_ (.B(_08768_),
    .A(_08674_),
    .X(_08769_));
 sg13g2_nor2_1 _14302_ (.A(net148),
    .B(_08769_),
    .Y(_00011_));
 sg13g2_nand3_1 _14303_ (.B(_08762_),
    .C(_08767_),
    .A(_08674_),
    .Y(_08770_));
 sg13g2_xor2_1 _14304_ (.B(_08770_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .X(_08771_));
 sg13g2_nor2_1 _14305_ (.A(net148),
    .B(_08771_),
    .Y(_00012_));
 sg13g2_inv_1 _14306_ (.Y(_08772_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ));
 sg13g2_nand4_1 _14307_ (.B(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ),
    .C(_08762_),
    .A(_08674_),
    .Y(_08773_),
    .D(_08767_));
 sg13g2_xnor2_1 _14308_ (.Y(_08774_),
    .A(_08772_),
    .B(_08773_));
 sg13g2_nor2_1 _14309_ (.A(net148),
    .B(_08774_),
    .Y(_00013_));
 sg13g2_nor2_1 _14310_ (.A(_08772_),
    .B(_08773_),
    .Y(_08775_));
 sg13g2_buf_8 _14311_ (.A(_08775_),
    .X(_08776_));
 sg13g2_xnor2_1 _14312_ (.Y(_08777_),
    .A(_08679_),
    .B(_08776_));
 sg13g2_nor2_1 _14313_ (.A(net148),
    .B(_08777_),
    .Y(_00014_));
 sg13g2_nand2_1 _14314_ (.Y(_08778_),
    .A(_08679_),
    .B(_08776_));
 sg13g2_xor2_1 _14315_ (.B(_08778_),
    .A(_08678_),
    .X(_08779_));
 sg13g2_nor2_1 _14316_ (.A(_08753_),
    .B(_08779_),
    .Y(_00015_));
 sg13g2_buf_1 _14317_ (.A(_08731_),
    .X(_08780_));
 sg13g2_nand3_1 _14318_ (.B(_08679_),
    .C(_08776_),
    .A(_08678_),
    .Y(_08781_));
 sg13g2_xor2_1 _14319_ (.B(_08781_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ),
    .X(_08782_));
 sg13g2_nor2_1 _14320_ (.A(net147),
    .B(_08782_),
    .Y(_00017_));
 sg13g2_and3_1 _14321_ (.X(_08783_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ),
    .B(_08678_),
    .C(_08679_));
 sg13g2_buf_1 _14322_ (.A(_08783_),
    .X(_08784_));
 sg13g2_nand2_1 _14323_ (.Y(_08785_),
    .A(_08776_),
    .B(_08784_));
 sg13g2_xor2_1 _14324_ (.B(_08785_),
    .A(_08677_),
    .X(_08786_));
 sg13g2_nor2_1 _14325_ (.A(net147),
    .B(_08786_),
    .Y(_00018_));
 sg13g2_nand3_1 _14326_ (.B(_08776_),
    .C(_08784_),
    .A(_08677_),
    .Y(_08787_));
 sg13g2_xor2_1 _14327_ (.B(_08787_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .X(_08788_));
 sg13g2_nor2_1 _14328_ (.A(net147),
    .B(_08788_),
    .Y(_00019_));
 sg13g2_and4_1 _14329_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ),
    .B(_08677_),
    .C(_08776_),
    .D(_08784_),
    .X(_08789_));
 sg13g2_buf_8 _14330_ (.A(_08789_),
    .X(_08790_));
 sg13g2_xnor2_1 _14331_ (.Y(_08791_),
    .A(_08682_),
    .B(_08790_));
 sg13g2_nor2_1 _14332_ (.A(net147),
    .B(_08791_),
    .Y(_00020_));
 sg13g2_nand2_1 _14333_ (.Y(_08792_),
    .A(_08682_),
    .B(_08790_));
 sg13g2_xor2_1 _14334_ (.B(_08792_),
    .A(_08684_),
    .X(_08793_));
 sg13g2_nor2_1 _14335_ (.A(net147),
    .B(_08793_),
    .Y(_00021_));
 sg13g2_nand3_1 _14336_ (.B(_08682_),
    .C(_08790_),
    .A(_08684_),
    .Y(_08794_));
 sg13g2_xor2_1 _14337_ (.B(_08794_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ),
    .X(_08795_));
 sg13g2_nor2_1 _14338_ (.A(_08780_),
    .B(_08795_),
    .Y(_00022_));
 sg13g2_and4_1 _14339_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ),
    .B(_08684_),
    .C(_08682_),
    .D(_08790_),
    .X(_08796_));
 sg13g2_xnor2_1 _14340_ (.Y(_08797_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .B(_08796_));
 sg13g2_nor2_1 _14341_ (.A(_08780_),
    .B(_08797_),
    .Y(_00023_));
 sg13g2_and2_1 _14342_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ),
    .B(_08796_),
    .X(_08798_));
 sg13g2_buf_8 _14343_ (.A(_08798_),
    .X(_08799_));
 sg13g2_xnor2_1 _14344_ (.Y(_08800_),
    .A(_08681_),
    .B(_08799_));
 sg13g2_nor2_1 _14345_ (.A(net147),
    .B(_08800_),
    .Y(_00024_));
 sg13g2_nand2_1 _14346_ (.Y(_08801_),
    .A(_08681_),
    .B(_08799_));
 sg13g2_xor2_1 _14347_ (.B(_08801_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .X(_08802_));
 sg13g2_nor2_1 _14348_ (.A(net147),
    .B(_08802_),
    .Y(_00025_));
 sg13g2_and2_1 _14349_ (.A(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ),
    .B(_08681_),
    .X(_08803_));
 sg13g2_buf_1 _14350_ (.A(_08803_),
    .X(_08804_));
 sg13g2_nand2_1 _14351_ (.Y(_08805_),
    .A(_08799_),
    .B(_08804_));
 sg13g2_xor2_1 _14352_ (.B(_08805_),
    .A(_08687_),
    .X(_08806_));
 sg13g2_nor2_1 _14353_ (.A(net147),
    .B(_08806_),
    .Y(_00026_));
 sg13g2_nand3_1 _14354_ (.B(_08799_),
    .C(_08804_),
    .A(_08687_),
    .Y(_08807_));
 sg13g2_xor2_1 _14355_ (.B(_08807_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .X(_08808_));
 sg13g2_nor2_1 _14356_ (.A(_08731_),
    .B(_08808_),
    .Y(_00028_));
 sg13g2_nand4_1 _14357_ (.B(_08687_),
    .C(_08799_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ),
    .Y(_08809_),
    .D(_08804_));
 sg13g2_xor2_1 _14358_ (.B(_08809_),
    .A(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ),
    .X(_08810_));
 sg13g2_nor2_1 _14359_ (.A(_08731_),
    .B(_08810_),
    .Y(_00029_));
 sg13g2_nand3_1 _14360_ (.B(_08609_),
    .C(_08662_),
    .A(net831),
    .Y(_08811_));
 sg13g2_nand3_1 _14361_ (.B(_08662_),
    .C(_08665_),
    .A(net795),
    .Y(_08812_));
 sg13g2_o21ai_1 _14362_ (.B1(_08812_),
    .Y(_08813_),
    .A1(_08655_),
    .A2(_08811_));
 sg13g2_buf_1 _14363_ (.A(\top_ihp.wb_uart.uart_tx.state[1] ),
    .X(_08814_));
 sg13g2_buf_1 _14364_ (.A(\top_ihp.wb_uart.uart_tx.state[0] ),
    .X(_08815_));
 sg13g2_nor2_2 _14365_ (.A(_08814_),
    .B(_08815_),
    .Y(_08816_));
 sg13g2_nor2b_1 _14366_ (.A(_08813_),
    .B_N(_08816_),
    .Y(_08817_));
 sg13g2_buf_2 _14367_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ),
    .X(_08818_));
 sg13g2_buf_2 _14368_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ),
    .X(_08819_));
 sg13g2_buf_1 _14369_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ),
    .X(_08820_));
 sg13g2_buf_1 _14370_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ),
    .X(_08821_));
 sg13g2_buf_1 _14371_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ),
    .X(_08822_));
 sg13g2_nor4_1 _14372_ (.A(_08820_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .C(_08821_),
    .D(_08822_),
    .Y(_08823_));
 sg13g2_buf_1 _14373_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ),
    .X(_08824_));
 sg13g2_buf_1 _14374_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ),
    .X(_08825_));
 sg13g2_nor4_1 _14375_ (.A(_08824_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .D(_08825_),
    .Y(_08826_));
 sg13g2_buf_1 _14376_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ),
    .X(_08827_));
 sg13g2_nor4_1 _14377_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ),
    .C(_08827_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .Y(_08828_));
 sg13g2_buf_8 _14378_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ),
    .X(_08829_));
 sg13g2_buf_8 _14379_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ),
    .X(_08830_));
 sg13g2_inv_1 _14380_ (.Y(_08831_),
    .A(_08830_));
 sg13g2_buf_1 _14381_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ),
    .X(_08832_));
 sg13g2_nor4_1 _14382_ (.A(_08829_),
    .B(_08831_),
    .C(_08832_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .Y(_08833_));
 sg13g2_nand4_1 _14383_ (.B(_08826_),
    .C(_08828_),
    .A(_08823_),
    .Y(_08834_),
    .D(_08833_));
 sg13g2_buf_1 _14384_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ),
    .X(_08835_));
 sg13g2_inv_1 _14385_ (.Y(_08836_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_nor4_1 _14386_ (.A(_08835_),
    .B(_08836_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ),
    .Y(_08837_));
 sg13g2_buf_1 _14387_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ),
    .X(_08838_));
 sg13g2_inv_1 _14388_ (.Y(_08839_),
    .A(_08838_));
 sg13g2_nor4_1 _14389_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .D(_08839_),
    .Y(_08840_));
 sg13g2_buf_1 _14390_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ),
    .X(_08841_));
 sg13g2_buf_1 _14391_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ),
    .X(_08842_));
 sg13g2_nor4_1 _14392_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ),
    .B(_08841_),
    .C(_08842_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ),
    .Y(_08843_));
 sg13g2_buf_2 _14393_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ),
    .X(_08844_));
 sg13g2_nand2_1 _14394_ (.Y(_08845_),
    .A(_08844_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_nor3_1 _14395_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ),
    .C(_08845_),
    .Y(_08846_));
 sg13g2_nand4_1 _14396_ (.B(_08840_),
    .C(_08843_),
    .A(_08837_),
    .Y(_08847_),
    .D(_08846_));
 sg13g2_nor2_1 _14397_ (.A(_08834_),
    .B(_08847_),
    .Y(_08848_));
 sg13g2_buf_1 _14398_ (.A(_08848_),
    .X(_08849_));
 sg13g2_nand4_1 _14399_ (.B(_08819_),
    .C(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .A(_08818_),
    .Y(_08850_),
    .D(_08849_));
 sg13g2_nor2_1 _14400_ (.A(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .B(_08850_),
    .Y(_08851_));
 sg13g2_nand2b_1 _14401_ (.Y(_08852_),
    .B(_08814_),
    .A_N(_08815_));
 sg13g2_buf_1 _14402_ (.A(_08852_),
    .X(_08853_));
 sg13g2_nand2_1 _14403_ (.Y(_08854_),
    .A(_08815_),
    .B(_08849_));
 sg13g2_o21ai_1 _14404_ (.B1(_08854_),
    .Y(_08855_),
    .A1(_08851_),
    .A2(_08853_));
 sg13g2_nor2_1 _14405_ (.A(_08817_),
    .B(_08855_),
    .Y(\top_ihp.wb_uart.uart_tx.next_state[0] ));
 sg13g2_xnor2_1 _14406_ (.Y(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .A(_08814_),
    .B(_08854_));
 sg13g2_nand4_1 _14407_ (.B(_08609_),
    .C(_08662_),
    .A(net831),
    .Y(_08856_),
    .D(_08816_));
 sg13g2_nand4_1 _14408_ (.B(_08662_),
    .C(_08665_),
    .A(net831),
    .Y(_08857_),
    .D(_08816_));
 sg13g2_o21ai_1 _14409_ (.B1(_08857_),
    .Y(_08858_),
    .A1(_08655_),
    .A2(_08856_));
 sg13g2_buf_1 _14410_ (.A(_08858_),
    .X(_08859_));
 sg13g2_nand2b_1 _14411_ (.Y(_08860_),
    .B(_08849_),
    .A_N(_08816_));
 sg13g2_nand2b_1 _14412_ (.Y(_08861_),
    .B(_08860_),
    .A_N(net593));
 sg13g2_buf_2 _14413_ (.A(_08861_),
    .X(_08862_));
 sg13g2_buf_1 _14414_ (.A(_08862_),
    .X(_08863_));
 sg13g2_nor2_1 _14415_ (.A(_08829_),
    .B(net146),
    .Y(_00037_));
 sg13g2_xnor2_1 _14416_ (.Y(_08864_),
    .A(_08829_),
    .B(_08830_));
 sg13g2_nor2_1 _14417_ (.A(net146),
    .B(_08864_),
    .Y(_00048_));
 sg13g2_nand2_1 _14418_ (.Y(_08865_),
    .A(_08829_),
    .B(_08830_));
 sg13g2_xor2_1 _14419_ (.B(_08865_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ),
    .X(_08866_));
 sg13g2_nor2_1 _14420_ (.A(net146),
    .B(_08866_),
    .Y(_00059_));
 sg13g2_and3_1 _14421_ (.X(_08867_),
    .A(_08829_),
    .B(_08830_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ));
 sg13g2_buf_1 _14422_ (.A(_08867_),
    .X(_08868_));
 sg13g2_xnor2_1 _14423_ (.Y(_08869_),
    .A(_08844_),
    .B(_08868_));
 sg13g2_nor2_1 _14424_ (.A(net146),
    .B(_08869_),
    .Y(_00062_));
 sg13g2_nand2_1 _14425_ (.Y(_08870_),
    .A(_08844_),
    .B(_08868_));
 sg13g2_xor2_1 _14426_ (.B(_08870_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ),
    .X(_08871_));
 sg13g2_nor2_1 _14427_ (.A(_08863_),
    .B(_08871_),
    .Y(_00063_));
 sg13g2_nand2b_1 _14428_ (.Y(_08872_),
    .B(_08868_),
    .A_N(_08845_));
 sg13g2_xor2_1 _14429_ (.B(_08872_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .X(_08873_));
 sg13g2_nor2_1 _14430_ (.A(_08863_),
    .B(_08873_),
    .Y(_00064_));
 sg13g2_and3_1 _14431_ (.X(_08874_),
    .A(_08844_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_and2_1 _14432_ (.A(_08868_),
    .B(_08874_),
    .X(_08875_));
 sg13g2_xnor2_1 _14433_ (.Y(_08876_),
    .A(_08838_),
    .B(_08875_));
 sg13g2_nor2_1 _14434_ (.A(net146),
    .B(_08876_),
    .Y(_00065_));
 sg13g2_nand2_1 _14435_ (.Y(_08877_),
    .A(_08838_),
    .B(_08875_));
 sg13g2_xor2_1 _14436_ (.B(_08877_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .X(_08878_));
 sg13g2_nor2_1 _14437_ (.A(net146),
    .B(_08878_),
    .Y(_00066_));
 sg13g2_and4_1 _14438_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ),
    .B(_08838_),
    .C(_08868_),
    .D(_08874_),
    .X(_08879_));
 sg13g2_xnor2_1 _14439_ (.Y(_08880_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ),
    .B(_08879_));
 sg13g2_nor2_1 _14440_ (.A(net146),
    .B(_08880_),
    .Y(_00067_));
 sg13g2_and2_1 _14441_ (.A(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ),
    .B(_08879_),
    .X(_08881_));
 sg13g2_buf_1 _14442_ (.A(_08881_),
    .X(_08882_));
 sg13g2_xnor2_1 _14443_ (.Y(_08883_),
    .A(_08835_),
    .B(_08882_));
 sg13g2_nor2_1 _14444_ (.A(net146),
    .B(_08883_),
    .Y(_00068_));
 sg13g2_buf_1 _14445_ (.A(_08862_),
    .X(_08884_));
 sg13g2_nand2_1 _14446_ (.Y(_08885_),
    .A(_08835_),
    .B(_08882_));
 sg13g2_xor2_1 _14447_ (.B(_08885_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .X(_08886_));
 sg13g2_nor2_1 _14448_ (.A(net145),
    .B(_08886_),
    .Y(_00038_));
 sg13g2_inv_1 _14449_ (.Y(_08887_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ));
 sg13g2_nand3_1 _14450_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ),
    .C(_08882_),
    .A(_08835_),
    .Y(_08888_));
 sg13g2_buf_1 _14451_ (.A(_08888_),
    .X(_08889_));
 sg13g2_xnor2_1 _14452_ (.Y(_08890_),
    .A(_08887_),
    .B(_08889_));
 sg13g2_nor2_1 _14453_ (.A(net145),
    .B(_08890_),
    .Y(_00039_));
 sg13g2_nor2_1 _14454_ (.A(_08887_),
    .B(_08889_),
    .Y(_08891_));
 sg13g2_xnor2_1 _14455_ (.Y(_08892_),
    .A(_08841_),
    .B(_08891_));
 sg13g2_nor2_1 _14456_ (.A(net145),
    .B(_08892_),
    .Y(_00040_));
 sg13g2_inv_1 _14457_ (.Y(_08893_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ));
 sg13g2_nand2_1 _14458_ (.Y(_08894_),
    .A(_08841_),
    .B(_08891_));
 sg13g2_xnor2_1 _14459_ (.Y(_08895_),
    .A(_08893_),
    .B(_08894_));
 sg13g2_nor2_1 _14460_ (.A(net145),
    .B(_08895_),
    .Y(_00041_));
 sg13g2_inv_1 _14461_ (.Y(_08896_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ));
 sg13g2_inv_1 _14462_ (.Y(_08897_),
    .A(_08841_));
 sg13g2_or4_1 _14463_ (.A(_08887_),
    .B(_08893_),
    .C(_08897_),
    .D(_08889_),
    .X(_08898_));
 sg13g2_buf_1 _14464_ (.A(_08898_),
    .X(_08899_));
 sg13g2_xnor2_1 _14465_ (.Y(_08900_),
    .A(_08896_),
    .B(_08899_));
 sg13g2_nor2_1 _14466_ (.A(net145),
    .B(_08900_),
    .Y(_00042_));
 sg13g2_nor2_1 _14467_ (.A(_08896_),
    .B(_08899_),
    .Y(_08901_));
 sg13g2_xnor2_1 _14468_ (.Y(_08902_),
    .A(_08842_),
    .B(_08901_));
 sg13g2_nor2_1 _14469_ (.A(net145),
    .B(_08902_),
    .Y(_00043_));
 sg13g2_nand2_1 _14470_ (.Y(_08903_),
    .A(_08842_),
    .B(_08901_));
 sg13g2_xor2_1 _14471_ (.B(_08903_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ),
    .X(_08904_));
 sg13g2_nor2_1 _14472_ (.A(net145),
    .B(_08904_),
    .Y(_00044_));
 sg13g2_inv_1 _14473_ (.Y(_08905_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ));
 sg13g2_nand3_1 _14474_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ),
    .C(_08901_),
    .A(_08842_),
    .Y(_08906_));
 sg13g2_xnor2_1 _14475_ (.Y(_08907_),
    .A(_08905_),
    .B(_08906_));
 sg13g2_nor2_1 _14476_ (.A(net145),
    .B(_08907_),
    .Y(_00045_));
 sg13g2_nor2_2 _14477_ (.A(_08905_),
    .B(_08906_),
    .Y(_08908_));
 sg13g2_xnor2_1 _14478_ (.Y(_08909_),
    .A(_08824_),
    .B(_08908_));
 sg13g2_nor2_1 _14479_ (.A(_08884_),
    .B(_08909_),
    .Y(_00046_));
 sg13g2_nand2_1 _14480_ (.Y(_08910_),
    .A(_08824_),
    .B(_08908_));
 sg13g2_xor2_1 _14481_ (.B(_08910_),
    .A(_08820_),
    .X(_08911_));
 sg13g2_nor2_1 _14482_ (.A(_08884_),
    .B(_08911_),
    .Y(_00047_));
 sg13g2_buf_1 _14483_ (.A(_08862_),
    .X(_08912_));
 sg13g2_nand3_1 _14484_ (.B(_08824_),
    .C(_08908_),
    .A(_08820_),
    .Y(_08913_));
 sg13g2_xor2_1 _14485_ (.B(_08913_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .X(_08914_));
 sg13g2_nor2_1 _14486_ (.A(_08912_),
    .B(_08914_),
    .Y(_00049_));
 sg13g2_inv_1 _14487_ (.Y(_08915_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ));
 sg13g2_nand4_1 _14488_ (.B(_08824_),
    .C(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ),
    .A(_08820_),
    .Y(_08916_),
    .D(_08908_));
 sg13g2_buf_2 _14489_ (.A(_08916_),
    .X(_08917_));
 sg13g2_xnor2_1 _14490_ (.Y(_08918_),
    .A(_08915_),
    .B(_08917_));
 sg13g2_nor2_1 _14491_ (.A(net144),
    .B(_08918_),
    .Y(_00050_));
 sg13g2_nor2_1 _14492_ (.A(_08915_),
    .B(_08917_),
    .Y(_08919_));
 sg13g2_xnor2_1 _14493_ (.Y(_08920_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ),
    .B(_08919_));
 sg13g2_nor2_1 _14494_ (.A(net144),
    .B(_08920_),
    .Y(_00051_));
 sg13g2_nand2_1 _14495_ (.Y(_08921_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ));
 sg13g2_nor2_2 _14496_ (.A(_08917_),
    .B(_08921_),
    .Y(_08922_));
 sg13g2_xnor2_1 _14497_ (.Y(_08923_),
    .A(_08825_),
    .B(_08922_));
 sg13g2_nor2_1 _14498_ (.A(net144),
    .B(_08923_),
    .Y(_00052_));
 sg13g2_nand2_1 _14499_ (.Y(_08924_),
    .A(_08825_),
    .B(_08922_));
 sg13g2_xor2_1 _14500_ (.B(_08924_),
    .A(_08832_),
    .X(_08925_));
 sg13g2_nor2_1 _14501_ (.A(net144),
    .B(_08925_),
    .Y(_00053_));
 sg13g2_nand3_1 _14502_ (.B(_08832_),
    .C(_08922_),
    .A(_08825_),
    .Y(_08926_));
 sg13g2_xor2_1 _14503_ (.B(_08926_),
    .A(_08821_),
    .X(_08927_));
 sg13g2_nor2_1 _14504_ (.A(net144),
    .B(_08927_),
    .Y(_00054_));
 sg13g2_nand4_1 _14505_ (.B(_08821_),
    .C(_08832_),
    .A(_08825_),
    .Y(_08928_),
    .D(_08922_));
 sg13g2_xor2_1 _14506_ (.B(_08928_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ),
    .X(_08929_));
 sg13g2_nor2_1 _14507_ (.A(net144),
    .B(_08929_),
    .Y(_00055_));
 sg13g2_nand4_1 _14508_ (.B(_08821_),
    .C(_08832_),
    .A(_08825_),
    .Y(_08930_),
    .D(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ));
 sg13g2_nor3_2 _14509_ (.A(_08917_),
    .B(_08921_),
    .C(_08930_),
    .Y(_08931_));
 sg13g2_xnor2_1 _14510_ (.Y(_08932_),
    .A(_08822_),
    .B(_08931_));
 sg13g2_nor2_1 _14511_ (.A(net144),
    .B(_08932_),
    .Y(_00056_));
 sg13g2_nand2_1 _14512_ (.Y(_08933_),
    .A(_08822_),
    .B(_08931_));
 sg13g2_xor2_1 _14513_ (.B(_08933_),
    .A(_08827_),
    .X(_08934_));
 sg13g2_nor2_1 _14514_ (.A(_08912_),
    .B(_08934_),
    .Y(_00057_));
 sg13g2_nand3_1 _14515_ (.B(_08827_),
    .C(_08931_),
    .A(_08822_),
    .Y(_08935_));
 sg13g2_xor2_1 _14516_ (.B(_08935_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ),
    .X(_08936_));
 sg13g2_nor2_1 _14517_ (.A(net144),
    .B(_08936_),
    .Y(_00058_));
 sg13g2_and2_1 _14518_ (.A(_08822_),
    .B(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ),
    .X(_08937_));
 sg13g2_nand3_1 _14519_ (.B(_08931_),
    .C(_08937_),
    .A(_08827_),
    .Y(_08938_));
 sg13g2_xor2_1 _14520_ (.B(_08938_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .X(_08939_));
 sg13g2_nor2_1 _14521_ (.A(_08862_),
    .B(_08939_),
    .Y(_00060_));
 sg13g2_nand4_1 _14522_ (.B(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ),
    .C(_08931_),
    .A(_08827_),
    .Y(_08940_),
    .D(_08937_));
 sg13g2_xor2_1 _14523_ (.B(_08940_),
    .A(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ),
    .X(_08941_));
 sg13g2_nor2_1 _14524_ (.A(_08862_),
    .B(_08941_),
    .Y(_00061_));
 sg13g2_buf_1 _14525_ (.A(\top_ihp.wb_imem.state[1] ),
    .X(_08942_));
 sg13g2_nand3_1 _14526_ (.B(_08584_),
    .C(_08592_),
    .A(net1024),
    .Y(_08943_));
 sg13g2_buf_2 _14527_ (.A(_08943_),
    .X(_08944_));
 sg13g2_buf_8 _14528_ (.A(_08944_),
    .X(_08945_));
 sg13g2_nor2_1 _14529_ (.A(_00117_),
    .B(net861),
    .Y(_08946_));
 sg13g2_buf_1 _14530_ (.A(\top_ihp.wb_emem.last_bit ),
    .X(_08947_));
 sg13g2_buf_2 _14531_ (.A(\top_ihp.wb_emem.state[2] ),
    .X(_08948_));
 sg13g2_buf_1 _14532_ (.A(\top_ihp.wb_emem.state[3] ),
    .X(_08949_));
 sg13g2_nor2_1 _14533_ (.A(_08948_),
    .B(net1023),
    .Y(_08950_));
 sg13g2_buf_1 _14534_ (.A(_08950_),
    .X(_08951_));
 sg13g2_buf_1 _14535_ (.A(\top_ihp.wb_emem.state[0] ),
    .X(_08952_));
 sg13g2_buf_2 _14536_ (.A(\top_ihp.wb_emem.state[1] ),
    .X(_08953_));
 sg13g2_and2_1 _14537_ (.A(net1022),
    .B(_08953_),
    .X(_08954_));
 sg13g2_buf_1 _14538_ (.A(_08954_),
    .X(_08955_));
 sg13g2_nand3_1 _14539_ (.B(_08951_),
    .C(_08955_),
    .A(_08947_),
    .Y(_08956_));
 sg13g2_buf_2 _14540_ (.A(_08956_),
    .X(_08957_));
 sg13g2_buf_8 _14541_ (.A(_08957_),
    .X(_08958_));
 sg13g2_buf_2 _14542_ (.A(\top_ihp.wb_ack_spi ),
    .X(_08959_));
 sg13g2_inv_1 _14543_ (.Y(_08960_),
    .A(_00119_));
 sg13g2_nor2b_1 _14544_ (.A(_08959_),
    .B_N(_08598_),
    .Y(_08961_));
 sg13g2_buf_2 _14545_ (.A(_08961_),
    .X(_08962_));
 sg13g2_a22oi_1 _14546_ (.Y(_08963_),
    .B1(_08962_),
    .B2(\top_ihp.wb_coproc.dat_o[15] ),
    .A2(_08960_),
    .A1(_08959_));
 sg13g2_buf_1 _14547_ (.A(_08947_),
    .X(_08964_));
 sg13g2_buf_1 _14548_ (.A(_08955_),
    .X(_08965_));
 sg13g2_and4_1 _14549_ (.A(net1021),
    .B(_00118_),
    .C(_08951_),
    .D(net891),
    .X(_08966_));
 sg13g2_a221oi_1 _14550_ (.B2(_08963_),
    .C1(_08966_),
    .B1(net846),
    .A1(net1024),
    .Y(_08967_),
    .A2(_08594_));
 sg13g2_buf_1 _14551_ (.A(\top_ihp.wb_ack_gpio ),
    .X(_08968_));
 sg13g2_nor2b_1 _14552_ (.A(_08968_),
    .B_N(_00080_),
    .Y(_08969_));
 sg13g2_buf_2 _14553_ (.A(_08969_),
    .X(_08970_));
 sg13g2_o21ai_1 _14554_ (.B1(_08970_),
    .Y(_08971_),
    .A1(_08946_),
    .A2(_08967_));
 sg13g2_buf_2 _14555_ (.A(_08971_),
    .X(_08972_));
 sg13g2_buf_1 _14556_ (.A(\top_ihp.wb_ack_uart ),
    .X(_08973_));
 sg13g2_nor2_1 _14557_ (.A(_08968_),
    .B(_08973_),
    .Y(_08974_));
 sg13g2_buf_2 _14558_ (.A(_08974_),
    .X(_08975_));
 sg13g2_nor2_1 _14559_ (.A(_08598_),
    .B(_08959_),
    .Y(_08976_));
 sg13g2_nand4_1 _14560_ (.B(_08957_),
    .C(_08975_),
    .A(_08944_),
    .Y(_08977_),
    .D(_08976_));
 sg13g2_buf_1 _14561_ (.A(_08977_),
    .X(_08978_));
 sg13g2_nand2_1 _14562_ (.Y(_08979_),
    .A(_08412_),
    .B(_08978_));
 sg13g2_buf_1 _14563_ (.A(_08979_),
    .X(_08980_));
 sg13g2_buf_1 _14564_ (.A(net763),
    .X(_08981_));
 sg13g2_buf_1 _14565_ (.A(net763),
    .X(_08982_));
 sg13g2_nand2_1 _14566_ (.Y(_08983_),
    .A(\top_ihp.oisc.decoder.instruction[15] ),
    .B(_08982_));
 sg13g2_o21ai_1 _14567_ (.B1(_08983_),
    .Y(_00241_),
    .A1(_08972_),
    .A2(net751));
 sg13g2_buf_1 _14568_ (.A(\top_ihp.oisc.micro_op[9] ),
    .X(_08984_));
 sg13g2_buf_2 _14569_ (.A(_08984_),
    .X(_08985_));
 sg13g2_and2_1 _14570_ (.A(\top_ihp.oisc.micro_state[1] ),
    .B(_08199_),
    .X(_08986_));
 sg13g2_buf_2 _14571_ (.A(_08986_),
    .X(_08987_));
 sg13g2_and2_1 _14572_ (.A(net1020),
    .B(_08987_),
    .X(\top_ihp.oisc.reg_rb[1] ));
 sg13g2_buf_1 _14573_ (.A(\top_ihp.oisc.micro_op[8] ),
    .X(_08988_));
 sg13g2_nand2_2 _14574_ (.Y(_08989_),
    .A(_08988_),
    .B(_08987_));
 sg13g2_inv_2 _14575_ (.Y(\top_ihp.oisc.reg_rb[0] ),
    .A(_08989_));
 sg13g2_inv_1 _14576_ (.Y(_08990_),
    .A(\top_ihp.oisc.micro_op[11] ));
 sg13g2_nand2_2 _14577_ (.Y(_08991_),
    .A(\top_ihp.oisc.micro_state[1] ),
    .B(_08199_));
 sg13g2_nor2_1 _14578_ (.A(_08990_),
    .B(_08991_),
    .Y(_08992_));
 sg13g2_buf_2 _14579_ (.A(_08992_),
    .X(\top_ihp.oisc.reg_rb[3] ));
 sg13g2_buf_2 _14580_ (.A(\top_ihp.oisc.micro_op[10] ),
    .X(_08993_));
 sg13g2_nand4_1 _14581_ (.B(_08203_),
    .C(_08204_),
    .A(_08202_),
    .Y(_08994_),
    .D(_08208_));
 sg13g2_buf_1 _14582_ (.A(_08994_),
    .X(_08995_));
 sg13g2_nor2_1 _14583_ (.A(_08995_),
    .B(_08987_),
    .Y(_08996_));
 sg13g2_a21oi_2 _14584_ (.B1(_08996_),
    .Y(_08997_),
    .A2(_08987_),
    .A1(net1041));
 sg13g2_inv_1 _14585_ (.Y(_08998_),
    .A(_08997_));
 sg13g2_buf_1 _14586_ (.A(_08998_),
    .X(_08999_));
 sg13g2_buf_1 _14587_ (.A(net830),
    .X(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_buf_1 _14588_ (.A(_08615_),
    .X(_09000_));
 sg13g2_buf_2 _14589_ (.A(\top_ihp.oisc.state[6] ),
    .X(_09001_));
 sg13g2_inv_1 _14590_ (.Y(_09002_),
    .A(_09001_));
 sg13g2_buf_8 _14591_ (.A(_08978_),
    .X(_09003_));
 sg13g2_a21oi_1 _14592_ (.A1(net982),
    .A2(_09002_),
    .Y(_09004_),
    .B1(_09003_));
 sg13g2_or2_1 _14593_ (.X(_09005_),
    .B(_00093_),
    .A(net1032));
 sg13g2_buf_1 _14594_ (.A(_08995_),
    .X(_09006_));
 sg13g2_nand2_1 _14595_ (.Y(_09007_),
    .A(net1032),
    .B(net890));
 sg13g2_o21ai_1 _14596_ (.B1(_09007_),
    .Y(_00002_),
    .A1(_09004_),
    .A2(_09005_));
 sg13g2_xor2_1 _14597_ (.B(\top_ihp.wb_spi.spi_clk_cnt[0] ),
    .A(\top_ihp.spi_clk_o ),
    .X(_00266_));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_nand2_2 _14599_ (.Y(_09008_),
    .A(net1032),
    .B(\top_ihp.oisc.micro_state[0] ));
 sg13g2_and2_1 _14600_ (.A(net890),
    .B(_09008_),
    .X(_09009_));
 sg13g2_buf_1 _14601_ (.A(_09009_),
    .X(_09010_));
 sg13g2_buf_1 _14602_ (.A(_09010_),
    .X(_09011_));
 sg13g2_buf_2 _14603_ (.A(\top_ihp.oisc.micro_pc[7] ),
    .X(_09012_));
 sg13g2_buf_1 _14604_ (.A(_09012_),
    .X(_09013_));
 sg13g2_buf_1 _14605_ (.A(net1019),
    .X(_09014_));
 sg13g2_buf_1 _14606_ (.A(\top_ihp.oisc.micro_pc[5] ),
    .X(_09015_));
 sg13g2_inv_1 _14607_ (.Y(_09016_),
    .A(net1040));
 sg13g2_buf_1 _14608_ (.A(_09016_),
    .X(_09017_));
 sg13g2_buf_1 _14609_ (.A(net980),
    .X(_09018_));
 sg13g2_buf_1 _14610_ (.A(\top_ihp.oisc.micro_pc[6] ),
    .X(_09019_));
 sg13g2_buf_1 _14611_ (.A(net1039),
    .X(_09020_));
 sg13g2_buf_1 _14612_ (.A(\top_ihp.oisc.micro_pc[3] ),
    .X(_09021_));
 sg13g2_buf_1 _14613_ (.A(_09021_),
    .X(_09022_));
 sg13g2_buf_1 _14614_ (.A(net1017),
    .X(_09023_));
 sg13g2_buf_1 _14615_ (.A(net979),
    .X(_09024_));
 sg13g2_buf_1 _14616_ (.A(net932),
    .X(_09025_));
 sg13g2_buf_1 _14617_ (.A(\top_ihp.oisc.micro_pc[0] ),
    .X(_09026_));
 sg13g2_buf_1 _14618_ (.A(_09026_),
    .X(_09027_));
 sg13g2_buf_1 _14619_ (.A(\top_ihp.oisc.micro_pc[2] ),
    .X(_09028_));
 sg13g2_nor2_1 _14620_ (.A(net1016),
    .B(net1038),
    .Y(_09029_));
 sg13g2_buf_1 _14621_ (.A(_09029_),
    .X(_09030_));
 sg13g2_buf_1 _14622_ (.A(\top_ihp.oisc.micro_pc[1] ),
    .X(_09031_));
 sg13g2_inv_2 _14623_ (.Y(_09032_),
    .A(_09031_));
 sg13g2_buf_1 _14624_ (.A(_09032_),
    .X(_09033_));
 sg13g2_buf_1 _14625_ (.A(\top_ihp.oisc.micro_pc[4] ),
    .X(_09034_));
 sg13g2_buf_1 _14626_ (.A(_09034_),
    .X(_09035_));
 sg13g2_buf_1 _14627_ (.A(net1015),
    .X(_09036_));
 sg13g2_nor2_1 _14628_ (.A(_09033_),
    .B(net977),
    .Y(_09037_));
 sg13g2_buf_1 _14629_ (.A(net1038),
    .X(_09038_));
 sg13g2_buf_1 _14630_ (.A(net1014),
    .X(_09039_));
 sg13g2_inv_1 _14631_ (.Y(_09040_),
    .A(_09026_));
 sg13g2_buf_1 _14632_ (.A(_09040_),
    .X(_09041_));
 sg13g2_nand2_2 _14633_ (.Y(_09042_),
    .A(net975),
    .B(net978));
 sg13g2_nor2_1 _14634_ (.A(_09028_),
    .B(_09032_),
    .Y(_09043_));
 sg13g2_buf_1 _14635_ (.A(_09043_),
    .X(_09044_));
 sg13g2_inv_2 _14636_ (.Y(_09045_),
    .A(net1038));
 sg13g2_buf_1 _14637_ (.A(_09031_),
    .X(_09046_));
 sg13g2_nor2_2 _14638_ (.A(_09045_),
    .B(net1013),
    .Y(_09047_));
 sg13g2_buf_1 _14639_ (.A(net1016),
    .X(_09048_));
 sg13g2_o21ai_1 _14640_ (.B1(_09048_),
    .Y(_09049_),
    .A1(net930),
    .A2(_09047_));
 sg13g2_o21ai_1 _14641_ (.B1(_09049_),
    .Y(_09050_),
    .A1(net976),
    .A2(_09042_));
 sg13g2_buf_1 _14642_ (.A(_09036_),
    .X(_09051_));
 sg13g2_a22oi_1 _14643_ (.Y(_09052_),
    .B1(_09050_),
    .B2(net929),
    .A2(_09037_),
    .A1(net931));
 sg13g2_buf_1 _14644_ (.A(net975),
    .X(_09053_));
 sg13g2_buf_1 _14645_ (.A(net928),
    .X(_09054_));
 sg13g2_inv_1 _14646_ (.Y(_09055_),
    .A(_09021_));
 sg13g2_buf_1 _14647_ (.A(_09055_),
    .X(_09056_));
 sg13g2_inv_2 _14648_ (.Y(_09057_),
    .A(_09034_));
 sg13g2_nor2_1 _14649_ (.A(_09056_),
    .B(_09057_),
    .Y(_09058_));
 sg13g2_buf_1 _14650_ (.A(_09058_),
    .X(_09059_));
 sg13g2_nand3_1 _14651_ (.B(net930),
    .C(net887),
    .A(net888),
    .Y(_09060_));
 sg13g2_o21ai_1 _14652_ (.B1(_09060_),
    .Y(_09061_),
    .A1(net889),
    .A2(_09052_));
 sg13g2_buf_1 _14653_ (.A(net1013),
    .X(_09062_));
 sg13g2_buf_1 _14654_ (.A(net972),
    .X(_09063_));
 sg13g2_buf_1 _14655_ (.A(_09063_),
    .X(_09064_));
 sg13g2_buf_1 _14656_ (.A(_09019_),
    .X(_09065_));
 sg13g2_buf_1 _14657_ (.A(_00217_),
    .X(_09066_));
 sg13g2_buf_1 _14658_ (.A(_09066_),
    .X(_09067_));
 sg13g2_buf_1 _14659_ (.A(_09057_),
    .X(_09068_));
 sg13g2_nor2_2 _14660_ (.A(net1011),
    .B(net971),
    .Y(_09069_));
 sg13g2_inv_2 _14661_ (.Y(_09070_),
    .A(_09066_));
 sg13g2_nor2_1 _14662_ (.A(_09070_),
    .B(net1017),
    .Y(_09071_));
 sg13g2_buf_2 _14663_ (.A(_09071_),
    .X(_09072_));
 sg13g2_nor2_2 _14664_ (.A(_09041_),
    .B(net977),
    .Y(_09073_));
 sg13g2_a22oi_1 _14665_ (.Y(_09074_),
    .B1(_09072_),
    .B2(_09073_),
    .A2(_09069_),
    .A1(net928));
 sg13g2_nor3_1 _14666_ (.A(net886),
    .B(net1012),
    .C(_09074_),
    .Y(_09075_));
 sg13g2_a21o_1 _14667_ (.A2(_09061_),
    .A1(net1018),
    .B1(_09075_),
    .X(_09076_));
 sg13g2_buf_1 _14668_ (.A(net973),
    .X(_09077_));
 sg13g2_buf_1 _14669_ (.A(net1014),
    .X(_09078_));
 sg13g2_nor2_1 _14670_ (.A(_09040_),
    .B(_09032_),
    .Y(_09079_));
 sg13g2_buf_1 _14671_ (.A(_09079_),
    .X(_09080_));
 sg13g2_nand2_1 _14672_ (.Y(_09081_),
    .A(_09078_),
    .B(net925));
 sg13g2_nand2_1 _14673_ (.Y(_09082_),
    .A(net929),
    .B(_09081_));
 sg13g2_buf_1 _14674_ (.A(net1013),
    .X(_09083_));
 sg13g2_nand2_2 _14675_ (.Y(_09084_),
    .A(net969),
    .B(net926));
 sg13g2_nand2_2 _14676_ (.Y(_09085_),
    .A(_09070_),
    .B(net1017));
 sg13g2_inv_1 _14677_ (.Y(_09086_),
    .A(_09085_));
 sg13g2_nand2_1 _14678_ (.Y(_09087_),
    .A(net978),
    .B(_09086_));
 sg13g2_o21ai_1 _14679_ (.B1(_09087_),
    .Y(_09088_),
    .A1(net976),
    .A2(_09084_));
 sg13g2_a221oi_1 _14680_ (.B2(net888),
    .C1(net1012),
    .B1(_09088_),
    .A1(net926),
    .Y(_09089_),
    .A2(_09082_));
 sg13g2_nand2_1 _14681_ (.Y(_09090_),
    .A(_09056_),
    .B(_09057_));
 sg13g2_buf_2 _14682_ (.A(_09090_),
    .X(_09091_));
 sg13g2_buf_1 _14683_ (.A(_09045_),
    .X(_09092_));
 sg13g2_nor2_1 _14684_ (.A(_09027_),
    .B(net968),
    .Y(_09093_));
 sg13g2_buf_2 _14685_ (.A(_09093_),
    .X(_09094_));
 sg13g2_buf_1 _14686_ (.A(net974),
    .X(_09095_));
 sg13g2_buf_1 _14687_ (.A(net1011),
    .X(_09096_));
 sg13g2_nand2_1 _14688_ (.Y(_09097_),
    .A(_09046_),
    .B(_09068_));
 sg13g2_nand2_1 _14689_ (.Y(_09098_),
    .A(net978),
    .B(_09035_));
 sg13g2_nand2_1 _14690_ (.Y(_09099_),
    .A(_09097_),
    .B(_09098_));
 sg13g2_nand3_1 _14691_ (.B(net967),
    .C(_09099_),
    .A(_09095_),
    .Y(_09100_));
 sg13g2_nand3_1 _14692_ (.B(_09091_),
    .C(_09100_),
    .A(net1012),
    .Y(_09101_));
 sg13g2_o21ai_1 _14693_ (.B1(_09101_),
    .Y(_09102_),
    .A1(_09091_),
    .A2(_09094_));
 sg13g2_o21ai_1 _14694_ (.B1(net933),
    .Y(_09103_),
    .A1(_09089_),
    .A2(_09102_));
 sg13g2_o21ai_1 _14695_ (.B1(_09103_),
    .Y(_09104_),
    .A1(net933),
    .A2(_09076_));
 sg13g2_inv_1 _14696_ (.Y(_09105_),
    .A(\top_ihp.oisc.micro_pc[6] ));
 sg13g2_buf_1 _14697_ (.A(_09105_),
    .X(_09106_));
 sg13g2_buf_1 _14698_ (.A(net980),
    .X(_09107_));
 sg13g2_buf_1 _14699_ (.A(_09039_),
    .X(_09108_));
 sg13g2_buf_1 _14700_ (.A(_00216_),
    .X(_09109_));
 sg13g2_nor2_1 _14701_ (.A(_09057_),
    .B(_09109_),
    .Y(_09110_));
 sg13g2_buf_2 _14702_ (.A(_09110_),
    .X(_09111_));
 sg13g2_nor2_1 _14703_ (.A(_09021_),
    .B(_09034_),
    .Y(_09112_));
 sg13g2_buf_1 _14704_ (.A(_09112_),
    .X(_09113_));
 sg13g2_or2_1 _14705_ (.X(_09114_),
    .B(_09111_),
    .A(net966));
 sg13g2_buf_1 _14706_ (.A(_09114_),
    .X(_09115_));
 sg13g2_buf_1 _14707_ (.A(net1016),
    .X(_09116_));
 sg13g2_buf_1 _14708_ (.A(net965),
    .X(_09117_));
 sg13g2_a22oi_1 _14709_ (.Y(_09118_),
    .B1(_09115_),
    .B2(net921),
    .A2(_09111_),
    .A1(net927));
 sg13g2_buf_1 _14710_ (.A(net970),
    .X(_09119_));
 sg13g2_nor2_1 _14711_ (.A(net973),
    .B(_09034_),
    .Y(_09120_));
 sg13g2_buf_2 _14712_ (.A(_09120_),
    .X(_09121_));
 sg13g2_buf_1 _14713_ (.A(_09121_),
    .X(_09122_));
 sg13g2_nand3_1 _14714_ (.B(_09119_),
    .C(_09122_),
    .A(net921),
    .Y(_09123_));
 sg13g2_o21ai_1 _14715_ (.B1(_09123_),
    .Y(_09124_),
    .A1(net922),
    .A2(_09118_));
 sg13g2_nand2_1 _14716_ (.Y(_09125_),
    .A(net923),
    .B(_09124_));
 sg13g2_buf_1 _14717_ (.A(_09015_),
    .X(_09126_));
 sg13g2_buf_1 _14718_ (.A(net1009),
    .X(_09127_));
 sg13g2_buf_1 _14719_ (.A(net964),
    .X(_09128_));
 sg13g2_nand2_1 _14720_ (.Y(_09129_),
    .A(net1016),
    .B(net1013));
 sg13g2_buf_2 _14721_ (.A(_09129_),
    .X(_09130_));
 sg13g2_nor2_1 _14722_ (.A(_09066_),
    .B(net1017),
    .Y(_09131_));
 sg13g2_buf_2 _14723_ (.A(_09131_),
    .X(_09132_));
 sg13g2_nand4_1 _14724_ (.B(_09130_),
    .C(_09098_),
    .A(_09128_),
    .Y(_09133_),
    .D(_09132_));
 sg13g2_nand3_1 _14725_ (.B(_09125_),
    .C(_09133_),
    .A(net1010),
    .Y(_09134_));
 sg13g2_buf_2 _14726_ (.A(_00214_),
    .X(_09135_));
 sg13g2_nand2_1 _14727_ (.Y(_09136_),
    .A(_09019_),
    .B(_09135_));
 sg13g2_nand3_1 _14728_ (.B(_09134_),
    .C(_09136_),
    .A(net1019),
    .Y(_09137_));
 sg13g2_o21ai_1 _14729_ (.B1(_09137_),
    .Y(_09138_),
    .A1(net981),
    .A2(_09104_));
 sg13g2_buf_1 _14730_ (.A(_09010_),
    .X(_09139_));
 sg13g2_nand2_1 _14731_ (.Y(_09140_),
    .A(_08203_),
    .B(net828));
 sg13g2_o21ai_1 _14732_ (.B1(_09140_),
    .Y(_00395_),
    .A1(net829),
    .A2(_09138_));
 sg13g2_inv_2 _14733_ (.Y(_09141_),
    .A(net1041));
 sg13g2_buf_2 _14734_ (.A(net1012),
    .X(_09142_));
 sg13g2_buf_1 _14735_ (.A(net972),
    .X(_09143_));
 sg13g2_nand2_1 _14736_ (.Y(_09144_),
    .A(_09030_),
    .B(net860));
 sg13g2_nor2_1 _14737_ (.A(net1014),
    .B(_09130_),
    .Y(_09145_));
 sg13g2_nor3_1 _14738_ (.A(net974),
    .B(net968),
    .C(_09062_),
    .Y(_09146_));
 sg13g2_o21ai_1 _14739_ (.B1(_09115_),
    .Y(_09147_),
    .A1(_09145_),
    .A2(_09146_));
 sg13g2_o21ai_1 _14740_ (.B1(_09147_),
    .Y(_09148_),
    .A1(net918),
    .A2(_09144_));
 sg13g2_nor2_1 _14741_ (.A(net975),
    .B(net1014),
    .Y(_09149_));
 sg13g2_buf_2 _14742_ (.A(_09149_),
    .X(_09150_));
 sg13g2_nor2_1 _14743_ (.A(_09021_),
    .B(_09057_),
    .Y(_09151_));
 sg13g2_buf_1 _14744_ (.A(_09151_),
    .X(_09152_));
 sg13g2_buf_1 _14745_ (.A(_09152_),
    .X(_09153_));
 sg13g2_a22oi_1 _14746_ (.Y(_09154_),
    .B1(_09150_),
    .B2(net885),
    .A2(net860),
    .A1(net920));
 sg13g2_buf_1 _14747_ (.A(net978),
    .X(_09155_));
 sg13g2_nand2_1 _14748_ (.Y(_09156_),
    .A(_09155_),
    .B(_09016_));
 sg13g2_nor2_1 _14749_ (.A(_09154_),
    .B(_09156_),
    .Y(_09157_));
 sg13g2_a21oi_1 _14750_ (.A1(net919),
    .A2(_09148_),
    .Y(_09158_),
    .B1(_09157_));
 sg13g2_nor2_1 _14751_ (.A(net977),
    .B(net980),
    .Y(_09159_));
 sg13g2_nand2_1 _14752_ (.Y(_09160_),
    .A(_09070_),
    .B(net973));
 sg13g2_buf_2 _14753_ (.A(_09160_),
    .X(_09161_));
 sg13g2_nand2_1 _14754_ (.Y(_09162_),
    .A(net1038),
    .B(_09031_));
 sg13g2_buf_1 _14755_ (.A(_09162_),
    .X(_09163_));
 sg13g2_nand2_1 _14756_ (.Y(_09164_),
    .A(_09032_),
    .B(_09066_));
 sg13g2_nand4_1 _14757_ (.B(_09021_),
    .C(_09163_),
    .A(net975),
    .Y(_09165_),
    .D(_09164_));
 sg13g2_o21ai_1 _14758_ (.B1(_09165_),
    .Y(_09166_),
    .A1(_09130_),
    .A2(_09161_));
 sg13g2_nor2_1 _14759_ (.A(net978),
    .B(net971),
    .Y(_09167_));
 sg13g2_nor2_2 _14760_ (.A(net1011),
    .B(net1015),
    .Y(_09168_));
 sg13g2_nor2_1 _14761_ (.A(net1013),
    .B(_09057_),
    .Y(_09169_));
 sg13g2_buf_1 _14762_ (.A(_09169_),
    .X(_09170_));
 sg13g2_a21o_1 _14763_ (.A2(_09168_),
    .A1(net969),
    .B1(_09170_),
    .X(_09171_));
 sg13g2_a22oi_1 _14764_ (.Y(_09172_),
    .B1(_09171_),
    .B2(net924),
    .A2(_09167_),
    .A1(_09094_));
 sg13g2_nand2_1 _14765_ (.Y(_09173_),
    .A(net1015),
    .B(net1040));
 sg13g2_buf_1 _14766_ (.A(_09173_),
    .X(_09174_));
 sg13g2_buf_1 _14767_ (.A(_09070_),
    .X(_09175_));
 sg13g2_nor2_1 _14768_ (.A(_09027_),
    .B(net1013),
    .Y(_09176_));
 sg13g2_nand2_1 _14769_ (.Y(_09177_),
    .A(net962),
    .B(_09176_));
 sg13g2_or2_1 _14770_ (.X(_09178_),
    .B(_09177_),
    .A(_09174_));
 sg13g2_o21ai_1 _14771_ (.B1(_09178_),
    .Y(_09179_),
    .A1(net964),
    .A2(_09172_));
 sg13g2_inv_1 _14772_ (.Y(_09180_),
    .A(_09109_));
 sg13g2_a221oi_1 _14773_ (.B2(_09180_),
    .C1(net1018),
    .B1(_09179_),
    .A1(_09159_),
    .Y(_09181_),
    .A2(_09166_));
 sg13g2_a21o_1 _14774_ (.A2(_09158_),
    .A1(net963),
    .B1(_09181_),
    .X(_09182_));
 sg13g2_nor2_1 _14775_ (.A(net975),
    .B(_09031_),
    .Y(_09183_));
 sg13g2_buf_2 _14776_ (.A(_09183_),
    .X(_09184_));
 sg13g2_nor2_1 _14777_ (.A(_09035_),
    .B(_09085_),
    .Y(_09185_));
 sg13g2_a21oi_1 _14778_ (.A1(_09184_),
    .A2(_09185_),
    .Y(_09186_),
    .B1(net1040));
 sg13g2_and2_1 _14779_ (.A(net1010),
    .B(_09186_),
    .X(_09187_));
 sg13g2_nand2_1 _14780_ (.Y(_09188_),
    .A(net1016),
    .B(net973));
 sg13g2_buf_1 _14781_ (.A(_09188_),
    .X(_09189_));
 sg13g2_nand2_1 _14782_ (.Y(_09190_),
    .A(_09045_),
    .B(_09032_));
 sg13g2_nor2_1 _14783_ (.A(net1015),
    .B(_09190_),
    .Y(_09191_));
 sg13g2_a21oi_1 _14784_ (.A1(net927),
    .A2(_09069_),
    .Y(_09192_),
    .B1(_09191_));
 sg13g2_or2_1 _14785_ (.X(_09193_),
    .B(_09192_),
    .A(_09189_));
 sg13g2_nor2_1 _14786_ (.A(net1014),
    .B(net969),
    .Y(_09194_));
 sg13g2_nand2_1 _14787_ (.Y(_09195_),
    .A(_09194_),
    .B(net887));
 sg13g2_nand3_1 _14788_ (.B(_09193_),
    .C(_09195_),
    .A(_09187_),
    .Y(_09196_));
 sg13g2_a22oi_1 _14789_ (.Y(_09197_),
    .B1(net966),
    .B2(net962),
    .A2(net887),
    .A1(net976));
 sg13g2_buf_1 _14790_ (.A(net974),
    .X(_09198_));
 sg13g2_nand3_1 _14791_ (.B(net962),
    .C(net885),
    .A(net916),
    .Y(_09199_));
 sg13g2_o21ai_1 _14792_ (.B1(_09199_),
    .Y(_09200_),
    .A1(net921),
    .A2(_09197_));
 sg13g2_a22oi_1 _14793_ (.Y(_09201_),
    .B1(_09200_),
    .B2(net917),
    .A2(net887),
    .A1(net930));
 sg13g2_nand2_2 _14794_ (.Y(_09202_),
    .A(net974),
    .B(net968));
 sg13g2_a21oi_1 _14795_ (.A1(_09024_),
    .A2(_09202_),
    .Y(_09203_),
    .B1(_09097_));
 sg13g2_nand2b_1 _14796_ (.Y(_09204_),
    .B(net1039),
    .A_N(_09203_));
 sg13g2_buf_1 _14797_ (.A(net965),
    .X(_09205_));
 sg13g2_a21oi_1 _14798_ (.A1(_09084_),
    .A2(_09195_),
    .Y(_09206_),
    .B1(_09205_));
 sg13g2_o21ai_1 _14799_ (.B1(net923),
    .Y(_09207_),
    .A1(_09204_),
    .A2(_09206_));
 sg13g2_o21ai_1 _14800_ (.B1(_09207_),
    .Y(_09208_),
    .A1(net1018),
    .A2(_09201_));
 sg13g2_nand3_1 _14801_ (.B(_09196_),
    .C(_09208_),
    .A(net1019),
    .Y(_09209_));
 sg13g2_o21ai_1 _14802_ (.B1(_09209_),
    .Y(_09210_),
    .A1(net981),
    .A2(_09182_));
 sg13g2_nor2_1 _14803_ (.A(net828),
    .B(_09210_),
    .Y(_09211_));
 sg13g2_a21oi_1 _14804_ (.A1(_09141_),
    .A2(_09011_),
    .Y(_00396_),
    .B1(_09211_));
 sg13g2_buf_1 _14805_ (.A(_09176_),
    .X(_09212_));
 sg13g2_a22oi_1 _14806_ (.Y(_09213_),
    .B1(_09168_),
    .B2(net914),
    .A2(_09167_),
    .A1(_09150_));
 sg13g2_buf_1 _14807_ (.A(_00215_),
    .X(_09214_));
 sg13g2_inv_1 _14808_ (.Y(_09215_),
    .A(_09214_));
 sg13g2_nand4_1 _14809_ (.B(net1012),
    .C(_09215_),
    .A(net918),
    .Y(_09216_),
    .D(net931));
 sg13g2_o21ai_1 _14810_ (.B1(_09216_),
    .Y(_09217_),
    .A1(net1018),
    .A2(_09213_));
 sg13g2_nor2_1 _14811_ (.A(net979),
    .B(net1040),
    .Y(_09218_));
 sg13g2_nor3_1 _14812_ (.A(net975),
    .B(_09083_),
    .C(_09067_),
    .Y(_09219_));
 sg13g2_o21ai_1 _14813_ (.B1(_09049_),
    .Y(_09220_),
    .A1(_09198_),
    .A2(_09163_));
 sg13g2_a22oi_1 _14814_ (.Y(_09221_),
    .B1(_09220_),
    .B2(net966),
    .A2(_09219_),
    .A1(_09111_));
 sg13g2_nor2_1 _14815_ (.A(_09031_),
    .B(net973),
    .Y(_09222_));
 sg13g2_buf_1 _14816_ (.A(_09222_),
    .X(_09223_));
 sg13g2_nand4_1 _14817_ (.B(_09214_),
    .C(_09150_),
    .A(net1012),
    .Y(_09224_),
    .D(net884));
 sg13g2_o21ai_1 _14818_ (.B1(_09224_),
    .Y(_09225_),
    .A1(net1018),
    .A2(_09221_));
 sg13g2_buf_1 _14819_ (.A(_09127_),
    .X(_09226_));
 sg13g2_a22oi_1 _14820_ (.Y(_09227_),
    .B1(_09225_),
    .B2(net913),
    .A2(_09218_),
    .A1(_09217_));
 sg13g2_nor2_1 _14821_ (.A(_09046_),
    .B(_09022_),
    .Y(_09228_));
 sg13g2_buf_2 _14822_ (.A(_09228_),
    .X(_09229_));
 sg13g2_nor2_1 _14823_ (.A(_09032_),
    .B(_09021_),
    .Y(_09230_));
 sg13g2_buf_1 _14824_ (.A(_09230_),
    .X(_09231_));
 sg13g2_nor2_1 _14825_ (.A(net912),
    .B(net884),
    .Y(_09232_));
 sg13g2_inv_1 _14826_ (.Y(_09233_),
    .A(_09232_));
 sg13g2_a22oi_1 _14827_ (.Y(_09234_),
    .B1(_09233_),
    .B2(_09150_),
    .A2(_09229_),
    .A1(_09094_));
 sg13g2_nor3_1 _14828_ (.A(net1018),
    .B(_09174_),
    .C(_09234_),
    .Y(_09235_));
 sg13g2_and2_1 _14829_ (.A(net931),
    .B(_09229_),
    .X(_09236_));
 sg13g2_and4_1 _14830_ (.A(net1018),
    .B(_09135_),
    .C(_09214_),
    .D(_09236_),
    .X(_09237_));
 sg13g2_o21ai_1 _14831_ (.B1(net1019),
    .Y(_09238_),
    .A1(_09235_),
    .A2(_09237_));
 sg13g2_o21ai_1 _14832_ (.B1(_09238_),
    .Y(_09239_),
    .A1(net1019),
    .A2(_09227_));
 sg13g2_nor2_1 _14833_ (.A(net828),
    .B(_09239_),
    .Y(_09240_));
 sg13g2_a21oi_1 _14834_ (.A1(_08990_),
    .A2(_09011_),
    .Y(_00397_),
    .B1(_09240_));
 sg13g2_nor2_2 _14835_ (.A(_09045_),
    .B(_09034_),
    .Y(_09241_));
 sg13g2_nand2_1 _14836_ (.Y(_09242_),
    .A(_09189_),
    .B(_09241_));
 sg13g2_nor2_1 _14837_ (.A(_09038_),
    .B(net979),
    .Y(_09243_));
 sg13g2_buf_1 _14838_ (.A(_09243_),
    .X(_09244_));
 sg13g2_nand2_1 _14839_ (.Y(_09245_),
    .A(net1038),
    .B(net1017));
 sg13g2_buf_2 _14840_ (.A(_09245_),
    .X(_09246_));
 sg13g2_and2_1 _14841_ (.A(_09198_),
    .B(_09246_),
    .X(_09247_));
 sg13g2_buf_1 _14842_ (.A(_09036_),
    .X(_09248_));
 sg13g2_o21ai_1 _14843_ (.B1(net911),
    .Y(_09249_),
    .A1(_09244_),
    .A2(_09247_));
 sg13g2_a21oi_1 _14844_ (.A1(_09242_),
    .A2(_09249_),
    .Y(_09250_),
    .B1(net917));
 sg13g2_buf_1 _14845_ (.A(net970),
    .X(_09251_));
 sg13g2_nand2_1 _14846_ (.Y(_09252_),
    .A(_09251_),
    .B(_09184_));
 sg13g2_o21ai_1 _14847_ (.B1(_09226_),
    .Y(_09253_),
    .A1(_09091_),
    .A2(_09252_));
 sg13g2_buf_1 _14848_ (.A(_00219_),
    .X(_09254_));
 sg13g2_nor2_1 _14849_ (.A(_09038_),
    .B(net1015),
    .Y(_09255_));
 sg13g2_buf_1 _14850_ (.A(net968),
    .X(_09256_));
 sg13g2_nand2_1 _14851_ (.Y(_09257_),
    .A(net968),
    .B(_09170_));
 sg13g2_o21ai_1 _14852_ (.B1(_09257_),
    .Y(_09258_),
    .A1(net909),
    .A2(_09099_));
 sg13g2_buf_1 _14853_ (.A(_09095_),
    .X(_09259_));
 sg13g2_a22oi_1 _14854_ (.Y(_09260_),
    .B1(_09258_),
    .B2(net883),
    .A2(_09255_),
    .A1(_09254_));
 sg13g2_o21ai_1 _14855_ (.B1(_09186_),
    .Y(_09261_),
    .A1(net889),
    .A2(_09260_));
 sg13g2_o21ai_1 _14856_ (.B1(_09261_),
    .Y(_09262_),
    .A1(_09250_),
    .A2(_09253_));
 sg13g2_and2_1 _14857_ (.A(_09212_),
    .B(_09153_),
    .X(_09263_));
 sg13g2_a21oi_1 _14858_ (.A1(net915),
    .A2(net860),
    .Y(_09264_),
    .B1(_09263_));
 sg13g2_nand2_1 _14859_ (.Y(_09265_),
    .A(_09047_),
    .B(net860));
 sg13g2_o21ai_1 _14860_ (.B1(_09265_),
    .Y(_09266_),
    .A1(net922),
    .A2(_09264_));
 sg13g2_buf_1 _14861_ (.A(net971),
    .X(_09267_));
 sg13g2_nor2_1 _14862_ (.A(_09045_),
    .B(net978),
    .Y(_09268_));
 sg13g2_a221oi_1 _14863_ (.B2(net888),
    .C1(net885),
    .B1(_09268_),
    .A1(net908),
    .Y(_09269_),
    .A2(_09180_));
 sg13g2_nor2_1 _14864_ (.A(net968),
    .B(net971),
    .Y(_09270_));
 sg13g2_o21ai_1 _14865_ (.B1(net915),
    .Y(_09271_),
    .A1(net917),
    .A2(_09270_));
 sg13g2_and3_1 _14866_ (.X(_09272_),
    .A(net919),
    .B(_09269_),
    .C(_09271_));
 sg13g2_a21oi_1 _14867_ (.A1(net933),
    .A2(_09266_),
    .Y(_09273_),
    .B1(_09272_));
 sg13g2_nor2_1 _14868_ (.A(net1016),
    .B(_09032_),
    .Y(_09274_));
 sg13g2_buf_2 _14869_ (.A(_09274_),
    .X(_09275_));
 sg13g2_nor2_2 _14870_ (.A(_09184_),
    .B(_09275_),
    .Y(_09276_));
 sg13g2_nor2_1 _14871_ (.A(_09092_),
    .B(net1017),
    .Y(_09277_));
 sg13g2_nor2b_1 _14872_ (.A(_09276_),
    .B_N(_09277_),
    .Y(_09278_));
 sg13g2_nor2_1 _14873_ (.A(_09068_),
    .B(_09278_),
    .Y(_09279_));
 sg13g2_nor2_1 _14874_ (.A(net1038),
    .B(net973),
    .Y(_09280_));
 sg13g2_buf_2 _14875_ (.A(_09280_),
    .X(_09281_));
 sg13g2_nand2_1 _14876_ (.Y(_09282_),
    .A(net979),
    .B(_09268_));
 sg13g2_nand2_1 _14877_ (.Y(_09283_),
    .A(net978),
    .B(_09072_));
 sg13g2_a21oi_1 _14878_ (.A1(_09282_),
    .A2(_09283_),
    .Y(_09284_),
    .B1(net924));
 sg13g2_a221oi_1 _14879_ (.B2(_09254_),
    .C1(_09284_),
    .B1(_09281_),
    .A1(_09072_),
    .Y(_09285_),
    .A2(net925));
 sg13g2_buf_2 _14880_ (.A(_00218_),
    .X(_09286_));
 sg13g2_a221oi_1 _14881_ (.B2(_09286_),
    .C1(net911),
    .B1(_09244_),
    .A1(_09094_),
    .Y(_09287_),
    .A2(_09232_));
 sg13g2_nand2_1 _14882_ (.Y(_09288_),
    .A(_09033_),
    .B(_09023_));
 sg13g2_nand2_1 _14883_ (.Y(_09289_),
    .A(net976),
    .B(net912));
 sg13g2_o21ai_1 _14884_ (.B1(_09289_),
    .Y(_09290_),
    .A1(_09251_),
    .A2(_09288_));
 sg13g2_nand2_1 _14885_ (.Y(_09291_),
    .A(_09259_),
    .B(_09290_));
 sg13g2_a22oi_1 _14886_ (.Y(_09292_),
    .B1(_09287_),
    .B2(_09291_),
    .A2(_09285_),
    .A1(_09279_));
 sg13g2_nand2_2 _14887_ (.Y(_09293_),
    .A(net978),
    .B(net973));
 sg13g2_nand2_1 _14888_ (.Y(_09294_),
    .A(net1016),
    .B(net979));
 sg13g2_o21ai_1 _14889_ (.B1(_09294_),
    .Y(_09295_),
    .A1(_09116_),
    .A2(_09293_));
 sg13g2_buf_1 _14890_ (.A(net1015),
    .X(_09296_));
 sg13g2_nand2_1 _14891_ (.Y(_09297_),
    .A(net979),
    .B(net961));
 sg13g2_o21ai_1 _14892_ (.B1(_09297_),
    .Y(_09298_),
    .A1(_09063_),
    .A2(net966));
 sg13g2_a22oi_1 _14893_ (.Y(_09299_),
    .B1(_09298_),
    .B2(_09150_),
    .A2(_09295_),
    .A1(_09241_));
 sg13g2_o21ai_1 _14894_ (.B1(_09246_),
    .Y(_09300_),
    .A1(_09091_),
    .A2(_09202_));
 sg13g2_nand2_1 _14895_ (.Y(_09301_),
    .A(net918),
    .B(_09300_));
 sg13g2_a21oi_1 _14896_ (.A1(_09299_),
    .A2(_09301_),
    .Y(_09302_),
    .B1(_09107_));
 sg13g2_a21oi_1 _14897_ (.A1(_09018_),
    .A2(_09292_),
    .Y(_09303_),
    .B1(_09302_));
 sg13g2_nor2_1 _14898_ (.A(net927),
    .B(net967),
    .Y(_09304_));
 sg13g2_nand2_1 _14899_ (.Y(_09305_),
    .A(net970),
    .B(net971));
 sg13g2_nand2_1 _14900_ (.Y(_09306_),
    .A(net932),
    .B(_09305_));
 sg13g2_a22oi_1 _14901_ (.Y(_09307_),
    .B1(_09306_),
    .B2(net918),
    .A2(_09304_),
    .A1(net887));
 sg13g2_nand2_2 _14902_ (.Y(_09308_),
    .A(net1017),
    .B(_09057_));
 sg13g2_nand2_1 _14903_ (.Y(_09309_),
    .A(net1013),
    .B(net1015));
 sg13g2_o21ai_1 _14904_ (.B1(_09309_),
    .Y(_09310_),
    .A1(net972),
    .A2(_09308_));
 sg13g2_nand2_1 _14905_ (.Y(_09311_),
    .A(net909),
    .B(_09310_));
 sg13g2_a21oi_1 _14906_ (.A1(_09307_),
    .A2(_09311_),
    .Y(_09312_),
    .B1(net888));
 sg13g2_buf_1 _14907_ (.A(_09205_),
    .X(_09313_));
 sg13g2_nand2_1 _14908_ (.Y(_09314_),
    .A(_09083_),
    .B(net979));
 sg13g2_a21oi_1 _14909_ (.A1(net922),
    .A2(_09314_),
    .Y(_09315_),
    .B1(_09229_));
 sg13g2_nor3_1 _14910_ (.A(net882),
    .B(_09248_),
    .C(_09315_),
    .Y(_09316_));
 sg13g2_o21ai_1 _14911_ (.B1(_09135_),
    .Y(_09317_),
    .A1(_09312_),
    .A2(_09316_));
 sg13g2_mux4_1 _14912_ (.S0(_09142_),
    .A0(_09262_),
    .A1(_09273_),
    .A2(_09303_),
    .A3(_09317_),
    .S1(net981),
    .X(_09318_));
 sg13g2_nand2_1 _14913_ (.Y(_09319_),
    .A(\top_ihp.oisc.micro_op[12] ),
    .B(net828));
 sg13g2_o21ai_1 _14914_ (.B1(_09319_),
    .Y(_00398_),
    .A1(net829),
    .A2(_09318_));
 sg13g2_a21oi_1 _14915_ (.A1(_09087_),
    .A2(_09289_),
    .Y(_09320_),
    .B1(net882));
 sg13g2_nor3_1 _14916_ (.A(_09054_),
    .B(net922),
    .C(net912),
    .Y(_09321_));
 sg13g2_nor2_1 _14917_ (.A(_09320_),
    .B(_09321_),
    .Y(_09322_));
 sg13g2_nand2_1 _14918_ (.Y(_09323_),
    .A(_09259_),
    .B(_09223_));
 sg13g2_o21ai_1 _14919_ (.B1(_09323_),
    .Y(_09324_),
    .A1(net882),
    .A2(_09084_));
 sg13g2_nor2_2 _14920_ (.A(_09106_),
    .B(_09012_),
    .Y(_09325_));
 sg13g2_nand2_1 _14921_ (.Y(_09326_),
    .A(net933),
    .B(_09325_));
 sg13g2_a21oi_1 _14922_ (.A1(_09069_),
    .A2(_09324_),
    .Y(_09327_),
    .B1(_09326_));
 sg13g2_o21ai_1 _14923_ (.B1(_09327_),
    .Y(_09328_),
    .A1(net911),
    .A2(_09322_));
 sg13g2_nand2_1 _14924_ (.Y(_09329_),
    .A(net916),
    .B(_09244_));
 sg13g2_a21oi_1 _14925_ (.A1(_09246_),
    .A2(_09329_),
    .Y(_09330_),
    .B1(_09309_));
 sg13g2_a22oi_1 _14926_ (.Y(_09331_),
    .B1(net914),
    .B2(_09132_),
    .A2(_09254_),
    .A1(net932));
 sg13g2_nor2_1 _14927_ (.A(net929),
    .B(_09331_),
    .Y(_09332_));
 sg13g2_o21ai_1 _14928_ (.B1(net919),
    .Y(_09333_),
    .A1(_09330_),
    .A2(_09332_));
 sg13g2_a22oi_1 _14929_ (.Y(_09334_),
    .B1(_09167_),
    .B2(net916),
    .A2(net971),
    .A1(net967));
 sg13g2_nand2b_1 _14930_ (.Y(_09335_),
    .B(net889),
    .A_N(_09334_));
 sg13g2_o21ai_1 _14931_ (.B1(_09277_),
    .Y(_09336_),
    .A1(net929),
    .A2(_09275_));
 sg13g2_o21ai_1 _14932_ (.B1(_09288_),
    .Y(_09337_),
    .A1(net976),
    .A2(_09099_));
 sg13g2_nand2_1 _14933_ (.Y(_09338_),
    .A(net888),
    .B(_09337_));
 sg13g2_nand4_1 _14934_ (.B(_09335_),
    .C(_09336_),
    .A(_09107_),
    .Y(_09339_),
    .D(_09338_));
 sg13g2_a21oi_1 _14935_ (.A1(_09333_),
    .A2(_09339_),
    .Y(_09340_),
    .B1(net963));
 sg13g2_buf_1 _14936_ (.A(_09267_),
    .X(_09341_));
 sg13g2_o21ai_1 _14937_ (.B1(_09177_),
    .Y(_09342_),
    .A1(_09025_),
    .A2(_09220_));
 sg13g2_nand4_1 _14938_ (.B(net963),
    .C(_09135_),
    .A(net881),
    .Y(_09343_),
    .D(_09342_));
 sg13g2_nand3b_1 _14939_ (.B(_09343_),
    .C(_09013_),
    .Y(_09344_),
    .A_N(_09340_));
 sg13g2_a21oi_1 _14940_ (.A1(net920),
    .A2(net884),
    .Y(_09345_),
    .B1(_09231_));
 sg13g2_nor2_1 _14941_ (.A(_09078_),
    .B(_09314_),
    .Y(_09346_));
 sg13g2_nor3_1 _14942_ (.A(_09117_),
    .B(_09229_),
    .C(_09346_),
    .Y(_09347_));
 sg13g2_a21o_1 _14943_ (.A2(_09345_),
    .A1(net883),
    .B1(_09347_),
    .X(_09348_));
 sg13g2_or2_1 _14944_ (.X(_09349_),
    .B(_09012_),
    .A(net1039));
 sg13g2_buf_1 _14945_ (.A(_09349_),
    .X(_09350_));
 sg13g2_a21oi_1 _14946_ (.A1(_09132_),
    .A2(_09184_),
    .Y(_09351_),
    .B1(_09350_));
 sg13g2_o21ai_1 _14947_ (.B1(_09351_),
    .Y(_09352_),
    .A1(_09248_),
    .A2(_09348_));
 sg13g2_or2_1 _14948_ (.X(_09353_),
    .B(_09152_),
    .A(_09121_));
 sg13g2_buf_1 _14949_ (.A(_09353_),
    .X(_09354_));
 sg13g2_nor2_1 _14950_ (.A(_09184_),
    .B(_09354_),
    .Y(_09355_));
 sg13g2_a22oi_1 _14951_ (.Y(_09356_),
    .B1(_09355_),
    .B2(_09096_),
    .A2(_09354_),
    .A1(_09219_));
 sg13g2_o21ai_1 _14952_ (.B1(net970),
    .Y(_09357_),
    .A1(_09048_),
    .A2(_09067_));
 sg13g2_a21oi_1 _14953_ (.A1(net860),
    .A2(_09357_),
    .Y(_09358_),
    .B1(net885));
 sg13g2_nand2_1 _14954_ (.Y(_09359_),
    .A(net921),
    .B(_09229_));
 sg13g2_o21ai_1 _14955_ (.B1(_09359_),
    .Y(_09360_),
    .A1(_09155_),
    .A2(_09358_));
 sg13g2_a21oi_1 _14956_ (.A1(net919),
    .A2(_09360_),
    .Y(_09361_),
    .B1(_09350_));
 sg13g2_a21oi_1 _14957_ (.A1(_09325_),
    .A2(_09356_),
    .Y(_09362_),
    .B1(_09361_));
 sg13g2_a21o_1 _14958_ (.A2(_09352_),
    .A1(net933),
    .B1(_09362_),
    .X(_09363_));
 sg13g2_nand3_1 _14959_ (.B(_09344_),
    .C(_09363_),
    .A(_09328_),
    .Y(_09364_));
 sg13g2_nand2_1 _14960_ (.Y(_09365_),
    .A(\top_ihp.oisc.micro_op[13] ),
    .B(_09139_));
 sg13g2_o21ai_1 _14961_ (.B1(_09365_),
    .Y(_00399_),
    .A1(net829),
    .A2(_09364_));
 sg13g2_inv_1 _14962_ (.Y(_09366_),
    .A(\top_ihp.oisc.micro_op[14] ));
 sg13g2_nand2_1 _14963_ (.Y(_09367_),
    .A(net969),
    .B(net1040));
 sg13g2_or2_1 _14964_ (.X(_09368_),
    .B(_09367_),
    .A(_09297_));
 sg13g2_o21ai_1 _14965_ (.B1(_09368_),
    .Y(_09369_),
    .A1(_09091_),
    .A2(_09156_));
 sg13g2_a22oi_1 _14966_ (.Y(_09370_),
    .B1(_09369_),
    .B2(net883),
    .A2(_09263_),
    .A1(net964));
 sg13g2_inv_1 _14967_ (.Y(_09371_),
    .A(_09314_));
 sg13g2_nor2_1 _14968_ (.A(_09277_),
    .B(_09281_),
    .Y(_09372_));
 sg13g2_a22oi_1 _14969_ (.Y(_09373_),
    .B1(_09372_),
    .B2(net924),
    .A2(_09371_),
    .A1(net931));
 sg13g2_nor3_1 _14970_ (.A(net908),
    .B(net964),
    .C(_09373_),
    .Y(_09374_));
 sg13g2_a21oi_1 _14971_ (.A1(_09161_),
    .A2(_09246_),
    .Y(_09375_),
    .B1(net961));
 sg13g2_a22oi_1 _14972_ (.Y(_09376_),
    .B1(_09375_),
    .B2(net925),
    .A2(net884),
    .A1(_09094_));
 sg13g2_nor2_1 _14973_ (.A(net980),
    .B(_09376_),
    .Y(_09377_));
 sg13g2_nor2_1 _14974_ (.A(_09374_),
    .B(_09377_),
    .Y(_09378_));
 sg13g2_o21ai_1 _14975_ (.B1(_09378_),
    .Y(_09379_),
    .A1(_09108_),
    .A2(_09370_));
 sg13g2_nor2_1 _14976_ (.A(net967),
    .B(_09042_),
    .Y(_09380_));
 sg13g2_o21ai_1 _14977_ (.B1(_09081_),
    .Y(_09381_),
    .A1(_09042_),
    .A2(_09372_));
 sg13g2_a22oi_1 _14978_ (.Y(_09382_),
    .B1(_09381_),
    .B2(net881),
    .A2(_09380_),
    .A1(_09111_));
 sg13g2_a21o_1 _14979_ (.A2(net932),
    .A1(net928),
    .B1(_09244_),
    .X(_09383_));
 sg13g2_a221oi_1 _14980_ (.B2(_09383_),
    .C1(net919),
    .B1(_09170_),
    .A1(_09073_),
    .Y(_09384_),
    .A2(_09088_));
 sg13g2_a21oi_1 _14981_ (.A1(net913),
    .A2(_09382_),
    .Y(_09385_),
    .B1(_09384_));
 sg13g2_o21ai_1 _14982_ (.B1(_09202_),
    .Y(_09386_),
    .A1(net921),
    .A2(_09305_));
 sg13g2_a22oi_1 _14983_ (.Y(_09387_),
    .B1(net884),
    .B2(net909),
    .A2(_09163_),
    .A1(net916));
 sg13g2_nor2_1 _14984_ (.A(net908),
    .B(_09387_),
    .Y(_09388_));
 sg13g2_a21oi_1 _14985_ (.A1(net912),
    .A2(_09386_),
    .Y(_09389_),
    .B1(_09388_));
 sg13g2_nor2_1 _14986_ (.A(_09070_),
    .B(net971),
    .Y(_09390_));
 sg13g2_a21o_1 _14987_ (.A2(_09390_),
    .A1(net969),
    .B1(_09191_),
    .X(_09391_));
 sg13g2_a22oi_1 _14988_ (.Y(_09392_),
    .B1(_09391_),
    .B2(net916),
    .A2(_09390_),
    .A1(net914));
 sg13g2_a21o_1 _14989_ (.A2(_09170_),
    .A1(net974),
    .B1(_09275_),
    .X(_09393_));
 sg13g2_o21ai_1 _14990_ (.B1(_09309_),
    .Y(_09394_),
    .A1(net961),
    .A2(_09190_));
 sg13g2_a221oi_1 _14991_ (.B2(net928),
    .C1(net932),
    .B1(_09394_),
    .A1(_09039_),
    .Y(_09395_),
    .A2(_09393_));
 sg13g2_a21oi_1 _14992_ (.A1(net889),
    .A2(_09392_),
    .Y(_09396_),
    .B1(_09395_));
 sg13g2_nand2_1 _14993_ (.Y(_09397_),
    .A(net923),
    .B(_09396_));
 sg13g2_o21ai_1 _14994_ (.B1(_09397_),
    .Y(_09398_),
    .A1(net923),
    .A2(_09389_));
 sg13g2_nor2_1 _14995_ (.A(net976),
    .B(_09091_),
    .Y(_09399_));
 sg13g2_a21oi_1 _14996_ (.A1(net920),
    .A2(_09308_),
    .Y(_09400_),
    .B1(net928));
 sg13g2_o21ai_1 _14997_ (.B1(net886),
    .Y(_09401_),
    .A1(_09399_),
    .A2(_09400_));
 sg13g2_nor3_1 _14998_ (.A(net975),
    .B(_09092_),
    .C(net972),
    .Y(_09402_));
 sg13g2_nand2_1 _14999_ (.Y(_09403_),
    .A(net1013),
    .B(_09175_));
 sg13g2_o21ai_1 _15000_ (.B1(_09195_),
    .Y(_09404_),
    .A1(_09091_),
    .A2(_09403_));
 sg13g2_a22oi_1 _15001_ (.Y(_09405_),
    .B1(_09404_),
    .B2(net888),
    .A2(_09402_),
    .A1(net887));
 sg13g2_inv_1 _15002_ (.Y(_09406_),
    .A(_09135_));
 sg13g2_a21oi_1 _15003_ (.A1(_09401_),
    .A2(_09405_),
    .Y(_09407_),
    .B1(_09406_));
 sg13g2_mux4_1 _15004_ (.S0(_09142_),
    .A0(_09379_),
    .A1(_09385_),
    .A2(_09398_),
    .A3(_09407_),
    .S1(_09013_),
    .X(_09408_));
 sg13g2_nor2_1 _15005_ (.A(net828),
    .B(_09408_),
    .Y(_09409_));
 sg13g2_a21oi_1 _15006_ (.A1(_09366_),
    .A2(net829),
    .Y(_00400_),
    .B1(_09409_));
 sg13g2_nand2_1 _15007_ (.Y(_09410_),
    .A(_09286_),
    .B(_09281_));
 sg13g2_o21ai_1 _15008_ (.B1(_09410_),
    .Y(_09411_),
    .A1(_09130_),
    .A2(_09281_));
 sg13g2_nand3_1 _15009_ (.B(_09161_),
    .C(_09246_),
    .A(net974),
    .Y(_09412_));
 sg13g2_o21ai_1 _15010_ (.B1(_09412_),
    .Y(_09413_),
    .A1(net965),
    .A2(_09246_));
 sg13g2_a22oi_1 _15011_ (.Y(_09414_),
    .B1(_09413_),
    .B2(net918),
    .A2(net914),
    .A1(_09072_));
 sg13g2_nor2_1 _15012_ (.A(net881),
    .B(_09414_),
    .Y(_09415_));
 sg13g2_a21oi_1 _15013_ (.A1(net881),
    .A2(_09411_),
    .Y(_09416_),
    .B1(_09415_));
 sg13g2_nor2_2 _15014_ (.A(_09121_),
    .B(_09152_),
    .Y(_09417_));
 sg13g2_a21oi_1 _15015_ (.A1(net910),
    .A2(_09417_),
    .Y(_09418_),
    .B1(_09185_));
 sg13g2_nand2_1 _15016_ (.Y(_09419_),
    .A(net909),
    .B(net885));
 sg13g2_o21ai_1 _15017_ (.B1(_09419_),
    .Y(_09420_),
    .A1(net915),
    .A2(_09418_));
 sg13g2_nand2_1 _15018_ (.Y(_09421_),
    .A(net926),
    .B(net925));
 sg13g2_nand2_1 _15019_ (.Y(_09422_),
    .A(_09254_),
    .B(_09059_));
 sg13g2_a21oi_1 _15020_ (.A1(_09421_),
    .A2(_09422_),
    .Y(_09423_),
    .B1(net922));
 sg13g2_a21oi_1 _15021_ (.A1(net917),
    .A2(_09420_),
    .Y(_09424_),
    .B1(_09423_));
 sg13g2_mux2_1 _15022_ (.A0(_09416_),
    .A1(_09424_),
    .S(net933),
    .X(_09425_));
 sg13g2_a21oi_1 _15023_ (.A1(_09072_),
    .A2(_09042_),
    .Y(_09426_),
    .B1(net910));
 sg13g2_o21ai_1 _15024_ (.B1(_09410_),
    .Y(_09427_),
    .A1(net925),
    .A2(_09426_));
 sg13g2_nor2_1 _15025_ (.A(net980),
    .B(net1039),
    .Y(_09428_));
 sg13g2_a22oi_1 _15026_ (.Y(_09429_),
    .B1(net884),
    .B2(net970),
    .A2(_09072_),
    .A1(net972));
 sg13g2_nand2b_1 _15027_ (.Y(_09430_),
    .B(net924),
    .A_N(_09429_));
 sg13g2_inv_1 _15028_ (.Y(_09431_),
    .A(_09254_));
 sg13g2_nand2_1 _15029_ (.Y(_09432_),
    .A(_09293_),
    .B(_09282_));
 sg13g2_a22oi_1 _15030_ (.Y(_09433_),
    .B1(_09432_),
    .B2(net928),
    .A2(_09281_),
    .A1(_09431_));
 sg13g2_a21oi_1 _15031_ (.A1(_09430_),
    .A2(_09433_),
    .Y(_09434_),
    .B1(_09136_));
 sg13g2_a21oi_1 _15032_ (.A1(_09427_),
    .A2(_09428_),
    .Y(_09435_),
    .B1(_09434_));
 sg13g2_nor2_1 _15033_ (.A(net881),
    .B(_09435_),
    .Y(_09436_));
 sg13g2_a221oi_1 _15034_ (.B2(_09255_),
    .C1(net964),
    .B1(_09295_),
    .A1(net911),
    .Y(_09437_),
    .A2(_09109_));
 sg13g2_a21o_1 _15035_ (.A2(net980),
    .A1(net920),
    .B1(_09399_),
    .X(_09438_));
 sg13g2_a22oi_1 _15036_ (.Y(_09439_),
    .B1(_09438_),
    .B2(net883),
    .A2(net923),
    .A1(net908));
 sg13g2_nor3_1 _15037_ (.A(net1018),
    .B(_09437_),
    .C(_09439_),
    .Y(_09440_));
 sg13g2_nor3_1 _15038_ (.A(net883),
    .B(_09132_),
    .C(_09281_),
    .Y(_09441_));
 sg13g2_nor4_1 _15039_ (.A(_09097_),
    .B(_09136_),
    .C(_09247_),
    .D(_09441_),
    .Y(_09442_));
 sg13g2_nor3_1 _15040_ (.A(_09436_),
    .B(_09440_),
    .C(_09442_),
    .Y(_09443_));
 sg13g2_nor2_1 _15041_ (.A(net969),
    .B(net961),
    .Y(_09444_));
 sg13g2_nand2_1 _15042_ (.Y(_09445_),
    .A(_09098_),
    .B(_09305_));
 sg13g2_a22oi_1 _15043_ (.Y(_09446_),
    .B1(_09445_),
    .B2(net888),
    .A2(_09444_),
    .A1(net922));
 sg13g2_nor2_1 _15044_ (.A(net1038),
    .B(_09057_),
    .Y(_09447_));
 sg13g2_nor2_1 _15045_ (.A(_09241_),
    .B(_09447_),
    .Y(_09448_));
 sg13g2_nor2_1 _15046_ (.A(net965),
    .B(_09255_),
    .Y(_09449_));
 sg13g2_a21oi_1 _15047_ (.A1(net916),
    .A2(_09448_),
    .Y(_09450_),
    .B1(_09449_));
 sg13g2_a221oi_1 _15048_ (.B2(net927),
    .C1(net926),
    .B1(_09450_),
    .A1(_09286_),
    .Y(_09451_),
    .A2(_09270_));
 sg13g2_a21o_1 _15049_ (.A2(_09446_),
    .A1(net926),
    .B1(_09451_),
    .X(_09452_));
 sg13g2_a21oi_1 _15050_ (.A1(net922),
    .A2(_09309_),
    .Y(_09453_),
    .B1(_09189_));
 sg13g2_nor2_1 _15051_ (.A(net921),
    .B(net908),
    .Y(_09454_));
 sg13g2_nor3_1 _15052_ (.A(_09073_),
    .B(_09087_),
    .C(_09454_),
    .Y(_09455_));
 sg13g2_nor3_1 _15053_ (.A(net919),
    .B(_09453_),
    .C(_09455_),
    .Y(_09456_));
 sg13g2_a21oi_1 _15054_ (.A1(net913),
    .A2(_09452_),
    .Y(_09457_),
    .B1(_09456_));
 sg13g2_nor2_1 _15055_ (.A(_09350_),
    .B(_09457_),
    .Y(_09458_));
 sg13g2_a221oi_1 _15056_ (.B2(net981),
    .C1(_09458_),
    .B1(_09443_),
    .A1(_09325_),
    .Y(_09459_),
    .A2(_09425_));
 sg13g2_mux2_1 _15057_ (.A0(_09459_),
    .A1(\top_ihp.oisc.micro_op[15] ),
    .S(_09139_),
    .X(_00401_));
 sg13g2_nor3_1 _15058_ (.A(net915),
    .B(net967),
    .C(net929),
    .Y(_09460_));
 sg13g2_a22oi_1 _15059_ (.Y(_09461_),
    .B1(_09232_),
    .B2(_09460_),
    .A2(_09184_),
    .A1(_09111_));
 sg13g2_a21oi_1 _15060_ (.A1(_09175_),
    .A2(_09153_),
    .Y(_09462_),
    .B1(_09241_));
 sg13g2_o21ai_1 _15061_ (.B1(_09144_),
    .Y(_09463_),
    .A1(net928),
    .A2(_09462_));
 sg13g2_a221oi_1 _15062_ (.B2(_09143_),
    .C1(_09065_),
    .B1(_09463_),
    .A1(_09212_),
    .Y(_09464_),
    .A2(net966));
 sg13g2_a21oi_1 _15063_ (.A1(net963),
    .A2(_09461_),
    .Y(_09465_),
    .B1(_09464_));
 sg13g2_a21o_1 _15064_ (.A2(_09111_),
    .A1(net1040),
    .B1(net972),
    .X(_09466_));
 sg13g2_a21oi_1 _15065_ (.A1(_09094_),
    .A2(_09466_),
    .Y(_09467_),
    .B1(_09150_));
 sg13g2_a221oi_1 _15066_ (.B2(net918),
    .C1(_09467_),
    .B1(_09308_),
    .A1(_09051_),
    .Y(_09468_),
    .A2(_09109_));
 sg13g2_nor2_1 _15067_ (.A(net967),
    .B(_09354_),
    .Y(_09469_));
 sg13g2_a22oi_1 _15068_ (.Y(_09470_),
    .B1(_09469_),
    .B2(_09117_),
    .A2(_09354_),
    .A1(_09030_));
 sg13g2_nor3_1 _15069_ (.A(_09143_),
    .B(net1010),
    .C(_09470_),
    .Y(_09471_));
 sg13g2_a21oi_1 _15070_ (.A1(net1010),
    .A2(_09468_),
    .Y(_09472_),
    .B1(_09471_));
 sg13g2_nor2_1 _15071_ (.A(_09018_),
    .B(_09472_),
    .Y(_09473_));
 sg13g2_a21oi_1 _15072_ (.A1(net933),
    .A2(_09465_),
    .Y(_09474_),
    .B1(_09473_));
 sg13g2_a21oi_1 _15073_ (.A1(net962),
    .A2(_09275_),
    .Y(_09475_),
    .B1(net961));
 sg13g2_nand2_1 _15074_ (.Y(_09476_),
    .A(net1015),
    .B(_09165_));
 sg13g2_a21oi_1 _15075_ (.A1(_09029_),
    .A2(net912),
    .Y(_09477_),
    .B1(_09476_));
 sg13g2_nor4_1 _15076_ (.A(net1040),
    .B(net1010),
    .C(_09475_),
    .D(_09477_),
    .Y(_09478_));
 sg13g2_nand2_1 _15077_ (.Y(_09479_),
    .A(net1014),
    .B(_09403_));
 sg13g2_o21ai_1 _15078_ (.B1(_09479_),
    .Y(_09480_),
    .A1(_09116_),
    .A2(_09164_));
 sg13g2_a22oi_1 _15079_ (.Y(_09481_),
    .B1(_09480_),
    .B2(_09077_),
    .A2(_09145_),
    .A1(_09161_));
 sg13g2_nand2_1 _15080_ (.Y(_09482_),
    .A(net968),
    .B(net971));
 sg13g2_nand3_1 _15081_ (.B(_09275_),
    .C(_09482_),
    .A(_09132_),
    .Y(_09483_));
 sg13g2_o21ai_1 _15082_ (.B1(_09483_),
    .Y(_09484_),
    .A1(net929),
    .A2(_09481_));
 sg13g2_nand2_1 _15083_ (.Y(_09485_),
    .A(net1014),
    .B(_09276_));
 sg13g2_o21ai_1 _15084_ (.B1(_09485_),
    .Y(_09486_),
    .A1(net1014),
    .A2(_09286_));
 sg13g2_nor2_1 _15085_ (.A(net932),
    .B(_09486_),
    .Y(_09487_));
 sg13g2_nor3_1 _15086_ (.A(net908),
    .B(_09346_),
    .C(_09487_),
    .Y(_09488_));
 sg13g2_a21oi_1 _15087_ (.A1(_09403_),
    .A2(_09164_),
    .Y(_09489_),
    .B1(_09294_));
 sg13g2_nand2_1 _15088_ (.Y(_09490_),
    .A(net969),
    .B(net1011));
 sg13g2_a21oi_1 _15089_ (.A1(net932),
    .A2(_09490_),
    .Y(_09491_),
    .B1(net965));
 sg13g2_nor4_1 _15090_ (.A(net977),
    .B(_09244_),
    .C(_09489_),
    .D(_09491_),
    .Y(_09492_));
 sg13g2_nor3_1 _15091_ (.A(net964),
    .B(_09488_),
    .C(_09492_),
    .Y(_09493_));
 sg13g2_a21oi_1 _15092_ (.A1(net919),
    .A2(_09484_),
    .Y(_09494_),
    .B1(_09493_));
 sg13g2_nor2_1 _15093_ (.A(net963),
    .B(_09494_),
    .Y(_09495_));
 sg13g2_o21ai_1 _15094_ (.B1(net1019),
    .Y(_09496_),
    .A1(_09478_),
    .A2(_09495_));
 sg13g2_o21ai_1 _15095_ (.B1(_09496_),
    .Y(_09497_),
    .A1(net981),
    .A2(_09474_));
 sg13g2_mux2_1 _15096_ (.A0(_09497_),
    .A1(_08202_),
    .S(net828),
    .X(_00402_));
 sg13g2_nor2_1 _15097_ (.A(_09015_),
    .B(net1039),
    .Y(_09498_));
 sg13g2_a21o_1 _15098_ (.A2(net885),
    .A1(_09119_),
    .B1(net860),
    .X(_09499_));
 sg13g2_a22oi_1 _15099_ (.Y(_09500_),
    .B1(_09499_),
    .B2(net886),
    .A2(_09113_),
    .A1(_09194_));
 sg13g2_a21oi_1 _15100_ (.A1(net922),
    .A2(net887),
    .Y(_09501_),
    .B1(_09399_));
 sg13g2_nand2_1 _15101_ (.Y(_09502_),
    .A(_09184_),
    .B(_09501_));
 sg13g2_o21ai_1 _15102_ (.B1(_09502_),
    .Y(_09503_),
    .A1(net882),
    .A2(_09500_));
 sg13g2_nor2_1 _15103_ (.A(net1016),
    .B(_09109_),
    .Y(_09504_));
 sg13g2_a22oi_1 _15104_ (.Y(_09505_),
    .B1(_09504_),
    .B2(_09170_),
    .A2(_09121_),
    .A1(net925));
 sg13g2_nand3_1 _15105_ (.B(net966),
    .C(_09276_),
    .A(net1011),
    .Y(_09506_));
 sg13g2_o21ai_1 _15106_ (.B1(_09506_),
    .Y(_09507_),
    .A1(net976),
    .A2(_09505_));
 sg13g2_a21o_1 _15107_ (.A2(_09507_),
    .A1(_09428_),
    .B1(_09478_),
    .X(_09508_));
 sg13g2_a21oi_1 _15108_ (.A1(_09498_),
    .A2(_09503_),
    .Y(_09509_),
    .B1(_09508_));
 sg13g2_nor2_1 _15109_ (.A(net974),
    .B(_09023_),
    .Y(_09510_));
 sg13g2_a21oi_1 _15110_ (.A1(net883),
    .A2(_09281_),
    .Y(_09511_),
    .B1(_09510_));
 sg13g2_nor4_1 _15111_ (.A(_09064_),
    .B(net963),
    .C(_09174_),
    .D(_09511_),
    .Y(_09512_));
 sg13g2_a21oi_1 _15112_ (.A1(_09053_),
    .A2(_09044_),
    .Y(_09513_),
    .B1(_09402_));
 sg13g2_a22oi_1 _15113_ (.Y(_09514_),
    .B1(_09121_),
    .B2(net914),
    .A2(net912),
    .A1(_09296_));
 sg13g2_or2_1 _15114_ (.X(_09515_),
    .B(_09514_),
    .A(net910));
 sg13g2_o21ai_1 _15115_ (.B1(_09515_),
    .Y(_09516_),
    .A1(_09122_),
    .A2(_09513_));
 sg13g2_a22oi_1 _15116_ (.Y(_09517_),
    .B1(_09275_),
    .B2(_09086_),
    .A2(_09229_),
    .A1(_09150_));
 sg13g2_nor3_1 _15117_ (.A(net911),
    .B(net1012),
    .C(_09517_),
    .Y(_09518_));
 sg13g2_a21oi_1 _15118_ (.A1(_09065_),
    .A2(_09516_),
    .Y(_09519_),
    .B1(_09518_));
 sg13g2_nor2_1 _15119_ (.A(net930),
    .B(_09047_),
    .Y(_09520_));
 sg13g2_o21ai_1 _15120_ (.B1(_09485_),
    .Y(_09521_),
    .A1(net962),
    .A2(_09276_));
 sg13g2_a22oi_1 _15121_ (.Y(_09522_),
    .B1(_09521_),
    .B2(net932),
    .A2(_09510_),
    .A1(_09520_));
 sg13g2_nand2_1 _15122_ (.Y(_09523_),
    .A(net975),
    .B(net884));
 sg13g2_nand2_1 _15123_ (.Y(_09524_),
    .A(net962),
    .B(net961));
 sg13g2_a21o_1 _15124_ (.A2(_09523_),
    .A1(_09421_),
    .B1(_09524_),
    .X(_09525_));
 sg13g2_o21ai_1 _15125_ (.B1(_09525_),
    .Y(_09526_),
    .A1(net929),
    .A2(_09522_));
 sg13g2_nor2_1 _15126_ (.A(net917),
    .B(net1010),
    .Y(_09527_));
 sg13g2_o21ai_1 _15127_ (.B1(_09256_),
    .Y(_09528_),
    .A1(_09111_),
    .A2(net860));
 sg13g2_nand2_1 _15128_ (.Y(_09529_),
    .A(_09053_),
    .B(_09375_));
 sg13g2_o21ai_1 _15129_ (.B1(_09529_),
    .Y(_09530_),
    .A1(_09054_),
    .A2(_09528_));
 sg13g2_a221oi_1 _15130_ (.B2(_09530_),
    .C1(_09226_),
    .B1(_09527_),
    .A1(net1010),
    .Y(_09531_),
    .A2(_09526_));
 sg13g2_a21oi_1 _15131_ (.A1(net913),
    .A2(_09519_),
    .Y(_09532_),
    .B1(_09531_));
 sg13g2_nor3_1 _15132_ (.A(net1019),
    .B(_09512_),
    .C(_09532_),
    .Y(_09533_));
 sg13g2_a21oi_1 _15133_ (.A1(net981),
    .A2(_09509_),
    .Y(_09534_),
    .B1(_09533_));
 sg13g2_mux2_1 _15134_ (.A0(_09534_),
    .A1(_08205_),
    .S(net828),
    .X(_00403_));
 sg13g2_inv_1 _15135_ (.Y(_09535_),
    .A(_08204_));
 sg13g2_nor2_1 _15136_ (.A(_09070_),
    .B(net973),
    .Y(_09536_));
 sg13g2_nand2_1 _15137_ (.Y(_09537_),
    .A(net969),
    .B(_09536_));
 sg13g2_o21ai_1 _15138_ (.B1(_09537_),
    .Y(_09538_),
    .A1(net970),
    .A2(_09293_));
 sg13g2_a221oi_1 _15139_ (.B2(net928),
    .C1(net977),
    .B1(_09538_),
    .A1(_09184_),
    .Y(_09539_),
    .A2(_09536_));
 sg13g2_nor4_1 _15140_ (.A(net964),
    .B(net1039),
    .C(_09279_),
    .D(_09539_),
    .Y(_09540_));
 sg13g2_o21ai_1 _15141_ (.B1(_09012_),
    .Y(_09541_),
    .A1(_09508_),
    .A2(_09540_));
 sg13g2_nor2b_1 _15142_ (.A(_09010_),
    .B_N(_09541_),
    .Y(_09542_));
 sg13g2_and3_1 _15143_ (.X(_09543_),
    .A(_09180_),
    .B(_09168_),
    .C(_09275_));
 sg13g2_inv_1 _15144_ (.Y(_09544_),
    .A(_09543_));
 sg13g2_nand2_1 _15145_ (.Y(_09545_),
    .A(net1009),
    .B(_09236_));
 sg13g2_a221oi_1 _15146_ (.B2(net931),
    .C1(net1009),
    .B1(_09229_),
    .A1(net925),
    .Y(_09546_),
    .A2(_09086_));
 sg13g2_a221oi_1 _15147_ (.B2(net911),
    .C1(_09546_),
    .B1(_09545_),
    .A1(_09159_),
    .Y(_09547_),
    .A2(_09544_));
 sg13g2_or2_1 _15148_ (.X(_09548_),
    .B(_09547_),
    .A(_09020_));
 sg13g2_nor3_1 _15149_ (.A(_09202_),
    .B(_09174_),
    .C(_09288_),
    .Y(_09549_));
 sg13g2_nand3_1 _15150_ (.B(_09159_),
    .C(net884),
    .A(net931),
    .Y(_09550_));
 sg13g2_nand3_1 _15151_ (.B(_09115_),
    .C(_09219_),
    .A(net1009),
    .Y(_09551_));
 sg13g2_o21ai_1 _15152_ (.B1(_09551_),
    .Y(_09552_),
    .A1(_09127_),
    .A2(_09544_));
 sg13g2_nor2_1 _15153_ (.A(net1010),
    .B(_09552_),
    .Y(_09553_));
 sg13g2_a21oi_1 _15154_ (.A1(_09550_),
    .A2(_09553_),
    .Y(_09554_),
    .B1(_09014_));
 sg13g2_o21ai_1 _15155_ (.B1(_09554_),
    .Y(_09555_),
    .A1(_09548_),
    .A2(_09549_));
 sg13g2_a22oi_1 _15156_ (.Y(_00404_),
    .B1(_09542_),
    .B2(_09555_),
    .A2(net829),
    .A1(_09535_));
 sg13g2_inv_1 _15157_ (.Y(_09556_),
    .A(_08206_));
 sg13g2_nor2_1 _15158_ (.A(net926),
    .B(_09016_),
    .Y(_09557_));
 sg13g2_nor2_1 _15159_ (.A(net927),
    .B(_09202_),
    .Y(_09558_));
 sg13g2_a22oi_1 _15160_ (.Y(_09559_),
    .B1(_09557_),
    .B2(_09047_),
    .A2(_09218_),
    .A1(net930));
 sg13g2_nor2_1 _15161_ (.A(net883),
    .B(_09559_),
    .Y(_09560_));
 sg13g2_a21oi_1 _15162_ (.A1(_09557_),
    .A2(_09558_),
    .Y(_09561_),
    .B1(_09560_));
 sg13g2_nor2_1 _15163_ (.A(net881),
    .B(_09561_),
    .Y(_09562_));
 sg13g2_nand4_1 _15164_ (.B(net923),
    .C(_09150_),
    .A(net911),
    .Y(_09563_),
    .D(_09229_));
 sg13g2_a21oi_1 _15165_ (.A1(_09553_),
    .A2(_09563_),
    .Y(_09564_),
    .B1(_09012_));
 sg13g2_o21ai_1 _15166_ (.B1(_09564_),
    .Y(_09565_),
    .A1(_09548_),
    .A2(_09562_));
 sg13g2_and2_1 _15167_ (.A(_09542_),
    .B(_09565_),
    .X(_09566_));
 sg13g2_a21oi_1 _15168_ (.A1(_09556_),
    .A2(net829),
    .Y(_00405_),
    .B1(_09566_));
 sg13g2_inv_1 _15169_ (.Y(_09567_),
    .A(_08207_));
 sg13g2_nand4_1 _15170_ (.B(_09159_),
    .C(_09223_),
    .A(net931),
    .Y(_09568_),
    .D(_09325_));
 sg13g2_a22oi_1 _15171_ (.Y(_00406_),
    .B1(_09566_),
    .B2(_09568_),
    .A2(_09008_),
    .A1(_09567_));
 sg13g2_inv_1 _15172_ (.Y(_09569_),
    .A(_08988_));
 sg13g2_nand2_1 _15173_ (.Y(_09570_),
    .A(_09189_),
    .B(_09246_));
 sg13g2_a21o_1 _15174_ (.A2(_09536_),
    .A1(net917),
    .B1(_09132_),
    .X(_09571_));
 sg13g2_a21oi_1 _15175_ (.A1(_09293_),
    .A2(_09490_),
    .Y(_09572_),
    .B1(net916));
 sg13g2_a221oi_1 _15176_ (.B2(net921),
    .C1(_09572_),
    .B1(_09571_),
    .A1(net927),
    .Y(_09573_),
    .A2(_09570_));
 sg13g2_nand2_1 _15177_ (.Y(_09574_),
    .A(net979),
    .B(_09286_));
 sg13g2_a21oi_1 _15178_ (.A1(_09084_),
    .A2(_09574_),
    .Y(_09575_),
    .B1(net909));
 sg13g2_o21ai_1 _15179_ (.B1(_09189_),
    .Y(_09576_),
    .A1(net910),
    .A2(_09042_));
 sg13g2_nor3_1 _15180_ (.A(net908),
    .B(_09575_),
    .C(_09576_),
    .Y(_09577_));
 sg13g2_a21oi_1 _15181_ (.A1(net881),
    .A2(_09573_),
    .Y(_09578_),
    .B1(_09577_));
 sg13g2_a22oi_1 _15182_ (.Y(_09579_),
    .B1(_09152_),
    .B2(net1011),
    .A2(_09121_),
    .A1(net970));
 sg13g2_a22oi_1 _15183_ (.Y(_09580_),
    .B1(_09417_),
    .B2(net965),
    .A2(net887),
    .A1(net968));
 sg13g2_o21ai_1 _15184_ (.B1(_09580_),
    .Y(_09581_),
    .A1(net924),
    .A2(_09579_));
 sg13g2_nand2_1 _15185_ (.Y(_09582_),
    .A(net974),
    .B(_09308_));
 sg13g2_a21oi_1 _15186_ (.A1(net1011),
    .A2(net885),
    .Y(_09583_),
    .B1(_09582_));
 sg13g2_a21oi_1 _15187_ (.A1(net1011),
    .A2(net966),
    .Y(_09584_),
    .B1(net965));
 sg13g2_nor3_1 _15188_ (.A(net927),
    .B(_09583_),
    .C(_09584_),
    .Y(_09585_));
 sg13g2_a21oi_1 _15189_ (.A1(net918),
    .A2(_09581_),
    .Y(_09586_),
    .B1(_09585_));
 sg13g2_nand2_1 _15190_ (.Y(_09587_),
    .A(net913),
    .B(_09586_));
 sg13g2_o21ai_1 _15191_ (.B1(_09587_),
    .Y(_09588_),
    .A1(net913),
    .A2(_09578_));
 sg13g2_o21ai_1 _15192_ (.B1(_09482_),
    .Y(_09589_),
    .A1(net967),
    .A2(_09297_));
 sg13g2_nor3_1 _15193_ (.A(net924),
    .B(net977),
    .C(_09072_),
    .Y(_09590_));
 sg13g2_a21oi_1 _15194_ (.A1(net915),
    .A2(_09589_),
    .Y(_09591_),
    .B1(_09590_));
 sg13g2_nand2_1 _15195_ (.Y(_09592_),
    .A(net920),
    .B(_09308_));
 sg13g2_nand2_1 _15196_ (.Y(_09593_),
    .A(_09256_),
    .B(net860));
 sg13g2_nand3_1 _15197_ (.B(_09592_),
    .C(_09593_),
    .A(_09080_),
    .Y(_09594_));
 sg13g2_o21ai_1 _15198_ (.B1(_09594_),
    .Y(_09595_),
    .A1(net886),
    .A2(_09591_));
 sg13g2_nand2b_1 _15199_ (.Y(_09596_),
    .B(_09595_),
    .A_N(_09136_));
 sg13g2_o21ai_1 _15200_ (.B1(_09596_),
    .Y(_09597_),
    .A1(net963),
    .A2(_09588_));
 sg13g2_a21o_1 _15201_ (.A2(_09558_),
    .A1(_09390_),
    .B1(net923),
    .X(_09598_));
 sg13g2_a21o_1 _15202_ (.A2(_09168_),
    .A1(net972),
    .B1(_09447_),
    .X(_09599_));
 sg13g2_a22oi_1 _15203_ (.Y(_09600_),
    .B1(_09599_),
    .B2(net915),
    .A2(net914),
    .A1(_09069_));
 sg13g2_nor2_1 _15204_ (.A(net970),
    .B(_09390_),
    .Y(_09601_));
 sg13g2_a21oi_1 _15205_ (.A1(net965),
    .A2(_09255_),
    .Y(_09602_),
    .B1(_09270_));
 sg13g2_o21ai_1 _15206_ (.B1(_09602_),
    .Y(_09603_),
    .A1(net916),
    .A2(_09601_));
 sg13g2_a221oi_1 _15207_ (.B2(net918),
    .C1(net889),
    .B1(_09603_),
    .A1(_09524_),
    .Y(_09604_),
    .A2(_09402_));
 sg13g2_a21oi_1 _15208_ (.A1(net889),
    .A2(_09600_),
    .Y(_09605_),
    .B1(_09604_));
 sg13g2_nor2_1 _15209_ (.A(net909),
    .B(_09444_),
    .Y(_09606_));
 sg13g2_or2_1 _15210_ (.X(_09607_),
    .B(_09606_),
    .A(_09189_));
 sg13g2_nor2_1 _15211_ (.A(net914),
    .B(_09241_),
    .Y(_09608_));
 sg13g2_o21ai_1 _15212_ (.B1(net976),
    .Y(_09609_),
    .A1(net977),
    .A2(_09130_));
 sg13g2_a221oi_1 _15213_ (.B2(net962),
    .C1(net926),
    .B1(_09609_),
    .A1(_09081_),
    .Y(_09610_),
    .A2(_09608_));
 sg13g2_nor2_1 _15214_ (.A(net961),
    .B(_09130_),
    .Y(_09611_));
 sg13g2_a22oi_1 _15215_ (.Y(_09612_),
    .B1(_09611_),
    .B2(_09085_),
    .A2(_09294_),
    .A1(_09170_));
 sg13g2_o21ai_1 _15216_ (.B1(net1039),
    .Y(_09613_),
    .A1(net920),
    .A2(_09612_));
 sg13g2_nor2_1 _15217_ (.A(_09610_),
    .B(_09613_),
    .Y(_09614_));
 sg13g2_a221oi_1 _15218_ (.B2(_09607_),
    .C1(_09614_),
    .B1(_09187_),
    .A1(net919),
    .Y(_09615_),
    .A2(net1012));
 sg13g2_o21ai_1 _15219_ (.B1(_09615_),
    .Y(_09616_),
    .A1(_09598_),
    .A2(_09605_));
 sg13g2_nand2_1 _15220_ (.Y(_09617_),
    .A(_09161_),
    .B(_09305_));
 sg13g2_a22oi_1 _15221_ (.Y(_09618_),
    .B1(_09617_),
    .B2(net883),
    .A2(_09417_),
    .A1(net909));
 sg13g2_nand2_1 _15222_ (.Y(_09619_),
    .A(net886),
    .B(_09618_));
 sg13g2_nand2_1 _15223_ (.Y(_09620_),
    .A(_09108_),
    .B(_09417_));
 sg13g2_nand3_1 _15224_ (.B(_09144_),
    .C(_09620_),
    .A(net917),
    .Y(_09621_));
 sg13g2_nand4_1 _15225_ (.B(_09325_),
    .C(_09619_),
    .A(net913),
    .Y(_09622_),
    .D(_09621_));
 sg13g2_o21ai_1 _15226_ (.B1(_09622_),
    .Y(_09623_),
    .A1(net1019),
    .A2(_09616_));
 sg13g2_a221oi_1 _15227_ (.B2(net981),
    .C1(_09623_),
    .B1(_09597_),
    .A1(net890),
    .Y(_09624_),
    .A2(_09008_));
 sg13g2_a21oi_1 _15228_ (.A1(_09569_),
    .A2(net829),
    .Y(_00407_),
    .B1(_09624_));
 sg13g2_nor2_1 _15229_ (.A(_09077_),
    .B(_09194_),
    .Y(_09625_));
 sg13g2_nand3_1 _15230_ (.B(net930),
    .C(_09113_),
    .A(_09017_),
    .Y(_09626_));
 sg13g2_o21ai_1 _15231_ (.B1(_09626_),
    .Y(_09627_),
    .A1(_09174_),
    .A2(_09625_));
 sg13g2_o21ai_1 _15232_ (.B1(_09544_),
    .Y(_09628_),
    .A1(_09341_),
    .A2(_09084_));
 sg13g2_a21oi_1 _15233_ (.A1(net888),
    .A2(net885),
    .Y(_09629_),
    .B1(_09073_));
 sg13g2_nor4_1 _15234_ (.A(net886),
    .B(_09096_),
    .C(_09128_),
    .D(_09629_),
    .Y(_09630_));
 sg13g2_a221oi_1 _15235_ (.B2(net913),
    .C1(_09630_),
    .B1(_09628_),
    .A1(net882),
    .Y(_09631_),
    .A2(_09627_));
 sg13g2_nor2_1 _15236_ (.A(_09062_),
    .B(net1040),
    .Y(_09632_));
 sg13g2_a21oi_1 _15237_ (.A1(net1009),
    .A2(net930),
    .Y(_09633_),
    .B1(_09632_));
 sg13g2_nand4_1 _15238_ (.B(net910),
    .C(net972),
    .A(net924),
    .Y(_09634_),
    .D(net980));
 sg13g2_o21ai_1 _15239_ (.B1(_09634_),
    .Y(_09635_),
    .A1(net915),
    .A2(_09633_));
 sg13g2_a21oi_1 _15240_ (.A1(_09156_),
    .A2(_09367_),
    .Y(_09636_),
    .B1(_09161_));
 sg13g2_a22oi_1 _15241_ (.Y(_09637_),
    .B1(_09636_),
    .B2(net882),
    .A2(_09635_),
    .A1(net889));
 sg13g2_nand2_1 _15242_ (.Y(_09638_),
    .A(net910),
    .B(_09557_));
 sg13g2_o21ai_1 _15243_ (.B1(_09638_),
    .Y(_09639_),
    .A1(net962),
    .A2(net1009));
 sg13g2_nand2_1 _15244_ (.Y(_09640_),
    .A(net1009),
    .B(_09244_));
 sg13g2_o21ai_1 _15245_ (.B1(_09640_),
    .Y(_09641_),
    .A1(net1009),
    .A2(_09085_));
 sg13g2_nor3_1 _15246_ (.A(net889),
    .B(net980),
    .C(_09252_),
    .Y(_09642_));
 sg13g2_a221oi_1 _15247_ (.B2(_09275_),
    .C1(_09642_),
    .B1(_09641_),
    .A1(_09276_),
    .Y(_09643_),
    .A2(_09639_));
 sg13g2_mux2_1 _15248_ (.A0(_09637_),
    .A1(_09643_),
    .S(_09341_),
    .X(_09644_));
 sg13g2_a21oi_1 _15249_ (.A1(_09130_),
    .A2(_09293_),
    .Y(_09645_),
    .B1(_09448_));
 sg13g2_a21oi_1 _15250_ (.A1(net929),
    .A2(_09286_),
    .Y(_09646_),
    .B1(_09037_));
 sg13g2_a21oi_1 _15251_ (.A1(net930),
    .A2(net966),
    .Y(_09647_),
    .B1(net964));
 sg13g2_o21ai_1 _15252_ (.B1(_09647_),
    .Y(_09648_),
    .A1(_09246_),
    .A2(_09646_));
 sg13g2_o21ai_1 _15253_ (.B1(_09523_),
    .Y(_09649_),
    .A1(_09041_),
    .A2(_09233_));
 sg13g2_a22oi_1 _15254_ (.Y(_09650_),
    .B1(_09649_),
    .B2(net920),
    .A2(net912),
    .A1(net931));
 sg13g2_a221oi_1 _15255_ (.B2(net924),
    .C1(net977),
    .B1(_09281_),
    .A1(net910),
    .Y(_09651_),
    .A2(net912));
 sg13g2_a21oi_1 _15256_ (.A1(net911),
    .A2(_09650_),
    .Y(_09652_),
    .B1(_09651_));
 sg13g2_a21oi_1 _15257_ (.A1(net914),
    .A2(_09185_),
    .Y(_09653_),
    .B1(net923));
 sg13g2_nand2b_1 _15258_ (.Y(_09654_),
    .B(_09653_),
    .A_N(_09652_));
 sg13g2_o21ai_1 _15259_ (.B1(_09654_),
    .Y(_09655_),
    .A1(_09645_),
    .A2(_09648_));
 sg13g2_o21ai_1 _15260_ (.B1(_09412_),
    .Y(_09656_),
    .A1(net921),
    .A2(_09161_));
 sg13g2_a22oi_1 _15261_ (.Y(_09657_),
    .B1(_09072_),
    .B2(net927),
    .A2(_09024_),
    .A1(net910));
 sg13g2_o21ai_1 _15262_ (.B1(net908),
    .Y(_09658_),
    .A1(net915),
    .A2(_09657_));
 sg13g2_a21o_1 _15263_ (.A2(_09656_),
    .A1(net917),
    .B1(_09658_),
    .X(_09659_));
 sg13g2_nand3_1 _15264_ (.B(_09476_),
    .C(_09659_),
    .A(_09135_),
    .Y(_09660_));
 sg13g2_mux4_1 _15265_ (.S0(net963),
    .A0(_09631_),
    .A1(_09644_),
    .A2(_09655_),
    .A3(_09660_),
    .S1(_09014_),
    .X(_09661_));
 sg13g2_nand2_1 _15266_ (.Y(_09662_),
    .A(net1020),
    .B(net828));
 sg13g2_o21ai_1 _15267_ (.B1(_09662_),
    .Y(_00408_),
    .A1(net829),
    .A2(_09661_));
 sg13g2_buf_1 _15268_ (.A(net1101),
    .X(_09663_));
 sg13g2_nand2_2 _15269_ (.Y(_09664_),
    .A(_08199_),
    .B(\top_ihp.oisc.micro_state[2] ));
 sg13g2_nand3_1 _15270_ (.B(_09006_),
    .C(_09664_),
    .A(_00091_),
    .Y(_09665_));
 sg13g2_nand2_1 _15271_ (.Y(_09666_),
    .A(_09663_),
    .B(_09665_));
 sg13g2_buf_1 _15272_ (.A(_09666_),
    .X(_09667_));
 sg13g2_buf_1 _15273_ (.A(_09667_),
    .X(_09668_));
 sg13g2_buf_1 _15274_ (.A(\top_ihp.oisc.state[3] ),
    .X(_09669_));
 sg13g2_buf_1 _15275_ (.A(_09669_),
    .X(_09670_));
 sg13g2_buf_1 _15276_ (.A(_09670_),
    .X(_09671_));
 sg13g2_inv_1 _15277_ (.Y(_09672_),
    .A(\top_ihp.oisc.op_b[31] ));
 sg13g2_buf_4 _15278_ (.X(_09673_),
    .A(\top_ihp.oisc.op_a[31] ));
 sg13g2_nor2_1 _15279_ (.A(_09672_),
    .B(_09673_),
    .Y(_09674_));
 sg13g2_nand3_1 _15280_ (.B(_08306_),
    .C(_08483_),
    .A(_08352_),
    .Y(_09675_));
 sg13g2_buf_1 _15281_ (.A(_09675_),
    .X(_09676_));
 sg13g2_xnor2_1 _15282_ (.Y(_09677_),
    .A(net1058),
    .B(_08219_));
 sg13g2_nand2_1 _15283_ (.Y(_09678_),
    .A(_09677_),
    .B(_08492_));
 sg13g2_nor3_1 _15284_ (.A(_09678_),
    .B(_08491_),
    .C(_08499_),
    .Y(_09679_));
 sg13g2_nand3_1 _15285_ (.B(_08397_),
    .C(_09679_),
    .A(_08309_),
    .Y(_09680_));
 sg13g2_xor2_1 _15286_ (.B(_08545_),
    .A(\top_ihp.oisc.op_b[30] ),
    .X(_09681_));
 sg13g2_or3_1 _15287_ (.A(_08556_),
    .B(_08560_),
    .C(_09681_),
    .X(_09682_));
 sg13g2_nand2_1 _15288_ (.Y(_09683_),
    .A(_08323_),
    .B(_08614_));
 sg13g2_xor2_1 _15289_ (.B(_08319_),
    .A(_08317_),
    .X(_09684_));
 sg13g2_nor2_1 _15290_ (.A(_09683_),
    .B(_09684_),
    .Y(_09685_));
 sg13g2_xor2_1 _15291_ (.B(_08328_),
    .A(_08326_),
    .X(_09686_));
 sg13g2_nand2b_1 _15292_ (.Y(_09687_),
    .B(_08334_),
    .A_N(_08331_));
 sg13g2_xor2_1 _15293_ (.B(_09673_),
    .A(\top_ihp.oisc.op_b[31] ),
    .X(_09688_));
 sg13g2_nor3_1 _15294_ (.A(_09686_),
    .B(_09687_),
    .C(_09688_),
    .Y(_09689_));
 sg13g2_nand2_1 _15295_ (.Y(_09690_),
    .A(_09685_),
    .B(_09689_));
 sg13g2_or3_1 _15296_ (.A(_08348_),
    .B(_08505_),
    .C(_09690_),
    .X(_09691_));
 sg13g2_nor4_1 _15297_ (.A(_09676_),
    .B(_09680_),
    .C(_09682_),
    .D(_09691_),
    .Y(_09692_));
 sg13g2_inv_1 _15298_ (.Y(_09693_),
    .A(_08545_));
 sg13g2_nand3_1 _15299_ (.B(_08552_),
    .C(_08561_),
    .A(_09693_),
    .Y(_09694_));
 sg13g2_nand3_1 _15300_ (.B(_08552_),
    .C(_08561_),
    .A(\top_ihp.oisc.op_b[30] ),
    .Y(_09695_));
 sg13g2_a21oi_1 _15301_ (.A1(_09694_),
    .A2(_09695_),
    .Y(_09696_),
    .B1(_08550_));
 sg13g2_a21o_1 _15302_ (.A2(_08545_),
    .A1(_08549_),
    .B1(_08576_),
    .X(_09697_));
 sg13g2_o21ai_1 _15303_ (.B1(_09697_),
    .Y(_09698_),
    .A1(_08549_),
    .A2(net1026));
 sg13g2_nor3_1 _15304_ (.A(_09673_),
    .B(_09696_),
    .C(_09698_),
    .Y(_09699_));
 sg13g2_nor3_1 _15305_ (.A(_09672_),
    .B(_09696_),
    .C(_09698_),
    .Y(_09700_));
 sg13g2_nor4_2 _15306_ (.A(_09674_),
    .B(_09692_),
    .C(_09699_),
    .Y(_09701_),
    .D(_09700_));
 sg13g2_or2_1 _15307_ (.X(_09702_),
    .B(_09701_),
    .A(_08203_));
 sg13g2_or3_1 _15308_ (.A(net1008),
    .B(net892),
    .C(_09664_),
    .X(_09703_));
 sg13g2_buf_1 _15309_ (.A(_09703_),
    .X(_09704_));
 sg13g2_nor2_1 _15310_ (.A(net882),
    .B(_09704_),
    .Y(_09705_));
 sg13g2_a22oi_1 _15311_ (.Y(_09706_),
    .B1(_09702_),
    .B2(_09705_),
    .A2(\top_ihp.oisc.decoder.decoded[0] ),
    .A1(net960));
 sg13g2_nor2_1 _15312_ (.A(_09702_),
    .B(_09704_),
    .Y(_09707_));
 sg13g2_o21ai_1 _15313_ (.B1(net882),
    .Y(_09708_),
    .A1(_09667_),
    .A2(_09707_));
 sg13g2_o21ai_1 _15314_ (.B1(_09708_),
    .Y(_00409_),
    .A1(net792),
    .A2(_09706_));
 sg13g2_nor2b_1 _15315_ (.A(_08202_),
    .B_N(_08203_),
    .Y(_09709_));
 sg13g2_nand2_1 _15316_ (.Y(_09710_),
    .A(_08203_),
    .B(_09026_));
 sg13g2_and2_1 _15317_ (.A(_08202_),
    .B(_09710_),
    .X(_09711_));
 sg13g2_mux2_1 _15318_ (.A0(_09711_),
    .A1(_09313_),
    .S(_09701_),
    .X(_09712_));
 sg13g2_a21oi_1 _15319_ (.A1(_09313_),
    .A2(_09709_),
    .Y(_09713_),
    .B1(_09712_));
 sg13g2_or4_1 _15320_ (.A(net886),
    .B(_09667_),
    .C(_09704_),
    .D(_09713_),
    .X(_09714_));
 sg13g2_nor3_1 _15321_ (.A(net1008),
    .B(net892),
    .C(_09664_),
    .Y(_09715_));
 sg13g2_buf_2 _15322_ (.A(_09715_),
    .X(_09716_));
 sg13g2_nand3_1 _15323_ (.B(_09716_),
    .C(_09713_),
    .A(net886),
    .Y(_09717_));
 sg13g2_and4_1 _15324_ (.A(net1008),
    .B(_09663_),
    .C(\top_ihp.oisc.decoder.decoded[1] ),
    .D(_09665_),
    .X(_09718_));
 sg13g2_a21oi_1 _15325_ (.A1(_09064_),
    .A2(_09667_),
    .Y(_09719_),
    .B1(_09718_));
 sg13g2_nand3_1 _15326_ (.B(_09717_),
    .C(_09719_),
    .A(_09714_),
    .Y(_00410_));
 sg13g2_buf_1 _15327_ (.A(_09701_),
    .X(_09720_));
 sg13g2_xnor2_1 _15328_ (.Y(_09721_),
    .A(net967),
    .B(_09130_));
 sg13g2_nand2_1 _15329_ (.Y(_09722_),
    .A(_09032_),
    .B(_09710_));
 sg13g2_a22oi_1 _15330_ (.Y(_09723_),
    .B1(_09722_),
    .B2(_08202_),
    .A2(net925),
    .A1(_08203_));
 sg13g2_xor2_1 _15331_ (.B(net920),
    .A(_08205_),
    .X(_09724_));
 sg13g2_xnor2_1 _15332_ (.Y(_09725_),
    .A(_09723_),
    .B(_09724_));
 sg13g2_nor2_1 _15333_ (.A(net732),
    .B(_09725_),
    .Y(_09726_));
 sg13g2_a21oi_1 _15334_ (.A1(net732),
    .A2(_09721_),
    .Y(_09727_),
    .B1(_09726_));
 sg13g2_a221oi_1 _15335_ (.B2(_09727_),
    .C1(net792),
    .B1(_09716_),
    .A1(net960),
    .Y(_09728_),
    .A2(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_a21oi_1 _15336_ (.A1(net909),
    .A2(net792),
    .Y(_00411_),
    .B1(_09728_));
 sg13g2_nor2_1 _15337_ (.A(_09286_),
    .B(_09163_),
    .Y(_09729_));
 sg13g2_xnor2_1 _15338_ (.Y(_09730_),
    .A(_09180_),
    .B(_09729_));
 sg13g2_nand2_1 _15339_ (.Y(_09731_),
    .A(_08205_),
    .B(_09028_));
 sg13g2_nor2_1 _15340_ (.A(_08205_),
    .B(net1038),
    .Y(_09732_));
 sg13g2_a21oi_2 _15341_ (.B1(_09732_),
    .Y(_09733_),
    .A2(_09731_),
    .A1(_09723_));
 sg13g2_xnor2_1 _15342_ (.Y(_09734_),
    .A(_08204_),
    .B(_09025_));
 sg13g2_xnor2_1 _15343_ (.Y(_09735_),
    .A(_09733_),
    .B(_09734_));
 sg13g2_nor2_1 _15344_ (.A(net732),
    .B(_09735_),
    .Y(_09736_));
 sg13g2_a21oi_1 _15345_ (.A1(net732),
    .A2(_09730_),
    .Y(_09737_),
    .B1(_09736_));
 sg13g2_a221oi_1 _15346_ (.B2(_09737_),
    .C1(net792),
    .B1(_09716_),
    .A1(net960),
    .Y(_09738_),
    .A2(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_a21oi_1 _15347_ (.A1(net926),
    .A2(net792),
    .Y(_00412_),
    .B1(_09738_));
 sg13g2_or2_1 _15348_ (.X(_09739_),
    .B(_09294_),
    .A(_09163_));
 sg13g2_buf_1 _15349_ (.A(_09739_),
    .X(_09740_));
 sg13g2_xnor2_1 _15350_ (.Y(_09741_),
    .A(_09214_),
    .B(_09740_));
 sg13g2_nor2_1 _15351_ (.A(net1017),
    .B(_09733_),
    .Y(_09742_));
 sg13g2_a21oi_1 _15352_ (.A1(_09022_),
    .A2(_09733_),
    .Y(_09743_),
    .B1(_08204_));
 sg13g2_nor2_1 _15353_ (.A(_09742_),
    .B(_09743_),
    .Y(_09744_));
 sg13g2_xnor2_1 _15354_ (.Y(_09745_),
    .A(_08206_),
    .B(_09051_));
 sg13g2_xnor2_1 _15355_ (.Y(_09746_),
    .A(_09744_),
    .B(_09745_));
 sg13g2_nor2_1 _15356_ (.A(net732),
    .B(_09746_),
    .Y(_09747_));
 sg13g2_a21oi_1 _15357_ (.A1(net732),
    .A2(_09741_),
    .Y(_09748_),
    .B1(_09747_));
 sg13g2_a221oi_1 _15358_ (.B2(_09748_),
    .C1(_09667_),
    .B1(_09716_),
    .A1(net960),
    .Y(_09749_),
    .A2(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_a21oi_1 _15359_ (.A1(net881),
    .A2(net792),
    .Y(_00413_),
    .B1(_09749_));
 sg13g2_nor2_1 _15360_ (.A(_09296_),
    .B(_09744_),
    .Y(_09750_));
 sg13g2_a21oi_1 _15361_ (.A1(net961),
    .A2(_09744_),
    .Y(_09751_),
    .B1(_08206_));
 sg13g2_nor2_2 _15362_ (.A(_09750_),
    .B(_09751_),
    .Y(_09752_));
 sg13g2_nand2_1 _15363_ (.Y(_09753_),
    .A(_08207_),
    .B(_09017_));
 sg13g2_nand2_1 _15364_ (.Y(_09754_),
    .A(_09567_),
    .B(_09126_));
 sg13g2_and2_1 _15365_ (.A(_09753_),
    .B(_09754_),
    .X(_09755_));
 sg13g2_xnor2_1 _15366_ (.Y(_09756_),
    .A(_09752_),
    .B(_09755_));
 sg13g2_nor2_1 _15367_ (.A(_09267_),
    .B(_09740_),
    .Y(_09757_));
 sg13g2_xnor2_1 _15368_ (.Y(_09758_),
    .A(_09135_),
    .B(_09757_));
 sg13g2_mux2_1 _15369_ (.A0(_09756_),
    .A1(_09758_),
    .S(_09720_),
    .X(_09759_));
 sg13g2_a221oi_1 _15370_ (.B2(_09759_),
    .C1(_09667_),
    .B1(_09716_),
    .A1(net960),
    .Y(_09760_),
    .A2(\top_ihp.oisc.decoder.decoded[5] ));
 sg13g2_a21oi_1 _15371_ (.A1(net933),
    .A2(net792),
    .Y(_00414_),
    .B1(_09760_));
 sg13g2_mux2_1 _15372_ (.A0(_09753_),
    .A1(_09754_),
    .S(_09752_),
    .X(_09761_));
 sg13g2_xnor2_1 _15373_ (.Y(_09762_),
    .A(_09020_),
    .B(_09761_));
 sg13g2_nor2_1 _15374_ (.A(_09174_),
    .B(_09740_),
    .Y(_09763_));
 sg13g2_xnor2_1 _15375_ (.Y(_09764_),
    .A(_00213_),
    .B(_09763_));
 sg13g2_mux2_1 _15376_ (.A0(_09762_),
    .A1(_09764_),
    .S(net732),
    .X(_09765_));
 sg13g2_a221oi_1 _15377_ (.B2(_09765_),
    .C1(_09667_),
    .B1(_09716_),
    .A1(net960),
    .Y(_09766_),
    .A2(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_a21oi_1 _15378_ (.A1(_09106_),
    .A2(net792),
    .Y(_00415_),
    .B1(_09766_));
 sg13g2_and2_1 _15379_ (.A(_08207_),
    .B(_09498_),
    .X(_09767_));
 sg13g2_nand2_1 _15380_ (.Y(_09768_),
    .A(_09126_),
    .B(net1039));
 sg13g2_nor2_1 _15381_ (.A(_08207_),
    .B(_09768_),
    .Y(_09769_));
 sg13g2_mux2_1 _15382_ (.A0(_09767_),
    .A1(_09769_),
    .S(_09752_),
    .X(_09770_));
 sg13g2_xnor2_1 _15383_ (.Y(_09771_),
    .A(_09012_),
    .B(_09770_));
 sg13g2_nor4_1 _15384_ (.A(_09286_),
    .B(_09297_),
    .C(_09163_),
    .D(_09768_),
    .Y(_09772_));
 sg13g2_xnor2_1 _15385_ (.Y(_09773_),
    .A(_00212_),
    .B(_09772_));
 sg13g2_nand2_1 _15386_ (.Y(_09774_),
    .A(net732),
    .B(_09773_));
 sg13g2_o21ai_1 _15387_ (.B1(_09774_),
    .Y(_09775_),
    .A1(_09720_),
    .A2(_09771_));
 sg13g2_a22oi_1 _15388_ (.Y(_09776_),
    .B1(_09716_),
    .B2(_09775_),
    .A2(\top_ihp.oisc.decoder.decoded[7] ),
    .A1(net960));
 sg13g2_nand2_1 _15389_ (.Y(_09777_),
    .A(net981),
    .B(_09668_));
 sg13g2_o21ai_1 _15390_ (.B1(_09777_),
    .Y(_00416_),
    .A1(_09668_),
    .A2(_09776_));
 sg13g2_inv_1 _15391_ (.Y(_09778_),
    .A(\top_ihp.oisc.micro_state[2] ));
 sg13g2_buf_1 _15392_ (.A(net1032),
    .X(_09779_));
 sg13g2_mux2_1 _15393_ (.A0(_13698_),
    .A1(_09778_),
    .S(net959),
    .X(_00417_));
 sg13g2_nand2b_1 _15394_ (.Y(_09780_),
    .B(\top_ihp.oisc.micro_state[1] ),
    .A_N(net959));
 sg13g2_o21ai_1 _15395_ (.B1(_09780_),
    .Y(_00418_),
    .A1(_08211_),
    .A2(_09008_));
 sg13g2_nand2_1 _15396_ (.Y(_09781_),
    .A(_09006_),
    .B(_08987_));
 sg13g2_o21ai_1 _15397_ (.B1(_09781_),
    .Y(_00419_),
    .A1(net959),
    .A2(_09778_));
 sg13g2_buf_1 _15398_ (.A(\top_ihp.oisc.state[2] ),
    .X(_09782_));
 sg13g2_or2_1 _15399_ (.X(_09783_),
    .B(_09669_),
    .A(net1037));
 sg13g2_buf_2 _15400_ (.A(_09783_),
    .X(_09784_));
 sg13g2_buf_1 _15401_ (.A(_09784_),
    .X(_09785_));
 sg13g2_buf_1 _15402_ (.A(_09785_),
    .X(_09786_));
 sg13g2_buf_2 _15403_ (.A(\top_ihp.oisc.state[4] ),
    .X(_09787_));
 sg13g2_buf_1 _15404_ (.A(_09787_),
    .X(_09788_));
 sg13g2_buf_1 _15405_ (.A(net1007),
    .X(_09789_));
 sg13g2_buf_1 _15406_ (.A(\top_ihp.oisc.decoder.decoded[13] ),
    .X(_09790_));
 sg13g2_buf_1 _15407_ (.A(net1036),
    .X(_09791_));
 sg13g2_buf_2 _15408_ (.A(_00090_),
    .X(_09792_));
 sg13g2_buf_1 _15409_ (.A(_09792_),
    .X(_09793_));
 sg13g2_buf_1 _15410_ (.A(\top_ihp.oisc.decoder.instruction[7] ),
    .X(_09794_));
 sg13g2_nand3_1 _15411_ (.B(_09793_),
    .C(_09794_),
    .A(_09791_),
    .Y(_09795_));
 sg13g2_buf_1 _15412_ (.A(\top_ihp.oisc.decoder.instruction[20] ),
    .X(_09796_));
 sg13g2_buf_1 _15413_ (.A(\top_ihp.oisc.decoder.decoded[15] ),
    .X(_09797_));
 sg13g2_nand2_1 _15414_ (.Y(_09798_),
    .A(net1006),
    .B(_09797_));
 sg13g2_inv_2 _15415_ (.Y(_09799_),
    .A(_09790_));
 sg13g2_nand2_1 _15416_ (.Y(_09800_),
    .A(_09799_),
    .B(_09792_));
 sg13g2_o21ai_1 _15417_ (.B1(_09800_),
    .Y(_09801_),
    .A1(net1005),
    .A2(_09798_));
 sg13g2_nand2_1 _15418_ (.Y(_09802_),
    .A(_09796_),
    .B(_09801_));
 sg13g2_buf_1 _15419_ (.A(\top_ihp.oisc.decoder.decoded[14] ),
    .X(_09803_));
 sg13g2_buf_1 _15420_ (.A(_09803_),
    .X(_09804_));
 sg13g2_a21oi_1 _15421_ (.A1(_09795_),
    .A2(_09802_),
    .Y(_09805_),
    .B1(net1004));
 sg13g2_buf_1 _15422_ (.A(\top_ihp.oisc.mem_addr_lowbits[0] ),
    .X(_09806_));
 sg13g2_nor2_1 _15423_ (.A(_08656_),
    .B(_08657_),
    .Y(_09807_));
 sg13g2_and2_1 _15424_ (.A(_09806_),
    .B(_09807_),
    .X(_09808_));
 sg13g2_buf_1 _15425_ (.A(_09808_),
    .X(_09809_));
 sg13g2_buf_1 _15426_ (.A(\top_ihp.oisc.mem_addr_lowbits[1] ),
    .X(_09810_));
 sg13g2_buf_1 _15427_ (.A(_09810_),
    .X(_09811_));
 sg13g2_nand2b_1 _15428_ (.Y(_09812_),
    .B(_00080_),
    .A_N(_08968_));
 sg13g2_buf_1 _15429_ (.A(_09812_),
    .X(_09813_));
 sg13g2_buf_1 _15430_ (.A(net957),
    .X(_09814_));
 sg13g2_buf_8 _15431_ (.A(net861),
    .X(_09815_));
 sg13g2_buf_1 _15432_ (.A(net845),
    .X(_09816_));
 sg13g2_buf_1 _15433_ (.A(net827),
    .X(_09817_));
 sg13g2_buf_1 _15434_ (.A(_08951_),
    .X(_09818_));
 sg13g2_and3_1 _15435_ (.X(_09819_),
    .A(net1021),
    .B(net879),
    .C(net891));
 sg13g2_buf_1 _15436_ (.A(_09819_),
    .X(_09820_));
 sg13g2_buf_1 _15437_ (.A(_09820_),
    .X(_09821_));
 sg13g2_buf_1 _15438_ (.A(_09821_),
    .X(_09822_));
 sg13g2_buf_1 _15439_ (.A(_08959_),
    .X(_09823_));
 sg13g2_buf_1 _15440_ (.A(_09823_),
    .X(_09824_));
 sg13g2_buf_1 _15441_ (.A(net956),
    .X(_09825_));
 sg13g2_inv_1 _15442_ (.Y(_09826_),
    .A(_00161_));
 sg13g2_buf_1 _15443_ (.A(_08962_),
    .X(_09827_));
 sg13g2_buf_1 _15444_ (.A(_09827_),
    .X(_09828_));
 sg13g2_buf_1 _15445_ (.A(net878),
    .X(_09829_));
 sg13g2_buf_1 _15446_ (.A(_09820_),
    .X(_09830_));
 sg13g2_a221oi_1 _15447_ (.B2(\top_ihp.wb_coproc.dat_o[24] ),
    .C1(net825),
    .B1(_09829_),
    .A1(_09825_),
    .Y(_09831_),
    .A2(_09826_));
 sg13g2_a21oi_1 _15448_ (.A1(_00160_),
    .A2(net790),
    .Y(_09832_),
    .B1(_09831_));
 sg13g2_buf_1 _15449_ (.A(net845),
    .X(_09833_));
 sg13g2_nor2_1 _15450_ (.A(_00159_),
    .B(net824),
    .Y(_09834_));
 sg13g2_a21oi_1 _15451_ (.A1(_09817_),
    .A2(_09832_),
    .Y(_09835_),
    .B1(_09834_));
 sg13g2_nor2_2 _15452_ (.A(net906),
    .B(_09835_),
    .Y(_09836_));
 sg13g2_inv_1 _15453_ (.Y(_09837_),
    .A(_00137_));
 sg13g2_a221oi_1 _15454_ (.B2(\top_ihp.wb_coproc.dat_o[8] ),
    .C1(_09821_),
    .B1(net878),
    .A1(net956),
    .Y(_09838_),
    .A2(_09837_));
 sg13g2_a21oi_1 _15455_ (.A1(_00136_),
    .A2(net825),
    .Y(_09839_),
    .B1(_09838_));
 sg13g2_nor2_1 _15456_ (.A(_00135_),
    .B(net845),
    .Y(_09840_));
 sg13g2_a21oi_1 _15457_ (.A1(net827),
    .A2(_09839_),
    .Y(_09841_),
    .B1(_09840_));
 sg13g2_nand2b_1 _15458_ (.Y(_09842_),
    .B(_08970_),
    .A_N(_09841_));
 sg13g2_nor2_1 _15459_ (.A(net1035),
    .B(_09842_),
    .Y(_09843_));
 sg13g2_a21o_1 _15460_ (.A2(_09836_),
    .A1(net1003),
    .B1(_09843_),
    .X(_09844_));
 sg13g2_nor2b_1 _15461_ (.A(_08656_),
    .B_N(_09806_),
    .Y(_09845_));
 sg13g2_buf_1 _15462_ (.A(_09845_),
    .X(_09846_));
 sg13g2_inv_1 _15463_ (.Y(_09847_),
    .A(_08657_));
 sg13g2_buf_1 _15464_ (.A(_09847_),
    .X(_09848_));
 sg13g2_o21ai_1 _15465_ (.B1(net954),
    .Y(_09849_),
    .A1(net1035),
    .A2(net955));
 sg13g2_buf_1 _15466_ (.A(net1024),
    .X(_09850_));
 sg13g2_and2_1 _15467_ (.A(net953),
    .B(net862),
    .X(_09851_));
 sg13g2_buf_1 _15468_ (.A(_09851_),
    .X(_09852_));
 sg13g2_buf_1 _15469_ (.A(net846),
    .X(_09853_));
 sg13g2_nor2_1 _15470_ (.A(\top_ihp.wb_dati_ram[0] ),
    .B(net823),
    .Y(_09854_));
 sg13g2_a221oi_1 _15471_ (.B2(net859),
    .C1(net790),
    .B1(\top_ihp.wb_coproc.dat_o[0] ),
    .A1(net905),
    .Y(_09855_),
    .A2(\top_ihp.wb_dati_spi[0] ));
 sg13g2_nor3_1 _15472_ (.A(_09852_),
    .B(_09854_),
    .C(_09855_),
    .Y(_09856_));
 sg13g2_a21oi_1 _15473_ (.A1(\top_ihp.wb_dati_rom[0] ),
    .A2(_09852_),
    .Y(_09857_),
    .B1(_09856_));
 sg13g2_nand2_1 _15474_ (.Y(_09858_),
    .A(_08968_),
    .B(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_o21ai_1 _15475_ (.B1(_09858_),
    .Y(_09859_),
    .A1(_08968_),
    .A2(_09857_));
 sg13g2_buf_1 _15476_ (.A(_08973_),
    .X(_09860_));
 sg13g2_mux2_1 _15477_ (.A0(_09859_),
    .A1(\top_ihp.wb_dati_uart[0] ),
    .S(_09860_),
    .X(_09861_));
 sg13g2_nor2_1 _15478_ (.A(_00120_),
    .B(_08945_),
    .Y(_09862_));
 sg13g2_inv_1 _15479_ (.Y(_09863_),
    .A(_00122_));
 sg13g2_a22oi_1 _15480_ (.Y(_09864_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[16] ),
    .A2(_09863_),
    .A1(net1002));
 sg13g2_and4_1 _15481_ (.A(net1021),
    .B(_00121_),
    .C(net879),
    .D(net891),
    .X(_09865_));
 sg13g2_a221oi_1 _15482_ (.B2(_09864_),
    .C1(_09865_),
    .B1(net846),
    .A1(_08942_),
    .Y(_09866_),
    .A2(net862));
 sg13g2_o21ai_1 _15483_ (.B1(_08975_),
    .Y(_09867_),
    .A1(_09862_),
    .A2(_09866_));
 sg13g2_buf_2 _15484_ (.A(_09867_),
    .X(_09868_));
 sg13g2_nand2b_1 _15485_ (.Y(_09869_),
    .B(_09806_),
    .A_N(_08656_));
 sg13g2_inv_1 _15486_ (.Y(_09870_),
    .A(net1035));
 sg13g2_buf_1 _15487_ (.A(_09870_),
    .X(_09871_));
 sg13g2_nor2_1 _15488_ (.A(_08657_),
    .B(_09871_),
    .Y(_09872_));
 sg13g2_buf_1 _15489_ (.A(_09872_),
    .X(_09873_));
 sg13g2_nand2_1 _15490_ (.Y(_09874_),
    .A(_09869_),
    .B(net877));
 sg13g2_and2_1 _15491_ (.A(_08415_),
    .B(_09001_),
    .X(_09875_));
 sg13g2_buf_1 _15492_ (.A(_09875_),
    .X(_09876_));
 sg13g2_buf_1 _15493_ (.A(_09876_),
    .X(_09877_));
 sg13g2_o21ai_1 _15494_ (.B1(net903),
    .Y(_09878_),
    .A1(_09868_),
    .A2(_09874_));
 sg13g2_a221oi_1 _15495_ (.B2(_09861_),
    .C1(_09878_),
    .B1(_09849_),
    .A1(_09809_),
    .Y(_09879_),
    .A2(_09844_));
 sg13g2_inv_2 _15496_ (.Y(_09880_),
    .A(_09787_));
 sg13g2_o21ai_1 _15497_ (.B1(_09880_),
    .Y(_09881_),
    .A1(_09683_),
    .A2(net903));
 sg13g2_nor2_1 _15498_ (.A(_09879_),
    .B(_09881_),
    .Y(_09882_));
 sg13g2_a21oi_1 _15499_ (.A1(net958),
    .A2(_09805_),
    .Y(_09883_),
    .B1(_09882_));
 sg13g2_buf_1 _15500_ (.A(_09785_),
    .X(_09884_));
 sg13g2_nand2_1 _15501_ (.Y(_09885_),
    .A(_08321_),
    .B(net876));
 sg13g2_o21ai_1 _15502_ (.B1(_09885_),
    .Y(_09886_),
    .A1(net880),
    .A2(_09883_));
 sg13g2_buf_2 _15503_ (.A(_09886_),
    .X(_09887_));
 sg13g2_buf_1 _15504_ (.A(_09887_),
    .X(_09888_));
 sg13g2_buf_1 _15505_ (.A(net143),
    .X(_09889_));
 sg13g2_nor2b_1 _15506_ (.A(_09790_),
    .B_N(_09797_),
    .Y(_09890_));
 sg13g2_buf_1 _15507_ (.A(_09890_),
    .X(_09891_));
 sg13g2_nand2_1 _15508_ (.Y(_09892_),
    .A(net1004),
    .B(_09891_));
 sg13g2_buf_1 _15509_ (.A(\top_ihp.oisc.decoder.decoded[12] ),
    .X(_09893_));
 sg13g2_a221oi_1 _15510_ (.B2(_09893_),
    .C1(_09664_),
    .B1(_08210_),
    .A1(_08415_),
    .Y(_09894_),
    .A2(_09001_));
 sg13g2_buf_2 _15511_ (.A(_09894_),
    .X(_09895_));
 sg13g2_nand2_1 _15512_ (.Y(_09896_),
    .A(_08415_),
    .B(_09001_));
 sg13g2_buf_2 _15513_ (.A(_09896_),
    .X(_09897_));
 sg13g2_nand3_1 _15514_ (.B(_09893_),
    .C(_08210_),
    .A(_08199_),
    .Y(_09898_));
 sg13g2_xor2_1 _15515_ (.B(net1036),
    .A(_09803_),
    .X(_09899_));
 sg13g2_a22oi_1 _15516_ (.Y(_09900_),
    .B1(_09899_),
    .B2(_09792_),
    .A2(_09898_),
    .A1(_09897_));
 sg13g2_buf_2 _15517_ (.A(_09900_),
    .X(_09901_));
 sg13g2_buf_1 _15518_ (.A(\top_ihp.oisc.decoder.instruction[10] ),
    .X(_09902_));
 sg13g2_a22oi_1 _15519_ (.Y(_09903_),
    .B1(_09901_),
    .B2(_09902_),
    .A2(_09895_),
    .A1(\top_ihp.oisc.micro_res_addr[3] ));
 sg13g2_nor2_1 _15520_ (.A(_09787_),
    .B(_09903_),
    .Y(_09904_));
 sg13g2_a21oi_2 _15521_ (.B1(_09904_),
    .Y(_09905_),
    .A2(_09892_),
    .A1(net1007));
 sg13g2_buf_1 _15522_ (.A(\top_ihp.oisc.decoder.instruction[9] ),
    .X(_09906_));
 sg13g2_a221oi_1 _15523_ (.B2(_09906_),
    .C1(_09787_),
    .B1(_09901_),
    .A1(\top_ihp.oisc.micro_res_addr[2] ),
    .Y(_09907_),
    .A2(_09895_));
 sg13g2_a21oi_1 _15524_ (.A1(_09787_),
    .A2(_09892_),
    .Y(_09908_),
    .B1(_09907_));
 sg13g2_nor2_1 _15525_ (.A(net1008),
    .B(_09908_),
    .Y(_09909_));
 sg13g2_buf_2 _15526_ (.A(_09909_),
    .X(_09910_));
 sg13g2_and2_1 _15527_ (.A(_09905_),
    .B(_09910_),
    .X(_09911_));
 sg13g2_buf_1 _15528_ (.A(_09911_),
    .X(_09912_));
 sg13g2_buf_1 _15529_ (.A(_00092_),
    .X(_09913_));
 sg13g2_nand2b_1 _15530_ (.Y(_09914_),
    .B(_09913_),
    .A_N(_09912_));
 sg13g2_buf_1 _15531_ (.A(_09914_),
    .X(_09915_));
 sg13g2_nand2b_1 _15532_ (.Y(_09916_),
    .B(_09913_),
    .A_N(_09669_));
 sg13g2_nor2_1 _15533_ (.A(_09787_),
    .B(_09916_),
    .Y(_09917_));
 sg13g2_nor2b_1 _15534_ (.A(_09895_),
    .B_N(_09917_),
    .Y(_09918_));
 sg13g2_buf_1 _15535_ (.A(\top_ihp.oisc.decoder.instruction[11] ),
    .X(_09919_));
 sg13g2_nand3_1 _15536_ (.B(_09901_),
    .C(_09917_),
    .A(_09919_),
    .Y(_09920_));
 sg13g2_buf_1 _15537_ (.A(_09920_),
    .X(_09921_));
 sg13g2_nor2_2 _15538_ (.A(_09787_),
    .B(_09784_),
    .Y(_09922_));
 sg13g2_buf_2 _15539_ (.A(\top_ihp.oisc.state[0] ),
    .X(_09923_));
 sg13g2_buf_2 _15540_ (.A(_09923_),
    .X(_09924_));
 sg13g2_a21oi_1 _15541_ (.A1(_09893_),
    .A2(_09001_),
    .Y(_09925_),
    .B1(net1000));
 sg13g2_nand3_1 _15542_ (.B(_09922_),
    .C(_09925_),
    .A(_09664_),
    .Y(_09926_));
 sg13g2_nand2_1 _15543_ (.Y(_09927_),
    .A(_09921_),
    .B(_09926_));
 sg13g2_nor2_1 _15544_ (.A(_09918_),
    .B(_09927_),
    .Y(_09928_));
 sg13g2_buf_2 _15545_ (.A(_09928_),
    .X(_09929_));
 sg13g2_buf_1 _15546_ (.A(\top_ihp.oisc.decoder.instruction[8] ),
    .X(_09930_));
 sg13g2_a22oi_1 _15547_ (.Y(_09931_),
    .B1(_09901_),
    .B2(_09930_),
    .A2(_09895_),
    .A1(\top_ihp.oisc.micro_res_addr[1] ));
 sg13g2_nand2b_1 _15548_ (.Y(_09932_),
    .B(_00091_),
    .A_N(_09931_));
 sg13g2_inv_1 _15549_ (.Y(_09933_),
    .A(\top_ihp.oisc.state[2] ));
 sg13g2_o21ai_1 _15550_ (.B1(_09933_),
    .Y(_09934_),
    .A1(net1007),
    .A2(_09932_));
 sg13g2_a22oi_1 _15551_ (.Y(_09935_),
    .B1(_09901_),
    .B2(_09794_),
    .A2(_09895_),
    .A1(\top_ihp.oisc.micro_res_addr[0] ));
 sg13g2_nand2b_1 _15552_ (.Y(_09936_),
    .B(_09922_),
    .A_N(_09935_));
 sg13g2_buf_1 _15553_ (.A(_09936_),
    .X(_09937_));
 sg13g2_nor2b_1 _15554_ (.A(_09934_),
    .B_N(_09937_),
    .Y(_09938_));
 sg13g2_buf_2 _15555_ (.A(_09938_),
    .X(_09939_));
 sg13g2_and2_1 _15556_ (.A(_09929_),
    .B(_09939_),
    .X(_09940_));
 sg13g2_buf_1 _15557_ (.A(_09940_),
    .X(_09941_));
 sg13g2_nand2_1 _15558_ (.Y(_09942_),
    .A(net692),
    .B(_09941_));
 sg13g2_buf_1 _15559_ (.A(_09942_),
    .X(_09943_));
 sg13g2_buf_1 _15560_ (.A(_09943_),
    .X(_09944_));
 sg13g2_mux2_1 _15561_ (.A0(net64),
    .A1(\top_ihp.oisc.regs[0][0] ),
    .S(net409),
    .X(_00484_));
 sg13g2_inv_1 _15562_ (.Y(_09945_),
    .A(_09803_));
 sg13g2_o21ai_1 _15563_ (.B1(_09945_),
    .Y(_09946_),
    .A1(_09792_),
    .A2(_09891_));
 sg13g2_a21oi_1 _15564_ (.A1(_09800_),
    .A2(_09946_),
    .Y(_09947_),
    .B1(_09880_));
 sg13g2_buf_2 _15565_ (.A(_09947_),
    .X(_09948_));
 sg13g2_inv_1 _15566_ (.Y(_09949_),
    .A(_09807_));
 sg13g2_nand2_1 _15567_ (.Y(_09950_),
    .A(_08973_),
    .B(\top_ihp.wb_dati_uart[7] ));
 sg13g2_nor2_1 _15568_ (.A(_00132_),
    .B(net861),
    .Y(_09951_));
 sg13g2_inv_1 _15569_ (.Y(_09952_),
    .A(_00134_));
 sg13g2_a22oi_1 _15570_ (.Y(_09953_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[7] ),
    .A2(_09952_),
    .A1(_08959_));
 sg13g2_and4_1 _15571_ (.A(net1021),
    .B(_00133_),
    .C(_08951_),
    .D(net891),
    .X(_09954_));
 sg13g2_a221oi_1 _15572_ (.B2(_09953_),
    .C1(_09954_),
    .B1(net846),
    .A1(net1024),
    .Y(_09955_),
    .A2(_08594_));
 sg13g2_nor2b_1 _15573_ (.A(_08973_),
    .B_N(_08543_),
    .Y(_09956_));
 sg13g2_buf_1 _15574_ (.A(_09956_),
    .X(_09957_));
 sg13g2_o21ai_1 _15575_ (.B1(_09957_),
    .Y(_09958_),
    .A1(_09951_),
    .A2(_09955_));
 sg13g2_nand3_1 _15576_ (.B(_09950_),
    .C(_09958_),
    .A(_09870_),
    .Y(_09959_));
 sg13g2_buf_1 _15577_ (.A(_09959_),
    .X(_09960_));
 sg13g2_nor2_1 _15578_ (.A(_00156_),
    .B(net861),
    .Y(_09961_));
 sg13g2_inv_1 _15579_ (.Y(_09962_),
    .A(_00158_));
 sg13g2_a22oi_1 _15580_ (.Y(_09963_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[23] ),
    .A2(_09962_),
    .A1(_08959_));
 sg13g2_and4_1 _15581_ (.A(net1021),
    .B(_00157_),
    .C(net879),
    .D(net891),
    .X(_09964_));
 sg13g2_a221oi_1 _15582_ (.B2(_09963_),
    .C1(_09964_),
    .B1(net846),
    .A1(net1024),
    .Y(_09965_),
    .A2(net862));
 sg13g2_o21ai_1 _15583_ (.B1(_08970_),
    .Y(_09966_),
    .A1(_09961_),
    .A2(_09965_));
 sg13g2_buf_1 _15584_ (.A(_09966_),
    .X(_09967_));
 sg13g2_buf_1 _15585_ (.A(\top_ihp.oisc.decoder.instruction[14] ),
    .X(_09968_));
 sg13g2_or3_1 _15586_ (.A(_09806_),
    .B(_09968_),
    .C(_09949_),
    .X(_09969_));
 sg13g2_a21oi_1 _15587_ (.A1(net1035),
    .A2(_09967_),
    .Y(_09970_),
    .B1(_09969_));
 sg13g2_a21o_1 _15588_ (.A2(_08963_),
    .A1(net846),
    .B1(_08966_),
    .X(_09971_));
 sg13g2_inv_1 _15589_ (.Y(_09972_),
    .A(_00179_));
 sg13g2_a22oi_1 _15590_ (.Y(_09973_),
    .B1(_09827_),
    .B2(\top_ihp.wb_coproc.dat_o[31] ),
    .A2(_09972_),
    .A1(net1002));
 sg13g2_mux2_1 _15591_ (.A0(_00178_),
    .A1(_09973_),
    .S(_08958_),
    .X(_09974_));
 sg13g2_mux4_1 _15592_ (.S0(net1035),
    .A0(_00117_),
    .A1(_00177_),
    .A2(_09971_),
    .A3(_09974_),
    .S1(net861),
    .X(_09975_));
 sg13g2_nor2_2 _15593_ (.A(net957),
    .B(_09975_),
    .Y(_09976_));
 sg13g2_nor2b_1 _15594_ (.A(_09968_),
    .B_N(_09806_),
    .Y(_09977_));
 sg13g2_a22oi_1 _15595_ (.Y(_09978_),
    .B1(_09976_),
    .B2(_09977_),
    .A2(_09970_),
    .A1(_09960_));
 sg13g2_o21ai_1 _15596_ (.B1(_09876_),
    .Y(_09979_),
    .A1(_09949_),
    .A2(_09978_));
 sg13g2_buf_1 _15597_ (.A(_09979_),
    .X(_09980_));
 sg13g2_inv_1 _15598_ (.Y(_09981_),
    .A(_09980_));
 sg13g2_buf_1 _15599_ (.A(net1025),
    .X(_09982_));
 sg13g2_nor2_1 _15600_ (.A(_00141_),
    .B(net845),
    .Y(_09983_));
 sg13g2_inv_1 _15601_ (.Y(_09984_),
    .A(_00143_));
 sg13g2_a221oi_1 _15602_ (.B2(\top_ihp.wb_coproc.dat_o[10] ),
    .C1(_09820_),
    .B1(net878),
    .A1(net956),
    .Y(_09985_),
    .A2(_09984_));
 sg13g2_a221oi_1 _15603_ (.B2(_00142_),
    .C1(_09985_),
    .B1(net826),
    .A1(_09850_),
    .Y(_09986_),
    .A2(_08595_));
 sg13g2_o21ai_1 _15604_ (.B1(_08970_),
    .Y(_09987_),
    .A1(_09983_),
    .A2(_09986_));
 sg13g2_inv_1 _15605_ (.Y(_09988_),
    .A(_09987_));
 sg13g2_nand2_1 _15606_ (.Y(_09989_),
    .A(net954),
    .B(net1035));
 sg13g2_nand2_1 _15607_ (.Y(_09990_),
    .A(_00166_),
    .B(net825));
 sg13g2_inv_1 _15608_ (.Y(_09991_),
    .A(_00167_));
 sg13g2_a22oi_1 _15609_ (.Y(_09992_),
    .B1(net878),
    .B2(\top_ihp.wb_coproc.dat_o[26] ),
    .A2(_09991_),
    .A1(net956));
 sg13g2_nand2_1 _15610_ (.Y(_09993_),
    .A(net823),
    .B(_09992_));
 sg13g2_nand3_1 _15611_ (.B(_09990_),
    .C(_09993_),
    .A(_09816_),
    .Y(_09994_));
 sg13g2_o21ai_1 _15612_ (.B1(_09994_),
    .Y(_09995_),
    .A1(_00165_),
    .A2(_09833_));
 sg13g2_nand2_2 _15613_ (.Y(_09996_),
    .A(_08970_),
    .B(_09995_));
 sg13g2_nand2b_1 _15614_ (.Y(_09997_),
    .B(net952),
    .A_N(_09987_));
 sg13g2_o21ai_1 _15615_ (.B1(_09997_),
    .Y(_09998_),
    .A1(_09989_),
    .A2(_09996_));
 sg13g2_buf_1 _15616_ (.A(_08656_),
    .X(_09999_));
 sg13g2_a22oi_1 _15617_ (.Y(_10000_),
    .B1(_09998_),
    .B2(net999),
    .A2(_09988_),
    .A1(net951));
 sg13g2_nand2_1 _15618_ (.Y(_10001_),
    .A(_08358_),
    .B(_08375_));
 sg13g2_xnor2_1 _15619_ (.Y(_10002_),
    .A(_08301_),
    .B(_10001_));
 sg13g2_buf_1 _15620_ (.A(_09897_),
    .X(_10003_));
 sg13g2_a221oi_1 _15621_ (.B2(net902),
    .C1(net1007),
    .B1(_10002_),
    .A1(_09981_),
    .Y(_10004_),
    .A2(_10000_));
 sg13g2_a21oi_1 _15622_ (.A1(\top_ihp.oisc.decoder.instruction[30] ),
    .A2(_09948_),
    .Y(_10005_),
    .B1(_10004_));
 sg13g2_nand2_1 _15623_ (.Y(_10006_),
    .A(net1053),
    .B(net876));
 sg13g2_o21ai_1 _15624_ (.B1(_10006_),
    .Y(_10007_),
    .A1(net880),
    .A2(_10005_));
 sg13g2_buf_1 _15625_ (.A(_10007_),
    .X(_10008_));
 sg13g2_buf_2 _15626_ (.A(_10008_),
    .X(_10009_));
 sg13g2_buf_2 _15627_ (.A(net142),
    .X(_10010_));
 sg13g2_mux2_1 _15628_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[0][10] ),
    .S(net409),
    .X(_00485_));
 sg13g2_buf_1 _15629_ (.A(net592),
    .X(_10011_));
 sg13g2_or2_1 _15630_ (.X(_10012_),
    .B(_09815_),
    .A(_00144_));
 sg13g2_nand2_1 _15631_ (.Y(_10013_),
    .A(_00145_),
    .B(net826));
 sg13g2_inv_1 _15632_ (.Y(_10014_),
    .A(_00146_));
 sg13g2_a22oi_1 _15633_ (.Y(_10015_),
    .B1(net878),
    .B2(\top_ihp.wb_coproc.dat_o[11] ),
    .A2(_10014_),
    .A1(net956));
 sg13g2_nand2_1 _15634_ (.Y(_10016_),
    .A(net823),
    .B(_10015_));
 sg13g2_nand3_1 _15635_ (.B(_10013_),
    .C(_10016_),
    .A(_09816_),
    .Y(_10017_));
 sg13g2_a21oi_1 _15636_ (.A1(_10012_),
    .A2(_10017_),
    .Y(_10018_),
    .B1(_09813_));
 sg13g2_or2_1 _15637_ (.X(_10019_),
    .B(net827),
    .A(_00168_));
 sg13g2_nand2_1 _15638_ (.Y(_10020_),
    .A(_00169_),
    .B(net826));
 sg13g2_inv_1 _15639_ (.Y(_10021_),
    .A(_00170_));
 sg13g2_a22oi_1 _15640_ (.Y(_10022_),
    .B1(_09828_),
    .B2(\top_ihp.wb_coproc.dat_o[27] ),
    .A2(_10021_),
    .A1(_09824_));
 sg13g2_nand2_1 _15641_ (.Y(_10023_),
    .A(net823),
    .B(_10022_));
 sg13g2_nand3_1 _15642_ (.B(_10020_),
    .C(_10023_),
    .A(net827),
    .Y(_10024_));
 sg13g2_a21oi_2 _15643_ (.B1(net957),
    .Y(_10025_),
    .A2(_10024_),
    .A1(_10019_));
 sg13g2_nand2_1 _15644_ (.Y(_10026_),
    .A(_09872_),
    .B(_10025_));
 sg13g2_nand2_1 _15645_ (.Y(_10027_),
    .A(net952),
    .B(_10018_));
 sg13g2_nand2_1 _15646_ (.Y(_10028_),
    .A(_10026_),
    .B(_10027_));
 sg13g2_a22oi_1 _15647_ (.Y(_10029_),
    .B1(_10028_),
    .B2(_08656_),
    .A2(_10018_),
    .A1(net1025));
 sg13g2_nand2_1 _15648_ (.Y(_10030_),
    .A(_08301_),
    .B(_08355_));
 sg13g2_a21oi_1 _15649_ (.A1(_08478_),
    .A2(_08482_),
    .Y(_10031_),
    .B1(_10030_));
 sg13g2_nor2_1 _15650_ (.A(_08457_),
    .B(_10031_),
    .Y(_10032_));
 sg13g2_xor2_1 _15651_ (.B(_10032_),
    .A(net1054),
    .X(_10033_));
 sg13g2_and2_1 _15652_ (.A(net1030),
    .B(_09897_),
    .X(_10034_));
 sg13g2_a221oi_1 _15653_ (.B2(_10034_),
    .C1(net1007),
    .B1(_10033_),
    .A1(_09981_),
    .Y(_10035_),
    .A2(_10029_));
 sg13g2_nor2_1 _15654_ (.A(_09782_),
    .B(net1008),
    .Y(_10036_));
 sg13g2_buf_1 _15655_ (.A(_10036_),
    .X(_10037_));
 sg13g2_o21ai_1 _15656_ (.B1(_10037_),
    .Y(_10038_),
    .A1(net903),
    .A2(_10033_));
 sg13g2_nand2b_1 _15657_ (.Y(_10039_),
    .B(_10038_),
    .A_N(net1030));
 sg13g2_o21ai_1 _15658_ (.B1(_10039_),
    .Y(_10040_),
    .A1(net907),
    .A2(_10035_));
 sg13g2_buf_2 _15659_ (.A(_10040_),
    .X(_10041_));
 sg13g2_buf_1 _15660_ (.A(_10037_),
    .X(_10042_));
 sg13g2_buf_1 _15661_ (.A(\top_ihp.oisc.decoder.instruction[31] ),
    .X(_10043_));
 sg13g2_nor2b_1 _15662_ (.A(net1005),
    .B_N(_09796_),
    .Y(_10044_));
 sg13g2_a22oi_1 _15663_ (.Y(_10045_),
    .B1(_09891_),
    .B2(_10044_),
    .A2(_10043_),
    .A1(net1005));
 sg13g2_nand4_1 _15664_ (.B(_09799_),
    .C(net1005),
    .A(_09804_),
    .Y(_10046_),
    .D(_09794_));
 sg13g2_o21ai_1 _15665_ (.B1(_10046_),
    .Y(_10047_),
    .A1(_09804_),
    .A2(_10045_));
 sg13g2_nand3_1 _15666_ (.B(net875),
    .C(_10047_),
    .A(net958),
    .Y(_10048_));
 sg13g2_and2_1 _15667_ (.A(_10041_),
    .B(_10048_),
    .X(_10049_));
 sg13g2_buf_2 _15668_ (.A(_10049_),
    .X(_10050_));
 sg13g2_buf_8 _15669_ (.A(_10050_),
    .X(_10051_));
 sg13g2_buf_1 _15670_ (.A(_09942_),
    .X(_10052_));
 sg13g2_nand2_1 _15671_ (.Y(_10053_),
    .A(\top_ihp.oisc.regs[0][11] ),
    .B(net591));
 sg13g2_o21ai_1 _15672_ (.B1(_10053_),
    .Y(_00486_),
    .A1(net408),
    .A2(net62));
 sg13g2_buf_1 _15673_ (.A(net907),
    .X(_10054_));
 sg13g2_nor2_1 _15674_ (.A(_09945_),
    .B(_09799_),
    .Y(_10055_));
 sg13g2_and2_1 _15675_ (.A(_09792_),
    .B(_10055_),
    .X(_10056_));
 sg13g2_buf_2 _15676_ (.A(_10056_),
    .X(_10057_));
 sg13g2_nor2_1 _15677_ (.A(net1004),
    .B(_09792_),
    .Y(_10058_));
 sg13g2_nand2_1 _15678_ (.Y(_10059_),
    .A(_09891_),
    .B(_10058_));
 sg13g2_buf_1 _15679_ (.A(_10059_),
    .X(_10060_));
 sg13g2_nand2b_1 _15680_ (.Y(_10061_),
    .B(_10060_),
    .A_N(_10057_));
 sg13g2_nand2_1 _15681_ (.Y(_10062_),
    .A(_09792_),
    .B(_10043_));
 sg13g2_o21ai_1 _15682_ (.B1(net1007),
    .Y(_10063_),
    .A1(_10062_),
    .A2(_10055_));
 sg13g2_buf_1 _15683_ (.A(_10063_),
    .X(_10064_));
 sg13g2_a21oi_1 _15684_ (.A1(net999),
    .A2(_10061_),
    .Y(_10065_),
    .B1(_10064_));
 sg13g2_a21oi_1 _15685_ (.A1(\top_ihp.wb_coproc.dat_o[12] ),
    .A2(_08598_),
    .Y(_10066_),
    .B1(net1002));
 sg13g2_a21o_1 _15686_ (.A2(_09823_),
    .A1(_00083_),
    .B1(_10066_),
    .X(_10067_));
 sg13g2_mux2_1 _15687_ (.A0(_00082_),
    .A1(_10067_),
    .S(_09853_),
    .X(_10068_));
 sg13g2_mux2_1 _15688_ (.A0(_00081_),
    .A1(_10068_),
    .S(net845),
    .X(_10069_));
 sg13g2_nor2_1 _15689_ (.A(net957),
    .B(_10069_),
    .Y(_10070_));
 sg13g2_buf_2 _15690_ (.A(_10070_),
    .X(_10071_));
 sg13g2_or2_1 _15691_ (.X(_10072_),
    .B(net827),
    .A(_00171_));
 sg13g2_inv_1 _15692_ (.Y(_10073_),
    .A(_00173_));
 sg13g2_a221oi_1 _15693_ (.B2(\top_ihp.wb_coproc.dat_o[28] ),
    .C1(net826),
    .B1(net878),
    .A1(net956),
    .Y(_10074_),
    .A2(_10073_));
 sg13g2_a21oi_1 _15694_ (.A1(_00172_),
    .A2(net825),
    .Y(_10075_),
    .B1(_10074_));
 sg13g2_nand2_1 _15695_ (.Y(_10076_),
    .A(net824),
    .B(_10075_));
 sg13g2_a21oi_2 _15696_ (.B1(net957),
    .Y(_10077_),
    .A2(_10076_),
    .A1(_10072_));
 sg13g2_nor3_1 _15697_ (.A(_09810_),
    .B(net957),
    .C(_10069_),
    .Y(_10078_));
 sg13g2_a21o_1 _15698_ (.A2(_10077_),
    .A1(net877),
    .B1(_10078_),
    .X(_10079_));
 sg13g2_a22oi_1 _15699_ (.Y(_10080_),
    .B1(_10079_),
    .B2(net999),
    .A2(_10071_),
    .A1(net951));
 sg13g2_o21ai_1 _15700_ (.B1(net1054),
    .Y(_10081_),
    .A1(_08457_),
    .A2(_10031_));
 sg13g2_nor3_1 _15701_ (.A(net1054),
    .B(_08457_),
    .C(_10031_),
    .Y(_10082_));
 sg13g2_a21oi_1 _15702_ (.A1(net1030),
    .A2(_10081_),
    .Y(_10083_),
    .B1(_10082_));
 sg13g2_xor2_1 _15703_ (.B(_10083_),
    .A(_08296_),
    .X(_10084_));
 sg13g2_a22oi_1 _15704_ (.Y(_10085_),
    .B1(_10084_),
    .B2(net902),
    .A2(_10080_),
    .A1(_09981_));
 sg13g2_nor2_1 _15705_ (.A(net958),
    .B(_10085_),
    .Y(_10086_));
 sg13g2_nor3_2 _15706_ (.A(net876),
    .B(_10065_),
    .C(_10086_),
    .Y(_10087_));
 sg13g2_a21oi_1 _15707_ (.A1(_08252_),
    .A2(net874),
    .Y(_10088_),
    .B1(_10087_));
 sg13g2_buf_2 _15708_ (.A(_10088_),
    .X(_10089_));
 sg13g2_buf_1 _15709_ (.A(net141),
    .X(_10090_));
 sg13g2_nand2_1 _15710_ (.Y(_10091_),
    .A(\top_ihp.oisc.regs[0][12] ),
    .B(net591));
 sg13g2_o21ai_1 _15711_ (.B1(_10091_),
    .Y(_00487_),
    .A1(net408),
    .A2(net61));
 sg13g2_buf_1 _15712_ (.A(net1025),
    .X(_10092_));
 sg13g2_inv_1 _15713_ (.Y(_10093_),
    .A(_00089_));
 sg13g2_a221oi_1 _15714_ (.B2(\top_ihp.wb_coproc.dat_o[13] ),
    .C1(net826),
    .B1(net878),
    .A1(net956),
    .Y(_10094_),
    .A2(_10093_));
 sg13g2_a21oi_1 _15715_ (.A1(_00088_),
    .A2(net825),
    .Y(_10095_),
    .B1(_10094_));
 sg13g2_nor2_1 _15716_ (.A(_00087_),
    .B(net827),
    .Y(_10096_));
 sg13g2_a21oi_2 _15717_ (.B1(_10096_),
    .Y(_10097_),
    .A2(_10095_),
    .A1(_09833_));
 sg13g2_nor2_1 _15718_ (.A(net906),
    .B(_10097_),
    .Y(_10098_));
 sg13g2_nand2b_1 _15719_ (.Y(_10099_),
    .B(_08970_),
    .A_N(_10097_));
 sg13g2_buf_1 _15720_ (.A(_10099_),
    .X(_10100_));
 sg13g2_inv_1 _15721_ (.Y(_10101_),
    .A(_00176_));
 sg13g2_a221oi_1 _15722_ (.B2(\top_ihp.wb_coproc.dat_o[29] ),
    .C1(net825),
    .B1(net859),
    .A1(net905),
    .Y(_10102_),
    .A2(_10101_));
 sg13g2_a21oi_1 _15723_ (.A1(_00175_),
    .A2(net790),
    .Y(_10103_),
    .B1(_10102_));
 sg13g2_nor2_1 _15724_ (.A(_00174_),
    .B(_09817_),
    .Y(_10104_));
 sg13g2_a21oi_1 _15725_ (.A1(net791),
    .A2(_10103_),
    .Y(_10105_),
    .B1(_10104_));
 sg13g2_nor2_2 _15726_ (.A(net906),
    .B(_10105_),
    .Y(_10106_));
 sg13g2_nand2_1 _15727_ (.Y(_10107_),
    .A(_09873_),
    .B(_10106_));
 sg13g2_o21ai_1 _15728_ (.B1(_10107_),
    .Y(_10108_),
    .A1(_09811_),
    .A2(net731));
 sg13g2_a221oi_1 _15729_ (.B2(net999),
    .C1(_09980_),
    .B1(_10108_),
    .A1(net950),
    .Y(_10109_),
    .A2(_10098_));
 sg13g2_buf_1 _15730_ (.A(net903),
    .X(_10110_));
 sg13g2_nor3_1 _15731_ (.A(_08296_),
    .B(_08298_),
    .C(_08299_),
    .Y(_10111_));
 sg13g2_inv_1 _15732_ (.Y(_10112_),
    .A(_10032_));
 sg13g2_a21oi_1 _15733_ (.A1(_10111_),
    .A2(_10112_),
    .Y(_10113_),
    .B1(_08460_));
 sg13g2_xor2_1 _15734_ (.B(_10113_),
    .A(_08295_),
    .X(_10114_));
 sg13g2_nor2_1 _15735_ (.A(net873),
    .B(_10114_),
    .Y(_10115_));
 sg13g2_buf_1 _15736_ (.A(_09880_),
    .X(_10116_));
 sg13g2_o21ai_1 _15737_ (.B1(net949),
    .Y(_10117_),
    .A1(_10109_),
    .A2(_10115_));
 sg13g2_a21oi_1 _15738_ (.A1(net950),
    .A2(_10061_),
    .Y(_10118_),
    .B1(_10064_));
 sg13g2_nor2_1 _15739_ (.A(net876),
    .B(_10118_),
    .Y(_10119_));
 sg13g2_a22oi_1 _15740_ (.Y(_10120_),
    .B1(_10117_),
    .B2(_10119_),
    .A2(net874),
    .A1(net1055));
 sg13g2_buf_1 _15741_ (.A(_10120_),
    .X(_10121_));
 sg13g2_buf_2 _15742_ (.A(_10121_),
    .X(_10122_));
 sg13g2_nand2_1 _15743_ (.Y(_10123_),
    .A(\top_ihp.oisc.regs[0][13] ),
    .B(net591));
 sg13g2_o21ai_1 _15744_ (.B1(_10123_),
    .Y(_00488_),
    .A1(net408),
    .A2(_10122_));
 sg13g2_or2_1 _15745_ (.X(_10124_),
    .B(net824),
    .A(_00084_));
 sg13g2_nand2_1 _15746_ (.Y(_10125_),
    .A(_00085_),
    .B(_09830_));
 sg13g2_inv_1 _15747_ (.Y(_10126_),
    .A(_00086_));
 sg13g2_a22oi_1 _15748_ (.Y(_10127_),
    .B1(net859),
    .B2(\top_ihp.wb_coproc.dat_o[14] ),
    .A2(_10126_),
    .A1(net905));
 sg13g2_nand2_1 _15749_ (.Y(_10128_),
    .A(_09853_),
    .B(_10127_));
 sg13g2_nand3_1 _15750_ (.B(_10125_),
    .C(_10128_),
    .A(net824),
    .Y(_10129_));
 sg13g2_a21oi_1 _15751_ (.A1(_10124_),
    .A2(_10129_),
    .Y(_10130_),
    .B1(net906));
 sg13g2_buf_2 _15752_ (.A(_10130_),
    .X(_10131_));
 sg13g2_a21o_1 _15753_ (.A2(_10129_),
    .A1(_10124_),
    .B1(net957),
    .X(_10132_));
 sg13g2_buf_1 _15754_ (.A(_10132_),
    .X(_10133_));
 sg13g2_inv_1 _15755_ (.Y(_10134_),
    .A(_00116_));
 sg13g2_a221oi_1 _15756_ (.B2(\top_ihp.wb_coproc.dat_o[30] ),
    .C1(net826),
    .B1(net859),
    .A1(net905),
    .Y(_10135_),
    .A2(_10134_));
 sg13g2_a21oi_1 _15757_ (.A1(_00115_),
    .A2(_09822_),
    .Y(_10136_),
    .B1(_10135_));
 sg13g2_nor2_1 _15758_ (.A(_00114_),
    .B(net824),
    .Y(_10137_));
 sg13g2_a21oi_1 _15759_ (.A1(net824),
    .A2(_10136_),
    .Y(_10138_),
    .B1(_10137_));
 sg13g2_nor2_2 _15760_ (.A(net906),
    .B(_10138_),
    .Y(_10139_));
 sg13g2_nand2_1 _15761_ (.Y(_10140_),
    .A(_09873_),
    .B(_10139_));
 sg13g2_o21ai_1 _15762_ (.B1(_10140_),
    .Y(_10141_),
    .A1(_09811_),
    .A2(_10133_));
 sg13g2_a221oi_1 _15763_ (.B2(net999),
    .C1(_09980_),
    .B1(_10141_),
    .A1(net950),
    .Y(_10142_),
    .A2(_10131_));
 sg13g2_nor2_1 _15764_ (.A(_08251_),
    .B(_08254_),
    .Y(_10143_));
 sg13g2_a21oi_1 _15765_ (.A1(net1055),
    .A2(_08257_),
    .Y(_10144_),
    .B1(_10143_));
 sg13g2_or2_1 _15766_ (.X(_10145_),
    .B(_10144_),
    .A(_08270_));
 sg13g2_a21o_1 _15767_ (.A2(_10001_),
    .A1(_08302_),
    .B1(_10145_),
    .X(_10146_));
 sg13g2_buf_1 _15768_ (.A(_10146_),
    .X(_10147_));
 sg13g2_xor2_1 _15769_ (.B(_08305_),
    .A(_10147_),
    .X(_10148_));
 sg13g2_nor2_1 _15770_ (.A(net873),
    .B(_10148_),
    .Y(_10149_));
 sg13g2_o21ai_1 _15771_ (.B1(net949),
    .Y(_10150_),
    .A1(_10142_),
    .A2(_10149_));
 sg13g2_inv_1 _15772_ (.Y(_10151_),
    .A(_10064_));
 sg13g2_buf_1 _15773_ (.A(_10057_),
    .X(_10152_));
 sg13g2_nor2_1 _15774_ (.A(_08659_),
    .B(_10060_),
    .Y(_10153_));
 sg13g2_a21oi_1 _15775_ (.A1(_09968_),
    .A2(net858),
    .Y(_10154_),
    .B1(_10153_));
 sg13g2_buf_1 _15776_ (.A(_09784_),
    .X(_10155_));
 sg13g2_a21oi_1 _15777_ (.A1(_10151_),
    .A2(_10154_),
    .Y(_10156_),
    .B1(net901));
 sg13g2_a22oi_1 _15778_ (.Y(_10157_),
    .B1(_10150_),
    .B2(_10156_),
    .A2(_09786_),
    .A1(net1051));
 sg13g2_buf_1 _15779_ (.A(_10157_),
    .X(_10158_));
 sg13g2_buf_2 _15780_ (.A(_10158_),
    .X(_10159_));
 sg13g2_nand2_1 _15781_ (.Y(_10160_),
    .A(\top_ihp.oisc.regs[0][14] ),
    .B(net591));
 sg13g2_o21ai_1 _15782_ (.B1(_10160_),
    .Y(_00489_),
    .A1(net408),
    .A2(net277));
 sg13g2_or2_1 _15783_ (.X(_10161_),
    .B(_09977_),
    .A(_08656_));
 sg13g2_a221oi_1 _15784_ (.B2(_10161_),
    .C1(_08657_),
    .B1(_09976_),
    .A1(_09960_),
    .Y(_10162_),
    .A2(_09970_));
 sg13g2_a21oi_1 _15785_ (.A1(net1025),
    .A2(_08972_),
    .Y(_10163_),
    .B1(_10162_));
 sg13g2_xor2_1 _15786_ (.B(_08487_),
    .A(_08304_),
    .X(_10164_));
 sg13g2_nand2_1 _15787_ (.Y(_10165_),
    .A(_09897_),
    .B(_10164_));
 sg13g2_o21ai_1 _15788_ (.B1(_10165_),
    .Y(_10166_),
    .A1(_09897_),
    .A2(_10163_));
 sg13g2_nand2_1 _15789_ (.Y(_10167_),
    .A(\top_ihp.oisc.decoder.instruction[15] ),
    .B(_10061_));
 sg13g2_a221oi_1 _15790_ (.B2(_10151_),
    .C1(_09784_),
    .B1(_10167_),
    .A1(_09880_),
    .Y(_10168_),
    .A2(_10166_));
 sg13g2_buf_1 _15791_ (.A(_10168_),
    .X(_10169_));
 sg13g2_a21oi_1 _15792_ (.A1(_08287_),
    .A2(_10054_),
    .Y(_10170_),
    .B1(net663));
 sg13g2_buf_2 _15793_ (.A(_10170_),
    .X(_10171_));
 sg13g2_nand2_1 _15794_ (.Y(_10172_),
    .A(\top_ihp.oisc.regs[0][15] ),
    .B(net591));
 sg13g2_o21ai_1 _15795_ (.B1(_10172_),
    .Y(_00490_),
    .A1(_10011_),
    .A2(net407));
 sg13g2_nor2_1 _15796_ (.A(_00237_),
    .B(_10060_),
    .Y(_10173_));
 sg13g2_a21oi_1 _15797_ (.A1(\top_ihp.oisc.decoder.instruction[16] ),
    .A2(net858),
    .Y(_10174_),
    .B1(_10173_));
 sg13g2_nor2_1 _15798_ (.A(_08362_),
    .B(_08364_),
    .Y(_10175_));
 sg13g2_nand2_1 _15799_ (.Y(_10176_),
    .A(_08340_),
    .B(_08343_));
 sg13g2_a221oi_1 _15800_ (.B2(_08337_),
    .C1(_10176_),
    .B1(_08335_),
    .A1(_08325_),
    .Y(_10177_),
    .A2(_08333_));
 sg13g2_buf_1 _15801_ (.A(_10177_),
    .X(_10178_));
 sg13g2_o21ai_1 _15802_ (.B1(net1029),
    .Y(_10179_),
    .A1(_10175_),
    .A2(_10178_));
 sg13g2_nor3_1 _15803_ (.A(_08366_),
    .B(_10175_),
    .C(_10178_),
    .Y(_10180_));
 sg13g2_a21oi_2 _15804_ (.B1(_10180_),
    .Y(_10181_),
    .A2(_10179_),
    .A1(_08345_));
 sg13g2_nor2b_1 _15805_ (.A(_09676_),
    .B_N(_08369_),
    .Y(_10182_));
 sg13g2_nand2b_1 _15806_ (.Y(_10183_),
    .B(net1030),
    .A_N(net1054));
 sg13g2_nor2_1 _15807_ (.A(_08372_),
    .B(_08373_),
    .Y(_10184_));
 sg13g2_nor3_1 _15808_ (.A(_08263_),
    .B(_10184_),
    .C(_08374_),
    .Y(_10185_));
 sg13g2_o21ai_1 _15809_ (.B1(_08263_),
    .Y(_10186_),
    .A1(_10184_),
    .A2(_08374_));
 sg13g2_o21ai_1 _15810_ (.B1(_10186_),
    .Y(_10187_),
    .A1(net1053),
    .A2(_10185_));
 sg13g2_a21o_1 _15811_ (.A2(_10187_),
    .A1(_10183_),
    .B1(_08298_),
    .X(_10188_));
 sg13g2_and3_1 _15812_ (.X(_10189_),
    .A(_08461_),
    .B(_08266_),
    .C(_08306_));
 sg13g2_nor2_1 _15813_ (.A(net1051),
    .B(_08452_),
    .Y(_10190_));
 sg13g2_a221oi_1 _15814_ (.B2(_08306_),
    .C1(_08288_),
    .B1(_10144_),
    .A1(_08279_),
    .Y(_10191_),
    .A2(_10190_));
 sg13g2_o21ai_1 _15815_ (.B1(_10191_),
    .Y(_10192_),
    .A1(_08479_),
    .A2(_09676_));
 sg13g2_a221oi_1 _15816_ (.B2(_10189_),
    .C1(_10192_),
    .B1(_10188_),
    .A1(_10181_),
    .Y(_10193_),
    .A2(_10182_));
 sg13g2_xor2_1 _15817_ (.B(_10193_),
    .A(_08307_),
    .X(_10194_));
 sg13g2_nor2_1 _15818_ (.A(_08656_),
    .B(_09806_),
    .Y(_10195_));
 sg13g2_nor3_1 _15819_ (.A(_08657_),
    .B(_09968_),
    .C(_10195_),
    .Y(_10196_));
 sg13g2_a22oi_1 _15820_ (.Y(_10197_),
    .B1(_09976_),
    .B2(_10196_),
    .A2(_09970_),
    .A1(_09960_));
 sg13g2_buf_2 _15821_ (.A(_10197_),
    .X(_10198_));
 sg13g2_o21ai_1 _15822_ (.B1(_10198_),
    .Y(_10199_),
    .A1(net954),
    .A2(_09868_));
 sg13g2_mux2_1 _15823_ (.A0(_10194_),
    .A1(_10199_),
    .S(net903),
    .X(_10200_));
 sg13g2_nor2_1 _15824_ (.A(net958),
    .B(_10200_),
    .Y(_10201_));
 sg13g2_a21oi_2 _15825_ (.B1(_10201_),
    .Y(_10202_),
    .A2(_10174_),
    .A1(_10151_));
 sg13g2_nor2_1 _15826_ (.A(_08291_),
    .B(_10042_),
    .Y(_10203_));
 sg13g2_a21oi_1 _15827_ (.A1(net875),
    .A2(_10202_),
    .Y(_10204_),
    .B1(_10203_));
 sg13g2_buf_1 _15828_ (.A(_10204_),
    .X(_10205_));
 sg13g2_buf_1 _15829_ (.A(net276),
    .X(_10206_));
 sg13g2_nand2_1 _15830_ (.Y(_10207_),
    .A(\top_ihp.oisc.regs[0][16] ),
    .B(net591));
 sg13g2_o21ai_1 _15831_ (.B1(_10207_),
    .Y(_00491_),
    .A1(net408),
    .A2(_10206_));
 sg13g2_nand2_1 _15832_ (.Y(_10208_),
    .A(net949),
    .B(_10037_));
 sg13g2_nor2_1 _15833_ (.A(_00123_),
    .B(_08944_),
    .Y(_10209_));
 sg13g2_inv_1 _15834_ (.Y(_10210_),
    .A(_00125_));
 sg13g2_a22oi_1 _15835_ (.Y(_10211_),
    .B1(_08962_),
    .B2(\top_ihp.wb_coproc.dat_o[17] ),
    .A2(_10210_),
    .A1(_08959_));
 sg13g2_and4_1 _15836_ (.A(_08947_),
    .B(_00124_),
    .C(_08951_),
    .D(_08955_),
    .X(_10212_));
 sg13g2_a221oi_1 _15837_ (.B2(_10211_),
    .C1(_10212_),
    .B1(_08957_),
    .A1(net1024),
    .Y(_10213_),
    .A2(_08594_));
 sg13g2_o21ai_1 _15838_ (.B1(_08975_),
    .Y(_10214_),
    .A1(_10209_),
    .A2(_10213_));
 sg13g2_buf_2 _15839_ (.A(_10214_),
    .X(_10215_));
 sg13g2_o21ai_1 _15840_ (.B1(_10198_),
    .Y(_10216_),
    .A1(net954),
    .A2(_10215_));
 sg13g2_xor2_1 _15841_ (.B(_08647_),
    .A(_08308_),
    .X(_10217_));
 sg13g2_mux2_1 _15842_ (.A0(_10216_),
    .A1(_10217_),
    .S(_10003_),
    .X(_10218_));
 sg13g2_a21oi_1 _15843_ (.A1(\top_ihp.oisc.decoder.instruction[17] ),
    .A2(_10057_),
    .Y(_10219_),
    .B1(_10064_));
 sg13g2_o21ai_1 _15844_ (.B1(_10219_),
    .Y(_10220_),
    .A1(_00238_),
    .A2(_10060_));
 sg13g2_mux2_1 _15845_ (.A0(net1052),
    .A1(_10220_),
    .S(_10037_),
    .X(_10221_));
 sg13g2_o21ai_1 _15846_ (.B1(_10221_),
    .Y(_10222_),
    .A1(_10208_),
    .A2(_10218_));
 sg13g2_buf_1 _15847_ (.A(_10222_),
    .X(_10223_));
 sg13g2_buf_1 _15848_ (.A(_10223_),
    .X(_10224_));
 sg13g2_nand2_1 _15849_ (.Y(_10225_),
    .A(\top_ihp.oisc.regs[0][17] ),
    .B(_10052_));
 sg13g2_o21ai_1 _15850_ (.B1(_10225_),
    .Y(_00492_),
    .A1(net408),
    .A2(net406));
 sg13g2_a22oi_1 _15851_ (.Y(_10226_),
    .B1(_10147_),
    .B2(_08310_),
    .A2(_08294_),
    .A1(_08290_));
 sg13g2_buf_1 _15852_ (.A(_10226_),
    .X(_10227_));
 sg13g2_xnor2_1 _15853_ (.Y(_10228_),
    .A(_08492_),
    .B(_10227_));
 sg13g2_buf_1 _15854_ (.A(net903),
    .X(_10229_));
 sg13g2_nor2_1 _15855_ (.A(_00126_),
    .B(_08944_),
    .Y(_10230_));
 sg13g2_inv_1 _15856_ (.Y(_10231_),
    .A(_00128_));
 sg13g2_a22oi_1 _15857_ (.Y(_10232_),
    .B1(_08962_),
    .B2(\top_ihp.wb_coproc.dat_o[18] ),
    .A2(_10231_),
    .A1(_08959_));
 sg13g2_and4_1 _15858_ (.A(_08964_),
    .B(_00127_),
    .C(_08951_),
    .D(net891),
    .X(_10233_));
 sg13g2_a221oi_1 _15859_ (.B2(_10232_),
    .C1(_10233_),
    .B1(_08957_),
    .A1(net1024),
    .Y(_10234_),
    .A2(_08594_));
 sg13g2_o21ai_1 _15860_ (.B1(_08975_),
    .Y(_10235_),
    .A1(_10230_),
    .A2(_10234_));
 sg13g2_inv_1 _15861_ (.Y(_10236_),
    .A(_10235_));
 sg13g2_nand2_1 _15862_ (.Y(_10237_),
    .A(net951),
    .B(_10236_));
 sg13g2_nand3_1 _15863_ (.B(_10198_),
    .C(_10237_),
    .A(_10229_),
    .Y(_10238_));
 sg13g2_o21ai_1 _15864_ (.B1(_10238_),
    .Y(_10239_),
    .A1(net873),
    .A2(_10228_));
 sg13g2_nand2_1 _15865_ (.Y(_10240_),
    .A(net949),
    .B(_10239_));
 sg13g2_nor2_1 _15866_ (.A(_00239_),
    .B(_10060_),
    .Y(_10241_));
 sg13g2_a21oi_1 _15867_ (.A1(\top_ihp.oisc.decoder.instruction[18] ),
    .A2(net858),
    .Y(_10242_),
    .B1(_10241_));
 sg13g2_a21oi_1 _15868_ (.A1(_10151_),
    .A2(_10242_),
    .Y(_10243_),
    .B1(net901));
 sg13g2_a22oi_1 _15869_ (.Y(_10244_),
    .B1(_10240_),
    .B2(_10243_),
    .A2(net880),
    .A1(net1059));
 sg13g2_buf_1 _15870_ (.A(_10244_),
    .X(_10245_));
 sg13g2_buf_2 _15871_ (.A(_10245_),
    .X(_10246_));
 sg13g2_nand2_1 _15872_ (.Y(_10247_),
    .A(\top_ihp.oisc.regs[0][18] ),
    .B(_10052_));
 sg13g2_o21ai_1 _15873_ (.B1(_10247_),
    .Y(_00493_),
    .A1(net408),
    .A2(_10246_));
 sg13g2_a21oi_1 _15874_ (.A1(\top_ihp.oisc.decoder.instruction[19] ),
    .A2(_10057_),
    .Y(_10248_),
    .B1(_10064_));
 sg13g2_o21ai_1 _15875_ (.B1(_10248_),
    .Y(_10249_),
    .A1(_00240_),
    .A2(_10060_));
 sg13g2_nand2_1 _15876_ (.Y(_10250_),
    .A(_10037_),
    .B(_10249_));
 sg13g2_nor2_1 _15877_ (.A(_00129_),
    .B(_08945_),
    .Y(_10251_));
 sg13g2_inv_1 _15878_ (.Y(_10252_),
    .A(_00131_));
 sg13g2_a22oi_1 _15879_ (.Y(_10253_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[19] ),
    .A2(_10252_),
    .A1(net1002));
 sg13g2_and4_1 _15880_ (.A(_08964_),
    .B(_00130_),
    .C(net879),
    .D(_08965_),
    .X(_10254_));
 sg13g2_a221oi_1 _15881_ (.B2(_10253_),
    .C1(_10254_),
    .B1(net846),
    .A1(net1024),
    .Y(_10255_),
    .A2(net862));
 sg13g2_o21ai_1 _15882_ (.B1(_08975_),
    .Y(_10256_),
    .A1(_10251_),
    .A2(_10255_));
 sg13g2_buf_2 _15883_ (.A(_10256_),
    .X(_10257_));
 sg13g2_inv_1 _15884_ (.Y(_10258_),
    .A(_10257_));
 sg13g2_nand3_1 _15885_ (.B(_09876_),
    .C(_10198_),
    .A(_09880_),
    .Y(_10259_));
 sg13g2_buf_2 _15886_ (.A(_10259_),
    .X(_10260_));
 sg13g2_a21oi_1 _15887_ (.A1(net951),
    .A2(_10258_),
    .Y(_10261_),
    .B1(_10260_));
 sg13g2_nand2_2 _15888_ (.Y(_10262_),
    .A(_09880_),
    .B(_09897_));
 sg13g2_nor4_1 _15889_ (.A(_08489_),
    .B(_08494_),
    .C(_08647_),
    .D(_10262_),
    .Y(_10263_));
 sg13g2_nor2_2 _15890_ (.A(net1007),
    .B(_09876_),
    .Y(_10264_));
 sg13g2_nand3_1 _15891_ (.B(_08494_),
    .C(_08639_),
    .A(_08489_),
    .Y(_10265_));
 sg13g2_o21ai_1 _15892_ (.B1(_10265_),
    .Y(_10266_),
    .A1(_08489_),
    .A2(_08639_));
 sg13g2_nand2_1 _15893_ (.Y(_10267_),
    .A(_10264_),
    .B(_10266_));
 sg13g2_nand4_1 _15894_ (.B(_08639_),
    .C(_08647_),
    .A(_08489_),
    .Y(_10268_),
    .D(_10264_));
 sg13g2_nand2_1 _15895_ (.Y(_10269_),
    .A(_10267_),
    .B(_10268_));
 sg13g2_nor4_1 _15896_ (.A(_10250_),
    .B(_10261_),
    .C(_10263_),
    .D(_10269_),
    .Y(_10270_));
 sg13g2_buf_2 _15897_ (.A(_10270_),
    .X(_10271_));
 sg13g2_a21oi_1 _15898_ (.A1(net1058),
    .A2(_10054_),
    .Y(_10272_),
    .B1(_10271_));
 sg13g2_buf_2 _15899_ (.A(_10272_),
    .X(_10273_));
 sg13g2_buf_1 _15900_ (.A(_10273_),
    .X(_10274_));
 sg13g2_buf_1 _15901_ (.A(net592),
    .X(_10275_));
 sg13g2_nand2_1 _15902_ (.Y(_10276_),
    .A(\top_ihp.oisc.regs[0][19] ),
    .B(net405));
 sg13g2_o21ai_1 _15903_ (.B1(_10276_),
    .Y(_00494_),
    .A1(net408),
    .A2(net60));
 sg13g2_buf_1 _15904_ (.A(net592),
    .X(_10277_));
 sg13g2_nor2_1 _15905_ (.A(_09945_),
    .B(net1036),
    .Y(_10278_));
 sg13g2_buf_1 _15906_ (.A(\top_ihp.oisc.decoder.instruction[21] ),
    .X(_10279_));
 sg13g2_mux2_1 _15907_ (.A0(_10279_),
    .A1(_09930_),
    .S(net1036),
    .X(_10280_));
 sg13g2_a22oi_1 _15908_ (.Y(_10281_),
    .B1(_10280_),
    .B2(_09945_),
    .A2(_10278_),
    .A1(_09930_));
 sg13g2_nor2b_1 _15909_ (.A(_10281_),
    .B_N(_09793_),
    .Y(_10282_));
 sg13g2_and2_1 _15910_ (.A(_09797_),
    .B(_10058_),
    .X(_10283_));
 sg13g2_buf_1 _15911_ (.A(_10283_),
    .X(_10284_));
 sg13g2_nand2_1 _15912_ (.Y(_10285_),
    .A(net1006),
    .B(_10279_));
 sg13g2_o21ai_1 _15913_ (.B1(_10285_),
    .Y(_10286_),
    .A1(net1006),
    .A2(_00233_));
 sg13g2_and2_1 _15914_ (.A(_10284_),
    .B(_10286_),
    .X(_10287_));
 sg13g2_o21ai_1 _15915_ (.B1(net958),
    .Y(_10288_),
    .A1(_10282_),
    .A2(_10287_));
 sg13g2_or2_1 _15916_ (.X(_10289_),
    .B(_09815_),
    .A(_00162_));
 sg13g2_nand2_1 _15917_ (.Y(_10290_),
    .A(_00163_),
    .B(net826));
 sg13g2_inv_1 _15918_ (.Y(_10291_),
    .A(_00164_));
 sg13g2_a22oi_1 _15919_ (.Y(_10292_),
    .B1(_09828_),
    .B2(\top_ihp.wb_coproc.dat_o[25] ),
    .A2(_10291_),
    .A1(_09824_));
 sg13g2_nand2_1 _15920_ (.Y(_10293_),
    .A(net823),
    .B(_10292_));
 sg13g2_nand3_1 _15921_ (.B(_10290_),
    .C(_10293_),
    .A(net827),
    .Y(_10294_));
 sg13g2_a21oi_2 _15922_ (.B1(net957),
    .Y(_10295_),
    .A2(_10294_),
    .A1(_10289_));
 sg13g2_nand2_1 _15923_ (.Y(_10296_),
    .A(net955),
    .B(_10295_));
 sg13g2_o21ai_1 _15924_ (.B1(_10296_),
    .Y(_10297_),
    .A1(net955),
    .A2(_10215_));
 sg13g2_nor2_1 _15925_ (.A(_00138_),
    .B(net827),
    .Y(_10298_));
 sg13g2_inv_1 _15926_ (.Y(_10299_),
    .A(_00140_));
 sg13g2_a221oi_1 _15927_ (.B2(\top_ihp.wb_coproc.dat_o[9] ),
    .C1(net826),
    .B1(net859),
    .A1(net905),
    .Y(_10300_),
    .A2(_10299_));
 sg13g2_a221oi_1 _15928_ (.B2(_00139_),
    .C1(_10300_),
    .B1(_09830_),
    .A1(_09850_),
    .Y(_10301_),
    .A2(_08595_));
 sg13g2_o21ai_1 _15929_ (.B1(_08970_),
    .Y(_10302_),
    .A1(_10298_),
    .A2(_10301_));
 sg13g2_buf_1 _15930_ (.A(_10302_),
    .X(_10303_));
 sg13g2_nand3_1 _15931_ (.B(_09846_),
    .C(_10303_),
    .A(net952),
    .Y(_10304_));
 sg13g2_o21ai_1 _15932_ (.B1(_10304_),
    .Y(_10305_),
    .A1(_09871_),
    .A2(_10297_));
 sg13g2_inv_1 _15933_ (.Y(_10306_),
    .A(_00232_));
 sg13g2_a221oi_1 _15934_ (.B2(\top_ihp.wb_coproc.dat_o[1] ),
    .C1(net790),
    .B1(net859),
    .A1(net905),
    .Y(_10307_),
    .A2(_10306_));
 sg13g2_a21oi_1 _15935_ (.A1(_00231_),
    .A2(net790),
    .Y(_10308_),
    .B1(_10307_));
 sg13g2_nand2_1 _15936_ (.Y(_10309_),
    .A(net791),
    .B(_10308_));
 sg13g2_o21ai_1 _15937_ (.B1(_10309_),
    .Y(_10310_),
    .A1(_00230_),
    .A2(net791));
 sg13g2_a22oi_1 _15938_ (.Y(_10311_),
    .B1(_09957_),
    .B2(_10310_),
    .A2(\top_ihp.wb_dati_uart[1] ),
    .A1(net1001));
 sg13g2_a221oi_1 _15939_ (.B2(_09849_),
    .C1(net902),
    .B1(_10311_),
    .A1(net954),
    .Y(_10312_),
    .A2(_10305_));
 sg13g2_xnor2_1 _15940_ (.Y(_10313_),
    .A(_08318_),
    .B(_08605_));
 sg13g2_nor2_1 _15941_ (.A(net872),
    .B(_10313_),
    .Y(_10314_));
 sg13g2_o21ai_1 _15942_ (.B1(net949),
    .Y(_10315_),
    .A1(_10312_),
    .A2(_10314_));
 sg13g2_a21oi_2 _15943_ (.B1(net876),
    .Y(_10316_),
    .A2(_10315_),
    .A1(_10288_));
 sg13g2_a21oi_1 _15944_ (.A1(_08317_),
    .A2(net874),
    .Y(_10317_),
    .B1(_10316_));
 sg13g2_buf_1 _15945_ (.A(_10317_),
    .X(_10318_));
 sg13g2_buf_1 _15946_ (.A(net274),
    .X(_10319_));
 sg13g2_nand2_1 _15947_ (.Y(_10320_),
    .A(\top_ihp.oisc.regs[0][1] ),
    .B(net405));
 sg13g2_o21ai_1 _15948_ (.B1(_10320_),
    .Y(_00495_),
    .A1(net404),
    .A2(net139));
 sg13g2_nor2_1 _15949_ (.A(_08245_),
    .B(_08246_),
    .Y(_10321_));
 sg13g2_or2_1 _15950_ (.X(_10322_),
    .B(_08247_),
    .A(_10321_));
 sg13g2_buf_1 _15951_ (.A(_10322_),
    .X(_10323_));
 sg13g2_nor2_1 _15952_ (.A(_09678_),
    .B(_10227_),
    .Y(_10324_));
 sg13g2_or2_1 _15953_ (.X(_10325_),
    .B(_10324_),
    .A(_10323_));
 sg13g2_xor2_1 _15954_ (.B(_10325_),
    .A(_08491_),
    .X(_10326_));
 sg13g2_nand2_1 _15955_ (.Y(_10327_),
    .A(_10264_),
    .B(_10326_));
 sg13g2_nand2_1 _15956_ (.Y(_10328_),
    .A(_09800_),
    .B(_09946_));
 sg13g2_a21o_1 _15957_ (.A2(_10328_),
    .A1(_10043_),
    .B1(_09880_),
    .X(_10329_));
 sg13g2_buf_1 _15958_ (.A(_10329_),
    .X(_10330_));
 sg13g2_buf_1 _15959_ (.A(_10330_),
    .X(_10331_));
 sg13g2_a21oi_1 _15960_ (.A1(_09796_),
    .A2(net858),
    .Y(_10332_),
    .B1(net822));
 sg13g2_inv_1 _15961_ (.Y(_10333_),
    .A(_00149_));
 sg13g2_a221oi_1 _15962_ (.B2(\top_ihp.wb_coproc.dat_o[20] ),
    .C1(net825),
    .B1(net859),
    .A1(net905),
    .Y(_10334_),
    .A2(_10333_));
 sg13g2_a21oi_1 _15963_ (.A1(_00148_),
    .A2(net790),
    .Y(_10335_),
    .B1(_10334_));
 sg13g2_nor2_1 _15964_ (.A(_00147_),
    .B(net824),
    .Y(_10336_));
 sg13g2_a21oi_1 _15965_ (.A1(net791),
    .A2(_10335_),
    .Y(_10337_),
    .B1(_10336_));
 sg13g2_nor2_1 _15966_ (.A(net906),
    .B(_10337_),
    .Y(_10338_));
 sg13g2_a21oi_1 _15967_ (.A1(net950),
    .A2(_10338_),
    .Y(_10339_),
    .B1(_10260_));
 sg13g2_nor3_1 _15968_ (.A(_10155_),
    .B(_10332_),
    .C(_10339_),
    .Y(_10340_));
 sg13g2_a22oi_1 _15969_ (.Y(_10341_),
    .B1(_10327_),
    .B2(_10340_),
    .A2(net880),
    .A1(net1056));
 sg13g2_buf_1 _15970_ (.A(_10341_),
    .X(_10342_));
 sg13g2_buf_2 _15971_ (.A(_10342_),
    .X(_10343_));
 sg13g2_nand2_1 _15972_ (.Y(_10344_),
    .A(\top_ihp.oisc.regs[0][20] ),
    .B(net405));
 sg13g2_o21ai_1 _15973_ (.B1(_10344_),
    .Y(_00496_),
    .A1(net404),
    .A2(net138));
 sg13g2_o21ai_1 _15974_ (.B1(_08644_),
    .Y(_10345_),
    .A1(_08496_),
    .A2(_08647_));
 sg13g2_xnor2_1 _15975_ (.Y(_10346_),
    .A(_08499_),
    .B(_10345_));
 sg13g2_inv_1 _15976_ (.Y(_10347_),
    .A(_00152_));
 sg13g2_a221oi_1 _15977_ (.B2(\top_ihp.wb_coproc.dat_o[21] ),
    .C1(net825),
    .B1(net859),
    .A1(net905),
    .Y(_10348_),
    .A2(_10347_));
 sg13g2_a21oi_1 _15978_ (.A1(_00151_),
    .A2(_09822_),
    .Y(_10349_),
    .B1(_10348_));
 sg13g2_nor2_1 _15979_ (.A(_00150_),
    .B(net824),
    .Y(_10350_));
 sg13g2_a21oi_1 _15980_ (.A1(net791),
    .A2(_10349_),
    .Y(_10351_),
    .B1(_10350_));
 sg13g2_nor2_1 _15981_ (.A(net906),
    .B(_10351_),
    .Y(_10352_));
 sg13g2_inv_1 _15982_ (.Y(_10353_),
    .A(_10198_));
 sg13g2_a21o_1 _15983_ (.A2(_10352_),
    .A1(net951),
    .B1(_10353_),
    .X(_10354_));
 sg13g2_mux2_1 _15984_ (.A0(_10346_),
    .A1(_10354_),
    .S(_10229_),
    .X(_10355_));
 sg13g2_buf_2 _15985_ (.A(_10355_),
    .X(_10356_));
 sg13g2_a21oi_1 _15986_ (.A1(_10279_),
    .A2(_10152_),
    .Y(_10357_),
    .B1(net822));
 sg13g2_nand2_1 _15987_ (.Y(_10358_),
    .A(_08235_),
    .B(net901));
 sg13g2_o21ai_1 _15988_ (.B1(_10358_),
    .Y(_10359_),
    .A1(_09786_),
    .A2(_10357_));
 sg13g2_o21ai_1 _15989_ (.B1(_10359_),
    .Y(_10360_),
    .A1(_10208_),
    .A2(_10356_));
 sg13g2_buf_1 _15990_ (.A(_10360_),
    .X(_10361_));
 sg13g2_buf_1 _15991_ (.A(net273),
    .X(_10362_));
 sg13g2_nand2_1 _15992_ (.Y(_10363_),
    .A(\top_ihp.oisc.regs[0][21] ),
    .B(net405));
 sg13g2_o21ai_1 _15993_ (.B1(_10363_),
    .Y(_00497_),
    .A1(net404),
    .A2(net137));
 sg13g2_xor2_1 _15994_ (.B(_08393_),
    .A(_08378_),
    .X(_10364_));
 sg13g2_inv_1 _15995_ (.Y(_10365_),
    .A(_00155_));
 sg13g2_a221oi_1 _15996_ (.B2(\top_ihp.wb_coproc.dat_o[22] ),
    .C1(net790),
    .B1(_09829_),
    .A1(_09825_),
    .Y(_10366_),
    .A2(_10365_));
 sg13g2_a21oi_1 _15997_ (.A1(_00154_),
    .A2(net790),
    .Y(_10367_),
    .B1(_10366_));
 sg13g2_nor2_1 _15998_ (.A(_00153_),
    .B(net791),
    .Y(_10368_));
 sg13g2_a21oi_1 _15999_ (.A1(net791),
    .A2(_10367_),
    .Y(_10369_),
    .B1(_10368_));
 sg13g2_nor2_1 _16000_ (.A(_09814_),
    .B(_10369_),
    .Y(_10370_));
 sg13g2_nand2_1 _16001_ (.Y(_10371_),
    .A(net950),
    .B(_10370_));
 sg13g2_nand3_1 _16002_ (.B(_10198_),
    .C(_10371_),
    .A(net873),
    .Y(_10372_));
 sg13g2_o21ai_1 _16003_ (.B1(_10372_),
    .Y(_10373_),
    .A1(_10110_),
    .A2(_10364_));
 sg13g2_buf_1 _16004_ (.A(\top_ihp.oisc.decoder.instruction[22] ),
    .X(_10374_));
 sg13g2_a21oi_1 _16005_ (.A1(_10374_),
    .A2(_10152_),
    .Y(_10375_),
    .B1(net822));
 sg13g2_nor2_1 _16006_ (.A(net907),
    .B(_10375_),
    .Y(_10376_));
 sg13g2_a21oi_1 _16007_ (.A1(_08391_),
    .A2(net901),
    .Y(_10377_),
    .B1(_10376_));
 sg13g2_a21o_1 _16008_ (.A2(_10373_),
    .A1(_09922_),
    .B1(_10377_),
    .X(_10378_));
 sg13g2_buf_1 _16009_ (.A(_10378_),
    .X(_10379_));
 sg13g2_buf_2 _16010_ (.A(_10379_),
    .X(_10380_));
 sg13g2_nand2_1 _16011_ (.Y(_10381_),
    .A(\top_ihp.oisc.regs[0][22] ),
    .B(net405));
 sg13g2_o21ai_1 _16012_ (.B1(_10381_),
    .Y(_00498_),
    .A1(net404),
    .A2(_10380_));
 sg13g2_nor2b_1 _16013_ (.A(_08526_),
    .B_N(_08599_),
    .Y(_10382_));
 sg13g2_xnor2_1 _16014_ (.Y(_10383_),
    .A(_08396_),
    .B(_10382_));
 sg13g2_nor2_1 _16015_ (.A(_09848_),
    .B(_09967_),
    .Y(_10384_));
 sg13g2_o21ai_1 _16016_ (.B1(net873),
    .Y(_10385_),
    .A1(_10353_),
    .A2(_10384_));
 sg13g2_o21ai_1 _16017_ (.B1(_10385_),
    .Y(_10386_),
    .A1(_10110_),
    .A2(_10383_));
 sg13g2_buf_1 _16018_ (.A(\top_ihp.oisc.decoder.instruction[23] ),
    .X(_10387_));
 sg13g2_a21oi_1 _16019_ (.A1(_10387_),
    .A2(net858),
    .Y(_10388_),
    .B1(net822));
 sg13g2_nand2_1 _16020_ (.Y(_10389_),
    .A(net1047),
    .B(net907));
 sg13g2_o21ai_1 _16021_ (.B1(_10389_),
    .Y(_10390_),
    .A1(_10155_),
    .A2(_10388_));
 sg13g2_o21ai_1 _16022_ (.B1(_10390_),
    .Y(_10391_),
    .A1(_10208_),
    .A2(_10386_));
 sg13g2_buf_1 _16023_ (.A(_10391_),
    .X(_10392_));
 sg13g2_buf_2 _16024_ (.A(_10392_),
    .X(_10393_));
 sg13g2_nand2_1 _16025_ (.Y(_10394_),
    .A(\top_ihp.oisc.regs[0][23] ),
    .B(net405));
 sg13g2_o21ai_1 _16026_ (.B1(_10394_),
    .Y(_00499_),
    .A1(net404),
    .A2(net271));
 sg13g2_buf_1 _16027_ (.A(\top_ihp.oisc.decoder.instruction[24] ),
    .X(_10395_));
 sg13g2_a21oi_1 _16028_ (.A1(_10395_),
    .A2(net858),
    .Y(_10396_),
    .B1(net822));
 sg13g2_a21oi_1 _16029_ (.A1(_08291_),
    .A2(_08272_),
    .Y(_10397_),
    .B1(_08275_));
 sg13g2_nand3b_1 _16030_ (.B(_08272_),
    .C(_08275_),
    .Y(_10398_),
    .A_N(_08282_));
 sg13g2_and2_1 _16031_ (.A(net1052),
    .B(_10398_),
    .X(_10399_));
 sg13g2_nor3_1 _16032_ (.A(_09678_),
    .B(_10397_),
    .C(_10399_),
    .Y(_10400_));
 sg13g2_nor3_1 _16033_ (.A(net1057),
    .B(_10323_),
    .C(_10400_),
    .Y(_10401_));
 sg13g2_o21ai_1 _16034_ (.B1(net1057),
    .Y(_10402_),
    .A1(_10323_),
    .A2(_10400_));
 sg13g2_o21ai_1 _16035_ (.B1(_10402_),
    .Y(_10403_),
    .A1(net1056),
    .A2(_10401_));
 sg13g2_nor2_1 _16036_ (.A(_08249_),
    .B(_08551_),
    .Y(_10404_));
 sg13g2_or2_1 _16037_ (.X(_10405_),
    .B(_08627_),
    .A(_08528_));
 sg13g2_a21oi_1 _16038_ (.A1(_10403_),
    .A2(_10404_),
    .Y(_10406_),
    .B1(_10405_));
 sg13g2_o21ai_1 _16039_ (.B1(_10406_),
    .Y(_10407_),
    .A1(_10193_),
    .A2(_09680_));
 sg13g2_xnor2_1 _16040_ (.Y(_10408_),
    .A(_08383_),
    .B(_10407_));
 sg13g2_nand2_1 _16041_ (.Y(_10409_),
    .A(_09982_),
    .B(_09836_));
 sg13g2_nand3_1 _16042_ (.B(_10198_),
    .C(_10409_),
    .A(net872),
    .Y(_10410_));
 sg13g2_o21ai_1 _16043_ (.B1(_10410_),
    .Y(_10411_),
    .A1(net873),
    .A2(_10408_));
 sg13g2_nor2_1 _16044_ (.A(net1048),
    .B(net875),
    .Y(_10412_));
 sg13g2_a221oi_1 _16045_ (.B2(_09922_),
    .C1(_10412_),
    .B1(_10411_),
    .A1(net875),
    .Y(_10413_),
    .A2(_10396_));
 sg13g2_buf_1 _16046_ (.A(_10413_),
    .X(_10414_));
 sg13g2_buf_2 _16047_ (.A(_10414_),
    .X(_10415_));
 sg13g2_buf_1 _16048_ (.A(net403),
    .X(_10416_));
 sg13g2_mux2_1 _16049_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[0][24] ),
    .S(net409),
    .X(_00500_));
 sg13g2_nand2_1 _16050_ (.Y(_10417_),
    .A(_08384_),
    .B(net874));
 sg13g2_buf_1 _16051_ (.A(\top_ihp.oisc.decoder.instruction[25] ),
    .X(_10418_));
 sg13g2_a21oi_1 _16052_ (.A1(_10418_),
    .A2(_10057_),
    .Y(_10419_),
    .B1(net822));
 sg13g2_a21oi_1 _16053_ (.A1(_10092_),
    .A2(_10295_),
    .Y(_10420_),
    .B1(_10260_));
 sg13g2_nor2_1 _16054_ (.A(net1048),
    .B(_08402_),
    .Y(_10421_));
 sg13g2_a21oi_1 _16055_ (.A1(_08381_),
    .A2(_10407_),
    .Y(_10422_),
    .B1(_10421_));
 sg13g2_xor2_1 _16056_ (.B(_10422_),
    .A(_08389_),
    .X(_10423_));
 sg13g2_nor2_2 _16057_ (.A(_10262_),
    .B(_10423_),
    .Y(_10424_));
 sg13g2_or4_1 _16058_ (.A(net907),
    .B(_10419_),
    .C(_10420_),
    .D(_10424_),
    .X(_10425_));
 sg13g2_buf_1 _16059_ (.A(_10425_),
    .X(_10426_));
 sg13g2_and2_1 _16060_ (.A(_10417_),
    .B(_10426_),
    .X(_10427_));
 sg13g2_buf_2 _16061_ (.A(_10427_),
    .X(_10428_));
 sg13g2_buf_8 _16062_ (.A(_10428_),
    .X(_10429_));
 sg13g2_nand2_1 _16063_ (.Y(_10430_),
    .A(\top_ihp.oisc.regs[0][25] ),
    .B(_10275_));
 sg13g2_o21ai_1 _16064_ (.B1(_10430_),
    .Y(_00501_),
    .A1(net404),
    .A2(net59));
 sg13g2_o21ai_1 _16065_ (.B1(_10198_),
    .Y(_10431_),
    .A1(net954),
    .A2(_09996_));
 sg13g2_nand2_1 _16066_ (.Y(_10432_),
    .A(_08502_),
    .B(_08503_));
 sg13g2_xnor2_1 _16067_ (.Y(_10433_),
    .A(_08410_),
    .B(_10432_));
 sg13g2_mux2_1 _16068_ (.A0(_10431_),
    .A1(_10433_),
    .S(net902),
    .X(_10434_));
 sg13g2_buf_1 _16069_ (.A(\top_ihp.oisc.decoder.instruction[26] ),
    .X(_10435_));
 sg13g2_a21oi_1 _16070_ (.A1(_10435_),
    .A2(net858),
    .Y(_10436_),
    .B1(net822));
 sg13g2_nand2_1 _16071_ (.Y(_10437_),
    .A(_08217_),
    .B(net907));
 sg13g2_o21ai_1 _16072_ (.B1(_10437_),
    .Y(_10438_),
    .A1(net901),
    .A2(_10436_));
 sg13g2_o21ai_1 _16073_ (.B1(_10438_),
    .Y(_10439_),
    .A1(_10208_),
    .A2(_10434_));
 sg13g2_buf_1 _16074_ (.A(_10439_),
    .X(_10440_));
 sg13g2_buf_2 _16075_ (.A(_10440_),
    .X(_10441_));
 sg13g2_nand2_1 _16076_ (.Y(_10442_),
    .A(\top_ihp.oisc.regs[0][26] ),
    .B(_10275_));
 sg13g2_o21ai_1 _16077_ (.B1(_10442_),
    .Y(_00502_),
    .A1(_10277_),
    .A2(net402));
 sg13g2_a21oi_1 _16078_ (.A1(\top_ihp.oisc.decoder.instruction[27] ),
    .A2(_10057_),
    .Y(_10443_),
    .B1(_10331_));
 sg13g2_a21oi_1 _16079_ (.A1(net1025),
    .A2(_10025_),
    .Y(_10444_),
    .B1(_10260_));
 sg13g2_or3_1 _16080_ (.A(_09784_),
    .B(_10443_),
    .C(_10444_),
    .X(_10445_));
 sg13g2_a21oi_1 _16081_ (.A1(_08602_),
    .A2(_10264_),
    .Y(_10446_),
    .B1(_10445_));
 sg13g2_buf_2 _16082_ (.A(_10446_),
    .X(_10447_));
 sg13g2_a21oi_1 _16083_ (.A1(net1046),
    .A2(net874),
    .Y(_10448_),
    .B1(_10447_));
 sg13g2_buf_2 _16084_ (.A(_10448_),
    .X(_10449_));
 sg13g2_buf_8 _16085_ (.A(_10449_),
    .X(_10450_));
 sg13g2_nand2_1 _16086_ (.Y(_10451_),
    .A(\top_ihp.oisc.regs[0][27] ),
    .B(net405));
 sg13g2_o21ai_1 _16087_ (.B1(_10451_),
    .Y(_00503_),
    .A1(net404),
    .A2(net31));
 sg13g2_a21oi_1 _16088_ (.A1(\top_ihp.oisc.decoder.instruction[28] ),
    .A2(_10057_),
    .Y(_10452_),
    .B1(_10331_));
 sg13g2_a21oi_1 _16089_ (.A1(_09982_),
    .A2(_10077_),
    .Y(_10453_),
    .B1(_10260_));
 sg13g2_nor3_1 _16090_ (.A(_09784_),
    .B(_10452_),
    .C(_10453_),
    .Y(_10454_));
 sg13g2_o21ai_1 _16091_ (.B1(_10454_),
    .Y(_10455_),
    .A1(_08540_),
    .A2(_10262_));
 sg13g2_buf_2 _16092_ (.A(_10455_),
    .X(_10456_));
 sg13g2_nand2_1 _16093_ (.Y(_10457_),
    .A(_08443_),
    .B(net874));
 sg13g2_and2_1 _16094_ (.A(_10456_),
    .B(_10457_),
    .X(_10458_));
 sg13g2_buf_8 _16095_ (.A(_10458_),
    .X(_10459_));
 sg13g2_buf_8 _16096_ (.A(_10459_),
    .X(_10460_));
 sg13g2_nand2_1 _16097_ (.Y(_10461_),
    .A(\top_ihp.oisc.regs[0][28] ),
    .B(net405));
 sg13g2_o21ai_1 _16098_ (.B1(_10461_),
    .Y(_00504_),
    .A1(net404),
    .A2(net30));
 sg13g2_a21oi_1 _16099_ (.A1(net950),
    .A2(_10106_),
    .Y(_10462_),
    .B1(_10260_));
 sg13g2_a21oi_1 _16100_ (.A1(\top_ihp.oisc.decoder.instruction[29] ),
    .A2(net858),
    .Y(_10463_),
    .B1(net822));
 sg13g2_a21oi_1 _16101_ (.A1(_08648_),
    .A2(_08654_),
    .Y(_10464_),
    .B1(_10262_));
 sg13g2_nor4_1 _16102_ (.A(_09884_),
    .B(_10462_),
    .C(_10463_),
    .D(_10464_),
    .Y(_10465_));
 sg13g2_a21oi_1 _16103_ (.A1(net1045),
    .A2(net874),
    .Y(_10466_),
    .B1(_10465_));
 sg13g2_buf_2 _16104_ (.A(_10466_),
    .X(_10467_));
 sg13g2_nand2_1 _16105_ (.Y(_10468_),
    .A(\top_ihp.oisc.regs[0][29] ),
    .B(net592));
 sg13g2_o21ai_1 _16106_ (.B1(_10468_),
    .Y(_00505_),
    .A1(_10277_),
    .A2(net269));
 sg13g2_nand2b_1 _16107_ (.Y(_10469_),
    .B(_08543_),
    .A_N(_08973_));
 sg13g2_buf_1 _16108_ (.A(_10469_),
    .X(_10470_));
 sg13g2_inv_1 _16109_ (.Y(_10471_),
    .A(_00101_));
 sg13g2_a22oi_1 _16110_ (.Y(_10472_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[2] ),
    .A2(_10471_),
    .A1(net1002));
 sg13g2_mux2_1 _16111_ (.A0(_00100_),
    .A1(_10472_),
    .S(_08958_),
    .X(_10473_));
 sg13g2_mux2_1 _16112_ (.A0(_00099_),
    .A1(_10473_),
    .S(net861),
    .X(_10474_));
 sg13g2_nand2_1 _16113_ (.Y(_10475_),
    .A(net1001),
    .B(\top_ihp.wb_dati_uart[2] ));
 sg13g2_o21ai_1 _16114_ (.B1(_10475_),
    .Y(_10476_),
    .A1(_10470_),
    .A2(_10474_));
 sg13g2_buf_1 _16115_ (.A(_10476_),
    .X(_10477_));
 sg13g2_o21ai_1 _16116_ (.B1(_09997_),
    .Y(_10478_),
    .A1(net952),
    .A2(_09996_));
 sg13g2_a22oi_1 _16117_ (.Y(_10479_),
    .B1(net749),
    .B2(net952),
    .A2(_10236_),
    .A1(_09872_));
 sg13g2_nor2_1 _16118_ (.A(net955),
    .B(_10479_),
    .Y(_10480_));
 sg13g2_a221oi_1 _16119_ (.B2(_09809_),
    .C1(_10480_),
    .B1(_10478_),
    .A1(_08658_),
    .Y(_10481_),
    .A2(_10477_));
 sg13g2_nor2_1 _16120_ (.A(_08319_),
    .B(_08323_),
    .Y(_10482_));
 sg13g2_a21oi_1 _16121_ (.A1(_08319_),
    .A2(_08323_),
    .Y(_10483_),
    .B1(_08318_));
 sg13g2_nor2_1 _16122_ (.A(_10482_),
    .B(_10483_),
    .Y(_10484_));
 sg13g2_xnor2_1 _16123_ (.Y(_10485_),
    .A(_09687_),
    .B(_10484_));
 sg13g2_nor2_1 _16124_ (.A(_09877_),
    .B(_10485_),
    .Y(_10486_));
 sg13g2_a21oi_1 _16125_ (.A1(net872),
    .A2(_10481_),
    .Y(_10487_),
    .B1(_10486_));
 sg13g2_and2_1 _16126_ (.A(net1036),
    .B(_09906_),
    .X(_10488_));
 sg13g2_a21oi_1 _16127_ (.A1(_09799_),
    .A2(_10374_),
    .Y(_10489_),
    .B1(_10488_));
 sg13g2_nand2_1 _16128_ (.Y(_10490_),
    .A(_09906_),
    .B(_10278_));
 sg13g2_o21ai_1 _16129_ (.B1(_10490_),
    .Y(_10491_),
    .A1(net1004),
    .A2(_10489_));
 sg13g2_nand2_1 _16130_ (.Y(_10492_),
    .A(net1006),
    .B(_10374_));
 sg13g2_o21ai_1 _16131_ (.B1(_10492_),
    .Y(_10493_),
    .A1(net1006),
    .A2(_00234_));
 sg13g2_a22oi_1 _16132_ (.Y(_10494_),
    .B1(_10493_),
    .B2(_10284_),
    .A2(_10491_),
    .A1(net1005));
 sg13g2_nand2_1 _16133_ (.Y(_10495_),
    .A(net1007),
    .B(_10494_));
 sg13g2_o21ai_1 _16134_ (.B1(_10495_),
    .Y(_10496_),
    .A1(_09788_),
    .A2(_10487_));
 sg13g2_nor2_1 _16135_ (.A(_09884_),
    .B(_10496_),
    .Y(_10497_));
 sg13g2_a21oi_1 _16136_ (.A1(net1050),
    .A2(net880),
    .Y(_10498_),
    .B1(_10497_));
 sg13g2_buf_1 _16137_ (.A(_10498_),
    .X(_10499_));
 sg13g2_buf_2 _16138_ (.A(_10499_),
    .X(_10500_));
 sg13g2_nand2_1 _16139_ (.Y(_10501_),
    .A(\top_ihp.oisc.regs[0][2] ),
    .B(net592));
 sg13g2_o21ai_1 _16140_ (.B1(_10501_),
    .Y(_00506_),
    .A1(net409),
    .A2(net136));
 sg13g2_a21oi_1 _16141_ (.A1(\top_ihp.oisc.decoder.instruction[30] ),
    .A2(_10057_),
    .Y(_10502_),
    .B1(_10330_));
 sg13g2_a21oi_1 _16142_ (.A1(net1025),
    .A2(_10139_),
    .Y(_10503_),
    .B1(_10260_));
 sg13g2_nor3_1 _16143_ (.A(_09784_),
    .B(_10502_),
    .C(_10503_),
    .Y(_10504_));
 sg13g2_o21ai_1 _16144_ (.B1(_10264_),
    .Y(_10505_),
    .A1(net1026),
    .A2(_08578_));
 sg13g2_a21o_1 _16145_ (.A2(_10504_),
    .A1(_08578_),
    .B1(net901),
    .X(_10506_));
 sg13g2_a22oi_1 _16146_ (.Y(_10507_),
    .B1(_10506_),
    .B2(net1026),
    .A2(_10505_),
    .A1(_10504_));
 sg13g2_buf_1 _16147_ (.A(_10507_),
    .X(_10508_));
 sg13g2_buf_2 _16148_ (.A(_10508_),
    .X(_10509_));
 sg13g2_nand2_1 _16149_ (.Y(_10510_),
    .A(\top_ihp.oisc.regs[0][30] ),
    .B(net592));
 sg13g2_o21ai_1 _16150_ (.B1(_10510_),
    .Y(_00507_),
    .A1(net409),
    .A2(net58));
 sg13g2_inv_1 _16151_ (.Y(_10511_),
    .A(\top_ihp.oisc.regs[0][31] ));
 sg13g2_mux2_1 _16152_ (.A0(_00177_),
    .A1(_09974_),
    .S(net791),
    .X(_10512_));
 sg13g2_nor3_1 _16153_ (.A(_09848_),
    .B(_09814_),
    .C(_10512_),
    .Y(_10513_));
 sg13g2_o21ai_1 _16154_ (.B1(net873),
    .Y(_10514_),
    .A1(_10353_),
    .A2(_10513_));
 sg13g2_nand2_1 _16155_ (.Y(_10515_),
    .A(_08444_),
    .B(_08538_));
 sg13g2_inv_1 _16156_ (.Y(_10516_),
    .A(_08443_));
 sg13g2_o21ai_1 _16157_ (.B1(_10516_),
    .Y(_10517_),
    .A1(_08444_),
    .A2(_08538_));
 sg13g2_nand3_1 _16158_ (.B(_10515_),
    .C(_10517_),
    .A(_08563_),
    .Y(_10518_));
 sg13g2_nand2b_1 _16159_ (.Y(_10519_),
    .B(_10518_),
    .A_N(_08567_));
 sg13g2_a21oi_1 _16160_ (.A1(net1026),
    .A2(_10519_),
    .Y(_10520_),
    .B1(_08549_));
 sg13g2_o21ai_1 _16161_ (.B1(_09688_),
    .Y(_10521_),
    .A1(net1026),
    .A2(_10519_));
 sg13g2_nor2_1 _16162_ (.A(_10520_),
    .B(_10521_),
    .Y(_10522_));
 sg13g2_o21ai_1 _16163_ (.B1(_10522_),
    .Y(_10523_),
    .A1(_08535_),
    .A2(_09682_));
 sg13g2_inv_1 _16164_ (.Y(_10524_),
    .A(_09688_));
 sg13g2_o21ai_1 _16165_ (.B1(_10524_),
    .Y(_10525_),
    .A1(_09696_),
    .A2(_09698_));
 sg13g2_nand3_1 _16166_ (.B(_10523_),
    .C(_10525_),
    .A(_10003_),
    .Y(_10526_));
 sg13g2_a21oi_1 _16167_ (.A1(_10514_),
    .A2(_10526_),
    .Y(_10527_),
    .B1(_09789_));
 sg13g2_inv_1 _16168_ (.Y(_10528_),
    .A(_10043_));
 sg13g2_a21oi_1 _16169_ (.A1(_09945_),
    .A2(_09891_),
    .Y(_10529_),
    .B1(net1005));
 sg13g2_nor3_1 _16170_ (.A(net949),
    .B(_10528_),
    .C(_10529_),
    .Y(_10530_));
 sg13g2_o21ai_1 _16171_ (.B1(_10042_),
    .Y(_10531_),
    .A1(_10527_),
    .A2(_10530_));
 sg13g2_buf_1 _16172_ (.A(_10531_),
    .X(_10532_));
 sg13g2_buf_2 _16173_ (.A(_10532_),
    .X(_10533_));
 sg13g2_and2_1 _16174_ (.A(_09673_),
    .B(net874),
    .X(_10534_));
 sg13g2_buf_2 _16175_ (.A(_10534_),
    .X(_10535_));
 sg13g2_buf_1 _16176_ (.A(_10535_),
    .X(_10536_));
 sg13g2_nor2_1 _16177_ (.A(_09943_),
    .B(net821),
    .Y(_10537_));
 sg13g2_a22oi_1 _16178_ (.Y(_00508_),
    .B1(net268),
    .B2(_10537_),
    .A2(_10011_),
    .A1(_10511_));
 sg13g2_inv_1 _16179_ (.Y(_10538_),
    .A(_00107_));
 sg13g2_a22oi_1 _16180_ (.Y(_10539_),
    .B1(net878),
    .B2(\top_ihp.wb_coproc.dat_o[3] ),
    .A2(_10538_),
    .A1(net956));
 sg13g2_mux2_1 _16181_ (.A0(_00106_),
    .A1(_10539_),
    .S(net823),
    .X(_10540_));
 sg13g2_mux2_1 _16182_ (.A0(_00105_),
    .A1(_10540_),
    .S(net845),
    .X(_10541_));
 sg13g2_nand2_1 _16183_ (.Y(_10542_),
    .A(net1001),
    .B(\top_ihp.wb_dati_uart[3] ));
 sg13g2_o21ai_1 _16184_ (.B1(_10542_),
    .Y(_10543_),
    .A1(_10470_),
    .A2(_10541_));
 sg13g2_buf_2 _16185_ (.A(_10543_),
    .X(_10544_));
 sg13g2_a22oi_1 _16186_ (.Y(_10545_),
    .B1(_10544_),
    .B2(net952),
    .A2(_10258_),
    .A1(net877));
 sg13g2_nand2_1 _16187_ (.Y(_10546_),
    .A(net1035),
    .B(_10025_));
 sg13g2_nand2_1 _16188_ (.Y(_10547_),
    .A(_10027_),
    .B(_10546_));
 sg13g2_a22oi_1 _16189_ (.Y(_10548_),
    .B1(_10547_),
    .B2(_09809_),
    .A2(_10544_),
    .A1(_08658_));
 sg13g2_o21ai_1 _16190_ (.B1(_10548_),
    .Y(_10549_),
    .A1(net955),
    .A2(_10545_));
 sg13g2_nor3_1 _16191_ (.A(net1050),
    .B(_10482_),
    .C(_10483_),
    .Y(_10550_));
 sg13g2_o21ai_1 _16192_ (.B1(net1050),
    .Y(_10551_),
    .A1(_10482_),
    .A2(_10483_));
 sg13g2_o21ai_1 _16193_ (.B1(_10551_),
    .Y(_10552_),
    .A1(_08330_),
    .A2(_10550_));
 sg13g2_xor2_1 _16194_ (.B(_10552_),
    .A(_09686_),
    .X(_10553_));
 sg13g2_mux2_1 _16195_ (.A0(_10549_),
    .A1(_10553_),
    .S(net902),
    .X(_10554_));
 sg13g2_and2_1 _16196_ (.A(net1036),
    .B(_09902_),
    .X(_10555_));
 sg13g2_a21oi_1 _16197_ (.A1(_09799_),
    .A2(_10387_),
    .Y(_10556_),
    .B1(_10555_));
 sg13g2_nand2_1 _16198_ (.Y(_10557_),
    .A(_09902_),
    .B(_10278_));
 sg13g2_o21ai_1 _16199_ (.B1(_10557_),
    .Y(_10558_),
    .A1(net1004),
    .A2(_10556_));
 sg13g2_nand2_1 _16200_ (.Y(_10559_),
    .A(net1006),
    .B(_10387_));
 sg13g2_o21ai_1 _16201_ (.B1(_10559_),
    .Y(_10560_),
    .A1(net1006),
    .A2(_00235_));
 sg13g2_a22oi_1 _16202_ (.Y(_10561_),
    .B1(_10560_),
    .B2(_10284_),
    .A2(_10558_),
    .A1(net1005));
 sg13g2_nand2_1 _16203_ (.Y(_10562_),
    .A(net958),
    .B(_10561_));
 sg13g2_o21ai_1 _16204_ (.B1(_10562_),
    .Y(_10563_),
    .A1(net958),
    .A2(_10554_));
 sg13g2_nand2_1 _16205_ (.Y(_10564_),
    .A(_08326_),
    .B(net876));
 sg13g2_o21ai_1 _16206_ (.B1(_10564_),
    .Y(_10565_),
    .A1(net880),
    .A2(_10563_));
 sg13g2_buf_1 _16207_ (.A(_10565_),
    .X(_10566_));
 sg13g2_buf_1 _16208_ (.A(_10566_),
    .X(_10567_));
 sg13g2_buf_1 _16209_ (.A(net135),
    .X(_10568_));
 sg13g2_mux2_1 _16210_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[0][3] ),
    .S(net409),
    .X(_00509_));
 sg13g2_and2_1 _16211_ (.A(net1036),
    .B(_09919_),
    .X(_10569_));
 sg13g2_a21oi_1 _16212_ (.A1(_09799_),
    .A2(_10395_),
    .Y(_10570_),
    .B1(_10569_));
 sg13g2_nand2_1 _16213_ (.Y(_10571_),
    .A(_09919_),
    .B(_10278_));
 sg13g2_o21ai_1 _16214_ (.B1(_10571_),
    .Y(_10572_),
    .A1(net1004),
    .A2(_10570_));
 sg13g2_nand2_1 _16215_ (.Y(_10573_),
    .A(net1006),
    .B(_10395_));
 sg13g2_o21ai_1 _16216_ (.B1(_10573_),
    .Y(_10574_),
    .A1(_09791_),
    .A2(_00236_));
 sg13g2_a22oi_1 _16217_ (.Y(_10575_),
    .B1(_10574_),
    .B2(_10284_),
    .A2(_10572_),
    .A1(net1005));
 sg13g2_inv_1 _16218_ (.Y(_10576_),
    .A(_00103_));
 sg13g2_nor2b_1 _16219_ (.A(_00104_),
    .B_N(net1002),
    .Y(_10577_));
 sg13g2_a21o_1 _16220_ (.A2(net904),
    .A1(\top_ihp.wb_coproc.dat_o[4] ),
    .B1(_10577_),
    .X(_10578_));
 sg13g2_mux2_1 _16221_ (.A0(_10576_),
    .A1(_10578_),
    .S(net846),
    .X(_10579_));
 sg13g2_nor2_1 _16222_ (.A(_00102_),
    .B(net861),
    .Y(_10580_));
 sg13g2_a21o_1 _16223_ (.A2(_10579_),
    .A1(net861),
    .B1(_10580_),
    .X(_10581_));
 sg13g2_a22oi_1 _16224_ (.Y(_10582_),
    .B1(_09957_),
    .B2(_10581_),
    .A2(\top_ihp.wb_dati_uart[4] ),
    .A1(net1001));
 sg13g2_buf_2 _16225_ (.A(_10582_),
    .X(_10583_));
 sg13g2_inv_1 _16226_ (.Y(_10584_),
    .A(_10583_));
 sg13g2_a22oi_1 _16227_ (.Y(_10585_),
    .B1(_10584_),
    .B2(net952),
    .A2(_10338_),
    .A1(net877));
 sg13g2_buf_1 _16228_ (.A(_10584_),
    .X(_10586_));
 sg13g2_a21o_1 _16229_ (.A2(_10077_),
    .A1(net1035),
    .B1(_10078_),
    .X(_10587_));
 sg13g2_a22oi_1 _16230_ (.Y(_10588_),
    .B1(_10587_),
    .B2(_09809_),
    .A2(_10586_),
    .A1(net1025));
 sg13g2_o21ai_1 _16231_ (.B1(_10588_),
    .Y(_10589_),
    .A1(net955),
    .A2(_10585_));
 sg13g2_a22oi_1 _16232_ (.Y(_10590_),
    .B1(_08335_),
    .B2(_08337_),
    .A2(_08333_),
    .A1(_08325_));
 sg13g2_xor2_1 _16233_ (.B(_10590_),
    .A(_08339_),
    .X(_10591_));
 sg13g2_xor2_1 _16234_ (.B(_10591_),
    .A(net1049),
    .X(_10592_));
 sg13g2_nor2_1 _16235_ (.A(_09877_),
    .B(_10592_),
    .Y(_10593_));
 sg13g2_a21oi_1 _16236_ (.A1(net872),
    .A2(_10589_),
    .Y(_10594_),
    .B1(_10593_));
 sg13g2_mux2_1 _16237_ (.A0(_10575_),
    .A1(_10594_),
    .S(net949),
    .X(_10595_));
 sg13g2_nand2_1 _16238_ (.Y(_10596_),
    .A(net1049),
    .B(net876));
 sg13g2_o21ai_1 _16239_ (.B1(_10596_),
    .Y(_10597_),
    .A1(net880),
    .A2(_10595_));
 sg13g2_buf_1 _16240_ (.A(_10597_),
    .X(_10598_));
 sg13g2_buf_2 _16241_ (.A(_10598_),
    .X(_10599_));
 sg13g2_buf_2 _16242_ (.A(net134),
    .X(_10600_));
 sg13g2_mux2_1 _16243_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[0][4] ),
    .S(net409),
    .X(_00510_));
 sg13g2_nor2_1 _16244_ (.A(_10590_),
    .B(_08361_),
    .Y(_10601_));
 sg13g2_nor2_1 _16245_ (.A(_08470_),
    .B(_10601_),
    .Y(_10602_));
 sg13g2_xor2_1 _16246_ (.B(_10602_),
    .A(_08342_),
    .X(_10603_));
 sg13g2_a21oi_1 _16247_ (.A1(_10418_),
    .A2(_09948_),
    .Y(_10604_),
    .B1(net872));
 sg13g2_a21o_1 _16248_ (.A2(_10604_),
    .A1(_10603_),
    .B1(net907),
    .X(_10605_));
 sg13g2_nor3_1 _16249_ (.A(_08363_),
    .B(net872),
    .C(_10603_),
    .Y(_10606_));
 sg13g2_buf_1 _16250_ (.A(\top_ihp.wb_dati_uart[5] ),
    .X(_10607_));
 sg13g2_inv_1 _16251_ (.Y(_10608_),
    .A(_00110_));
 sg13g2_a22oi_1 _16252_ (.Y(_10609_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[5] ),
    .A2(_10608_),
    .A1(net1002));
 sg13g2_mux2_1 _16253_ (.A0(_00109_),
    .A1(_10609_),
    .S(net823),
    .X(_10610_));
 sg13g2_mux2_1 _16254_ (.A0(_00108_),
    .A1(_10610_),
    .S(net845),
    .X(_10611_));
 sg13g2_inv_1 _16255_ (.Y(_10612_),
    .A(_10611_));
 sg13g2_a22oi_1 _16256_ (.Y(_10613_),
    .B1(_09957_),
    .B2(_10612_),
    .A2(_10607_),
    .A1(net1001));
 sg13g2_buf_1 _16257_ (.A(_10613_),
    .X(_10614_));
 sg13g2_nand2_1 _16258_ (.Y(_10615_),
    .A(net877),
    .B(_10352_));
 sg13g2_o21ai_1 _16259_ (.B1(_10615_),
    .Y(_10616_),
    .A1(net1003),
    .A2(_10614_));
 sg13g2_nand2_1 _16260_ (.Y(_10617_),
    .A(net1003),
    .B(_10106_));
 sg13g2_o21ai_1 _16261_ (.B1(_10617_),
    .Y(_10618_),
    .A1(net1003),
    .A2(_10100_));
 sg13g2_o21ai_1 _16262_ (.B1(net903),
    .Y(_10619_),
    .A1(net954),
    .A2(_10614_));
 sg13g2_a221oi_1 _16263_ (.B2(_09809_),
    .C1(_10619_),
    .B1(_10618_),
    .A1(_09869_),
    .Y(_10620_),
    .A2(_10616_));
 sg13g2_or3_1 _16264_ (.A(_09789_),
    .B(_10606_),
    .C(_10620_),
    .X(_10621_));
 sg13g2_a21oi_1 _16265_ (.A1(_10418_),
    .A2(_09948_),
    .Y(_10622_),
    .B1(net901));
 sg13g2_a22oi_1 _16266_ (.Y(_10623_),
    .B1(_10621_),
    .B2(_10622_),
    .A2(_10605_),
    .A1(_08363_));
 sg13g2_buf_1 _16267_ (.A(_10623_),
    .X(_10624_));
 sg13g2_buf_1 _16268_ (.A(_10624_),
    .X(_10625_));
 sg13g2_buf_1 _16269_ (.A(net267),
    .X(_10626_));
 sg13g2_mux2_1 _16270_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[0][5] ),
    .S(net409),
    .X(_00511_));
 sg13g2_or3_1 _16271_ (.A(net1029),
    .B(_10175_),
    .C(_10178_),
    .X(_10627_));
 sg13g2_nand2_1 _16272_ (.Y(_10628_),
    .A(_10179_),
    .B(_10627_));
 sg13g2_a21o_1 _16273_ (.A2(_09948_),
    .A1(_10435_),
    .B1(net872),
    .X(_10629_));
 sg13g2_o21ai_1 _16274_ (.B1(net875),
    .Y(_10630_),
    .A1(_10628_),
    .A2(_10629_));
 sg13g2_inv_1 _16275_ (.Y(_10631_),
    .A(_00113_));
 sg13g2_a22oi_1 _16276_ (.Y(_10632_),
    .B1(net904),
    .B2(\top_ihp.wb_coproc.dat_o[6] ),
    .A2(_10631_),
    .A1(net1002));
 sg13g2_mux2_1 _16277_ (.A0(_00112_),
    .A1(_10632_),
    .S(net823),
    .X(_10633_));
 sg13g2_mux2_1 _16278_ (.A0(_00111_),
    .A1(_10633_),
    .S(net845),
    .X(_10634_));
 sg13g2_nand2_1 _16279_ (.Y(_10635_),
    .A(net1001),
    .B(\top_ihp.wb_dati_uart[6] ));
 sg13g2_o21ai_1 _16280_ (.B1(_10635_),
    .Y(_10636_),
    .A1(_10470_),
    .A2(_10634_));
 sg13g2_buf_2 _16281_ (.A(_10636_),
    .X(_10637_));
 sg13g2_a22oi_1 _16282_ (.Y(_10638_),
    .B1(_10637_),
    .B2(net952),
    .A2(_10370_),
    .A1(net877));
 sg13g2_nand2_1 _16283_ (.Y(_10639_),
    .A(net1003),
    .B(_10139_));
 sg13g2_o21ai_1 _16284_ (.B1(_10639_),
    .Y(_10640_),
    .A1(net1003),
    .A2(_10133_));
 sg13g2_a221oi_1 _16285_ (.B2(_09809_),
    .C1(net902),
    .B1(_10640_),
    .A1(net951),
    .Y(_10641_),
    .A2(_10637_));
 sg13g2_o21ai_1 _16286_ (.B1(_10641_),
    .Y(_10642_),
    .A1(net955),
    .A2(_10638_));
 sg13g2_nand3_1 _16287_ (.B(net902),
    .C(_10628_),
    .A(_08345_),
    .Y(_10643_));
 sg13g2_nand3_1 _16288_ (.B(_10642_),
    .C(_10643_),
    .A(_10116_),
    .Y(_10644_));
 sg13g2_a21oi_1 _16289_ (.A1(_10435_),
    .A2(_09948_),
    .Y(_10645_),
    .B1(net901));
 sg13g2_a22oi_1 _16290_ (.Y(_10646_),
    .B1(_10644_),
    .B2(_10645_),
    .A2(_10630_),
    .A1(_08365_));
 sg13g2_buf_1 _16291_ (.A(_10646_),
    .X(_10647_));
 sg13g2_buf_2 _16292_ (.A(_10647_),
    .X(_10648_));
 sg13g2_buf_2 _16293_ (.A(net132),
    .X(_10649_));
 sg13g2_mux2_1 _16294_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[0][6] ),
    .S(net591),
    .X(_00512_));
 sg13g2_nand2_1 _16295_ (.Y(_10650_),
    .A(_09950_),
    .B(_09958_));
 sg13g2_nand2_1 _16296_ (.Y(_10651_),
    .A(net1003),
    .B(_09869_));
 sg13g2_nand2_1 _16297_ (.Y(_10652_),
    .A(net955),
    .B(_09976_));
 sg13g2_o21ai_1 _16298_ (.B1(_10652_),
    .Y(_10653_),
    .A1(_09967_),
    .A2(_10651_));
 sg13g2_a22oi_1 _16299_ (.Y(_10654_),
    .B1(_10653_),
    .B2(net954),
    .A2(_10650_),
    .A1(_09849_));
 sg13g2_xor2_1 _16300_ (.B(_10181_),
    .A(_08344_),
    .X(_10655_));
 sg13g2_nor2_1 _16301_ (.A(net903),
    .B(_10655_),
    .Y(_10656_));
 sg13g2_a21oi_1 _16302_ (.A1(net872),
    .A2(_10654_),
    .Y(_10657_),
    .B1(_10656_));
 sg13g2_a22oi_1 _16303_ (.Y(_10658_),
    .B1(_10657_),
    .B2(_10116_),
    .A2(_09948_),
    .A1(\top_ihp.oisc.decoder.instruction[27] ));
 sg13g2_nor2_1 _16304_ (.A(_08314_),
    .B(net875),
    .Y(_10659_));
 sg13g2_a21o_1 _16305_ (.A2(_10658_),
    .A1(net875),
    .B1(_10659_),
    .X(_10660_));
 sg13g2_buf_1 _16306_ (.A(_10660_),
    .X(_10661_));
 sg13g2_buf_1 _16307_ (.A(_10661_),
    .X(_10662_));
 sg13g2_nand2_1 _16308_ (.Y(_10663_),
    .A(\top_ihp.oisc.regs[0][7] ),
    .B(net592));
 sg13g2_o21ai_1 _16309_ (.B1(_10663_),
    .Y(_00513_),
    .A1(_09944_),
    .A2(net401));
 sg13g2_inv_1 _16310_ (.Y(_10664_),
    .A(_09842_));
 sg13g2_a21o_1 _16311_ (.A2(net877),
    .A1(_09836_),
    .B1(_09843_),
    .X(_10665_));
 sg13g2_a221oi_1 _16312_ (.B2(_09999_),
    .C1(_09980_),
    .B1(_10665_),
    .A1(net950),
    .Y(_10666_),
    .A2(_10664_));
 sg13g2_o21ai_1 _16313_ (.B1(_08369_),
    .Y(_10667_),
    .A1(_08316_),
    .A2(_10181_));
 sg13g2_xnor2_1 _16314_ (.Y(_10668_),
    .A(_08352_),
    .B(_10667_));
 sg13g2_o21ai_1 _16315_ (.B1(_09880_),
    .Y(_10669_),
    .A1(net873),
    .A2(_10668_));
 sg13g2_a21oi_1 _16316_ (.A1(\top_ihp.oisc.decoder.instruction[28] ),
    .A2(_09948_),
    .Y(_10670_),
    .B1(net907));
 sg13g2_o21ai_1 _16317_ (.B1(_10670_),
    .Y(_10671_),
    .A1(_10666_),
    .A2(_10669_));
 sg13g2_o21ai_1 _16318_ (.B1(_10671_),
    .Y(_10672_),
    .A1(_08350_),
    .A2(net875));
 sg13g2_buf_1 _16319_ (.A(_10672_),
    .X(_10673_));
 sg13g2_buf_2 _16320_ (.A(_10673_),
    .X(_10674_));
 sg13g2_nand2_1 _16321_ (.Y(_10675_),
    .A(\top_ihp.oisc.regs[0][8] ),
    .B(net592));
 sg13g2_o21ai_1 _16322_ (.B1(_10675_),
    .Y(_00514_),
    .A1(_09944_),
    .A2(_10674_));
 sg13g2_inv_1 _16323_ (.Y(_10676_),
    .A(_10303_));
 sg13g2_nand2_1 _16324_ (.Y(_10677_),
    .A(net877),
    .B(_10295_));
 sg13g2_o21ai_1 _16325_ (.B1(_10677_),
    .Y(_10678_),
    .A1(net1003),
    .A2(_10303_));
 sg13g2_a22oi_1 _16326_ (.Y(_10679_),
    .B1(_10678_),
    .B2(net999),
    .A2(_10676_),
    .A1(net951));
 sg13g2_nand2_1 _16327_ (.Y(_10680_),
    .A(_08478_),
    .B(_08482_));
 sg13g2_xnor2_1 _16328_ (.Y(_10681_),
    .A(_08355_),
    .B(_10680_));
 sg13g2_a221oi_1 _16329_ (.B2(net902),
    .C1(_09788_),
    .B1(_10681_),
    .A1(_09981_),
    .Y(_10682_),
    .A2(_10679_));
 sg13g2_a21oi_1 _16330_ (.A1(\top_ihp.oisc.decoder.instruction[29] ),
    .A2(_09948_),
    .Y(_10683_),
    .B1(_10682_));
 sg13g2_nand2_1 _16331_ (.Y(_10684_),
    .A(_08353_),
    .B(net876));
 sg13g2_o21ai_1 _16332_ (.B1(_10684_),
    .Y(_10685_),
    .A1(net880),
    .A2(_10683_));
 sg13g2_buf_1 _16333_ (.A(_10685_),
    .X(_10686_));
 sg13g2_buf_1 _16334_ (.A(_10686_),
    .X(_10687_));
 sg13g2_buf_1 _16335_ (.A(net131),
    .X(_10688_));
 sg13g2_mux2_1 _16336_ (.A0(_10688_),
    .A1(\top_ihp.oisc.regs[0][9] ),
    .S(net591),
    .X(_00515_));
 sg13g2_nand3_1 _16337_ (.B(net1004),
    .C(_09891_),
    .A(_09670_),
    .Y(_10689_));
 sg13g2_buf_1 _16338_ (.A(_10689_),
    .X(_10690_));
 sg13g2_nand2b_1 _16339_ (.Y(_10691_),
    .B(_09910_),
    .A_N(_09905_));
 sg13g2_inv_1 _16340_ (.Y(_10692_),
    .A(_09913_));
 sg13g2_a21oi_1 _16341_ (.A1(_10690_),
    .A2(_10691_),
    .Y(_10693_),
    .B1(_10692_));
 sg13g2_buf_2 _16342_ (.A(_10693_),
    .X(_10694_));
 sg13g2_and2_1 _16343_ (.A(_09937_),
    .B(_09934_),
    .X(_10695_));
 sg13g2_buf_1 _16344_ (.A(_10695_),
    .X(_10696_));
 sg13g2_and2_1 _16345_ (.A(_09929_),
    .B(net740),
    .X(_10697_));
 sg13g2_buf_1 _16346_ (.A(_10697_),
    .X(_10698_));
 sg13g2_nand2_1 _16347_ (.Y(_10699_),
    .A(_10694_),
    .B(_10698_));
 sg13g2_buf_1 _16348_ (.A(_10699_),
    .X(_10700_));
 sg13g2_buf_1 _16349_ (.A(_10700_),
    .X(_10701_));
 sg13g2_buf_1 _16350_ (.A(_10700_),
    .X(_10702_));
 sg13g2_nand2_1 _16351_ (.Y(_10703_),
    .A(_00267_),
    .B(net589));
 sg13g2_o21ai_1 _16352_ (.B1(_10703_),
    .Y(_00516_),
    .A1(net64),
    .A2(_10701_));
 sg13g2_buf_2 _16353_ (.A(_10008_),
    .X(_10704_));
 sg13g2_a21o_1 _16354_ (.A2(_10691_),
    .A1(_10690_),
    .B1(_10692_),
    .X(_10705_));
 sg13g2_buf_1 _16355_ (.A(_10705_),
    .X(_10706_));
 sg13g2_nand2_1 _16356_ (.Y(_10707_),
    .A(_09929_),
    .B(_10696_));
 sg13g2_nor2_1 _16357_ (.A(_10706_),
    .B(_10707_),
    .Y(_10708_));
 sg13g2_buf_2 _16358_ (.A(_10708_),
    .X(_10709_));
 sg13g2_mux2_1 _16359_ (.A0(\top_ihp.oisc.regs[10][10] ),
    .A1(net130),
    .S(_10709_),
    .X(_00517_));
 sg13g2_nand2_1 _16360_ (.Y(_10710_),
    .A(\top_ihp.oisc.regs[10][11] ),
    .B(net589));
 sg13g2_o21ai_1 _16361_ (.B1(_10710_),
    .Y(_00518_),
    .A1(net62),
    .A2(_10701_));
 sg13g2_nand2_1 _16362_ (.Y(_10711_),
    .A(\top_ihp.oisc.regs[10][12] ),
    .B(net589));
 sg13g2_o21ai_1 _16363_ (.B1(_10711_),
    .Y(_00519_),
    .A1(net61),
    .A2(net590));
 sg13g2_nand2_1 _16364_ (.Y(_10712_),
    .A(\top_ihp.oisc.regs[10][13] ),
    .B(_10702_));
 sg13g2_o21ai_1 _16365_ (.B1(_10712_),
    .Y(_00520_),
    .A1(net278),
    .A2(net590));
 sg13g2_nand2_1 _16366_ (.Y(_10713_),
    .A(\top_ihp.oisc.regs[10][14] ),
    .B(_10702_));
 sg13g2_o21ai_1 _16367_ (.B1(_10713_),
    .Y(_00521_),
    .A1(net277),
    .A2(net590));
 sg13g2_buf_1 _16368_ (.A(_10700_),
    .X(_10714_));
 sg13g2_nand2_1 _16369_ (.Y(_10715_),
    .A(\top_ihp.oisc.regs[10][15] ),
    .B(_10714_));
 sg13g2_o21ai_1 _16370_ (.B1(_10715_),
    .Y(_00522_),
    .A1(net407),
    .A2(net590));
 sg13g2_nand2_1 _16371_ (.Y(_10716_),
    .A(\top_ihp.oisc.regs[10][16] ),
    .B(net588));
 sg13g2_o21ai_1 _16372_ (.B1(_10716_),
    .Y(_00523_),
    .A1(net140),
    .A2(net590));
 sg13g2_nand2_1 _16373_ (.Y(_10717_),
    .A(\top_ihp.oisc.regs[10][17] ),
    .B(net588));
 sg13g2_o21ai_1 _16374_ (.B1(_10717_),
    .Y(_00524_),
    .A1(net406),
    .A2(net590));
 sg13g2_nand2_1 _16375_ (.Y(_10718_),
    .A(\top_ihp.oisc.regs[10][18] ),
    .B(net588));
 sg13g2_o21ai_1 _16376_ (.B1(_10718_),
    .Y(_00525_),
    .A1(net275),
    .A2(net590));
 sg13g2_buf_1 _16377_ (.A(_10700_),
    .X(_10719_));
 sg13g2_nand2_1 _16378_ (.Y(_10720_),
    .A(\top_ihp.oisc.regs[10][19] ),
    .B(net588));
 sg13g2_o21ai_1 _16379_ (.B1(_10720_),
    .Y(_00526_),
    .A1(net60),
    .A2(net587));
 sg13g2_nand2_1 _16380_ (.Y(_10721_),
    .A(\top_ihp.oisc.regs[10][1] ),
    .B(net588));
 sg13g2_o21ai_1 _16381_ (.B1(_10721_),
    .Y(_00527_),
    .A1(net139),
    .A2(net587));
 sg13g2_nand2_1 _16382_ (.Y(_10722_),
    .A(\top_ihp.oisc.regs[10][20] ),
    .B(net588));
 sg13g2_o21ai_1 _16383_ (.B1(_10722_),
    .Y(_00528_),
    .A1(net138),
    .A2(net587));
 sg13g2_nand2_1 _16384_ (.Y(_10723_),
    .A(\top_ihp.oisc.regs[10][21] ),
    .B(net588));
 sg13g2_o21ai_1 _16385_ (.B1(_10723_),
    .Y(_00529_),
    .A1(net137),
    .A2(net587));
 sg13g2_nand2_1 _16386_ (.Y(_10724_),
    .A(\top_ihp.oisc.regs[10][22] ),
    .B(_10714_));
 sg13g2_o21ai_1 _16387_ (.B1(_10724_),
    .Y(_00530_),
    .A1(net272),
    .A2(net587));
 sg13g2_nand2_1 _16388_ (.Y(_10725_),
    .A(\top_ihp.oisc.regs[10][23] ),
    .B(net588));
 sg13g2_o21ai_1 _16389_ (.B1(_10725_),
    .Y(_00531_),
    .A1(net271),
    .A2(net587));
 sg13g2_buf_2 _16390_ (.A(_10414_),
    .X(_10726_));
 sg13g2_mux2_1 _16391_ (.A0(\top_ihp.oisc.regs[10][24] ),
    .A1(net400),
    .S(_10709_),
    .X(_00532_));
 sg13g2_buf_1 _16392_ (.A(_10700_),
    .X(_10727_));
 sg13g2_nand2_1 _16393_ (.Y(_10728_),
    .A(\top_ihp.oisc.regs[10][25] ),
    .B(net586));
 sg13g2_o21ai_1 _16394_ (.B1(_10728_),
    .Y(_00533_),
    .A1(net59),
    .A2(net587));
 sg13g2_nand2_1 _16395_ (.Y(_10729_),
    .A(\top_ihp.oisc.regs[10][26] ),
    .B(net586));
 sg13g2_o21ai_1 _16396_ (.B1(_10729_),
    .Y(_00534_),
    .A1(net402),
    .A2(net587));
 sg13g2_nand2_1 _16397_ (.Y(_10730_),
    .A(\top_ihp.oisc.regs[10][27] ),
    .B(net586));
 sg13g2_o21ai_1 _16398_ (.B1(_10730_),
    .Y(_00535_),
    .A1(net31),
    .A2(_10719_));
 sg13g2_nand2_1 _16399_ (.Y(_10731_),
    .A(\top_ihp.oisc.regs[10][28] ),
    .B(net586));
 sg13g2_o21ai_1 _16400_ (.B1(_10731_),
    .Y(_00536_),
    .A1(net30),
    .A2(_10719_));
 sg13g2_nand2_1 _16401_ (.Y(_10732_),
    .A(\top_ihp.oisc.regs[10][29] ),
    .B(net586));
 sg13g2_o21ai_1 _16402_ (.B1(_10732_),
    .Y(_00537_),
    .A1(net269),
    .A2(net589));
 sg13g2_nand2_1 _16403_ (.Y(_10733_),
    .A(\top_ihp.oisc.regs[10][2] ),
    .B(_10727_));
 sg13g2_o21ai_1 _16404_ (.B1(_10733_),
    .Y(_00538_),
    .A1(net136),
    .A2(net589));
 sg13g2_nand2_1 _16405_ (.Y(_10734_),
    .A(\top_ihp.oisc.regs[10][30] ),
    .B(net586));
 sg13g2_o21ai_1 _16406_ (.B1(_10734_),
    .Y(_00539_),
    .A1(net58),
    .A2(net589));
 sg13g2_inv_1 _16407_ (.Y(_10735_),
    .A(\top_ihp.oisc.regs[10][31] ));
 sg13g2_nor2_1 _16408_ (.A(net821),
    .B(net586),
    .Y(_10736_));
 sg13g2_buf_1 _16409_ (.A(_10532_),
    .X(_10737_));
 sg13g2_buf_1 _16410_ (.A(net265),
    .X(_10738_));
 sg13g2_a22oi_1 _16411_ (.Y(_00540_),
    .B1(_10736_),
    .B2(net129),
    .A2(net590),
    .A1(_10735_));
 sg13g2_buf_2 _16412_ (.A(_10566_),
    .X(_10739_));
 sg13g2_mux2_1 _16413_ (.A0(\top_ihp.oisc.regs[10][3] ),
    .A1(net128),
    .S(_10709_),
    .X(_00541_));
 sg13g2_buf_2 _16414_ (.A(_10598_),
    .X(_10740_));
 sg13g2_mux2_1 _16415_ (.A0(\top_ihp.oisc.regs[10][4] ),
    .A1(net127),
    .S(_10709_),
    .X(_00542_));
 sg13g2_buf_2 _16416_ (.A(_10624_),
    .X(_10741_));
 sg13g2_mux2_1 _16417_ (.A0(\top_ihp.oisc.regs[10][5] ),
    .A1(net264),
    .S(_10709_),
    .X(_00543_));
 sg13g2_buf_2 _16418_ (.A(_10647_),
    .X(_10742_));
 sg13g2_mux2_1 _16419_ (.A0(\top_ihp.oisc.regs[10][6] ),
    .A1(net126),
    .S(_10709_),
    .X(_00544_));
 sg13g2_nand2_1 _16420_ (.Y(_10743_),
    .A(\top_ihp.oisc.regs[10][7] ),
    .B(_10727_));
 sg13g2_o21ai_1 _16421_ (.B1(_10743_),
    .Y(_00545_),
    .A1(net401),
    .A2(net589));
 sg13g2_nand2_1 _16422_ (.Y(_10744_),
    .A(\top_ihp.oisc.regs[10][8] ),
    .B(net586));
 sg13g2_o21ai_1 _16423_ (.B1(_10744_),
    .Y(_00546_),
    .A1(net266),
    .A2(net589));
 sg13g2_buf_2 _16424_ (.A(_10686_),
    .X(_10745_));
 sg13g2_mux2_1 _16425_ (.A0(\top_ihp.oisc.regs[10][9] ),
    .A1(net125),
    .S(_10709_),
    .X(_00547_));
 sg13g2_nor2_1 _16426_ (.A(_09937_),
    .B(_09932_),
    .Y(_10746_));
 sg13g2_buf_2 _16427_ (.A(_10746_),
    .X(_10747_));
 sg13g2_and2_1 _16428_ (.A(_09929_),
    .B(_10747_),
    .X(_10748_));
 sg13g2_buf_2 _16429_ (.A(_10748_),
    .X(_10749_));
 sg13g2_nand2_1 _16430_ (.Y(_10750_),
    .A(_10694_),
    .B(_10749_));
 sg13g2_buf_1 _16431_ (.A(_10750_),
    .X(_10751_));
 sg13g2_buf_1 _16432_ (.A(net662),
    .X(_10752_));
 sg13g2_buf_1 _16433_ (.A(_10750_),
    .X(_10753_));
 sg13g2_nand2_1 _16434_ (.Y(_10754_),
    .A(_00268_),
    .B(net661));
 sg13g2_o21ai_1 _16435_ (.B1(_10754_),
    .Y(_00548_),
    .A1(net64),
    .A2(net585));
 sg13g2_buf_2 _16436_ (.A(net662),
    .X(_10755_));
 sg13g2_mux2_1 _16437_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[11][10] ),
    .S(net584),
    .X(_00549_));
 sg13g2_nand2_1 _16438_ (.Y(_10756_),
    .A(\top_ihp.oisc.regs[11][11] ),
    .B(net661));
 sg13g2_o21ai_1 _16439_ (.B1(_10756_),
    .Y(_00550_),
    .A1(net62),
    .A2(net585));
 sg13g2_nand2_1 _16440_ (.Y(_10757_),
    .A(\top_ihp.oisc.regs[11][12] ),
    .B(net661));
 sg13g2_o21ai_1 _16441_ (.B1(_10757_),
    .Y(_00551_),
    .A1(net61),
    .A2(net585));
 sg13g2_nand2_1 _16442_ (.Y(_10758_),
    .A(\top_ihp.oisc.regs[11][13] ),
    .B(_10753_));
 sg13g2_o21ai_1 _16443_ (.B1(_10758_),
    .Y(_00552_),
    .A1(net278),
    .A2(net585));
 sg13g2_nand2_1 _16444_ (.Y(_10759_),
    .A(\top_ihp.oisc.regs[11][14] ),
    .B(net661));
 sg13g2_o21ai_1 _16445_ (.B1(_10759_),
    .Y(_00553_),
    .A1(net277),
    .A2(_10752_));
 sg13g2_nand2_1 _16446_ (.Y(_10760_),
    .A(\top_ihp.oisc.regs[11][15] ),
    .B(net661));
 sg13g2_o21ai_1 _16447_ (.B1(_10760_),
    .Y(_00554_),
    .A1(net407),
    .A2(net585));
 sg13g2_nand2_1 _16448_ (.Y(_10761_),
    .A(\top_ihp.oisc.regs[11][16] ),
    .B(net661));
 sg13g2_o21ai_1 _16449_ (.B1(_10761_),
    .Y(_00555_),
    .A1(net140),
    .A2(net585));
 sg13g2_nand2_1 _16450_ (.Y(_10762_),
    .A(\top_ihp.oisc.regs[11][17] ),
    .B(_10753_));
 sg13g2_o21ai_1 _16451_ (.B1(_10762_),
    .Y(_00556_),
    .A1(net406),
    .A2(net585));
 sg13g2_buf_1 _16452_ (.A(net662),
    .X(_10763_));
 sg13g2_nand2_1 _16453_ (.Y(_10764_),
    .A(\top_ihp.oisc.regs[11][18] ),
    .B(net583));
 sg13g2_o21ai_1 _16454_ (.B1(_10764_),
    .Y(_00557_),
    .A1(net275),
    .A2(_10752_));
 sg13g2_buf_2 _16455_ (.A(_10271_),
    .X(_10765_));
 sg13g2_mux2_1 _16456_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[11][19] ),
    .S(net584),
    .X(_00558_));
 sg13g2_nand2_1 _16457_ (.Y(_10766_),
    .A(_00269_),
    .B(net583));
 sg13g2_o21ai_1 _16458_ (.B1(_10766_),
    .Y(_00559_),
    .A1(_10316_),
    .A2(net585));
 sg13g2_buf_1 _16459_ (.A(net662),
    .X(_10767_));
 sg13g2_nand2_1 _16460_ (.Y(_10768_),
    .A(\top_ihp.oisc.regs[11][20] ),
    .B(net583));
 sg13g2_o21ai_1 _16461_ (.B1(_10768_),
    .Y(_00560_),
    .A1(net138),
    .A2(_10767_));
 sg13g2_nand2_1 _16462_ (.Y(_10769_),
    .A(\top_ihp.oisc.regs[11][21] ),
    .B(_10763_));
 sg13g2_o21ai_1 _16463_ (.B1(_10769_),
    .Y(_00561_),
    .A1(net137),
    .A2(net582));
 sg13g2_nand2_1 _16464_ (.Y(_10770_),
    .A(\top_ihp.oisc.regs[11][22] ),
    .B(net583));
 sg13g2_o21ai_1 _16465_ (.B1(_10770_),
    .Y(_00562_),
    .A1(net272),
    .A2(net582));
 sg13g2_nand2_1 _16466_ (.Y(_10771_),
    .A(\top_ihp.oisc.regs[11][23] ),
    .B(net583));
 sg13g2_o21ai_1 _16467_ (.B1(_10771_),
    .Y(_00563_),
    .A1(net271),
    .A2(net582));
 sg13g2_mux2_1 _16468_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[11][24] ),
    .S(net584),
    .X(_00564_));
 sg13g2_buf_8 _16469_ (.A(_10426_),
    .X(_10772_));
 sg13g2_buf_1 _16470_ (.A(net262),
    .X(_10773_));
 sg13g2_nand2_1 _16471_ (.Y(_10774_),
    .A(\top_ihp.oisc.regs[11][25] ),
    .B(net583));
 sg13g2_o21ai_1 _16472_ (.B1(_10774_),
    .Y(_00565_),
    .A1(net124),
    .A2(net582));
 sg13g2_nand2_1 _16473_ (.Y(_10775_),
    .A(\top_ihp.oisc.regs[11][26] ),
    .B(_10763_));
 sg13g2_o21ai_1 _16474_ (.B1(_10775_),
    .Y(_00566_),
    .A1(net402),
    .A2(net582));
 sg13g2_buf_2 _16475_ (.A(_10447_),
    .X(_10776_));
 sg13g2_mux2_1 _16476_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[11][27] ),
    .S(net584),
    .X(_00567_));
 sg13g2_nand2_1 _16477_ (.Y(_10777_),
    .A(\top_ihp.oisc.regs[11][28] ),
    .B(net583));
 sg13g2_o21ai_1 _16478_ (.B1(_10777_),
    .Y(_00568_),
    .A1(net30),
    .A2(_10767_));
 sg13g2_nand2_1 _16479_ (.Y(_10778_),
    .A(\top_ihp.oisc.regs[11][29] ),
    .B(net583));
 sg13g2_o21ai_1 _16480_ (.B1(_10778_),
    .Y(_00569_),
    .A1(net269),
    .A2(net582));
 sg13g2_buf_2 _16481_ (.A(_10499_),
    .X(_10779_));
 sg13g2_mux2_1 _16482_ (.A0(net122),
    .A1(_00270_),
    .S(net584),
    .X(_00570_));
 sg13g2_nand2_1 _16483_ (.Y(_10780_),
    .A(\top_ihp.oisc.regs[11][30] ),
    .B(net662));
 sg13g2_o21ai_1 _16484_ (.B1(_10780_),
    .Y(_00571_),
    .A1(net58),
    .A2(net582));
 sg13g2_nand2_1 _16485_ (.Y(_10781_),
    .A(\top_ihp.oisc.regs[11][31] ),
    .B(net662));
 sg13g2_o21ai_1 _16486_ (.B1(_10781_),
    .Y(_00572_),
    .A1(net268),
    .A2(net582));
 sg13g2_nand2_1 _16487_ (.Y(_10782_),
    .A(_00271_),
    .B(net662));
 sg13g2_o21ai_1 _16488_ (.B1(_10782_),
    .Y(_00573_),
    .A1(net57),
    .A2(net584));
 sg13g2_nand2_1 _16489_ (.Y(_10783_),
    .A(_00272_),
    .B(net662));
 sg13g2_o21ai_1 _16490_ (.B1(_10783_),
    .Y(_00574_),
    .A1(net56),
    .A2(net584));
 sg13g2_mux2_1 _16491_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[11][5] ),
    .S(net584),
    .X(_00575_));
 sg13g2_mux2_1 _16492_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[11][6] ),
    .S(net661),
    .X(_00576_));
 sg13g2_nand2_1 _16493_ (.Y(_10784_),
    .A(\top_ihp.oisc.regs[11][7] ),
    .B(_10751_));
 sg13g2_o21ai_1 _16494_ (.B1(_10784_),
    .Y(_00577_),
    .A1(net401),
    .A2(_10755_));
 sg13g2_nand2_1 _16495_ (.Y(_10785_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(_10751_));
 sg13g2_o21ai_1 _16496_ (.B1(_10785_),
    .Y(_00578_),
    .A1(net266),
    .A2(_10755_));
 sg13g2_mux2_1 _16497_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[11][9] ),
    .S(net661),
    .X(_00579_));
 sg13g2_nor3_1 _16498_ (.A(_09905_),
    .B(_09910_),
    .C(_09916_),
    .Y(_10786_));
 sg13g2_buf_2 _16499_ (.A(_10786_),
    .X(_10787_));
 sg13g2_nand2_1 _16500_ (.Y(_10788_),
    .A(_09941_),
    .B(_10787_));
 sg13g2_buf_1 _16501_ (.A(_10788_),
    .X(_10789_));
 sg13g2_buf_1 _16502_ (.A(net660),
    .X(_10790_));
 sg13g2_buf_2 _16503_ (.A(net660),
    .X(_10791_));
 sg13g2_nand2_1 _16504_ (.Y(_10792_),
    .A(_00273_),
    .B(net580));
 sg13g2_o21ai_1 _16505_ (.B1(_10792_),
    .Y(_00580_),
    .A1(net64),
    .A2(net581));
 sg13g2_nand2_1 _16506_ (.Y(_10793_),
    .A(_00274_),
    .B(net580));
 sg13g2_o21ai_1 _16507_ (.B1(_10793_),
    .Y(_00581_),
    .A1(net63),
    .A2(net581));
 sg13g2_buf_2 _16508_ (.A(net660),
    .X(_10794_));
 sg13g2_mux2_1 _16509_ (.A0(_10041_),
    .A1(_00275_),
    .S(net579),
    .X(_00582_));
 sg13g2_nand2_1 _16510_ (.Y(_10795_),
    .A(_00276_),
    .B(net580));
 sg13g2_o21ai_1 _16511_ (.B1(_10795_),
    .Y(_00583_),
    .A1(_10087_),
    .A2(net581));
 sg13g2_buf_1 _16512_ (.A(_10121_),
    .X(_10796_));
 sg13g2_mux2_1 _16513_ (.A0(net261),
    .A1(_00277_),
    .S(net579),
    .X(_00584_));
 sg13g2_buf_1 _16514_ (.A(_10158_),
    .X(_10797_));
 sg13g2_mux2_1 _16515_ (.A0(net260),
    .A1(_00278_),
    .S(_10794_),
    .X(_00585_));
 sg13g2_buf_2 _16516_ (.A(_10170_),
    .X(_10798_));
 sg13g2_mux2_1 _16517_ (.A0(net399),
    .A1(_00279_),
    .S(net579),
    .X(_00586_));
 sg13g2_nand2_1 _16518_ (.Y(_10799_),
    .A(_00280_),
    .B(net580));
 sg13g2_o21ai_1 _16519_ (.B1(_10799_),
    .Y(_00587_),
    .A1(_10202_),
    .A2(net581));
 sg13g2_buf_1 _16520_ (.A(_10223_),
    .X(_10800_));
 sg13g2_mux2_1 _16521_ (.A0(net398),
    .A1(_00281_),
    .S(net579),
    .X(_00588_));
 sg13g2_buf_1 _16522_ (.A(_10245_),
    .X(_10801_));
 sg13g2_mux2_1 _16523_ (.A0(net259),
    .A1(_00282_),
    .S(_10794_),
    .X(_00589_));
 sg13g2_nand2_1 _16524_ (.Y(_10802_),
    .A(_00283_),
    .B(net580));
 sg13g2_o21ai_1 _16525_ (.B1(_10802_),
    .Y(_00590_),
    .A1(net263),
    .A2(net581));
 sg13g2_nand2_1 _16526_ (.Y(_10803_),
    .A(_00284_),
    .B(net580));
 sg13g2_o21ai_1 _16527_ (.B1(_10803_),
    .Y(_00591_),
    .A1(_10316_),
    .A2(net581));
 sg13g2_buf_2 _16528_ (.A(_10342_),
    .X(_10804_));
 sg13g2_buf_2 _16529_ (.A(_10789_),
    .X(_10805_));
 sg13g2_mux2_1 _16530_ (.A0(net121),
    .A1(_00285_),
    .S(net578),
    .X(_00592_));
 sg13g2_nand2_1 _16531_ (.Y(_10806_),
    .A(_00286_),
    .B(net580));
 sg13g2_o21ai_1 _16532_ (.B1(_10806_),
    .Y(_00593_),
    .A1(_10356_),
    .A2(net581));
 sg13g2_buf_2 _16533_ (.A(_10379_),
    .X(_10807_));
 sg13g2_mux2_1 _16534_ (.A0(net258),
    .A1(_00287_),
    .S(net578),
    .X(_00594_));
 sg13g2_buf_1 _16535_ (.A(_10392_),
    .X(_10808_));
 sg13g2_mux2_1 _16536_ (.A0(net257),
    .A1(_00288_),
    .S(net578),
    .X(_00595_));
 sg13g2_nand2_1 _16537_ (.Y(_10809_),
    .A(_00289_),
    .B(net580));
 sg13g2_o21ai_1 _16538_ (.B1(_10809_),
    .Y(_00596_),
    .A1(net270),
    .A2(_10790_));
 sg13g2_mux2_1 _16539_ (.A0(_10424_),
    .A1(_00290_),
    .S(net578),
    .X(_00597_));
 sg13g2_buf_2 _16540_ (.A(_10440_),
    .X(_10810_));
 sg13g2_mux2_1 _16541_ (.A0(net397),
    .A1(_00291_),
    .S(net578),
    .X(_00598_));
 sg13g2_nand2_1 _16542_ (.Y(_10811_),
    .A(_00292_),
    .B(_10789_));
 sg13g2_o21ai_1 _16543_ (.B1(_10811_),
    .Y(_00599_),
    .A1(net123),
    .A2(_10790_));
 sg13g2_mux2_1 _16544_ (.A0(_10456_),
    .A1(_00293_),
    .S(_10805_),
    .X(_00600_));
 sg13g2_buf_2 _16545_ (.A(_10466_),
    .X(_10812_));
 sg13g2_mux2_1 _16546_ (.A0(net256),
    .A1(_00294_),
    .S(_10805_),
    .X(_00601_));
 sg13g2_mux2_1 _16547_ (.A0(net122),
    .A1(_00295_),
    .S(net578),
    .X(_00602_));
 sg13g2_buf_8 _16548_ (.A(_10508_),
    .X(_10813_));
 sg13g2_mux2_1 _16549_ (.A0(net53),
    .A1(_00296_),
    .S(net578),
    .X(_00603_));
 sg13g2_mux2_1 _16550_ (.A0(net265),
    .A1(_00297_),
    .S(net578),
    .X(_00604_));
 sg13g2_nand2_1 _16551_ (.Y(_10814_),
    .A(_00298_),
    .B(net660));
 sg13g2_o21ai_1 _16552_ (.B1(_10814_),
    .Y(_00605_),
    .A1(net57),
    .A2(net581));
 sg13g2_nand2_1 _16553_ (.Y(_10815_),
    .A(_00299_),
    .B(net660));
 sg13g2_o21ai_1 _16554_ (.B1(_10815_),
    .Y(_00606_),
    .A1(net56),
    .A2(net579));
 sg13g2_nand2_1 _16555_ (.Y(_10816_),
    .A(_00300_),
    .B(net660));
 sg13g2_o21ai_1 _16556_ (.B1(_10816_),
    .Y(_00607_),
    .A1(net133),
    .A2(net579));
 sg13g2_nand2_1 _16557_ (.Y(_10817_),
    .A(_00301_),
    .B(net660));
 sg13g2_o21ai_1 _16558_ (.B1(_10817_),
    .Y(_00608_),
    .A1(net55),
    .A2(net579));
 sg13g2_buf_2 _16559_ (.A(_10661_),
    .X(_10818_));
 sg13g2_mux2_1 _16560_ (.A0(net396),
    .A1(_00302_),
    .S(_10791_),
    .X(_00609_));
 sg13g2_buf_2 _16561_ (.A(_10673_),
    .X(_10819_));
 sg13g2_mux2_1 _16562_ (.A0(net255),
    .A1(_00303_),
    .S(_10791_),
    .X(_00610_));
 sg13g2_nand2_1 _16563_ (.Y(_10820_),
    .A(_00304_),
    .B(net660));
 sg13g2_o21ai_1 _16564_ (.B1(_10820_),
    .Y(_00611_),
    .A1(net54),
    .A2(net579));
 sg13g2_nor2b_1 _16565_ (.A(_09937_),
    .B_N(_09932_),
    .Y(_10821_));
 sg13g2_buf_2 _16566_ (.A(_10821_),
    .X(_10822_));
 sg13g2_and2_1 _16567_ (.A(_09929_),
    .B(_10822_),
    .X(_10823_));
 sg13g2_buf_1 _16568_ (.A(_10823_),
    .X(_10824_));
 sg13g2_nand2_1 _16569_ (.Y(_10825_),
    .A(_10787_),
    .B(_10824_));
 sg13g2_buf_1 _16570_ (.A(_10825_),
    .X(_10826_));
 sg13g2_buf_2 _16571_ (.A(net659),
    .X(_10827_));
 sg13g2_mux2_1 _16572_ (.A0(_09889_),
    .A1(\top_ihp.oisc.regs[13][0] ),
    .S(net577),
    .X(_00612_));
 sg13g2_buf_1 _16573_ (.A(net659),
    .X(_10828_));
 sg13g2_buf_2 _16574_ (.A(net659),
    .X(_10829_));
 sg13g2_nand2_1 _16575_ (.Y(_10830_),
    .A(_00305_),
    .B(net575));
 sg13g2_o21ai_1 _16576_ (.B1(_10830_),
    .Y(_00613_),
    .A1(_10010_),
    .A2(net576));
 sg13g2_mux2_1 _16577_ (.A0(_10041_),
    .A1(_00306_),
    .S(net577),
    .X(_00614_));
 sg13g2_nand2_1 _16578_ (.Y(_10831_),
    .A(_00307_),
    .B(net575));
 sg13g2_o21ai_1 _16579_ (.B1(_10831_),
    .Y(_00615_),
    .A1(_10087_),
    .A2(net576));
 sg13g2_mux2_1 _16580_ (.A0(net261),
    .A1(_00308_),
    .S(net577),
    .X(_00616_));
 sg13g2_mux2_1 _16581_ (.A0(net260),
    .A1(_00309_),
    .S(_10827_),
    .X(_00617_));
 sg13g2_mux2_1 _16582_ (.A0(net399),
    .A1(_00310_),
    .S(net577),
    .X(_00618_));
 sg13g2_nand2_1 _16583_ (.Y(_10832_),
    .A(_00311_),
    .B(net575));
 sg13g2_o21ai_1 _16584_ (.B1(_10832_),
    .Y(_00619_),
    .A1(_10202_),
    .A2(net576));
 sg13g2_mux2_1 _16585_ (.A0(net398),
    .A1(_00312_),
    .S(net577),
    .X(_00620_));
 sg13g2_mux2_1 _16586_ (.A0(net259),
    .A1(_00313_),
    .S(_10827_),
    .X(_00621_));
 sg13g2_nand2_1 _16587_ (.Y(_10833_),
    .A(_00314_),
    .B(net575));
 sg13g2_o21ai_1 _16588_ (.B1(_10833_),
    .Y(_00622_),
    .A1(_10765_),
    .A2(net576));
 sg13g2_buf_1 _16589_ (.A(net274),
    .X(_10834_));
 sg13g2_nand2_1 _16590_ (.Y(_10835_),
    .A(\top_ihp.oisc.regs[13][1] ),
    .B(net575));
 sg13g2_o21ai_1 _16591_ (.B1(_10835_),
    .Y(_00623_),
    .A1(net120),
    .A2(net576));
 sg13g2_buf_2 _16592_ (.A(net659),
    .X(_10836_));
 sg13g2_mux2_1 _16593_ (.A0(net121),
    .A1(_00315_),
    .S(net574),
    .X(_00624_));
 sg13g2_nand2_1 _16594_ (.Y(_10837_),
    .A(_00316_),
    .B(net575));
 sg13g2_o21ai_1 _16595_ (.B1(_10837_),
    .Y(_00625_),
    .A1(_10356_),
    .A2(net576));
 sg13g2_mux2_1 _16596_ (.A0(net258),
    .A1(_00317_),
    .S(net574),
    .X(_00626_));
 sg13g2_mux2_1 _16597_ (.A0(net257),
    .A1(_00318_),
    .S(net574),
    .X(_00627_));
 sg13g2_nand2_1 _16598_ (.Y(_10838_),
    .A(_00319_),
    .B(net575));
 sg13g2_o21ai_1 _16599_ (.B1(_10838_),
    .Y(_00628_),
    .A1(_10416_),
    .A2(_10828_));
 sg13g2_mux2_1 _16600_ (.A0(_10424_),
    .A1(_00320_),
    .S(net574),
    .X(_00629_));
 sg13g2_mux2_1 _16601_ (.A0(net397),
    .A1(_00321_),
    .S(net574),
    .X(_00630_));
 sg13g2_nand2_1 _16602_ (.Y(_10839_),
    .A(_00322_),
    .B(net575));
 sg13g2_o21ai_1 _16603_ (.B1(_10839_),
    .Y(_00631_),
    .A1(net123),
    .A2(_10828_));
 sg13g2_mux2_1 _16604_ (.A0(_10456_),
    .A1(_00323_),
    .S(_10836_),
    .X(_00632_));
 sg13g2_mux2_1 _16605_ (.A0(net256),
    .A1(_00324_),
    .S(_10836_),
    .X(_00633_));
 sg13g2_mux2_1 _16606_ (.A0(net122),
    .A1(_00325_),
    .S(net574),
    .X(_00634_));
 sg13g2_mux2_1 _16607_ (.A0(net53),
    .A1(_00326_),
    .S(net574),
    .X(_00635_));
 sg13g2_mux2_1 _16608_ (.A0(net265),
    .A1(_00327_),
    .S(net574),
    .X(_00636_));
 sg13g2_nand2_1 _16609_ (.Y(_10840_),
    .A(_00328_),
    .B(net659));
 sg13g2_o21ai_1 _16610_ (.B1(_10840_),
    .Y(_00637_),
    .A1(_10568_),
    .A2(net576));
 sg13g2_nand2_1 _16611_ (.Y(_10841_),
    .A(_00329_),
    .B(net659));
 sg13g2_o21ai_1 _16612_ (.B1(_10841_),
    .Y(_00638_),
    .A1(_10600_),
    .A2(net576));
 sg13g2_nand2_1 _16613_ (.Y(_10842_),
    .A(_00330_),
    .B(net659));
 sg13g2_o21ai_1 _16614_ (.B1(_10842_),
    .Y(_00639_),
    .A1(_10626_),
    .A2(net577));
 sg13g2_nand2_1 _16615_ (.Y(_10843_),
    .A(_00331_),
    .B(net659));
 sg13g2_o21ai_1 _16616_ (.B1(_10843_),
    .Y(_00640_),
    .A1(_10649_),
    .A2(net577));
 sg13g2_mux2_1 _16617_ (.A0(net396),
    .A1(_00332_),
    .S(_10829_),
    .X(_00641_));
 sg13g2_mux2_1 _16618_ (.A0(net255),
    .A1(_00333_),
    .S(_10829_),
    .X(_00642_));
 sg13g2_nand2_1 _16619_ (.Y(_10844_),
    .A(_00334_),
    .B(_10826_));
 sg13g2_o21ai_1 _16620_ (.B1(_10844_),
    .Y(_00643_),
    .A1(net54),
    .A2(net577));
 sg13g2_buf_2 _16621_ (.A(_09887_),
    .X(_10845_));
 sg13g2_or3_1 _16622_ (.A(_09905_),
    .B(_09910_),
    .C(_09916_),
    .X(_10846_));
 sg13g2_buf_2 _16623_ (.A(_10846_),
    .X(_10847_));
 sg13g2_nor2_1 _16624_ (.A(_10707_),
    .B(_10847_),
    .Y(_10848_));
 sg13g2_buf_2 _16625_ (.A(_10848_),
    .X(_10849_));
 sg13g2_mux2_1 _16626_ (.A0(\top_ihp.oisc.regs[14][0] ),
    .A1(net119),
    .S(net691),
    .X(_00644_));
 sg13g2_mux2_1 _16627_ (.A0(\top_ihp.oisc.regs[14][10] ),
    .A1(net130),
    .S(net691),
    .X(_00645_));
 sg13g2_nand2_1 _16628_ (.Y(_10850_),
    .A(_10698_),
    .B(_10787_));
 sg13g2_buf_2 _16629_ (.A(_10850_),
    .X(_10851_));
 sg13g2_buf_1 _16630_ (.A(_10851_),
    .X(_10852_));
 sg13g2_buf_1 _16631_ (.A(_10851_),
    .X(_10853_));
 sg13g2_nand2_1 _16632_ (.Y(_10854_),
    .A(\top_ihp.oisc.regs[14][11] ),
    .B(net572));
 sg13g2_o21ai_1 _16633_ (.B1(_10854_),
    .Y(_00646_),
    .A1(net62),
    .A2(net573));
 sg13g2_buf_1 _16634_ (.A(net141),
    .X(_10855_));
 sg13g2_nor2_1 _16635_ (.A(\top_ihp.oisc.regs[14][12] ),
    .B(_10848_),
    .Y(_10856_));
 sg13g2_a21oi_1 _16636_ (.A1(_10855_),
    .A2(net691),
    .Y(_00647_),
    .B1(_10856_));
 sg13g2_nand2_1 _16637_ (.Y(_10857_),
    .A(\top_ihp.oisc.regs[14][13] ),
    .B(net572));
 sg13g2_o21ai_1 _16638_ (.B1(_10857_),
    .Y(_00648_),
    .A1(net278),
    .A2(net573));
 sg13g2_nand2_1 _16639_ (.Y(_10858_),
    .A(\top_ihp.oisc.regs[14][14] ),
    .B(net572));
 sg13g2_o21ai_1 _16640_ (.B1(_10858_),
    .Y(_00649_),
    .A1(net277),
    .A2(_10852_));
 sg13g2_nand2_1 _16641_ (.Y(_10859_),
    .A(\top_ihp.oisc.regs[14][15] ),
    .B(net572));
 sg13g2_o21ai_1 _16642_ (.B1(_10859_),
    .Y(_00650_),
    .A1(net407),
    .A2(net573));
 sg13g2_nand2_1 _16643_ (.Y(_10860_),
    .A(\top_ihp.oisc.regs[14][16] ),
    .B(net572));
 sg13g2_o21ai_1 _16644_ (.B1(_10860_),
    .Y(_00651_),
    .A1(net140),
    .A2(net573));
 sg13g2_nand2_1 _16645_ (.Y(_10861_),
    .A(\top_ihp.oisc.regs[14][17] ),
    .B(net572));
 sg13g2_o21ai_1 _16646_ (.B1(_10861_),
    .Y(_00652_),
    .A1(net406),
    .A2(net573));
 sg13g2_nand2_1 _16647_ (.Y(_10862_),
    .A(\top_ihp.oisc.regs[14][18] ),
    .B(net572));
 sg13g2_o21ai_1 _16648_ (.B1(_10862_),
    .Y(_00653_),
    .A1(net275),
    .A2(net573));
 sg13g2_nand2_1 _16649_ (.Y(_10863_),
    .A(\top_ihp.oisc.regs[14][19] ),
    .B(net572));
 sg13g2_o21ai_1 _16650_ (.B1(_10863_),
    .Y(_00654_),
    .A1(net60),
    .A2(net573));
 sg13g2_buf_1 _16651_ (.A(_10851_),
    .X(_10864_));
 sg13g2_nand2_1 _16652_ (.Y(_10865_),
    .A(\top_ihp.oisc.regs[14][1] ),
    .B(net571));
 sg13g2_o21ai_1 _16653_ (.B1(_10865_),
    .Y(_00655_),
    .A1(net120),
    .A2(_10852_));
 sg13g2_buf_1 _16654_ (.A(_10851_),
    .X(_10866_));
 sg13g2_nand2_1 _16655_ (.Y(_10867_),
    .A(\top_ihp.oisc.regs[14][20] ),
    .B(net571));
 sg13g2_o21ai_1 _16656_ (.B1(_10867_),
    .Y(_00656_),
    .A1(net138),
    .A2(net570));
 sg13g2_nand2_1 _16657_ (.Y(_10868_),
    .A(\top_ihp.oisc.regs[14][21] ),
    .B(net571));
 sg13g2_o21ai_1 _16658_ (.B1(_10868_),
    .Y(_00657_),
    .A1(net137),
    .A2(net570));
 sg13g2_nand2_1 _16659_ (.Y(_10869_),
    .A(\top_ihp.oisc.regs[14][22] ),
    .B(net571));
 sg13g2_o21ai_1 _16660_ (.B1(_10869_),
    .Y(_00658_),
    .A1(net272),
    .A2(net570));
 sg13g2_nand2_1 _16661_ (.Y(_10870_),
    .A(\top_ihp.oisc.regs[14][23] ),
    .B(_10864_));
 sg13g2_o21ai_1 _16662_ (.B1(_10870_),
    .Y(_00659_),
    .A1(net271),
    .A2(net570));
 sg13g2_mux2_1 _16663_ (.A0(\top_ihp.oisc.regs[14][24] ),
    .A1(net400),
    .S(net691),
    .X(_00660_));
 sg13g2_nor2_1 _16664_ (.A(\top_ihp.oisc.regs[14][25] ),
    .B(_10848_),
    .Y(_10871_));
 sg13g2_a21oi_1 _16665_ (.A1(_10429_),
    .A2(net691),
    .Y(_00661_),
    .B1(_10871_));
 sg13g2_nand2_1 _16666_ (.Y(_10872_),
    .A(\top_ihp.oisc.regs[14][26] ),
    .B(net571));
 sg13g2_o21ai_1 _16667_ (.B1(_10872_),
    .Y(_00662_),
    .A1(net402),
    .A2(_10866_));
 sg13g2_nand2_1 _16668_ (.Y(_10873_),
    .A(\top_ihp.oisc.regs[14][27] ),
    .B(net571));
 sg13g2_o21ai_1 _16669_ (.B1(_10873_),
    .Y(_00663_),
    .A1(net31),
    .A2(net570));
 sg13g2_nand2_1 _16670_ (.Y(_10874_),
    .A(\top_ihp.oisc.regs[14][28] ),
    .B(net571));
 sg13g2_o21ai_1 _16671_ (.B1(_10874_),
    .Y(_00664_),
    .A1(_10460_),
    .A2(net570));
 sg13g2_nand2_1 _16672_ (.Y(_10875_),
    .A(\top_ihp.oisc.regs[14][29] ),
    .B(net571));
 sg13g2_o21ai_1 _16673_ (.B1(_10875_),
    .Y(_00665_),
    .A1(net269),
    .A2(net570));
 sg13g2_nand2_1 _16674_ (.Y(_10876_),
    .A(\top_ihp.oisc.regs[14][2] ),
    .B(_10864_));
 sg13g2_o21ai_1 _16675_ (.B1(_10876_),
    .Y(_00666_),
    .A1(net136),
    .A2(_10866_));
 sg13g2_nand2_1 _16676_ (.Y(_10877_),
    .A(\top_ihp.oisc.regs[14][30] ),
    .B(_10851_));
 sg13g2_o21ai_1 _16677_ (.B1(_10877_),
    .Y(_00667_),
    .A1(net58),
    .A2(net570));
 sg13g2_inv_1 _16678_ (.Y(_10878_),
    .A(\top_ihp.oisc.regs[14][31] ));
 sg13g2_nor2_1 _16679_ (.A(net821),
    .B(_10851_),
    .Y(_10879_));
 sg13g2_a22oi_1 _16680_ (.Y(_00668_),
    .B1(_10879_),
    .B2(net129),
    .A2(net573),
    .A1(_10878_));
 sg13g2_mux2_1 _16681_ (.A0(\top_ihp.oisc.regs[14][3] ),
    .A1(net128),
    .S(net691),
    .X(_00669_));
 sg13g2_mux2_1 _16682_ (.A0(\top_ihp.oisc.regs[14][4] ),
    .A1(net127),
    .S(_10849_),
    .X(_00670_));
 sg13g2_mux2_1 _16683_ (.A0(\top_ihp.oisc.regs[14][5] ),
    .A1(net264),
    .S(net691),
    .X(_00671_));
 sg13g2_mux2_1 _16684_ (.A0(\top_ihp.oisc.regs[14][6] ),
    .A1(net126),
    .S(net691),
    .X(_00672_));
 sg13g2_nand2_1 _16685_ (.Y(_10880_),
    .A(\top_ihp.oisc.regs[14][7] ),
    .B(_10851_));
 sg13g2_o21ai_1 _16686_ (.B1(_10880_),
    .Y(_00673_),
    .A1(net401),
    .A2(_10853_));
 sg13g2_nand2_1 _16687_ (.Y(_10881_),
    .A(\top_ihp.oisc.regs[14][8] ),
    .B(_10851_));
 sg13g2_o21ai_1 _16688_ (.B1(_10881_),
    .Y(_00674_),
    .A1(net266),
    .A2(_10853_));
 sg13g2_mux2_1 _16689_ (.A0(\top_ihp.oisc.regs[14][9] ),
    .A1(net125),
    .S(_10849_),
    .X(_00675_));
 sg13g2_nand2_1 _16690_ (.Y(_10882_),
    .A(_10749_),
    .B(_10787_));
 sg13g2_buf_1 _16691_ (.A(_10882_),
    .X(_10883_));
 sg13g2_buf_2 _16692_ (.A(_10883_),
    .X(_10884_));
 sg13g2_mux2_1 _16693_ (.A0(_09889_),
    .A1(\top_ihp.oisc.regs[15][0] ),
    .S(_10884_),
    .X(_00676_));
 sg13g2_mux2_1 _16694_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[15][10] ),
    .S(_10884_),
    .X(_00677_));
 sg13g2_buf_2 _16695_ (.A(net658),
    .X(_10885_));
 sg13g2_buf_1 _16696_ (.A(net658),
    .X(_10886_));
 sg13g2_nand2_1 _16697_ (.Y(_10887_),
    .A(\top_ihp.oisc.regs[15][11] ),
    .B(net567));
 sg13g2_o21ai_1 _16698_ (.B1(_10887_),
    .Y(_00678_),
    .A1(net62),
    .A2(net568));
 sg13g2_buf_1 _16699_ (.A(_10089_),
    .X(_10888_));
 sg13g2_nand2_1 _16700_ (.Y(_10889_),
    .A(\top_ihp.oisc.regs[15][12] ),
    .B(net567));
 sg13g2_o21ai_1 _16701_ (.B1(_10889_),
    .Y(_00679_),
    .A1(net51),
    .A2(net568));
 sg13g2_nand2_1 _16702_ (.Y(_10890_),
    .A(\top_ihp.oisc.regs[15][13] ),
    .B(net567));
 sg13g2_o21ai_1 _16703_ (.B1(_10890_),
    .Y(_00680_),
    .A1(net278),
    .A2(net568));
 sg13g2_nand2_1 _16704_ (.Y(_10891_),
    .A(\top_ihp.oisc.regs[15][14] ),
    .B(_10886_));
 sg13g2_o21ai_1 _16705_ (.B1(_10891_),
    .Y(_00681_),
    .A1(net277),
    .A2(net568));
 sg13g2_nand2_1 _16706_ (.Y(_10892_),
    .A(\top_ihp.oisc.regs[15][15] ),
    .B(net567));
 sg13g2_o21ai_1 _16707_ (.B1(_10892_),
    .Y(_00682_),
    .A1(net407),
    .A2(net568));
 sg13g2_nand2_1 _16708_ (.Y(_10893_),
    .A(\top_ihp.oisc.regs[15][16] ),
    .B(net567));
 sg13g2_o21ai_1 _16709_ (.B1(_10893_),
    .Y(_00683_),
    .A1(net140),
    .A2(_10885_));
 sg13g2_nand2_1 _16710_ (.Y(_10894_),
    .A(\top_ihp.oisc.regs[15][17] ),
    .B(net567));
 sg13g2_o21ai_1 _16711_ (.B1(_10894_),
    .Y(_00684_),
    .A1(net406),
    .A2(net568));
 sg13g2_nand2_1 _16712_ (.Y(_10895_),
    .A(\top_ihp.oisc.regs[15][18] ),
    .B(_10886_));
 sg13g2_o21ai_1 _16713_ (.B1(_10895_),
    .Y(_00685_),
    .A1(net275),
    .A2(_10885_));
 sg13g2_mux2_1 _16714_ (.A0(_10765_),
    .A1(\top_ihp.oisc.regs[15][19] ),
    .S(net569),
    .X(_00686_));
 sg13g2_buf_1 _16715_ (.A(net658),
    .X(_10896_));
 sg13g2_nand2_1 _16716_ (.Y(_10897_),
    .A(\top_ihp.oisc.regs[15][1] ),
    .B(net566));
 sg13g2_o21ai_1 _16717_ (.B1(_10897_),
    .Y(_00687_),
    .A1(_10834_),
    .A2(net568));
 sg13g2_nand2_1 _16718_ (.Y(_10898_),
    .A(\top_ihp.oisc.regs[15][20] ),
    .B(net566));
 sg13g2_o21ai_1 _16719_ (.B1(_10898_),
    .Y(_00688_),
    .A1(net138),
    .A2(net568));
 sg13g2_buf_1 _16720_ (.A(net658),
    .X(_10899_));
 sg13g2_nand2_1 _16721_ (.Y(_10900_),
    .A(\top_ihp.oisc.regs[15][21] ),
    .B(net566));
 sg13g2_o21ai_1 _16722_ (.B1(_10900_),
    .Y(_00689_),
    .A1(net137),
    .A2(net565));
 sg13g2_nand2_1 _16723_ (.Y(_10901_),
    .A(\top_ihp.oisc.regs[15][22] ),
    .B(net566));
 sg13g2_o21ai_1 _16724_ (.B1(_10901_),
    .Y(_00690_),
    .A1(net272),
    .A2(net565));
 sg13g2_nand2_1 _16725_ (.Y(_10902_),
    .A(\top_ihp.oisc.regs[15][23] ),
    .B(_10896_));
 sg13g2_o21ai_1 _16726_ (.B1(_10902_),
    .Y(_00691_),
    .A1(net271),
    .A2(_10899_));
 sg13g2_mux2_1 _16727_ (.A0(_10416_),
    .A1(\top_ihp.oisc.regs[15][24] ),
    .S(net569),
    .X(_00692_));
 sg13g2_nand2_1 _16728_ (.Y(_10903_),
    .A(\top_ihp.oisc.regs[15][25] ),
    .B(_10896_));
 sg13g2_o21ai_1 _16729_ (.B1(_10903_),
    .Y(_00693_),
    .A1(_10424_),
    .A2(net565));
 sg13g2_nand2_1 _16730_ (.Y(_10904_),
    .A(\top_ihp.oisc.regs[15][26] ),
    .B(net566));
 sg13g2_o21ai_1 _16731_ (.B1(_10904_),
    .Y(_00694_),
    .A1(net402),
    .A2(_10899_));
 sg13g2_mux2_1 _16732_ (.A0(_10776_),
    .A1(\top_ihp.oisc.regs[15][27] ),
    .S(net569),
    .X(_00695_));
 sg13g2_nand2_1 _16733_ (.Y(_10905_),
    .A(\top_ihp.oisc.regs[15][28] ),
    .B(net566));
 sg13g2_o21ai_1 _16734_ (.B1(_10905_),
    .Y(_00696_),
    .A1(_10460_),
    .A2(net565));
 sg13g2_nand2_1 _16735_ (.Y(_10906_),
    .A(\top_ihp.oisc.regs[15][29] ),
    .B(net566));
 sg13g2_o21ai_1 _16736_ (.B1(_10906_),
    .Y(_00697_),
    .A1(net269),
    .A2(net565));
 sg13g2_nand2_1 _16737_ (.Y(_10907_),
    .A(\top_ihp.oisc.regs[15][2] ),
    .B(net566));
 sg13g2_o21ai_1 _16738_ (.B1(_10907_),
    .Y(_00698_),
    .A1(net136),
    .A2(net565));
 sg13g2_nand2_1 _16739_ (.Y(_10908_),
    .A(\top_ihp.oisc.regs[15][30] ),
    .B(net658));
 sg13g2_o21ai_1 _16740_ (.B1(_10908_),
    .Y(_00699_),
    .A1(_10509_),
    .A2(net565));
 sg13g2_nand2_1 _16741_ (.Y(_10909_),
    .A(\top_ihp.oisc.regs[15][31] ),
    .B(net658));
 sg13g2_o21ai_1 _16742_ (.B1(_10909_),
    .Y(_00700_),
    .A1(net268),
    .A2(net565));
 sg13g2_mux2_1 _16743_ (.A0(_10568_),
    .A1(\top_ihp.oisc.regs[15][3] ),
    .S(net569),
    .X(_00701_));
 sg13g2_mux2_1 _16744_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[15][4] ),
    .S(net569),
    .X(_00702_));
 sg13g2_mux2_1 _16745_ (.A0(_10626_),
    .A1(\top_ihp.oisc.regs[15][5] ),
    .S(net569),
    .X(_00703_));
 sg13g2_mux2_1 _16746_ (.A0(_10649_),
    .A1(\top_ihp.oisc.regs[15][6] ),
    .S(net567),
    .X(_00704_));
 sg13g2_nand2_1 _16747_ (.Y(_10910_),
    .A(\top_ihp.oisc.regs[15][7] ),
    .B(net658));
 sg13g2_o21ai_1 _16748_ (.B1(_10910_),
    .Y(_00705_),
    .A1(net401),
    .A2(net569));
 sg13g2_nand2_1 _16749_ (.Y(_10911_),
    .A(\top_ihp.oisc.regs[15][8] ),
    .B(net658));
 sg13g2_o21ai_1 _16750_ (.B1(_10911_),
    .Y(_00706_),
    .A1(net266),
    .A2(net569));
 sg13g2_mux2_1 _16751_ (.A0(_10688_),
    .A1(\top_ihp.oisc.regs[15][9] ),
    .S(net567),
    .X(_00707_));
 sg13g2_buf_1 _16752_ (.A(\top_ihp.oisc.regs[16][0] ),
    .X(_00708_));
 sg13g2_buf_1 _16753_ (.A(\top_ihp.oisc.regs[16][10] ),
    .X(_00709_));
 sg13g2_buf_1 _16754_ (.A(\top_ihp.oisc.regs[16][11] ),
    .X(_00710_));
 sg13g2_buf_1 _16755_ (.A(\top_ihp.oisc.regs[16][12] ),
    .X(_00711_));
 sg13g2_buf_1 _16756_ (.A(\top_ihp.oisc.regs[16][13] ),
    .X(_00712_));
 sg13g2_buf_1 _16757_ (.A(\top_ihp.oisc.regs[16][14] ),
    .X(_00713_));
 sg13g2_buf_1 _16758_ (.A(\top_ihp.oisc.regs[16][15] ),
    .X(_00714_));
 sg13g2_buf_1 _16759_ (.A(\top_ihp.oisc.regs[16][16] ),
    .X(_00715_));
 sg13g2_buf_1 _16760_ (.A(\top_ihp.oisc.regs[16][17] ),
    .X(_00716_));
 sg13g2_buf_1 _16761_ (.A(\top_ihp.oisc.regs[16][18] ),
    .X(_00717_));
 sg13g2_buf_1 _16762_ (.A(\top_ihp.oisc.regs[16][19] ),
    .X(_00718_));
 sg13g2_buf_1 _16763_ (.A(\top_ihp.oisc.regs[16][1] ),
    .X(_00719_));
 sg13g2_buf_1 _16764_ (.A(\top_ihp.oisc.regs[16][20] ),
    .X(_00720_));
 sg13g2_buf_1 _16765_ (.A(\top_ihp.oisc.regs[16][21] ),
    .X(_00721_));
 sg13g2_buf_1 _16766_ (.A(\top_ihp.oisc.regs[16][22] ),
    .X(_00722_));
 sg13g2_buf_1 _16767_ (.A(\top_ihp.oisc.regs[16][23] ),
    .X(_00723_));
 sg13g2_buf_1 _16768_ (.A(\top_ihp.oisc.regs[16][24] ),
    .X(_00724_));
 sg13g2_buf_1 _16769_ (.A(\top_ihp.oisc.regs[16][25] ),
    .X(_00725_));
 sg13g2_buf_1 _16770_ (.A(\top_ihp.oisc.regs[16][26] ),
    .X(_00726_));
 sg13g2_buf_1 _16771_ (.A(\top_ihp.oisc.regs[16][27] ),
    .X(_00727_));
 sg13g2_buf_1 _16772_ (.A(\top_ihp.oisc.regs[16][28] ),
    .X(_00728_));
 sg13g2_buf_1 _16773_ (.A(\top_ihp.oisc.regs[16][29] ),
    .X(_00729_));
 sg13g2_buf_1 _16774_ (.A(\top_ihp.oisc.regs[16][2] ),
    .X(_00730_));
 sg13g2_buf_1 _16775_ (.A(\top_ihp.oisc.regs[16][30] ),
    .X(_00731_));
 sg13g2_buf_1 _16776_ (.A(\top_ihp.oisc.regs[16][31] ),
    .X(_00732_));
 sg13g2_buf_1 _16777_ (.A(\top_ihp.oisc.regs[16][3] ),
    .X(_00733_));
 sg13g2_buf_1 _16778_ (.A(\top_ihp.oisc.regs[16][4] ),
    .X(_00734_));
 sg13g2_buf_1 _16779_ (.A(\top_ihp.oisc.regs[16][5] ),
    .X(_00735_));
 sg13g2_buf_1 _16780_ (.A(\top_ihp.oisc.regs[16][6] ),
    .X(_00736_));
 sg13g2_buf_1 _16781_ (.A(\top_ihp.oisc.regs[16][7] ),
    .X(_00737_));
 sg13g2_buf_1 _16782_ (.A(\top_ihp.oisc.regs[16][8] ),
    .X(_00738_));
 sg13g2_buf_1 _16783_ (.A(\top_ihp.oisc.regs[16][9] ),
    .X(_00739_));
 sg13g2_buf_1 _16784_ (.A(\top_ihp.oisc.regs[17][0] ),
    .X(_00740_));
 sg13g2_buf_1 _16785_ (.A(\top_ihp.oisc.regs[17][10] ),
    .X(_00741_));
 sg13g2_buf_1 _16786_ (.A(\top_ihp.oisc.regs[17][11] ),
    .X(_00742_));
 sg13g2_buf_1 _16787_ (.A(\top_ihp.oisc.regs[17][12] ),
    .X(_00743_));
 sg13g2_buf_1 _16788_ (.A(\top_ihp.oisc.regs[17][13] ),
    .X(_00744_));
 sg13g2_buf_1 _16789_ (.A(\top_ihp.oisc.regs[17][14] ),
    .X(_00745_));
 sg13g2_buf_1 _16790_ (.A(\top_ihp.oisc.regs[17][15] ),
    .X(_00746_));
 sg13g2_buf_1 _16791_ (.A(\top_ihp.oisc.regs[17][16] ),
    .X(_00747_));
 sg13g2_buf_1 _16792_ (.A(\top_ihp.oisc.regs[17][17] ),
    .X(_00748_));
 sg13g2_buf_1 _16793_ (.A(\top_ihp.oisc.regs[17][18] ),
    .X(_00749_));
 sg13g2_buf_1 _16794_ (.A(\top_ihp.oisc.regs[17][19] ),
    .X(_00750_));
 sg13g2_buf_1 _16795_ (.A(\top_ihp.oisc.regs[17][1] ),
    .X(_00751_));
 sg13g2_buf_1 _16796_ (.A(\top_ihp.oisc.regs[17][20] ),
    .X(_00752_));
 sg13g2_buf_1 _16797_ (.A(\top_ihp.oisc.regs[17][21] ),
    .X(_00753_));
 sg13g2_buf_1 _16798_ (.A(\top_ihp.oisc.regs[17][22] ),
    .X(_00754_));
 sg13g2_buf_1 _16799_ (.A(\top_ihp.oisc.regs[17][23] ),
    .X(_00755_));
 sg13g2_buf_1 _16800_ (.A(\top_ihp.oisc.regs[17][24] ),
    .X(_00756_));
 sg13g2_buf_1 _16801_ (.A(\top_ihp.oisc.regs[17][25] ),
    .X(_00757_));
 sg13g2_buf_1 _16802_ (.A(\top_ihp.oisc.regs[17][26] ),
    .X(_00758_));
 sg13g2_buf_1 _16803_ (.A(\top_ihp.oisc.regs[17][27] ),
    .X(_00759_));
 sg13g2_buf_1 _16804_ (.A(\top_ihp.oisc.regs[17][28] ),
    .X(_00760_));
 sg13g2_buf_1 _16805_ (.A(\top_ihp.oisc.regs[17][29] ),
    .X(_00761_));
 sg13g2_buf_1 _16806_ (.A(\top_ihp.oisc.regs[17][2] ),
    .X(_00762_));
 sg13g2_buf_1 _16807_ (.A(\top_ihp.oisc.regs[17][30] ),
    .X(_00763_));
 sg13g2_buf_1 _16808_ (.A(\top_ihp.oisc.regs[17][31] ),
    .X(_00764_));
 sg13g2_buf_1 _16809_ (.A(\top_ihp.oisc.regs[17][3] ),
    .X(_00765_));
 sg13g2_buf_1 _16810_ (.A(\top_ihp.oisc.regs[17][4] ),
    .X(_00766_));
 sg13g2_buf_1 _16811_ (.A(\top_ihp.oisc.regs[17][5] ),
    .X(_00767_));
 sg13g2_buf_1 _16812_ (.A(\top_ihp.oisc.regs[17][6] ),
    .X(_00768_));
 sg13g2_buf_1 _16813_ (.A(\top_ihp.oisc.regs[17][7] ),
    .X(_00769_));
 sg13g2_buf_1 _16814_ (.A(\top_ihp.oisc.regs[17][8] ),
    .X(_00770_));
 sg13g2_buf_1 _16815_ (.A(\top_ihp.oisc.regs[17][9] ),
    .X(_00771_));
 sg13g2_buf_1 _16816_ (.A(\top_ihp.oisc.regs[18][0] ),
    .X(_00772_));
 sg13g2_buf_1 _16817_ (.A(\top_ihp.oisc.regs[18][10] ),
    .X(_00773_));
 sg13g2_buf_1 _16818_ (.A(\top_ihp.oisc.regs[18][11] ),
    .X(_00774_));
 sg13g2_buf_1 _16819_ (.A(\top_ihp.oisc.regs[18][12] ),
    .X(_00775_));
 sg13g2_buf_1 _16820_ (.A(\top_ihp.oisc.regs[18][13] ),
    .X(_00776_));
 sg13g2_buf_1 _16821_ (.A(\top_ihp.oisc.regs[18][14] ),
    .X(_00777_));
 sg13g2_buf_1 _16822_ (.A(\top_ihp.oisc.regs[18][15] ),
    .X(_00778_));
 sg13g2_buf_1 _16823_ (.A(\top_ihp.oisc.regs[18][16] ),
    .X(_00779_));
 sg13g2_buf_1 _16824_ (.A(\top_ihp.oisc.regs[18][17] ),
    .X(_00780_));
 sg13g2_buf_1 _16825_ (.A(\top_ihp.oisc.regs[18][18] ),
    .X(_00781_));
 sg13g2_buf_1 _16826_ (.A(\top_ihp.oisc.regs[18][19] ),
    .X(_00782_));
 sg13g2_buf_1 _16827_ (.A(\top_ihp.oisc.regs[18][1] ),
    .X(_00783_));
 sg13g2_buf_1 _16828_ (.A(\top_ihp.oisc.regs[18][20] ),
    .X(_00784_));
 sg13g2_buf_1 _16829_ (.A(\top_ihp.oisc.regs[18][21] ),
    .X(_00785_));
 sg13g2_buf_1 _16830_ (.A(\top_ihp.oisc.regs[18][22] ),
    .X(_00786_));
 sg13g2_buf_1 _16831_ (.A(\top_ihp.oisc.regs[18][23] ),
    .X(_00787_));
 sg13g2_buf_1 _16832_ (.A(\top_ihp.oisc.regs[18][24] ),
    .X(_00788_));
 sg13g2_buf_1 _16833_ (.A(\top_ihp.oisc.regs[18][25] ),
    .X(_00789_));
 sg13g2_buf_1 _16834_ (.A(\top_ihp.oisc.regs[18][26] ),
    .X(_00790_));
 sg13g2_buf_1 _16835_ (.A(\top_ihp.oisc.regs[18][27] ),
    .X(_00791_));
 sg13g2_buf_1 _16836_ (.A(\top_ihp.oisc.regs[18][28] ),
    .X(_00792_));
 sg13g2_buf_1 _16837_ (.A(\top_ihp.oisc.regs[18][29] ),
    .X(_00793_));
 sg13g2_buf_1 _16838_ (.A(\top_ihp.oisc.regs[18][2] ),
    .X(_00794_));
 sg13g2_buf_1 _16839_ (.A(\top_ihp.oisc.regs[18][30] ),
    .X(_00795_));
 sg13g2_buf_1 _16840_ (.A(\top_ihp.oisc.regs[18][31] ),
    .X(_00796_));
 sg13g2_buf_1 _16841_ (.A(\top_ihp.oisc.regs[18][3] ),
    .X(_00797_));
 sg13g2_buf_1 _16842_ (.A(\top_ihp.oisc.regs[18][4] ),
    .X(_00798_));
 sg13g2_buf_1 _16843_ (.A(\top_ihp.oisc.regs[18][5] ),
    .X(_00799_));
 sg13g2_buf_1 _16844_ (.A(\top_ihp.oisc.regs[18][6] ),
    .X(_00800_));
 sg13g2_buf_1 _16845_ (.A(\top_ihp.oisc.regs[18][7] ),
    .X(_00801_));
 sg13g2_buf_1 _16846_ (.A(\top_ihp.oisc.regs[18][8] ),
    .X(_00802_));
 sg13g2_buf_1 _16847_ (.A(\top_ihp.oisc.regs[18][9] ),
    .X(_00803_));
 sg13g2_buf_1 _16848_ (.A(\top_ihp.oisc.regs[19][0] ),
    .X(_00804_));
 sg13g2_buf_1 _16849_ (.A(\top_ihp.oisc.regs[19][10] ),
    .X(_00805_));
 sg13g2_buf_1 _16850_ (.A(\top_ihp.oisc.regs[19][11] ),
    .X(_00806_));
 sg13g2_buf_1 _16851_ (.A(\top_ihp.oisc.regs[19][12] ),
    .X(_00807_));
 sg13g2_buf_1 _16852_ (.A(\top_ihp.oisc.regs[19][13] ),
    .X(_00808_));
 sg13g2_buf_1 _16853_ (.A(\top_ihp.oisc.regs[19][14] ),
    .X(_00809_));
 sg13g2_buf_1 _16854_ (.A(\top_ihp.oisc.regs[19][15] ),
    .X(_00810_));
 sg13g2_buf_1 _16855_ (.A(\top_ihp.oisc.regs[19][16] ),
    .X(_00811_));
 sg13g2_buf_1 _16856_ (.A(\top_ihp.oisc.regs[19][17] ),
    .X(_00812_));
 sg13g2_buf_1 _16857_ (.A(\top_ihp.oisc.regs[19][18] ),
    .X(_00813_));
 sg13g2_buf_1 _16858_ (.A(\top_ihp.oisc.regs[19][19] ),
    .X(_00814_));
 sg13g2_buf_1 _16859_ (.A(\top_ihp.oisc.regs[19][1] ),
    .X(_00815_));
 sg13g2_buf_1 _16860_ (.A(\top_ihp.oisc.regs[19][20] ),
    .X(_00816_));
 sg13g2_buf_1 _16861_ (.A(\top_ihp.oisc.regs[19][21] ),
    .X(_00817_));
 sg13g2_buf_1 _16862_ (.A(\top_ihp.oisc.regs[19][22] ),
    .X(_00818_));
 sg13g2_buf_1 _16863_ (.A(\top_ihp.oisc.regs[19][23] ),
    .X(_00819_));
 sg13g2_buf_1 _16864_ (.A(\top_ihp.oisc.regs[19][24] ),
    .X(_00820_));
 sg13g2_buf_1 _16865_ (.A(\top_ihp.oisc.regs[19][25] ),
    .X(_00821_));
 sg13g2_buf_1 _16866_ (.A(\top_ihp.oisc.regs[19][26] ),
    .X(_00822_));
 sg13g2_buf_1 _16867_ (.A(\top_ihp.oisc.regs[19][27] ),
    .X(_00823_));
 sg13g2_buf_1 _16868_ (.A(\top_ihp.oisc.regs[19][28] ),
    .X(_00824_));
 sg13g2_buf_1 _16869_ (.A(\top_ihp.oisc.regs[19][29] ),
    .X(_00825_));
 sg13g2_buf_1 _16870_ (.A(\top_ihp.oisc.regs[19][2] ),
    .X(_00826_));
 sg13g2_buf_1 _16871_ (.A(\top_ihp.oisc.regs[19][30] ),
    .X(_00827_));
 sg13g2_buf_1 _16872_ (.A(\top_ihp.oisc.regs[19][31] ),
    .X(_00828_));
 sg13g2_buf_1 _16873_ (.A(\top_ihp.oisc.regs[19][3] ),
    .X(_00829_));
 sg13g2_buf_1 _16874_ (.A(\top_ihp.oisc.regs[19][4] ),
    .X(_00830_));
 sg13g2_buf_1 _16875_ (.A(\top_ihp.oisc.regs[19][5] ),
    .X(_00831_));
 sg13g2_buf_1 _16876_ (.A(\top_ihp.oisc.regs[19][6] ),
    .X(_00832_));
 sg13g2_buf_1 _16877_ (.A(\top_ihp.oisc.regs[19][7] ),
    .X(_00833_));
 sg13g2_buf_1 _16878_ (.A(\top_ihp.oisc.regs[19][8] ),
    .X(_00834_));
 sg13g2_buf_1 _16879_ (.A(\top_ihp.oisc.regs[19][9] ),
    .X(_00835_));
 sg13g2_nor2_2 _16880_ (.A(_10692_),
    .B(_09912_),
    .Y(_10912_));
 sg13g2_nand2_1 _16881_ (.Y(_10913_),
    .A(_09929_),
    .B(_10822_));
 sg13g2_nor2_1 _16882_ (.A(_10912_),
    .B(_10913_),
    .Y(_10914_));
 sg13g2_buf_2 _16883_ (.A(_10914_),
    .X(_10915_));
 sg13g2_buf_1 _16884_ (.A(_10915_),
    .X(_10916_));
 sg13g2_mux2_1 _16885_ (.A0(\top_ihp.oisc.regs[1][0] ),
    .A1(net119),
    .S(net564),
    .X(_00836_));
 sg13g2_mux2_1 _16886_ (.A0(\top_ihp.oisc.regs[1][10] ),
    .A1(net130),
    .S(net564),
    .X(_00837_));
 sg13g2_buf_1 _16887_ (.A(_10050_),
    .X(_10917_));
 sg13g2_nor2_1 _16888_ (.A(\top_ihp.oisc.regs[1][11] ),
    .B(_10915_),
    .Y(_10918_));
 sg13g2_a21oi_1 _16889_ (.A1(_10917_),
    .A2(_10916_),
    .Y(_00838_),
    .B1(_10918_));
 sg13g2_nand2_1 _16890_ (.Y(_10919_),
    .A(net692),
    .B(_10824_));
 sg13g2_buf_1 _16891_ (.A(_10919_),
    .X(_10920_));
 sg13g2_buf_1 _16892_ (.A(net563),
    .X(_10921_));
 sg13g2_buf_1 _16893_ (.A(net563),
    .X(_10922_));
 sg13g2_nand2_1 _16894_ (.Y(_10923_),
    .A(\top_ihp.oisc.regs[1][12] ),
    .B(net394));
 sg13g2_o21ai_1 _16895_ (.B1(_10923_),
    .Y(_00839_),
    .A1(_10888_),
    .A2(net395));
 sg13g2_nand2_1 _16896_ (.Y(_10924_),
    .A(\top_ihp.oisc.regs[1][13] ),
    .B(net394));
 sg13g2_o21ai_1 _16897_ (.B1(_10924_),
    .Y(_00840_),
    .A1(_10122_),
    .A2(net395));
 sg13g2_buf_1 _16898_ (.A(net563),
    .X(_10925_));
 sg13g2_nand2_1 _16899_ (.Y(_10926_),
    .A(\top_ihp.oisc.regs[1][14] ),
    .B(net393));
 sg13g2_o21ai_1 _16900_ (.B1(_10926_),
    .Y(_00841_),
    .A1(_10159_),
    .A2(net395));
 sg13g2_nand2_1 _16901_ (.Y(_10927_),
    .A(\top_ihp.oisc.regs[1][15] ),
    .B(net393));
 sg13g2_o21ai_1 _16902_ (.B1(_10927_),
    .Y(_00842_),
    .A1(_10171_),
    .A2(net395));
 sg13g2_nand2_1 _16903_ (.Y(_10928_),
    .A(\top_ihp.oisc.regs[1][16] ),
    .B(net393));
 sg13g2_o21ai_1 _16904_ (.B1(_10928_),
    .Y(_00843_),
    .A1(_10206_),
    .A2(net395));
 sg13g2_nand2_1 _16905_ (.Y(_10929_),
    .A(\top_ihp.oisc.regs[1][17] ),
    .B(net393));
 sg13g2_o21ai_1 _16906_ (.B1(_10929_),
    .Y(_00844_),
    .A1(_10224_),
    .A2(net395));
 sg13g2_nand2_1 _16907_ (.Y(_10930_),
    .A(\top_ihp.oisc.regs[1][18] ),
    .B(net393));
 sg13g2_o21ai_1 _16908_ (.B1(_10930_),
    .Y(_00845_),
    .A1(_10246_),
    .A2(net395));
 sg13g2_buf_2 _16909_ (.A(_10271_),
    .X(_10931_));
 sg13g2_mux2_1 _16910_ (.A0(\top_ihp.oisc.regs[1][19] ),
    .A1(_10931_),
    .S(net564),
    .X(_00846_));
 sg13g2_buf_1 _16911_ (.A(_10318_),
    .X(_10932_));
 sg13g2_nor2_1 _16912_ (.A(\top_ihp.oisc.regs[1][1] ),
    .B(_10915_),
    .Y(_10933_));
 sg13g2_a21oi_1 _16913_ (.A1(net118),
    .A2(net564),
    .Y(_00847_),
    .B1(_10933_));
 sg13g2_nand2_1 _16914_ (.Y(_10934_),
    .A(\top_ihp.oisc.regs[1][20] ),
    .B(net393));
 sg13g2_o21ai_1 _16915_ (.B1(_10934_),
    .Y(_00848_),
    .A1(_10343_),
    .A2(_10921_));
 sg13g2_nand2_1 _16916_ (.Y(_10935_),
    .A(\top_ihp.oisc.regs[1][21] ),
    .B(net393));
 sg13g2_o21ai_1 _16917_ (.B1(_10935_),
    .Y(_00849_),
    .A1(_10362_),
    .A2(net395));
 sg13g2_nand2_1 _16918_ (.Y(_10936_),
    .A(\top_ihp.oisc.regs[1][22] ),
    .B(_10925_));
 sg13g2_o21ai_1 _16919_ (.B1(_10936_),
    .Y(_00850_),
    .A1(_10380_),
    .A2(_10921_));
 sg13g2_nand2_1 _16920_ (.Y(_10937_),
    .A(\top_ihp.oisc.regs[1][23] ),
    .B(_10925_));
 sg13g2_o21ai_1 _16921_ (.B1(_10937_),
    .Y(_00851_),
    .A1(_10393_),
    .A2(_10922_));
 sg13g2_mux2_1 _16922_ (.A0(\top_ihp.oisc.regs[1][24] ),
    .A1(net400),
    .S(net564),
    .X(_00852_));
 sg13g2_nand2_1 _16923_ (.Y(_10938_),
    .A(\top_ihp.oisc.regs[1][25] ),
    .B(net393));
 sg13g2_o21ai_1 _16924_ (.B1(_10938_),
    .Y(_00853_),
    .A1(_10773_),
    .A2(net394));
 sg13g2_nand2_1 _16925_ (.Y(_10939_),
    .A(\top_ihp.oisc.regs[1][26] ),
    .B(net563));
 sg13g2_o21ai_1 _16926_ (.B1(_10939_),
    .Y(_00854_),
    .A1(_10441_),
    .A2(net394));
 sg13g2_buf_1 _16927_ (.A(_10447_),
    .X(_10940_));
 sg13g2_mux2_1 _16928_ (.A0(\top_ihp.oisc.regs[1][27] ),
    .A1(net117),
    .S(net564),
    .X(_00855_));
 sg13g2_buf_1 _16929_ (.A(_10456_),
    .X(_10941_));
 sg13g2_nor2_1 _16930_ (.A(\top_ihp.oisc.regs[1][28] ),
    .B(_10915_),
    .Y(_10942_));
 sg13g2_a21oi_1 _16931_ (.A1(net116),
    .A2(_10916_),
    .Y(_00856_),
    .B1(_10942_));
 sg13g2_nand2_1 _16932_ (.Y(_10943_),
    .A(\top_ihp.oisc.regs[1][29] ),
    .B(net563));
 sg13g2_o21ai_1 _16933_ (.B1(_10943_),
    .Y(_00857_),
    .A1(_10467_),
    .A2(_10922_));
 sg13g2_nand2_1 _16934_ (.Y(_10944_),
    .A(\top_ihp.oisc.regs[1][2] ),
    .B(net563));
 sg13g2_o21ai_1 _16935_ (.B1(_10944_),
    .Y(_00858_),
    .A1(_10500_),
    .A2(net394));
 sg13g2_mux2_1 _16936_ (.A0(_00335_),
    .A1(net53),
    .S(net564),
    .X(_00859_));
 sg13g2_nand2_1 _16937_ (.Y(_10945_),
    .A(\top_ihp.oisc.regs[1][31] ),
    .B(net563));
 sg13g2_o21ai_1 _16938_ (.B1(_10945_),
    .Y(_00860_),
    .A1(net268),
    .A2(net394));
 sg13g2_mux2_1 _16939_ (.A0(\top_ihp.oisc.regs[1][3] ),
    .A1(net128),
    .S(net564),
    .X(_00861_));
 sg13g2_mux2_1 _16940_ (.A0(\top_ihp.oisc.regs[1][4] ),
    .A1(net127),
    .S(_10915_),
    .X(_00862_));
 sg13g2_mux2_1 _16941_ (.A0(\top_ihp.oisc.regs[1][5] ),
    .A1(net264),
    .S(_10915_),
    .X(_00863_));
 sg13g2_mux2_1 _16942_ (.A0(\top_ihp.oisc.regs[1][6] ),
    .A1(net126),
    .S(_10915_),
    .X(_00864_));
 sg13g2_nand2_1 _16943_ (.Y(_10946_),
    .A(\top_ihp.oisc.regs[1][7] ),
    .B(net563));
 sg13g2_o21ai_1 _16944_ (.B1(_10946_),
    .Y(_00865_),
    .A1(_10662_),
    .A2(net394));
 sg13g2_nand2_1 _16945_ (.Y(_10947_),
    .A(\top_ihp.oisc.regs[1][8] ),
    .B(_10920_));
 sg13g2_o21ai_1 _16946_ (.B1(_10947_),
    .Y(_00866_),
    .A1(_10674_),
    .A2(net394));
 sg13g2_mux2_1 _16947_ (.A0(\top_ihp.oisc.regs[1][9] ),
    .A1(net125),
    .S(_10915_),
    .X(_00867_));
 sg13g2_buf_1 _16948_ (.A(\top_ihp.oisc.regs[20][0] ),
    .X(_00868_));
 sg13g2_buf_1 _16949_ (.A(\top_ihp.oisc.regs[20][10] ),
    .X(_00869_));
 sg13g2_buf_1 _16950_ (.A(\top_ihp.oisc.regs[20][11] ),
    .X(_00870_));
 sg13g2_buf_1 _16951_ (.A(\top_ihp.oisc.regs[20][12] ),
    .X(_00871_));
 sg13g2_buf_1 _16952_ (.A(\top_ihp.oisc.regs[20][13] ),
    .X(_00872_));
 sg13g2_buf_1 _16953_ (.A(\top_ihp.oisc.regs[20][14] ),
    .X(_00873_));
 sg13g2_buf_1 _16954_ (.A(\top_ihp.oisc.regs[20][15] ),
    .X(_00874_));
 sg13g2_buf_1 _16955_ (.A(\top_ihp.oisc.regs[20][16] ),
    .X(_00875_));
 sg13g2_buf_1 _16956_ (.A(\top_ihp.oisc.regs[20][17] ),
    .X(_00876_));
 sg13g2_buf_1 _16957_ (.A(\top_ihp.oisc.regs[20][18] ),
    .X(_00877_));
 sg13g2_buf_1 _16958_ (.A(\top_ihp.oisc.regs[20][19] ),
    .X(_00878_));
 sg13g2_buf_1 _16959_ (.A(\top_ihp.oisc.regs[20][1] ),
    .X(_00879_));
 sg13g2_buf_1 _16960_ (.A(\top_ihp.oisc.regs[20][20] ),
    .X(_00880_));
 sg13g2_buf_1 _16961_ (.A(\top_ihp.oisc.regs[20][21] ),
    .X(_00881_));
 sg13g2_buf_1 _16962_ (.A(\top_ihp.oisc.regs[20][22] ),
    .X(_00882_));
 sg13g2_buf_1 _16963_ (.A(\top_ihp.oisc.regs[20][23] ),
    .X(_00883_));
 sg13g2_buf_1 _16964_ (.A(\top_ihp.oisc.regs[20][24] ),
    .X(_00884_));
 sg13g2_buf_1 _16965_ (.A(\top_ihp.oisc.regs[20][25] ),
    .X(_00885_));
 sg13g2_buf_1 _16966_ (.A(\top_ihp.oisc.regs[20][26] ),
    .X(_00886_));
 sg13g2_buf_1 _16967_ (.A(\top_ihp.oisc.regs[20][27] ),
    .X(_00887_));
 sg13g2_buf_1 _16968_ (.A(\top_ihp.oisc.regs[20][28] ),
    .X(_00888_));
 sg13g2_buf_1 _16969_ (.A(\top_ihp.oisc.regs[20][29] ),
    .X(_00889_));
 sg13g2_buf_1 _16970_ (.A(\top_ihp.oisc.regs[20][2] ),
    .X(_00890_));
 sg13g2_buf_1 _16971_ (.A(\top_ihp.oisc.regs[20][30] ),
    .X(_00891_));
 sg13g2_buf_1 _16972_ (.A(\top_ihp.oisc.regs[20][31] ),
    .X(_00892_));
 sg13g2_buf_1 _16973_ (.A(\top_ihp.oisc.regs[20][3] ),
    .X(_00893_));
 sg13g2_buf_1 _16974_ (.A(\top_ihp.oisc.regs[20][4] ),
    .X(_00894_));
 sg13g2_buf_1 _16975_ (.A(\top_ihp.oisc.regs[20][5] ),
    .X(_00895_));
 sg13g2_buf_1 _16976_ (.A(\top_ihp.oisc.regs[20][6] ),
    .X(_00896_));
 sg13g2_buf_1 _16977_ (.A(\top_ihp.oisc.regs[20][7] ),
    .X(_00897_));
 sg13g2_buf_1 _16978_ (.A(\top_ihp.oisc.regs[20][8] ),
    .X(_00898_));
 sg13g2_buf_1 _16979_ (.A(\top_ihp.oisc.regs[20][9] ),
    .X(_00899_));
 sg13g2_buf_1 _16980_ (.A(\top_ihp.oisc.regs[21][0] ),
    .X(_00900_));
 sg13g2_buf_1 _16981_ (.A(\top_ihp.oisc.regs[21][10] ),
    .X(_00901_));
 sg13g2_buf_1 _16982_ (.A(\top_ihp.oisc.regs[21][11] ),
    .X(_00902_));
 sg13g2_buf_1 _16983_ (.A(\top_ihp.oisc.regs[21][12] ),
    .X(_00903_));
 sg13g2_buf_1 _16984_ (.A(\top_ihp.oisc.regs[21][13] ),
    .X(_00904_));
 sg13g2_buf_1 _16985_ (.A(\top_ihp.oisc.regs[21][14] ),
    .X(_00905_));
 sg13g2_buf_1 _16986_ (.A(\top_ihp.oisc.regs[21][15] ),
    .X(_00906_));
 sg13g2_buf_1 _16987_ (.A(\top_ihp.oisc.regs[21][16] ),
    .X(_00907_));
 sg13g2_buf_1 _16988_ (.A(\top_ihp.oisc.regs[21][17] ),
    .X(_00908_));
 sg13g2_buf_1 _16989_ (.A(\top_ihp.oisc.regs[21][18] ),
    .X(_00909_));
 sg13g2_buf_1 _16990_ (.A(\top_ihp.oisc.regs[21][19] ),
    .X(_00910_));
 sg13g2_buf_1 _16991_ (.A(\top_ihp.oisc.regs[21][1] ),
    .X(_00911_));
 sg13g2_buf_1 _16992_ (.A(\top_ihp.oisc.regs[21][20] ),
    .X(_00912_));
 sg13g2_buf_1 _16993_ (.A(\top_ihp.oisc.regs[21][21] ),
    .X(_00913_));
 sg13g2_buf_1 _16994_ (.A(\top_ihp.oisc.regs[21][22] ),
    .X(_00914_));
 sg13g2_buf_1 _16995_ (.A(\top_ihp.oisc.regs[21][23] ),
    .X(_00915_));
 sg13g2_buf_1 _16996_ (.A(\top_ihp.oisc.regs[21][24] ),
    .X(_00916_));
 sg13g2_buf_1 _16997_ (.A(\top_ihp.oisc.regs[21][25] ),
    .X(_00917_));
 sg13g2_buf_1 _16998_ (.A(\top_ihp.oisc.regs[21][26] ),
    .X(_00918_));
 sg13g2_buf_1 _16999_ (.A(\top_ihp.oisc.regs[21][27] ),
    .X(_00919_));
 sg13g2_buf_1 _17000_ (.A(\top_ihp.oisc.regs[21][28] ),
    .X(_00920_));
 sg13g2_buf_1 _17001_ (.A(\top_ihp.oisc.regs[21][29] ),
    .X(_00921_));
 sg13g2_buf_1 _17002_ (.A(\top_ihp.oisc.regs[21][2] ),
    .X(_00922_));
 sg13g2_buf_1 _17003_ (.A(\top_ihp.oisc.regs[21][30] ),
    .X(_00923_));
 sg13g2_buf_1 _17004_ (.A(\top_ihp.oisc.regs[21][31] ),
    .X(_00924_));
 sg13g2_buf_1 _17005_ (.A(\top_ihp.oisc.regs[21][3] ),
    .X(_00925_));
 sg13g2_buf_1 _17006_ (.A(\top_ihp.oisc.regs[21][4] ),
    .X(_00926_));
 sg13g2_buf_1 _17007_ (.A(\top_ihp.oisc.regs[21][5] ),
    .X(_00927_));
 sg13g2_buf_1 _17008_ (.A(\top_ihp.oisc.regs[21][6] ),
    .X(_00928_));
 sg13g2_buf_1 _17009_ (.A(\top_ihp.oisc.regs[21][7] ),
    .X(_00929_));
 sg13g2_buf_1 _17010_ (.A(\top_ihp.oisc.regs[21][8] ),
    .X(_00930_));
 sg13g2_buf_1 _17011_ (.A(\top_ihp.oisc.regs[21][9] ),
    .X(_00931_));
 sg13g2_buf_1 _17012_ (.A(\top_ihp.oisc.regs[22][0] ),
    .X(_00932_));
 sg13g2_buf_1 _17013_ (.A(\top_ihp.oisc.regs[22][10] ),
    .X(_00933_));
 sg13g2_buf_1 _17014_ (.A(\top_ihp.oisc.regs[22][11] ),
    .X(_00934_));
 sg13g2_buf_1 _17015_ (.A(\top_ihp.oisc.regs[22][12] ),
    .X(_00935_));
 sg13g2_buf_1 _17016_ (.A(\top_ihp.oisc.regs[22][13] ),
    .X(_00936_));
 sg13g2_buf_1 _17017_ (.A(\top_ihp.oisc.regs[22][14] ),
    .X(_00937_));
 sg13g2_buf_1 _17018_ (.A(\top_ihp.oisc.regs[22][15] ),
    .X(_00938_));
 sg13g2_buf_1 _17019_ (.A(\top_ihp.oisc.regs[22][16] ),
    .X(_00939_));
 sg13g2_buf_1 _17020_ (.A(\top_ihp.oisc.regs[22][17] ),
    .X(_00940_));
 sg13g2_buf_1 _17021_ (.A(\top_ihp.oisc.regs[22][18] ),
    .X(_00941_));
 sg13g2_buf_1 _17022_ (.A(\top_ihp.oisc.regs[22][19] ),
    .X(_00942_));
 sg13g2_buf_1 _17023_ (.A(\top_ihp.oisc.regs[22][1] ),
    .X(_00943_));
 sg13g2_buf_1 _17024_ (.A(\top_ihp.oisc.regs[22][20] ),
    .X(_00944_));
 sg13g2_buf_1 _17025_ (.A(\top_ihp.oisc.regs[22][21] ),
    .X(_00945_));
 sg13g2_buf_1 _17026_ (.A(\top_ihp.oisc.regs[22][22] ),
    .X(_00946_));
 sg13g2_buf_1 _17027_ (.A(\top_ihp.oisc.regs[22][23] ),
    .X(_00947_));
 sg13g2_buf_1 _17028_ (.A(\top_ihp.oisc.regs[22][24] ),
    .X(_00948_));
 sg13g2_buf_1 _17029_ (.A(\top_ihp.oisc.regs[22][25] ),
    .X(_00949_));
 sg13g2_buf_1 _17030_ (.A(\top_ihp.oisc.regs[22][26] ),
    .X(_00950_));
 sg13g2_buf_1 _17031_ (.A(\top_ihp.oisc.regs[22][27] ),
    .X(_00951_));
 sg13g2_buf_1 _17032_ (.A(\top_ihp.oisc.regs[22][28] ),
    .X(_00952_));
 sg13g2_buf_1 _17033_ (.A(\top_ihp.oisc.regs[22][29] ),
    .X(_00953_));
 sg13g2_buf_1 _17034_ (.A(\top_ihp.oisc.regs[22][2] ),
    .X(_00954_));
 sg13g2_buf_1 _17035_ (.A(\top_ihp.oisc.regs[22][30] ),
    .X(_00955_));
 sg13g2_buf_1 _17036_ (.A(\top_ihp.oisc.regs[22][31] ),
    .X(_00956_));
 sg13g2_buf_1 _17037_ (.A(\top_ihp.oisc.regs[22][3] ),
    .X(_00957_));
 sg13g2_buf_1 _17038_ (.A(\top_ihp.oisc.regs[22][4] ),
    .X(_00958_));
 sg13g2_buf_1 _17039_ (.A(\top_ihp.oisc.regs[22][5] ),
    .X(_00959_));
 sg13g2_buf_1 _17040_ (.A(\top_ihp.oisc.regs[22][6] ),
    .X(_00960_));
 sg13g2_buf_1 _17041_ (.A(\top_ihp.oisc.regs[22][7] ),
    .X(_00961_));
 sg13g2_buf_1 _17042_ (.A(\top_ihp.oisc.regs[22][8] ),
    .X(_00962_));
 sg13g2_buf_1 _17043_ (.A(\top_ihp.oisc.regs[22][9] ),
    .X(_00963_));
 sg13g2_buf_1 _17044_ (.A(\top_ihp.oisc.regs[23][0] ),
    .X(_00964_));
 sg13g2_buf_1 _17045_ (.A(\top_ihp.oisc.regs[23][10] ),
    .X(_00965_));
 sg13g2_buf_1 _17046_ (.A(\top_ihp.oisc.regs[23][11] ),
    .X(_00966_));
 sg13g2_buf_1 _17047_ (.A(\top_ihp.oisc.regs[23][12] ),
    .X(_00967_));
 sg13g2_buf_1 _17048_ (.A(\top_ihp.oisc.regs[23][13] ),
    .X(_00968_));
 sg13g2_buf_1 _17049_ (.A(\top_ihp.oisc.regs[23][14] ),
    .X(_00969_));
 sg13g2_buf_1 _17050_ (.A(\top_ihp.oisc.regs[23][15] ),
    .X(_00970_));
 sg13g2_buf_1 _17051_ (.A(\top_ihp.oisc.regs[23][16] ),
    .X(_00971_));
 sg13g2_buf_1 _17052_ (.A(\top_ihp.oisc.regs[23][17] ),
    .X(_00972_));
 sg13g2_buf_1 _17053_ (.A(\top_ihp.oisc.regs[23][18] ),
    .X(_00973_));
 sg13g2_buf_1 _17054_ (.A(\top_ihp.oisc.regs[23][19] ),
    .X(_00974_));
 sg13g2_buf_1 _17055_ (.A(\top_ihp.oisc.regs[23][1] ),
    .X(_00975_));
 sg13g2_buf_1 _17056_ (.A(\top_ihp.oisc.regs[23][20] ),
    .X(_00976_));
 sg13g2_buf_1 _17057_ (.A(\top_ihp.oisc.regs[23][21] ),
    .X(_00977_));
 sg13g2_buf_1 _17058_ (.A(\top_ihp.oisc.regs[23][22] ),
    .X(_00978_));
 sg13g2_buf_1 _17059_ (.A(\top_ihp.oisc.regs[23][23] ),
    .X(_00979_));
 sg13g2_buf_1 _17060_ (.A(\top_ihp.oisc.regs[23][24] ),
    .X(_00980_));
 sg13g2_buf_1 _17061_ (.A(\top_ihp.oisc.regs[23][25] ),
    .X(_00981_));
 sg13g2_buf_1 _17062_ (.A(\top_ihp.oisc.regs[23][26] ),
    .X(_00982_));
 sg13g2_buf_1 _17063_ (.A(\top_ihp.oisc.regs[23][27] ),
    .X(_00983_));
 sg13g2_buf_1 _17064_ (.A(\top_ihp.oisc.regs[23][28] ),
    .X(_00984_));
 sg13g2_buf_1 _17065_ (.A(\top_ihp.oisc.regs[23][29] ),
    .X(_00985_));
 sg13g2_buf_1 _17066_ (.A(\top_ihp.oisc.regs[23][2] ),
    .X(_00986_));
 sg13g2_buf_1 _17067_ (.A(\top_ihp.oisc.regs[23][30] ),
    .X(_00987_));
 sg13g2_buf_1 _17068_ (.A(\top_ihp.oisc.regs[23][31] ),
    .X(_00988_));
 sg13g2_buf_1 _17069_ (.A(\top_ihp.oisc.regs[23][3] ),
    .X(_00989_));
 sg13g2_buf_1 _17070_ (.A(\top_ihp.oisc.regs[23][4] ),
    .X(_00990_));
 sg13g2_buf_1 _17071_ (.A(\top_ihp.oisc.regs[23][5] ),
    .X(_00991_));
 sg13g2_buf_1 _17072_ (.A(\top_ihp.oisc.regs[23][6] ),
    .X(_00992_));
 sg13g2_buf_1 _17073_ (.A(\top_ihp.oisc.regs[23][7] ),
    .X(_00993_));
 sg13g2_buf_1 _17074_ (.A(\top_ihp.oisc.regs[23][8] ),
    .X(_00994_));
 sg13g2_buf_1 _17075_ (.A(\top_ihp.oisc.regs[23][9] ),
    .X(_00995_));
 sg13g2_buf_1 _17076_ (.A(\top_ihp.oisc.regs[24][0] ),
    .X(_00996_));
 sg13g2_buf_1 _17077_ (.A(\top_ihp.oisc.regs[24][10] ),
    .X(_00997_));
 sg13g2_buf_1 _17078_ (.A(\top_ihp.oisc.regs[24][11] ),
    .X(_00998_));
 sg13g2_buf_1 _17079_ (.A(\top_ihp.oisc.regs[24][12] ),
    .X(_00999_));
 sg13g2_buf_1 _17080_ (.A(\top_ihp.oisc.regs[24][13] ),
    .X(_01000_));
 sg13g2_buf_1 _17081_ (.A(\top_ihp.oisc.regs[24][14] ),
    .X(_01001_));
 sg13g2_buf_1 _17082_ (.A(\top_ihp.oisc.regs[24][15] ),
    .X(_01002_));
 sg13g2_buf_1 _17083_ (.A(\top_ihp.oisc.regs[24][16] ),
    .X(_01003_));
 sg13g2_buf_1 _17084_ (.A(\top_ihp.oisc.regs[24][17] ),
    .X(_01004_));
 sg13g2_buf_1 _17085_ (.A(\top_ihp.oisc.regs[24][18] ),
    .X(_01005_));
 sg13g2_buf_1 _17086_ (.A(\top_ihp.oisc.regs[24][19] ),
    .X(_01006_));
 sg13g2_buf_1 _17087_ (.A(\top_ihp.oisc.regs[24][1] ),
    .X(_01007_));
 sg13g2_buf_1 _17088_ (.A(\top_ihp.oisc.regs[24][20] ),
    .X(_01008_));
 sg13g2_buf_1 _17089_ (.A(\top_ihp.oisc.regs[24][21] ),
    .X(_01009_));
 sg13g2_buf_1 _17090_ (.A(\top_ihp.oisc.regs[24][22] ),
    .X(_01010_));
 sg13g2_buf_1 _17091_ (.A(\top_ihp.oisc.regs[24][23] ),
    .X(_01011_));
 sg13g2_buf_1 _17092_ (.A(\top_ihp.oisc.regs[24][24] ),
    .X(_01012_));
 sg13g2_buf_1 _17093_ (.A(\top_ihp.oisc.regs[24][25] ),
    .X(_01013_));
 sg13g2_buf_1 _17094_ (.A(\top_ihp.oisc.regs[24][26] ),
    .X(_01014_));
 sg13g2_buf_1 _17095_ (.A(\top_ihp.oisc.regs[24][27] ),
    .X(_01015_));
 sg13g2_buf_1 _17096_ (.A(\top_ihp.oisc.regs[24][28] ),
    .X(_01016_));
 sg13g2_buf_1 _17097_ (.A(\top_ihp.oisc.regs[24][29] ),
    .X(_01017_));
 sg13g2_buf_1 _17098_ (.A(\top_ihp.oisc.regs[24][2] ),
    .X(_01018_));
 sg13g2_buf_1 _17099_ (.A(\top_ihp.oisc.regs[24][30] ),
    .X(_01019_));
 sg13g2_buf_1 _17100_ (.A(\top_ihp.oisc.regs[24][31] ),
    .X(_01020_));
 sg13g2_buf_1 _17101_ (.A(\top_ihp.oisc.regs[24][3] ),
    .X(_01021_));
 sg13g2_buf_1 _17102_ (.A(\top_ihp.oisc.regs[24][4] ),
    .X(_01022_));
 sg13g2_buf_1 _17103_ (.A(\top_ihp.oisc.regs[24][5] ),
    .X(_01023_));
 sg13g2_buf_1 _17104_ (.A(\top_ihp.oisc.regs[24][6] ),
    .X(_01024_));
 sg13g2_buf_1 _17105_ (.A(\top_ihp.oisc.regs[24][7] ),
    .X(_01025_));
 sg13g2_buf_1 _17106_ (.A(\top_ihp.oisc.regs[24][8] ),
    .X(_01026_));
 sg13g2_buf_1 _17107_ (.A(\top_ihp.oisc.regs[24][9] ),
    .X(_01027_));
 sg13g2_buf_1 _17108_ (.A(\top_ihp.oisc.regs[25][0] ),
    .X(_01028_));
 sg13g2_buf_1 _17109_ (.A(\top_ihp.oisc.regs[25][10] ),
    .X(_01029_));
 sg13g2_buf_1 _17110_ (.A(\top_ihp.oisc.regs[25][11] ),
    .X(_01030_));
 sg13g2_buf_1 _17111_ (.A(\top_ihp.oisc.regs[25][12] ),
    .X(_01031_));
 sg13g2_buf_1 _17112_ (.A(\top_ihp.oisc.regs[25][13] ),
    .X(_01032_));
 sg13g2_buf_1 _17113_ (.A(\top_ihp.oisc.regs[25][14] ),
    .X(_01033_));
 sg13g2_buf_1 _17114_ (.A(\top_ihp.oisc.regs[25][15] ),
    .X(_01034_));
 sg13g2_buf_1 _17115_ (.A(\top_ihp.oisc.regs[25][16] ),
    .X(_01035_));
 sg13g2_buf_1 _17116_ (.A(\top_ihp.oisc.regs[25][17] ),
    .X(_01036_));
 sg13g2_buf_1 _17117_ (.A(\top_ihp.oisc.regs[25][18] ),
    .X(_01037_));
 sg13g2_buf_1 _17118_ (.A(\top_ihp.oisc.regs[25][19] ),
    .X(_01038_));
 sg13g2_buf_1 _17119_ (.A(\top_ihp.oisc.regs[25][1] ),
    .X(_01039_));
 sg13g2_buf_1 _17120_ (.A(\top_ihp.oisc.regs[25][20] ),
    .X(_01040_));
 sg13g2_buf_1 _17121_ (.A(\top_ihp.oisc.regs[25][21] ),
    .X(_01041_));
 sg13g2_buf_1 _17122_ (.A(\top_ihp.oisc.regs[25][22] ),
    .X(_01042_));
 sg13g2_buf_1 _17123_ (.A(\top_ihp.oisc.regs[25][23] ),
    .X(_01043_));
 sg13g2_buf_1 _17124_ (.A(\top_ihp.oisc.regs[25][24] ),
    .X(_01044_));
 sg13g2_buf_1 _17125_ (.A(\top_ihp.oisc.regs[25][25] ),
    .X(_01045_));
 sg13g2_buf_1 _17126_ (.A(\top_ihp.oisc.regs[25][26] ),
    .X(_01046_));
 sg13g2_buf_1 _17127_ (.A(\top_ihp.oisc.regs[25][27] ),
    .X(_01047_));
 sg13g2_buf_1 _17128_ (.A(\top_ihp.oisc.regs[25][28] ),
    .X(_01048_));
 sg13g2_buf_1 _17129_ (.A(\top_ihp.oisc.regs[25][29] ),
    .X(_01049_));
 sg13g2_buf_1 _17130_ (.A(\top_ihp.oisc.regs[25][2] ),
    .X(_01050_));
 sg13g2_buf_1 _17131_ (.A(\top_ihp.oisc.regs[25][30] ),
    .X(_01051_));
 sg13g2_buf_1 _17132_ (.A(\top_ihp.oisc.regs[25][31] ),
    .X(_01052_));
 sg13g2_buf_1 _17133_ (.A(\top_ihp.oisc.regs[25][3] ),
    .X(_01053_));
 sg13g2_buf_1 _17134_ (.A(\top_ihp.oisc.regs[25][4] ),
    .X(_01054_));
 sg13g2_buf_1 _17135_ (.A(\top_ihp.oisc.regs[25][5] ),
    .X(_01055_));
 sg13g2_buf_1 _17136_ (.A(\top_ihp.oisc.regs[25][6] ),
    .X(_01056_));
 sg13g2_buf_1 _17137_ (.A(\top_ihp.oisc.regs[25][7] ),
    .X(_01057_));
 sg13g2_buf_1 _17138_ (.A(\top_ihp.oisc.regs[25][8] ),
    .X(_01058_));
 sg13g2_buf_1 _17139_ (.A(\top_ihp.oisc.regs[25][9] ),
    .X(_01059_));
 sg13g2_buf_1 _17140_ (.A(\top_ihp.oisc.regs[26][0] ),
    .X(_01060_));
 sg13g2_buf_1 _17141_ (.A(\top_ihp.oisc.regs[26][10] ),
    .X(_01061_));
 sg13g2_buf_1 _17142_ (.A(\top_ihp.oisc.regs[26][11] ),
    .X(_01062_));
 sg13g2_buf_1 _17143_ (.A(\top_ihp.oisc.regs[26][12] ),
    .X(_01063_));
 sg13g2_buf_1 _17144_ (.A(\top_ihp.oisc.regs[26][13] ),
    .X(_01064_));
 sg13g2_buf_1 _17145_ (.A(\top_ihp.oisc.regs[26][14] ),
    .X(_01065_));
 sg13g2_buf_1 _17146_ (.A(\top_ihp.oisc.regs[26][15] ),
    .X(_01066_));
 sg13g2_buf_1 _17147_ (.A(\top_ihp.oisc.regs[26][16] ),
    .X(_01067_));
 sg13g2_buf_1 _17148_ (.A(\top_ihp.oisc.regs[26][17] ),
    .X(_01068_));
 sg13g2_buf_1 _17149_ (.A(\top_ihp.oisc.regs[26][18] ),
    .X(_01069_));
 sg13g2_buf_1 _17150_ (.A(\top_ihp.oisc.regs[26][19] ),
    .X(_01070_));
 sg13g2_buf_1 _17151_ (.A(\top_ihp.oisc.regs[26][1] ),
    .X(_01071_));
 sg13g2_buf_1 _17152_ (.A(\top_ihp.oisc.regs[26][20] ),
    .X(_01072_));
 sg13g2_buf_1 _17153_ (.A(\top_ihp.oisc.regs[26][21] ),
    .X(_01073_));
 sg13g2_buf_1 _17154_ (.A(\top_ihp.oisc.regs[26][22] ),
    .X(_01074_));
 sg13g2_buf_1 _17155_ (.A(\top_ihp.oisc.regs[26][23] ),
    .X(_01075_));
 sg13g2_buf_1 _17156_ (.A(\top_ihp.oisc.regs[26][24] ),
    .X(_01076_));
 sg13g2_buf_1 _17157_ (.A(\top_ihp.oisc.regs[26][25] ),
    .X(_01077_));
 sg13g2_buf_1 _17158_ (.A(\top_ihp.oisc.regs[26][26] ),
    .X(_01078_));
 sg13g2_buf_1 _17159_ (.A(\top_ihp.oisc.regs[26][27] ),
    .X(_01079_));
 sg13g2_buf_1 _17160_ (.A(\top_ihp.oisc.regs[26][28] ),
    .X(_01080_));
 sg13g2_buf_1 _17161_ (.A(\top_ihp.oisc.regs[26][29] ),
    .X(_01081_));
 sg13g2_buf_1 _17162_ (.A(\top_ihp.oisc.regs[26][2] ),
    .X(_01082_));
 sg13g2_buf_1 _17163_ (.A(\top_ihp.oisc.regs[26][30] ),
    .X(_01083_));
 sg13g2_buf_1 _17164_ (.A(\top_ihp.oisc.regs[26][31] ),
    .X(_01084_));
 sg13g2_buf_1 _17165_ (.A(\top_ihp.oisc.regs[26][3] ),
    .X(_01085_));
 sg13g2_buf_1 _17166_ (.A(\top_ihp.oisc.regs[26][4] ),
    .X(_01086_));
 sg13g2_buf_1 _17167_ (.A(\top_ihp.oisc.regs[26][5] ),
    .X(_01087_));
 sg13g2_buf_1 _17168_ (.A(\top_ihp.oisc.regs[26][6] ),
    .X(_01088_));
 sg13g2_buf_1 _17169_ (.A(\top_ihp.oisc.regs[26][7] ),
    .X(_01089_));
 sg13g2_buf_1 _17170_ (.A(\top_ihp.oisc.regs[26][8] ),
    .X(_01090_));
 sg13g2_buf_1 _17171_ (.A(\top_ihp.oisc.regs[26][9] ),
    .X(_01091_));
 sg13g2_buf_1 _17172_ (.A(\top_ihp.oisc.regs[27][0] ),
    .X(_01092_));
 sg13g2_buf_1 _17173_ (.A(\top_ihp.oisc.regs[27][10] ),
    .X(_01093_));
 sg13g2_buf_1 _17174_ (.A(\top_ihp.oisc.regs[27][11] ),
    .X(_01094_));
 sg13g2_buf_1 _17175_ (.A(\top_ihp.oisc.regs[27][12] ),
    .X(_01095_));
 sg13g2_buf_1 _17176_ (.A(\top_ihp.oisc.regs[27][13] ),
    .X(_01096_));
 sg13g2_buf_1 _17177_ (.A(\top_ihp.oisc.regs[27][14] ),
    .X(_01097_));
 sg13g2_buf_1 _17178_ (.A(\top_ihp.oisc.regs[27][15] ),
    .X(_01098_));
 sg13g2_buf_1 _17179_ (.A(\top_ihp.oisc.regs[27][16] ),
    .X(_01099_));
 sg13g2_buf_1 _17180_ (.A(\top_ihp.oisc.regs[27][17] ),
    .X(_01100_));
 sg13g2_buf_1 _17181_ (.A(\top_ihp.oisc.regs[27][18] ),
    .X(_01101_));
 sg13g2_buf_1 _17182_ (.A(\top_ihp.oisc.regs[27][19] ),
    .X(_01102_));
 sg13g2_buf_1 _17183_ (.A(\top_ihp.oisc.regs[27][1] ),
    .X(_01103_));
 sg13g2_buf_1 _17184_ (.A(\top_ihp.oisc.regs[27][20] ),
    .X(_01104_));
 sg13g2_buf_1 _17185_ (.A(\top_ihp.oisc.regs[27][21] ),
    .X(_01105_));
 sg13g2_buf_1 _17186_ (.A(\top_ihp.oisc.regs[27][22] ),
    .X(_01106_));
 sg13g2_buf_1 _17187_ (.A(\top_ihp.oisc.regs[27][23] ),
    .X(_01107_));
 sg13g2_buf_1 _17188_ (.A(\top_ihp.oisc.regs[27][24] ),
    .X(_01108_));
 sg13g2_buf_1 _17189_ (.A(\top_ihp.oisc.regs[27][25] ),
    .X(_01109_));
 sg13g2_buf_1 _17190_ (.A(\top_ihp.oisc.regs[27][26] ),
    .X(_01110_));
 sg13g2_buf_1 _17191_ (.A(\top_ihp.oisc.regs[27][27] ),
    .X(_01111_));
 sg13g2_buf_1 _17192_ (.A(\top_ihp.oisc.regs[27][28] ),
    .X(_01112_));
 sg13g2_buf_1 _17193_ (.A(\top_ihp.oisc.regs[27][29] ),
    .X(_01113_));
 sg13g2_buf_1 _17194_ (.A(\top_ihp.oisc.regs[27][2] ),
    .X(_01114_));
 sg13g2_buf_1 _17195_ (.A(\top_ihp.oisc.regs[27][30] ),
    .X(_01115_));
 sg13g2_buf_1 _17196_ (.A(\top_ihp.oisc.regs[27][31] ),
    .X(_01116_));
 sg13g2_buf_1 _17197_ (.A(\top_ihp.oisc.regs[27][3] ),
    .X(_01117_));
 sg13g2_buf_1 _17198_ (.A(\top_ihp.oisc.regs[27][4] ),
    .X(_01118_));
 sg13g2_buf_1 _17199_ (.A(\top_ihp.oisc.regs[27][5] ),
    .X(_01119_));
 sg13g2_buf_1 _17200_ (.A(\top_ihp.oisc.regs[27][6] ),
    .X(_01120_));
 sg13g2_buf_1 _17201_ (.A(\top_ihp.oisc.regs[27][7] ),
    .X(_01121_));
 sg13g2_buf_1 _17202_ (.A(\top_ihp.oisc.regs[27][8] ),
    .X(_01122_));
 sg13g2_buf_1 _17203_ (.A(\top_ihp.oisc.regs[27][9] ),
    .X(_01123_));
 sg13g2_buf_1 _17204_ (.A(\top_ihp.oisc.regs[28][0] ),
    .X(_01124_));
 sg13g2_buf_1 _17205_ (.A(\top_ihp.oisc.regs[28][10] ),
    .X(_01125_));
 sg13g2_buf_1 _17206_ (.A(\top_ihp.oisc.regs[28][11] ),
    .X(_01126_));
 sg13g2_buf_1 _17207_ (.A(\top_ihp.oisc.regs[28][12] ),
    .X(_01127_));
 sg13g2_buf_1 _17208_ (.A(\top_ihp.oisc.regs[28][13] ),
    .X(_01128_));
 sg13g2_buf_1 _17209_ (.A(\top_ihp.oisc.regs[28][14] ),
    .X(_01129_));
 sg13g2_buf_1 _17210_ (.A(\top_ihp.oisc.regs[28][15] ),
    .X(_01130_));
 sg13g2_buf_1 _17211_ (.A(\top_ihp.oisc.regs[28][16] ),
    .X(_01131_));
 sg13g2_buf_1 _17212_ (.A(\top_ihp.oisc.regs[28][17] ),
    .X(_01132_));
 sg13g2_buf_1 _17213_ (.A(\top_ihp.oisc.regs[28][18] ),
    .X(_01133_));
 sg13g2_buf_1 _17214_ (.A(\top_ihp.oisc.regs[28][19] ),
    .X(_01134_));
 sg13g2_buf_1 _17215_ (.A(\top_ihp.oisc.regs[28][1] ),
    .X(_01135_));
 sg13g2_buf_1 _17216_ (.A(\top_ihp.oisc.regs[28][20] ),
    .X(_01136_));
 sg13g2_buf_1 _17217_ (.A(\top_ihp.oisc.regs[28][21] ),
    .X(_01137_));
 sg13g2_buf_1 _17218_ (.A(\top_ihp.oisc.regs[28][22] ),
    .X(_01138_));
 sg13g2_buf_1 _17219_ (.A(\top_ihp.oisc.regs[28][23] ),
    .X(_01139_));
 sg13g2_buf_1 _17220_ (.A(\top_ihp.oisc.regs[28][24] ),
    .X(_01140_));
 sg13g2_buf_1 _17221_ (.A(\top_ihp.oisc.regs[28][25] ),
    .X(_01141_));
 sg13g2_buf_1 _17222_ (.A(\top_ihp.oisc.regs[28][26] ),
    .X(_01142_));
 sg13g2_buf_1 _17223_ (.A(\top_ihp.oisc.regs[28][27] ),
    .X(_01143_));
 sg13g2_buf_1 _17224_ (.A(\top_ihp.oisc.regs[28][28] ),
    .X(_01144_));
 sg13g2_buf_1 _17225_ (.A(\top_ihp.oisc.regs[28][29] ),
    .X(_01145_));
 sg13g2_buf_1 _17226_ (.A(\top_ihp.oisc.regs[28][2] ),
    .X(_01146_));
 sg13g2_buf_1 _17227_ (.A(\top_ihp.oisc.regs[28][30] ),
    .X(_01147_));
 sg13g2_buf_1 _17228_ (.A(\top_ihp.oisc.regs[28][31] ),
    .X(_01148_));
 sg13g2_buf_1 _17229_ (.A(\top_ihp.oisc.regs[28][3] ),
    .X(_01149_));
 sg13g2_buf_1 _17230_ (.A(\top_ihp.oisc.regs[28][4] ),
    .X(_01150_));
 sg13g2_buf_1 _17231_ (.A(\top_ihp.oisc.regs[28][5] ),
    .X(_01151_));
 sg13g2_buf_1 _17232_ (.A(\top_ihp.oisc.regs[28][6] ),
    .X(_01152_));
 sg13g2_buf_1 _17233_ (.A(\top_ihp.oisc.regs[28][7] ),
    .X(_01153_));
 sg13g2_buf_1 _17234_ (.A(\top_ihp.oisc.regs[28][8] ),
    .X(_01154_));
 sg13g2_buf_1 _17235_ (.A(\top_ihp.oisc.regs[28][9] ),
    .X(_01155_));
 sg13g2_buf_1 _17236_ (.A(\top_ihp.oisc.regs[29][0] ),
    .X(_01156_));
 sg13g2_buf_1 _17237_ (.A(\top_ihp.oisc.regs[29][10] ),
    .X(_01157_));
 sg13g2_buf_1 _17238_ (.A(\top_ihp.oisc.regs[29][11] ),
    .X(_01158_));
 sg13g2_buf_1 _17239_ (.A(\top_ihp.oisc.regs[29][12] ),
    .X(_01159_));
 sg13g2_buf_1 _17240_ (.A(\top_ihp.oisc.regs[29][13] ),
    .X(_01160_));
 sg13g2_buf_1 _17241_ (.A(\top_ihp.oisc.regs[29][14] ),
    .X(_01161_));
 sg13g2_buf_1 _17242_ (.A(\top_ihp.oisc.regs[29][15] ),
    .X(_01162_));
 sg13g2_buf_1 _17243_ (.A(\top_ihp.oisc.regs[29][16] ),
    .X(_01163_));
 sg13g2_buf_1 _17244_ (.A(\top_ihp.oisc.regs[29][17] ),
    .X(_01164_));
 sg13g2_buf_1 _17245_ (.A(\top_ihp.oisc.regs[29][18] ),
    .X(_01165_));
 sg13g2_buf_1 _17246_ (.A(\top_ihp.oisc.regs[29][19] ),
    .X(_01166_));
 sg13g2_buf_1 _17247_ (.A(\top_ihp.oisc.regs[29][1] ),
    .X(_01167_));
 sg13g2_buf_1 _17248_ (.A(\top_ihp.oisc.regs[29][20] ),
    .X(_01168_));
 sg13g2_buf_1 _17249_ (.A(\top_ihp.oisc.regs[29][21] ),
    .X(_01169_));
 sg13g2_buf_1 _17250_ (.A(\top_ihp.oisc.regs[29][22] ),
    .X(_01170_));
 sg13g2_buf_1 _17251_ (.A(\top_ihp.oisc.regs[29][23] ),
    .X(_01171_));
 sg13g2_buf_1 _17252_ (.A(\top_ihp.oisc.regs[29][24] ),
    .X(_01172_));
 sg13g2_buf_1 _17253_ (.A(\top_ihp.oisc.regs[29][25] ),
    .X(_01173_));
 sg13g2_buf_1 _17254_ (.A(\top_ihp.oisc.regs[29][26] ),
    .X(_01174_));
 sg13g2_buf_1 _17255_ (.A(\top_ihp.oisc.regs[29][27] ),
    .X(_01175_));
 sg13g2_buf_1 _17256_ (.A(\top_ihp.oisc.regs[29][28] ),
    .X(_01176_));
 sg13g2_buf_1 _17257_ (.A(\top_ihp.oisc.regs[29][29] ),
    .X(_01177_));
 sg13g2_buf_1 _17258_ (.A(\top_ihp.oisc.regs[29][2] ),
    .X(_01178_));
 sg13g2_buf_1 _17259_ (.A(\top_ihp.oisc.regs[29][30] ),
    .X(_01179_));
 sg13g2_buf_1 _17260_ (.A(\top_ihp.oisc.regs[29][31] ),
    .X(_01180_));
 sg13g2_buf_1 _17261_ (.A(\top_ihp.oisc.regs[29][3] ),
    .X(_01181_));
 sg13g2_buf_1 _17262_ (.A(\top_ihp.oisc.regs[29][4] ),
    .X(_01182_));
 sg13g2_buf_1 _17263_ (.A(\top_ihp.oisc.regs[29][5] ),
    .X(_01183_));
 sg13g2_buf_1 _17264_ (.A(\top_ihp.oisc.regs[29][6] ),
    .X(_01184_));
 sg13g2_buf_1 _17265_ (.A(\top_ihp.oisc.regs[29][7] ),
    .X(_01185_));
 sg13g2_buf_1 _17266_ (.A(\top_ihp.oisc.regs[29][8] ),
    .X(_01186_));
 sg13g2_buf_1 _17267_ (.A(\top_ihp.oisc.regs[29][9] ),
    .X(_01187_));
 sg13g2_nor2_1 _17268_ (.A(_10912_),
    .B(_10707_),
    .Y(_10948_));
 sg13g2_buf_4 _17269_ (.X(_10949_),
    .A(_10948_));
 sg13g2_mux2_1 _17270_ (.A0(\top_ihp.oisc.regs[2][0] ),
    .A1(net119),
    .S(_10949_),
    .X(_01188_));
 sg13g2_mux2_1 _17271_ (.A0(\top_ihp.oisc.regs[2][10] ),
    .A1(net130),
    .S(_10949_),
    .X(_01189_));
 sg13g2_nand2_1 _17272_ (.Y(_10950_),
    .A(net692),
    .B(_10698_));
 sg13g2_buf_1 _17273_ (.A(_10950_),
    .X(_10951_));
 sg13g2_buf_1 _17274_ (.A(_10951_),
    .X(_10952_));
 sg13g2_buf_1 _17275_ (.A(net392),
    .X(_10953_));
 sg13g2_buf_1 _17276_ (.A(_10951_),
    .X(_10954_));
 sg13g2_nand2_1 _17277_ (.Y(_10955_),
    .A(\top_ihp.oisc.regs[2][11] ),
    .B(_10954_));
 sg13g2_o21ai_1 _17278_ (.B1(_10955_),
    .Y(_01190_),
    .A1(net62),
    .A2(_10953_));
 sg13g2_nand2_1 _17279_ (.Y(_10956_),
    .A(\top_ihp.oisc.regs[2][12] ),
    .B(net391));
 sg13g2_o21ai_1 _17280_ (.B1(_10956_),
    .Y(_01191_),
    .A1(_10888_),
    .A2(net253));
 sg13g2_nand2_1 _17281_ (.Y(_10957_),
    .A(\top_ihp.oisc.regs[2][13] ),
    .B(net391));
 sg13g2_o21ai_1 _17282_ (.B1(_10957_),
    .Y(_01192_),
    .A1(net278),
    .A2(net253));
 sg13g2_nand2_1 _17283_ (.Y(_10958_),
    .A(\top_ihp.oisc.regs[2][14] ),
    .B(net391));
 sg13g2_o21ai_1 _17284_ (.B1(_10958_),
    .Y(_01193_),
    .A1(_10159_),
    .A2(net253));
 sg13g2_nand2_1 _17285_ (.Y(_10959_),
    .A(\top_ihp.oisc.regs[2][15] ),
    .B(net391));
 sg13g2_o21ai_1 _17286_ (.B1(_10959_),
    .Y(_01194_),
    .A1(_10171_),
    .A2(net253));
 sg13g2_nand2_1 _17287_ (.Y(_10960_),
    .A(\top_ihp.oisc.regs[2][16] ),
    .B(net391));
 sg13g2_o21ai_1 _17288_ (.B1(_10960_),
    .Y(_01195_),
    .A1(net140),
    .A2(net253));
 sg13g2_buf_1 _17289_ (.A(_10951_),
    .X(_10961_));
 sg13g2_nand2_1 _17290_ (.Y(_10962_),
    .A(\top_ihp.oisc.regs[2][17] ),
    .B(net390));
 sg13g2_o21ai_1 _17291_ (.B1(_10962_),
    .Y(_01196_),
    .A1(_10224_),
    .A2(net253));
 sg13g2_nand2_1 _17292_ (.Y(_10963_),
    .A(\top_ihp.oisc.regs[2][18] ),
    .B(net390));
 sg13g2_o21ai_1 _17293_ (.B1(_10963_),
    .Y(_01197_),
    .A1(net275),
    .A2(_10953_));
 sg13g2_nand2_1 _17294_ (.Y(_10964_),
    .A(\top_ihp.oisc.regs[2][19] ),
    .B(net390));
 sg13g2_o21ai_1 _17295_ (.B1(_10964_),
    .Y(_01198_),
    .A1(_10274_),
    .A2(net253));
 sg13g2_buf_1 _17296_ (.A(net392),
    .X(_10965_));
 sg13g2_nand2_1 _17297_ (.Y(_10966_),
    .A(\top_ihp.oisc.regs[2][1] ),
    .B(net390));
 sg13g2_o21ai_1 _17298_ (.B1(_10966_),
    .Y(_01199_),
    .A1(_10834_),
    .A2(net252));
 sg13g2_nand2_1 _17299_ (.Y(_10967_),
    .A(\top_ihp.oisc.regs[2][20] ),
    .B(net390));
 sg13g2_o21ai_1 _17300_ (.B1(_10967_),
    .Y(_01200_),
    .A1(_10343_),
    .A2(net252));
 sg13g2_nand2_1 _17301_ (.Y(_10968_),
    .A(\top_ihp.oisc.regs[2][21] ),
    .B(net390));
 sg13g2_o21ai_1 _17302_ (.B1(_10968_),
    .Y(_01201_),
    .A1(_10362_),
    .A2(net252));
 sg13g2_nand2_1 _17303_ (.Y(_10969_),
    .A(\top_ihp.oisc.regs[2][22] ),
    .B(net390));
 sg13g2_o21ai_1 _17304_ (.B1(_10969_),
    .Y(_01202_),
    .A1(net272),
    .A2(net252));
 sg13g2_nand2_1 _17305_ (.Y(_10970_),
    .A(\top_ihp.oisc.regs[2][23] ),
    .B(_10961_));
 sg13g2_o21ai_1 _17306_ (.B1(_10970_),
    .Y(_01203_),
    .A1(_10393_),
    .A2(net252));
 sg13g2_mux2_1 _17307_ (.A0(\top_ihp.oisc.regs[2][24] ),
    .A1(net400),
    .S(_10949_),
    .X(_01204_));
 sg13g2_nand2_1 _17308_ (.Y(_10971_),
    .A(\top_ihp.oisc.regs[2][25] ),
    .B(net390));
 sg13g2_o21ai_1 _17309_ (.B1(_10971_),
    .Y(_01205_),
    .A1(_10429_),
    .A2(net252));
 sg13g2_nand2_1 _17310_ (.Y(_10972_),
    .A(\top_ihp.oisc.regs[2][26] ),
    .B(_10961_));
 sg13g2_o21ai_1 _17311_ (.B1(_10972_),
    .Y(_01206_),
    .A1(_10441_),
    .A2(_10965_));
 sg13g2_nand2_1 _17312_ (.Y(_10973_),
    .A(\top_ihp.oisc.regs[2][27] ),
    .B(net392));
 sg13g2_o21ai_1 _17313_ (.B1(_10973_),
    .Y(_01207_),
    .A1(_10450_),
    .A2(net252));
 sg13g2_buf_8 _17314_ (.A(_10459_),
    .X(_10974_));
 sg13g2_nand2_1 _17315_ (.Y(_10975_),
    .A(\top_ihp.oisc.regs[2][28] ),
    .B(net392));
 sg13g2_o21ai_1 _17316_ (.B1(_10975_),
    .Y(_01208_),
    .A1(_10974_),
    .A2(net252));
 sg13g2_nand2_1 _17317_ (.Y(_10976_),
    .A(\top_ihp.oisc.regs[2][29] ),
    .B(net392));
 sg13g2_o21ai_1 _17318_ (.B1(_10976_),
    .Y(_01209_),
    .A1(_10467_),
    .A2(_10965_));
 sg13g2_nand2_1 _17319_ (.Y(_10977_),
    .A(\top_ihp.oisc.regs[2][2] ),
    .B(net392));
 sg13g2_o21ai_1 _17320_ (.B1(_10977_),
    .Y(_01210_),
    .A1(_10500_),
    .A2(net391));
 sg13g2_nand2_1 _17321_ (.Y(_10978_),
    .A(\top_ihp.oisc.regs[2][30] ),
    .B(net392));
 sg13g2_o21ai_1 _17322_ (.B1(_10978_),
    .Y(_01211_),
    .A1(_10509_),
    .A2(net391));
 sg13g2_inv_1 _17323_ (.Y(_10979_),
    .A(\top_ihp.oisc.regs[2][31] ));
 sg13g2_nor2_1 _17324_ (.A(_10536_),
    .B(net392),
    .Y(_10980_));
 sg13g2_a22oi_1 _17325_ (.Y(_01212_),
    .B1(_10980_),
    .B2(_10738_),
    .A2(net253),
    .A1(_10979_));
 sg13g2_mux2_1 _17326_ (.A0(\top_ihp.oisc.regs[2][3] ),
    .A1(net128),
    .S(_10949_),
    .X(_01213_));
 sg13g2_mux2_1 _17327_ (.A0(\top_ihp.oisc.regs[2][4] ),
    .A1(net127),
    .S(_10949_),
    .X(_01214_));
 sg13g2_mux2_1 _17328_ (.A0(\top_ihp.oisc.regs[2][5] ),
    .A1(net264),
    .S(_10949_),
    .X(_01215_));
 sg13g2_mux2_1 _17329_ (.A0(\top_ihp.oisc.regs[2][6] ),
    .A1(net126),
    .S(_10949_),
    .X(_01216_));
 sg13g2_nand2_1 _17330_ (.Y(_10981_),
    .A(\top_ihp.oisc.regs[2][7] ),
    .B(_10952_));
 sg13g2_o21ai_1 _17331_ (.B1(_10981_),
    .Y(_01217_),
    .A1(_10662_),
    .A2(net391));
 sg13g2_nand2_1 _17332_ (.Y(_10982_),
    .A(\top_ihp.oisc.regs[2][8] ),
    .B(_10952_));
 sg13g2_o21ai_1 _17333_ (.B1(_10982_),
    .Y(_01218_),
    .A1(net266),
    .A2(_10954_));
 sg13g2_mux2_1 _17334_ (.A0(\top_ihp.oisc.regs[2][9] ),
    .A1(net125),
    .S(_10949_),
    .X(_01219_));
 sg13g2_buf_1 _17335_ (.A(\top_ihp.oisc.regs[30][0] ),
    .X(_01220_));
 sg13g2_buf_1 _17336_ (.A(\top_ihp.oisc.regs[30][10] ),
    .X(_01221_));
 sg13g2_buf_1 _17337_ (.A(\top_ihp.oisc.regs[30][11] ),
    .X(_01222_));
 sg13g2_buf_1 _17338_ (.A(\top_ihp.oisc.regs[30][12] ),
    .X(_01223_));
 sg13g2_buf_1 _17339_ (.A(\top_ihp.oisc.regs[30][13] ),
    .X(_01224_));
 sg13g2_buf_1 _17340_ (.A(\top_ihp.oisc.regs[30][14] ),
    .X(_01225_));
 sg13g2_buf_1 _17341_ (.A(\top_ihp.oisc.regs[30][15] ),
    .X(_01226_));
 sg13g2_buf_1 _17342_ (.A(\top_ihp.oisc.regs[30][16] ),
    .X(_01227_));
 sg13g2_buf_1 _17343_ (.A(\top_ihp.oisc.regs[30][17] ),
    .X(_01228_));
 sg13g2_buf_1 _17344_ (.A(\top_ihp.oisc.regs[30][18] ),
    .X(_01229_));
 sg13g2_buf_1 _17345_ (.A(\top_ihp.oisc.regs[30][19] ),
    .X(_01230_));
 sg13g2_buf_1 _17346_ (.A(\top_ihp.oisc.regs[30][1] ),
    .X(_01231_));
 sg13g2_buf_1 _17347_ (.A(\top_ihp.oisc.regs[30][20] ),
    .X(_01232_));
 sg13g2_buf_1 _17348_ (.A(\top_ihp.oisc.regs[30][21] ),
    .X(_01233_));
 sg13g2_buf_1 _17349_ (.A(\top_ihp.oisc.regs[30][22] ),
    .X(_01234_));
 sg13g2_buf_1 _17350_ (.A(\top_ihp.oisc.regs[30][23] ),
    .X(_01235_));
 sg13g2_buf_1 _17351_ (.A(\top_ihp.oisc.regs[30][24] ),
    .X(_01236_));
 sg13g2_buf_1 _17352_ (.A(\top_ihp.oisc.regs[30][25] ),
    .X(_01237_));
 sg13g2_buf_1 _17353_ (.A(\top_ihp.oisc.regs[30][26] ),
    .X(_01238_));
 sg13g2_buf_1 _17354_ (.A(\top_ihp.oisc.regs[30][27] ),
    .X(_01239_));
 sg13g2_buf_1 _17355_ (.A(\top_ihp.oisc.regs[30][28] ),
    .X(_01240_));
 sg13g2_buf_1 _17356_ (.A(\top_ihp.oisc.regs[30][29] ),
    .X(_01241_));
 sg13g2_buf_1 _17357_ (.A(\top_ihp.oisc.regs[30][2] ),
    .X(_01242_));
 sg13g2_buf_1 _17358_ (.A(\top_ihp.oisc.regs[30][30] ),
    .X(_01243_));
 sg13g2_buf_1 _17359_ (.A(\top_ihp.oisc.regs[30][31] ),
    .X(_01244_));
 sg13g2_buf_1 _17360_ (.A(\top_ihp.oisc.regs[30][3] ),
    .X(_01245_));
 sg13g2_buf_1 _17361_ (.A(\top_ihp.oisc.regs[30][4] ),
    .X(_01246_));
 sg13g2_buf_1 _17362_ (.A(\top_ihp.oisc.regs[30][5] ),
    .X(_01247_));
 sg13g2_buf_1 _17363_ (.A(\top_ihp.oisc.regs[30][6] ),
    .X(_01248_));
 sg13g2_buf_1 _17364_ (.A(\top_ihp.oisc.regs[30][7] ),
    .X(_01249_));
 sg13g2_buf_1 _17365_ (.A(\top_ihp.oisc.regs[30][8] ),
    .X(_01250_));
 sg13g2_buf_1 _17366_ (.A(\top_ihp.oisc.regs[30][9] ),
    .X(_01251_));
 sg13g2_buf_1 _17367_ (.A(\top_ihp.oisc.regs[31][0] ),
    .X(_01252_));
 sg13g2_buf_1 _17368_ (.A(\top_ihp.oisc.regs[31][10] ),
    .X(_01253_));
 sg13g2_buf_1 _17369_ (.A(\top_ihp.oisc.regs[31][11] ),
    .X(_01254_));
 sg13g2_buf_1 _17370_ (.A(\top_ihp.oisc.regs[31][12] ),
    .X(_01255_));
 sg13g2_buf_1 _17371_ (.A(\top_ihp.oisc.regs[31][13] ),
    .X(_01256_));
 sg13g2_buf_1 _17372_ (.A(\top_ihp.oisc.regs[31][14] ),
    .X(_01257_));
 sg13g2_buf_1 _17373_ (.A(\top_ihp.oisc.regs[31][15] ),
    .X(_01258_));
 sg13g2_buf_1 _17374_ (.A(\top_ihp.oisc.regs[31][16] ),
    .X(_01259_));
 sg13g2_buf_1 _17375_ (.A(\top_ihp.oisc.regs[31][17] ),
    .X(_01260_));
 sg13g2_buf_1 _17376_ (.A(\top_ihp.oisc.regs[31][18] ),
    .X(_01261_));
 sg13g2_buf_1 _17377_ (.A(\top_ihp.oisc.regs[31][19] ),
    .X(_01262_));
 sg13g2_buf_1 _17378_ (.A(\top_ihp.oisc.regs[31][1] ),
    .X(_01263_));
 sg13g2_buf_1 _17379_ (.A(\top_ihp.oisc.regs[31][20] ),
    .X(_01264_));
 sg13g2_buf_1 _17380_ (.A(\top_ihp.oisc.regs[31][21] ),
    .X(_01265_));
 sg13g2_buf_1 _17381_ (.A(\top_ihp.oisc.regs[31][22] ),
    .X(_01266_));
 sg13g2_buf_1 _17382_ (.A(\top_ihp.oisc.regs[31][23] ),
    .X(_01267_));
 sg13g2_buf_1 _17383_ (.A(\top_ihp.oisc.regs[31][24] ),
    .X(_01268_));
 sg13g2_buf_1 _17384_ (.A(\top_ihp.oisc.regs[31][25] ),
    .X(_01269_));
 sg13g2_buf_1 _17385_ (.A(\top_ihp.oisc.regs[31][26] ),
    .X(_01270_));
 sg13g2_buf_1 _17386_ (.A(\top_ihp.oisc.regs[31][27] ),
    .X(_01271_));
 sg13g2_buf_1 _17387_ (.A(\top_ihp.oisc.regs[31][28] ),
    .X(_01272_));
 sg13g2_buf_1 _17388_ (.A(\top_ihp.oisc.regs[31][29] ),
    .X(_01273_));
 sg13g2_buf_1 _17389_ (.A(\top_ihp.oisc.regs[31][2] ),
    .X(_01274_));
 sg13g2_buf_1 _17390_ (.A(\top_ihp.oisc.regs[31][30] ),
    .X(_01275_));
 sg13g2_buf_1 _17391_ (.A(\top_ihp.oisc.regs[31][31] ),
    .X(_01276_));
 sg13g2_buf_1 _17392_ (.A(\top_ihp.oisc.regs[31][3] ),
    .X(_01277_));
 sg13g2_buf_1 _17393_ (.A(\top_ihp.oisc.regs[31][4] ),
    .X(_01278_));
 sg13g2_buf_1 _17394_ (.A(\top_ihp.oisc.regs[31][5] ),
    .X(_01279_));
 sg13g2_buf_1 _17395_ (.A(\top_ihp.oisc.regs[31][6] ),
    .X(_01280_));
 sg13g2_buf_1 _17396_ (.A(\top_ihp.oisc.regs[31][7] ),
    .X(_01281_));
 sg13g2_buf_1 _17397_ (.A(\top_ihp.oisc.regs[31][8] ),
    .X(_01282_));
 sg13g2_buf_1 _17398_ (.A(\top_ihp.oisc.regs[31][9] ),
    .X(_01283_));
 sg13g2_buf_1 _17399_ (.A(\top_ihp.oisc.regs[32][0] ),
    .X(_01284_));
 sg13g2_buf_1 _17400_ (.A(\top_ihp.oisc.regs[32][10] ),
    .X(_01285_));
 sg13g2_buf_1 _17401_ (.A(\top_ihp.oisc.regs[32][11] ),
    .X(_01286_));
 sg13g2_buf_1 _17402_ (.A(\top_ihp.oisc.regs[32][12] ),
    .X(_01287_));
 sg13g2_buf_1 _17403_ (.A(\top_ihp.oisc.regs[32][13] ),
    .X(_01288_));
 sg13g2_buf_1 _17404_ (.A(\top_ihp.oisc.regs[32][14] ),
    .X(_01289_));
 sg13g2_buf_1 _17405_ (.A(\top_ihp.oisc.regs[32][15] ),
    .X(_01290_));
 sg13g2_buf_1 _17406_ (.A(\top_ihp.oisc.regs[32][16] ),
    .X(_01291_));
 sg13g2_buf_1 _17407_ (.A(\top_ihp.oisc.regs[32][17] ),
    .X(_01292_));
 sg13g2_buf_1 _17408_ (.A(\top_ihp.oisc.regs[32][18] ),
    .X(_01293_));
 sg13g2_buf_1 _17409_ (.A(\top_ihp.oisc.regs[32][19] ),
    .X(_01294_));
 sg13g2_buf_1 _17410_ (.A(\top_ihp.oisc.regs[32][1] ),
    .X(_01295_));
 sg13g2_buf_1 _17411_ (.A(\top_ihp.oisc.regs[32][20] ),
    .X(_01296_));
 sg13g2_buf_1 _17412_ (.A(\top_ihp.oisc.regs[32][21] ),
    .X(_01297_));
 sg13g2_buf_1 _17413_ (.A(\top_ihp.oisc.regs[32][22] ),
    .X(_01298_));
 sg13g2_buf_1 _17414_ (.A(\top_ihp.oisc.regs[32][23] ),
    .X(_01299_));
 sg13g2_buf_1 _17415_ (.A(\top_ihp.oisc.regs[32][24] ),
    .X(_01300_));
 sg13g2_buf_1 _17416_ (.A(\top_ihp.oisc.regs[32][25] ),
    .X(_01301_));
 sg13g2_buf_1 _17417_ (.A(\top_ihp.oisc.regs[32][26] ),
    .X(_01302_));
 sg13g2_buf_1 _17418_ (.A(\top_ihp.oisc.regs[32][27] ),
    .X(_01303_));
 sg13g2_buf_1 _17419_ (.A(\top_ihp.oisc.regs[32][28] ),
    .X(_01304_));
 sg13g2_buf_1 _17420_ (.A(\top_ihp.oisc.regs[32][29] ),
    .X(_01305_));
 sg13g2_buf_1 _17421_ (.A(\top_ihp.oisc.regs[32][2] ),
    .X(_01306_));
 sg13g2_buf_1 _17422_ (.A(\top_ihp.oisc.regs[32][30] ),
    .X(_01307_));
 sg13g2_buf_1 _17423_ (.A(\top_ihp.oisc.regs[32][31] ),
    .X(_01308_));
 sg13g2_buf_1 _17424_ (.A(\top_ihp.oisc.regs[32][3] ),
    .X(_01309_));
 sg13g2_buf_1 _17425_ (.A(\top_ihp.oisc.regs[32][4] ),
    .X(_01310_));
 sg13g2_buf_1 _17426_ (.A(\top_ihp.oisc.regs[32][5] ),
    .X(_01311_));
 sg13g2_buf_1 _17427_ (.A(\top_ihp.oisc.regs[32][6] ),
    .X(_01312_));
 sg13g2_buf_1 _17428_ (.A(\top_ihp.oisc.regs[32][7] ),
    .X(_01313_));
 sg13g2_buf_1 _17429_ (.A(\top_ihp.oisc.regs[32][8] ),
    .X(_01314_));
 sg13g2_buf_1 _17430_ (.A(\top_ihp.oisc.regs[32][9] ),
    .X(_01315_));
 sg13g2_nand3_1 _17431_ (.B(_09921_),
    .C(_09926_),
    .A(_09918_),
    .Y(_10983_));
 sg13g2_buf_1 _17432_ (.A(_10983_),
    .X(_10984_));
 sg13g2_a21oi_1 _17433_ (.A1(_09912_),
    .A2(_09939_),
    .Y(_10985_),
    .B1(_10984_));
 sg13g2_and2_1 _17434_ (.A(_09914_),
    .B(_10985_),
    .X(_10986_));
 sg13g2_buf_1 _17435_ (.A(_10986_),
    .X(_10987_));
 sg13g2_nand2_1 _17436_ (.Y(_10988_),
    .A(_10822_),
    .B(_10987_));
 sg13g2_buf_1 _17437_ (.A(_10988_),
    .X(_10989_));
 sg13g2_buf_2 _17438_ (.A(net389),
    .X(_10990_));
 sg13g2_mux2_1 _17439_ (.A0(net64),
    .A1(\top_ihp.oisc.regs[33][0] ),
    .S(net251),
    .X(_01316_));
 sg13g2_mux2_1 _17440_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[33][10] ),
    .S(net251),
    .X(_01317_));
 sg13g2_buf_1 _17441_ (.A(_10050_),
    .X(_10991_));
 sg13g2_buf_1 _17442_ (.A(net389),
    .X(_10992_));
 sg13g2_buf_1 _17443_ (.A(net389),
    .X(_10993_));
 sg13g2_nand2_1 _17444_ (.Y(_10994_),
    .A(\top_ihp.oisc.regs[33][11] ),
    .B(net249));
 sg13g2_o21ai_1 _17445_ (.B1(_10994_),
    .Y(_01318_),
    .A1(net49),
    .A2(net250));
 sg13g2_nand2_1 _17446_ (.Y(_10995_),
    .A(\top_ihp.oisc.regs[33][12] ),
    .B(net249));
 sg13g2_o21ai_1 _17447_ (.B1(_10995_),
    .Y(_01319_),
    .A1(net51),
    .A2(net250));
 sg13g2_nand2_1 _17448_ (.Y(_10996_),
    .A(\top_ihp.oisc.regs[33][13] ),
    .B(_10993_));
 sg13g2_o21ai_1 _17449_ (.B1(_10996_),
    .Y(_01320_),
    .A1(net278),
    .A2(net250));
 sg13g2_nand2_1 _17450_ (.Y(_10997_),
    .A(\top_ihp.oisc.regs[33][14] ),
    .B(net249));
 sg13g2_o21ai_1 _17451_ (.B1(_10997_),
    .Y(_01321_),
    .A1(net277),
    .A2(_10992_));
 sg13g2_nand2_1 _17452_ (.Y(_10998_),
    .A(\top_ihp.oisc.regs[33][15] ),
    .B(_10993_));
 sg13g2_o21ai_1 _17453_ (.B1(_10998_),
    .Y(_01322_),
    .A1(net407),
    .A2(net250));
 sg13g2_nand2_1 _17454_ (.Y(_10999_),
    .A(\top_ihp.oisc.regs[33][16] ),
    .B(net249));
 sg13g2_o21ai_1 _17455_ (.B1(_10999_),
    .Y(_01323_),
    .A1(net140),
    .A2(net250));
 sg13g2_nand2_1 _17456_ (.Y(_11000_),
    .A(\top_ihp.oisc.regs[33][17] ),
    .B(net249));
 sg13g2_o21ai_1 _17457_ (.B1(_11000_),
    .Y(_01324_),
    .A1(net406),
    .A2(net250));
 sg13g2_nand2_1 _17458_ (.Y(_11001_),
    .A(\top_ihp.oisc.regs[33][18] ),
    .B(net249));
 sg13g2_o21ai_1 _17459_ (.B1(_11001_),
    .Y(_01325_),
    .A1(net275),
    .A2(_10992_));
 sg13g2_mux2_1 _17460_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[33][19] ),
    .S(net251),
    .X(_01326_));
 sg13g2_buf_1 _17461_ (.A(net389),
    .X(_11002_));
 sg13g2_nand2_1 _17462_ (.Y(_11003_),
    .A(\top_ihp.oisc.regs[33][1] ),
    .B(net248));
 sg13g2_o21ai_1 _17463_ (.B1(_11003_),
    .Y(_01327_),
    .A1(net120),
    .A2(net250));
 sg13g2_nand2_1 _17464_ (.Y(_11004_),
    .A(\top_ihp.oisc.regs[33][20] ),
    .B(_11002_));
 sg13g2_o21ai_1 _17465_ (.B1(_11004_),
    .Y(_01328_),
    .A1(net138),
    .A2(net250));
 sg13g2_buf_1 _17466_ (.A(net389),
    .X(_11005_));
 sg13g2_nand2_1 _17467_ (.Y(_11006_),
    .A(\top_ihp.oisc.regs[33][21] ),
    .B(net248));
 sg13g2_o21ai_1 _17468_ (.B1(_11006_),
    .Y(_01329_),
    .A1(net137),
    .A2(net247));
 sg13g2_nand2_1 _17469_ (.Y(_11007_),
    .A(\top_ihp.oisc.regs[33][22] ),
    .B(net248));
 sg13g2_o21ai_1 _17470_ (.B1(_11007_),
    .Y(_01330_),
    .A1(net272),
    .A2(net247));
 sg13g2_nand2_1 _17471_ (.Y(_11008_),
    .A(\top_ihp.oisc.regs[33][23] ),
    .B(net248));
 sg13g2_o21ai_1 _17472_ (.B1(_11008_),
    .Y(_01331_),
    .A1(net271),
    .A2(net247));
 sg13g2_mux2_1 _17473_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[33][24] ),
    .S(net251),
    .X(_01332_));
 sg13g2_nand2_1 _17474_ (.Y(_11009_),
    .A(\top_ihp.oisc.regs[33][25] ),
    .B(net248));
 sg13g2_o21ai_1 _17475_ (.B1(_11009_),
    .Y(_01333_),
    .A1(net124),
    .A2(net247));
 sg13g2_nand2_1 _17476_ (.Y(_11010_),
    .A(\top_ihp.oisc.regs[33][26] ),
    .B(net248));
 sg13g2_o21ai_1 _17477_ (.B1(_11010_),
    .Y(_01334_),
    .A1(net402),
    .A2(net247));
 sg13g2_mux2_1 _17478_ (.A0(_10776_),
    .A1(\top_ihp.oisc.regs[33][27] ),
    .S(net251),
    .X(_01335_));
 sg13g2_nand2_1 _17479_ (.Y(_11011_),
    .A(\top_ihp.oisc.regs[33][28] ),
    .B(_11002_));
 sg13g2_o21ai_1 _17480_ (.B1(_11011_),
    .Y(_01336_),
    .A1(net29),
    .A2(_11005_));
 sg13g2_nand2_1 _17481_ (.Y(_11012_),
    .A(\top_ihp.oisc.regs[33][29] ),
    .B(net248));
 sg13g2_o21ai_1 _17482_ (.B1(_11012_),
    .Y(_01337_),
    .A1(net269),
    .A2(net247));
 sg13g2_nand2_1 _17483_ (.Y(_11013_),
    .A(\top_ihp.oisc.regs[33][2] ),
    .B(net248));
 sg13g2_o21ai_1 _17484_ (.B1(_11013_),
    .Y(_01338_),
    .A1(net136),
    .A2(net247));
 sg13g2_nand2_1 _17485_ (.Y(_11014_),
    .A(\top_ihp.oisc.regs[33][30] ),
    .B(net389));
 sg13g2_o21ai_1 _17486_ (.B1(_11014_),
    .Y(_01339_),
    .A1(net58),
    .A2(net247));
 sg13g2_nand2_1 _17487_ (.Y(_11015_),
    .A(\top_ihp.oisc.regs[33][31] ),
    .B(_10989_));
 sg13g2_o21ai_1 _17488_ (.B1(_11015_),
    .Y(_01340_),
    .A1(net268),
    .A2(_11005_));
 sg13g2_mux2_1 _17489_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[33][3] ),
    .S(_10990_),
    .X(_01341_));
 sg13g2_mux2_1 _17490_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[33][4] ),
    .S(net251),
    .X(_01342_));
 sg13g2_mux2_1 _17491_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[33][5] ),
    .S(_10990_),
    .X(_01343_));
 sg13g2_mux2_1 _17492_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[33][6] ),
    .S(net249),
    .X(_01344_));
 sg13g2_nand2_1 _17493_ (.Y(_11016_),
    .A(\top_ihp.oisc.regs[33][7] ),
    .B(net389));
 sg13g2_o21ai_1 _17494_ (.B1(_11016_),
    .Y(_01345_),
    .A1(net401),
    .A2(net251));
 sg13g2_nand2_1 _17495_ (.Y(_11017_),
    .A(\top_ihp.oisc.regs[33][8] ),
    .B(net389));
 sg13g2_o21ai_1 _17496_ (.B1(_11017_),
    .Y(_01346_),
    .A1(net266),
    .A2(net251));
 sg13g2_mux2_1 _17497_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[33][9] ),
    .S(net249),
    .X(_01347_));
 sg13g2_nand2_1 _17498_ (.Y(_11018_),
    .A(net740),
    .B(_10987_));
 sg13g2_buf_1 _17499_ (.A(_11018_),
    .X(_11019_));
 sg13g2_buf_2 _17500_ (.A(net388),
    .X(_11020_));
 sg13g2_mux2_1 _17501_ (.A0(net64),
    .A1(\top_ihp.oisc.regs[34][0] ),
    .S(_11020_),
    .X(_01348_));
 sg13g2_mux2_1 _17502_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[34][10] ),
    .S(net246),
    .X(_01349_));
 sg13g2_buf_2 _17503_ (.A(net388),
    .X(_11021_));
 sg13g2_buf_2 _17504_ (.A(net388),
    .X(_11022_));
 sg13g2_nand2_1 _17505_ (.Y(_11023_),
    .A(\top_ihp.oisc.regs[34][11] ),
    .B(net244));
 sg13g2_o21ai_1 _17506_ (.B1(_11023_),
    .Y(_01350_),
    .A1(net49),
    .A2(net245));
 sg13g2_nand2_1 _17507_ (.Y(_11024_),
    .A(\top_ihp.oisc.regs[34][12] ),
    .B(net244));
 sg13g2_o21ai_1 _17508_ (.B1(_11024_),
    .Y(_01351_),
    .A1(net51),
    .A2(net245));
 sg13g2_nand2_1 _17509_ (.Y(_11025_),
    .A(\top_ihp.oisc.regs[34][13] ),
    .B(net244));
 sg13g2_o21ai_1 _17510_ (.B1(_11025_),
    .Y(_01352_),
    .A1(net278),
    .A2(net245));
 sg13g2_nand2_1 _17511_ (.Y(_11026_),
    .A(\top_ihp.oisc.regs[34][14] ),
    .B(net244));
 sg13g2_o21ai_1 _17512_ (.B1(_11026_),
    .Y(_01353_),
    .A1(net277),
    .A2(_11021_));
 sg13g2_mux2_1 _17513_ (.A0(net399),
    .A1(_00336_),
    .S(net246),
    .X(_01354_));
 sg13g2_nand2_1 _17514_ (.Y(_11027_),
    .A(\top_ihp.oisc.regs[34][16] ),
    .B(net244));
 sg13g2_o21ai_1 _17515_ (.B1(_11027_),
    .Y(_01355_),
    .A1(net140),
    .A2(net245));
 sg13g2_nand2_1 _17516_ (.Y(_11028_),
    .A(\top_ihp.oisc.regs[34][17] ),
    .B(_11022_));
 sg13g2_o21ai_1 _17517_ (.B1(_11028_),
    .Y(_01356_),
    .A1(net406),
    .A2(net245));
 sg13g2_nand2_1 _17518_ (.Y(_11029_),
    .A(\top_ihp.oisc.regs[34][18] ),
    .B(_11022_));
 sg13g2_o21ai_1 _17519_ (.B1(_11029_),
    .Y(_01357_),
    .A1(net275),
    .A2(_11021_));
 sg13g2_nand2_1 _17520_ (.Y(_11030_),
    .A(\top_ihp.oisc.regs[34][19] ),
    .B(net244));
 sg13g2_o21ai_1 _17521_ (.B1(_11030_),
    .Y(_01358_),
    .A1(net60),
    .A2(net245));
 sg13g2_buf_2 _17522_ (.A(net388),
    .X(_11031_));
 sg13g2_nand2_1 _17523_ (.Y(_11032_),
    .A(\top_ihp.oisc.regs[34][1] ),
    .B(net243));
 sg13g2_o21ai_1 _17524_ (.B1(_11032_),
    .Y(_01359_),
    .A1(net120),
    .A2(net245));
 sg13g2_buf_1 _17525_ (.A(net388),
    .X(_11033_));
 sg13g2_nand2_1 _17526_ (.Y(_11034_),
    .A(\top_ihp.oisc.regs[34][20] ),
    .B(_11031_));
 sg13g2_o21ai_1 _17527_ (.B1(_11034_),
    .Y(_01360_),
    .A1(net138),
    .A2(_11033_));
 sg13g2_nand2_1 _17528_ (.Y(_11035_),
    .A(\top_ihp.oisc.regs[34][21] ),
    .B(net243));
 sg13g2_o21ai_1 _17529_ (.B1(_11035_),
    .Y(_01361_),
    .A1(net137),
    .A2(_11033_));
 sg13g2_nand2_1 _17530_ (.Y(_11036_),
    .A(\top_ihp.oisc.regs[34][22] ),
    .B(net243));
 sg13g2_o21ai_1 _17531_ (.B1(_11036_),
    .Y(_01362_),
    .A1(net272),
    .A2(net242));
 sg13g2_nand2_1 _17532_ (.Y(_11037_),
    .A(\top_ihp.oisc.regs[34][23] ),
    .B(net243));
 sg13g2_o21ai_1 _17533_ (.B1(_11037_),
    .Y(_01363_),
    .A1(net271),
    .A2(net242));
 sg13g2_mux2_1 _17534_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[34][24] ),
    .S(net246),
    .X(_01364_));
 sg13g2_nand2_1 _17535_ (.Y(_11038_),
    .A(\top_ihp.oisc.regs[34][25] ),
    .B(net243));
 sg13g2_o21ai_1 _17536_ (.B1(_11038_),
    .Y(_01365_),
    .A1(net59),
    .A2(net242));
 sg13g2_nand2_1 _17537_ (.Y(_11039_),
    .A(\top_ihp.oisc.regs[34][26] ),
    .B(net243));
 sg13g2_o21ai_1 _17538_ (.B1(_11039_),
    .Y(_01366_),
    .A1(net402),
    .A2(net242));
 sg13g2_mux2_1 _17539_ (.A0(_10449_),
    .A1(_00337_),
    .S(net246),
    .X(_01367_));
 sg13g2_nand2_1 _17540_ (.Y(_11040_),
    .A(\top_ihp.oisc.regs[34][28] ),
    .B(_11031_));
 sg13g2_o21ai_1 _17541_ (.B1(_11040_),
    .Y(_01368_),
    .A1(net29),
    .A2(net242));
 sg13g2_nand2_1 _17542_ (.Y(_11041_),
    .A(\top_ihp.oisc.regs[34][29] ),
    .B(net243));
 sg13g2_o21ai_1 _17543_ (.B1(_11041_),
    .Y(_01369_),
    .A1(net269),
    .A2(net242));
 sg13g2_nand2_1 _17544_ (.Y(_11042_),
    .A(\top_ihp.oisc.regs[34][2] ),
    .B(net243));
 sg13g2_o21ai_1 _17545_ (.B1(_11042_),
    .Y(_01370_),
    .A1(net136),
    .A2(net242));
 sg13g2_nand2_1 _17546_ (.Y(_11043_),
    .A(\top_ihp.oisc.regs[34][30] ),
    .B(net388));
 sg13g2_o21ai_1 _17547_ (.B1(_11043_),
    .Y(_01371_),
    .A1(net58),
    .A2(net242));
 sg13g2_inv_1 _17548_ (.Y(_11044_),
    .A(\top_ihp.oisc.regs[34][31] ));
 sg13g2_nor2_1 _17549_ (.A(net821),
    .B(_11019_),
    .Y(_11045_));
 sg13g2_a22oi_1 _17550_ (.Y(_01372_),
    .B1(_11045_),
    .B2(net129),
    .A2(net245),
    .A1(_11044_));
 sg13g2_mux2_1 _17551_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[34][3] ),
    .S(_11020_),
    .X(_01373_));
 sg13g2_mux2_1 _17552_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[34][4] ),
    .S(net246),
    .X(_01374_));
 sg13g2_mux2_1 _17553_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[34][5] ),
    .S(net246),
    .X(_01375_));
 sg13g2_mux2_1 _17554_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[34][6] ),
    .S(net244),
    .X(_01376_));
 sg13g2_nand2_1 _17555_ (.Y(_11046_),
    .A(\top_ihp.oisc.regs[34][7] ),
    .B(net388));
 sg13g2_o21ai_1 _17556_ (.B1(_11046_),
    .Y(_01377_),
    .A1(net401),
    .A2(net246));
 sg13g2_nand2_1 _17557_ (.Y(_11047_),
    .A(\top_ihp.oisc.regs[34][8] ),
    .B(net388));
 sg13g2_o21ai_1 _17558_ (.B1(_11047_),
    .Y(_01378_),
    .A1(net266),
    .A2(net246));
 sg13g2_mux2_1 _17559_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[34][9] ),
    .S(net244),
    .X(_01379_));
 sg13g2_and2_1 _17560_ (.A(_10747_),
    .B(_10987_),
    .X(_11048_));
 sg13g2_buf_1 _17561_ (.A(_11048_),
    .X(_11049_));
 sg13g2_buf_2 _17562_ (.A(_11049_),
    .X(_11050_));
 sg13g2_mux2_1 _17563_ (.A0(\top_ihp.oisc.regs[35][0] ),
    .A1(net119),
    .S(net241),
    .X(_01380_));
 sg13g2_mux2_1 _17564_ (.A0(\top_ihp.oisc.regs[35][10] ),
    .A1(net130),
    .S(net241),
    .X(_01381_));
 sg13g2_mux2_1 _17565_ (.A0(_00338_),
    .A1(_10050_),
    .S(net241),
    .X(_01382_));
 sg13g2_nand2_1 _17566_ (.Y(_11051_),
    .A(_10747_),
    .B(_10987_));
 sg13g2_buf_1 _17567_ (.A(_11051_),
    .X(_11052_));
 sg13g2_buf_2 _17568_ (.A(_11052_),
    .X(_11053_));
 sg13g2_buf_2 _17569_ (.A(_11052_),
    .X(_11054_));
 sg13g2_nand2_1 _17570_ (.Y(_11055_),
    .A(\top_ihp.oisc.regs[35][12] ),
    .B(net239));
 sg13g2_o21ai_1 _17571_ (.B1(_11055_),
    .Y(_01383_),
    .A1(net51),
    .A2(net240));
 sg13g2_nand2_1 _17572_ (.Y(_11056_),
    .A(\top_ihp.oisc.regs[35][13] ),
    .B(net239));
 sg13g2_o21ai_1 _17573_ (.B1(_11056_),
    .Y(_01384_),
    .A1(net278),
    .A2(net240));
 sg13g2_nand2_1 _17574_ (.Y(_11057_),
    .A(\top_ihp.oisc.regs[35][14] ),
    .B(net239));
 sg13g2_o21ai_1 _17575_ (.B1(_11057_),
    .Y(_01385_),
    .A1(net277),
    .A2(_11053_));
 sg13g2_nand2_1 _17576_ (.Y(_11058_),
    .A(\top_ihp.oisc.regs[35][15] ),
    .B(_11054_));
 sg13g2_o21ai_1 _17577_ (.B1(_11058_),
    .Y(_01386_),
    .A1(net407),
    .A2(net240));
 sg13g2_nand2_1 _17578_ (.Y(_11059_),
    .A(\top_ihp.oisc.regs[35][16] ),
    .B(_11054_));
 sg13g2_o21ai_1 _17579_ (.B1(_11059_),
    .Y(_01387_),
    .A1(net140),
    .A2(_11053_));
 sg13g2_nand2_1 _17580_ (.Y(_11060_),
    .A(\top_ihp.oisc.regs[35][17] ),
    .B(net239));
 sg13g2_o21ai_1 _17581_ (.B1(_11060_),
    .Y(_01388_),
    .A1(net406),
    .A2(net240));
 sg13g2_nand2_1 _17582_ (.Y(_11061_),
    .A(\top_ihp.oisc.regs[35][18] ),
    .B(net239));
 sg13g2_o21ai_1 _17583_ (.B1(_11061_),
    .Y(_01389_),
    .A1(net275),
    .A2(net240));
 sg13g2_mux2_1 _17584_ (.A0(\top_ihp.oisc.regs[35][19] ),
    .A1(net254),
    .S(net241),
    .X(_01390_));
 sg13g2_nand2_1 _17585_ (.Y(_11062_),
    .A(\top_ihp.oisc.regs[35][1] ),
    .B(net239));
 sg13g2_o21ai_1 _17586_ (.B1(_11062_),
    .Y(_01391_),
    .A1(net120),
    .A2(net240));
 sg13g2_nand2_1 _17587_ (.Y(_11063_),
    .A(\top_ihp.oisc.regs[35][20] ),
    .B(net239));
 sg13g2_o21ai_1 _17588_ (.B1(_11063_),
    .Y(_01392_),
    .A1(net138),
    .A2(net240));
 sg13g2_nand2_1 _17589_ (.Y(_11064_),
    .A(\top_ihp.oisc.regs[35][21] ),
    .B(net239));
 sg13g2_o21ai_1 _17590_ (.B1(_11064_),
    .Y(_01393_),
    .A1(net137),
    .A2(net240));
 sg13g2_buf_1 _17591_ (.A(_11052_),
    .X(_11065_));
 sg13g2_buf_1 _17592_ (.A(_11052_),
    .X(_11066_));
 sg13g2_nand2_1 _17593_ (.Y(_11067_),
    .A(\top_ihp.oisc.regs[35][22] ),
    .B(net237));
 sg13g2_o21ai_1 _17594_ (.B1(_11067_),
    .Y(_01394_),
    .A1(net272),
    .A2(net238));
 sg13g2_nand2_1 _17595_ (.Y(_11068_),
    .A(\top_ihp.oisc.regs[35][23] ),
    .B(net237));
 sg13g2_o21ai_1 _17596_ (.B1(_11068_),
    .Y(_01395_),
    .A1(net271),
    .A2(net238));
 sg13g2_mux2_1 _17597_ (.A0(\top_ihp.oisc.regs[35][24] ),
    .A1(net400),
    .S(net241),
    .X(_01396_));
 sg13g2_nand2_1 _17598_ (.Y(_11069_),
    .A(\top_ihp.oisc.regs[35][25] ),
    .B(net237));
 sg13g2_o21ai_1 _17599_ (.B1(_11069_),
    .Y(_01397_),
    .A1(net124),
    .A2(net238));
 sg13g2_nand2_1 _17600_ (.Y(_11070_),
    .A(\top_ihp.oisc.regs[35][26] ),
    .B(net237));
 sg13g2_o21ai_1 _17601_ (.B1(_11070_),
    .Y(_01398_),
    .A1(net402),
    .A2(net238));
 sg13g2_mux2_1 _17602_ (.A0(\top_ihp.oisc.regs[35][27] ),
    .A1(net117),
    .S(net241),
    .X(_01399_));
 sg13g2_nand2_1 _17603_ (.Y(_11071_),
    .A(\top_ihp.oisc.regs[35][28] ),
    .B(_11066_));
 sg13g2_o21ai_1 _17604_ (.B1(_11071_),
    .Y(_01400_),
    .A1(net29),
    .A2(_11065_));
 sg13g2_nand2_1 _17605_ (.Y(_11072_),
    .A(\top_ihp.oisc.regs[35][29] ),
    .B(net237));
 sg13g2_o21ai_1 _17606_ (.B1(_11072_),
    .Y(_01401_),
    .A1(net269),
    .A2(net238));
 sg13g2_nand2_1 _17607_ (.Y(_11073_),
    .A(\top_ihp.oisc.regs[35][2] ),
    .B(net237));
 sg13g2_o21ai_1 _17608_ (.B1(_11073_),
    .Y(_01402_),
    .A1(net136),
    .A2(_11065_));
 sg13g2_nand2_1 _17609_ (.Y(_11074_),
    .A(\top_ihp.oisc.regs[35][30] ),
    .B(net237));
 sg13g2_o21ai_1 _17610_ (.B1(_11074_),
    .Y(_01403_),
    .A1(net58),
    .A2(net238));
 sg13g2_mux2_1 _17611_ (.A0(_00339_),
    .A1(net265),
    .S(net241),
    .X(_01404_));
 sg13g2_mux2_1 _17612_ (.A0(\top_ihp.oisc.regs[35][3] ),
    .A1(net128),
    .S(net241),
    .X(_01405_));
 sg13g2_mux2_1 _17613_ (.A0(\top_ihp.oisc.regs[35][4] ),
    .A1(_10740_),
    .S(_11050_),
    .X(_01406_));
 sg13g2_mux2_1 _17614_ (.A0(\top_ihp.oisc.regs[35][5] ),
    .A1(net264),
    .S(_11050_),
    .X(_01407_));
 sg13g2_mux2_1 _17615_ (.A0(\top_ihp.oisc.regs[35][6] ),
    .A1(net126),
    .S(_11049_),
    .X(_01408_));
 sg13g2_nand2_1 _17616_ (.Y(_11075_),
    .A(\top_ihp.oisc.regs[35][7] ),
    .B(_11066_));
 sg13g2_o21ai_1 _17617_ (.B1(_11075_),
    .Y(_01409_),
    .A1(net401),
    .A2(net238));
 sg13g2_nand2_1 _17618_ (.Y(_11076_),
    .A(\top_ihp.oisc.regs[35][8] ),
    .B(net237));
 sg13g2_o21ai_1 _17619_ (.B1(_11076_),
    .Y(_01410_),
    .A1(net266),
    .A2(net238));
 sg13g2_mux2_1 _17620_ (.A0(\top_ihp.oisc.regs[35][9] ),
    .A1(net125),
    .S(_11049_),
    .X(_01411_));
 sg13g2_nand2_1 _17621_ (.Y(_11077_),
    .A(_09913_),
    .B(_10690_));
 sg13g2_nor2_1 _17622_ (.A(net1008),
    .B(_09905_),
    .Y(_11078_));
 sg13g2_or3_1 _17623_ (.A(_09910_),
    .B(_11077_),
    .C(_11078_),
    .X(_11079_));
 sg13g2_buf_2 _17624_ (.A(_11079_),
    .X(_11080_));
 sg13g2_nor2_2 _17625_ (.A(_10984_),
    .B(_11080_),
    .Y(_11081_));
 sg13g2_nand2_1 _17626_ (.Y(_11082_),
    .A(_09939_),
    .B(_11081_));
 sg13g2_buf_1 _17627_ (.A(_11082_),
    .X(_11083_));
 sg13g2_buf_2 _17628_ (.A(net657),
    .X(_11084_));
 sg13g2_mux2_1 _17629_ (.A0(net64),
    .A1(\top_ihp.oisc.regs[36][0] ),
    .S(_11084_),
    .X(_01412_));
 sg13g2_mux2_1 _17630_ (.A0(_10010_),
    .A1(\top_ihp.oisc.regs[36][10] ),
    .S(_11084_),
    .X(_01413_));
 sg13g2_buf_2 _17631_ (.A(net657),
    .X(_11085_));
 sg13g2_buf_2 _17632_ (.A(net657),
    .X(_11086_));
 sg13g2_nand2_1 _17633_ (.Y(_11087_),
    .A(\top_ihp.oisc.regs[36][11] ),
    .B(net560));
 sg13g2_o21ai_1 _17634_ (.B1(_11087_),
    .Y(_01414_),
    .A1(net49),
    .A2(net561));
 sg13g2_nand2_1 _17635_ (.Y(_11088_),
    .A(\top_ihp.oisc.regs[36][12] ),
    .B(net560));
 sg13g2_o21ai_1 _17636_ (.B1(_11088_),
    .Y(_01415_),
    .A1(net51),
    .A2(net561));
 sg13g2_buf_1 _17637_ (.A(net261),
    .X(_11089_));
 sg13g2_nand2_1 _17638_ (.Y(_11090_),
    .A(\top_ihp.oisc.regs[36][13] ),
    .B(net560));
 sg13g2_o21ai_1 _17639_ (.B1(_11090_),
    .Y(_01416_),
    .A1(net115),
    .A2(net561));
 sg13g2_buf_1 _17640_ (.A(net260),
    .X(_11091_));
 sg13g2_nand2_1 _17641_ (.Y(_11092_),
    .A(\top_ihp.oisc.regs[36][14] ),
    .B(net560));
 sg13g2_o21ai_1 _17642_ (.B1(_11092_),
    .Y(_01417_),
    .A1(net114),
    .A2(net561));
 sg13g2_nand2_1 _17643_ (.Y(_11093_),
    .A(\top_ihp.oisc.regs[36][15] ),
    .B(net560));
 sg13g2_o21ai_1 _17644_ (.B1(_11093_),
    .Y(_01418_),
    .A1(net407),
    .A2(net561));
 sg13g2_buf_1 _17645_ (.A(net276),
    .X(_11094_));
 sg13g2_nand2_1 _17646_ (.Y(_11095_),
    .A(\top_ihp.oisc.regs[36][16] ),
    .B(_11086_));
 sg13g2_o21ai_1 _17647_ (.B1(_11095_),
    .Y(_01419_),
    .A1(net113),
    .A2(net561));
 sg13g2_buf_1 _17648_ (.A(net398),
    .X(_11096_));
 sg13g2_nand2_1 _17649_ (.Y(_11097_),
    .A(\top_ihp.oisc.regs[36][17] ),
    .B(net560));
 sg13g2_o21ai_1 _17650_ (.B1(_11097_),
    .Y(_01420_),
    .A1(net236),
    .A2(_11085_));
 sg13g2_buf_1 _17651_ (.A(net259),
    .X(_11098_));
 sg13g2_nand2_1 _17652_ (.Y(_11099_),
    .A(\top_ihp.oisc.regs[36][18] ),
    .B(_11086_));
 sg13g2_o21ai_1 _17653_ (.B1(_11099_),
    .Y(_01421_),
    .A1(net112),
    .A2(net561));
 sg13g2_mux2_1 _17654_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[36][19] ),
    .S(net562),
    .X(_01422_));
 sg13g2_buf_2 _17655_ (.A(net657),
    .X(_11100_));
 sg13g2_nand2_1 _17656_ (.Y(_11101_),
    .A(\top_ihp.oisc.regs[36][1] ),
    .B(_11100_));
 sg13g2_o21ai_1 _17657_ (.B1(_11101_),
    .Y(_01423_),
    .A1(net120),
    .A2(net561));
 sg13g2_buf_1 _17658_ (.A(_10804_),
    .X(_11102_));
 sg13g2_nand2_1 _17659_ (.Y(_11103_),
    .A(\top_ihp.oisc.regs[36][20] ),
    .B(net559));
 sg13g2_o21ai_1 _17660_ (.B1(_11103_),
    .Y(_01424_),
    .A1(net48),
    .A2(_11085_));
 sg13g2_buf_1 _17661_ (.A(net273),
    .X(_11104_));
 sg13g2_buf_1 _17662_ (.A(net657),
    .X(_11105_));
 sg13g2_nand2_1 _17663_ (.Y(_11106_),
    .A(\top_ihp.oisc.regs[36][21] ),
    .B(_11100_));
 sg13g2_o21ai_1 _17664_ (.B1(_11106_),
    .Y(_01425_),
    .A1(net111),
    .A2(net558));
 sg13g2_buf_2 _17665_ (.A(_10807_),
    .X(_11107_));
 sg13g2_nand2_1 _17666_ (.Y(_11108_),
    .A(\top_ihp.oisc.regs[36][22] ),
    .B(net559));
 sg13g2_o21ai_1 _17667_ (.B1(_11108_),
    .Y(_01426_),
    .A1(net110),
    .A2(net558));
 sg13g2_buf_1 _17668_ (.A(_10808_),
    .X(_11109_));
 sg13g2_nand2_1 _17669_ (.Y(_11110_),
    .A(\top_ihp.oisc.regs[36][23] ),
    .B(net559));
 sg13g2_o21ai_1 _17670_ (.B1(_11110_),
    .Y(_01427_),
    .A1(net109),
    .A2(net558));
 sg13g2_mux2_1 _17671_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[36][24] ),
    .S(net562),
    .X(_01428_));
 sg13g2_nand2_1 _17672_ (.Y(_11111_),
    .A(\top_ihp.oisc.regs[36][25] ),
    .B(net559));
 sg13g2_o21ai_1 _17673_ (.B1(_11111_),
    .Y(_01429_),
    .A1(net124),
    .A2(net558));
 sg13g2_buf_2 _17674_ (.A(net397),
    .X(_11112_));
 sg13g2_nand2_1 _17675_ (.Y(_11113_),
    .A(\top_ihp.oisc.regs[36][26] ),
    .B(net559));
 sg13g2_o21ai_1 _17676_ (.B1(_11113_),
    .Y(_01430_),
    .A1(net235),
    .A2(_11105_));
 sg13g2_mux2_1 _17677_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[36][27] ),
    .S(net562),
    .X(_01431_));
 sg13g2_nand2_1 _17678_ (.Y(_11114_),
    .A(\top_ihp.oisc.regs[36][28] ),
    .B(net559));
 sg13g2_o21ai_1 _17679_ (.B1(_11114_),
    .Y(_01432_),
    .A1(net29),
    .A2(net558));
 sg13g2_buf_1 _17680_ (.A(net256),
    .X(_11115_));
 sg13g2_nand2_1 _17681_ (.Y(_11116_),
    .A(\top_ihp.oisc.regs[36][29] ),
    .B(net559));
 sg13g2_o21ai_1 _17682_ (.B1(_11116_),
    .Y(_01433_),
    .A1(net108),
    .A2(_11105_));
 sg13g2_nand2_1 _17683_ (.Y(_11117_),
    .A(\top_ihp.oisc.regs[36][2] ),
    .B(net559));
 sg13g2_o21ai_1 _17684_ (.B1(_11117_),
    .Y(_01434_),
    .A1(net136),
    .A2(net558));
 sg13g2_nand2_1 _17685_ (.Y(_11118_),
    .A(\top_ihp.oisc.regs[36][30] ),
    .B(net657));
 sg13g2_o21ai_1 _17686_ (.B1(_11118_),
    .Y(_01435_),
    .A1(net58),
    .A2(net558));
 sg13g2_nand2_1 _17687_ (.Y(_11119_),
    .A(\top_ihp.oisc.regs[36][31] ),
    .B(_11083_));
 sg13g2_o21ai_1 _17688_ (.B1(_11119_),
    .Y(_01436_),
    .A1(net268),
    .A2(net558));
 sg13g2_mux2_1 _17689_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[36][3] ),
    .S(net562),
    .X(_01437_));
 sg13g2_mux2_1 _17690_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[36][4] ),
    .S(net562),
    .X(_01438_));
 sg13g2_mux2_1 _17691_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[36][5] ),
    .S(net562),
    .X(_01439_));
 sg13g2_mux2_1 _17692_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[36][6] ),
    .S(net560),
    .X(_01440_));
 sg13g2_buf_1 _17693_ (.A(_10818_),
    .X(_11120_));
 sg13g2_nand2_1 _17694_ (.Y(_11121_),
    .A(\top_ihp.oisc.regs[36][7] ),
    .B(net657));
 sg13g2_o21ai_1 _17695_ (.B1(_11121_),
    .Y(_01441_),
    .A1(net234),
    .A2(net562));
 sg13g2_buf_2 _17696_ (.A(_10819_),
    .X(_11122_));
 sg13g2_nand2_1 _17697_ (.Y(_11123_),
    .A(\top_ihp.oisc.regs[36][8] ),
    .B(net657));
 sg13g2_o21ai_1 _17698_ (.B1(_11123_),
    .Y(_01442_),
    .A1(net107),
    .A2(net562));
 sg13g2_mux2_1 _17699_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[36][9] ),
    .S(net560),
    .X(_01443_));
 sg13g2_nand2_1 _17700_ (.Y(_11124_),
    .A(_10822_),
    .B(_11081_));
 sg13g2_buf_2 _17701_ (.A(_11124_),
    .X(_11125_));
 sg13g2_buf_2 _17702_ (.A(_11125_),
    .X(_11126_));
 sg13g2_mux2_1 _17703_ (.A0(net64),
    .A1(\top_ihp.oisc.regs[37][0] ),
    .S(net557),
    .X(_01444_));
 sg13g2_mux2_1 _17704_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[37][10] ),
    .S(net557),
    .X(_01445_));
 sg13g2_buf_2 _17705_ (.A(_11125_),
    .X(_11127_));
 sg13g2_buf_1 _17706_ (.A(_11125_),
    .X(_11128_));
 sg13g2_nand2_1 _17707_ (.Y(_11129_),
    .A(\top_ihp.oisc.regs[37][11] ),
    .B(net555));
 sg13g2_o21ai_1 _17708_ (.B1(_11129_),
    .Y(_01446_),
    .A1(net49),
    .A2(net556));
 sg13g2_nand2_1 _17709_ (.Y(_11130_),
    .A(\top_ihp.oisc.regs[37][12] ),
    .B(_11128_));
 sg13g2_o21ai_1 _17710_ (.B1(_11130_),
    .Y(_01447_),
    .A1(net51),
    .A2(net556));
 sg13g2_nand2_1 _17711_ (.Y(_11131_),
    .A(\top_ihp.oisc.regs[37][13] ),
    .B(net555));
 sg13g2_o21ai_1 _17712_ (.B1(_11131_),
    .Y(_01448_),
    .A1(_11089_),
    .A2(net556));
 sg13g2_nand2_1 _17713_ (.Y(_11132_),
    .A(\top_ihp.oisc.regs[37][14] ),
    .B(_11128_));
 sg13g2_o21ai_1 _17714_ (.B1(_11132_),
    .Y(_01449_),
    .A1(net114),
    .A2(_11127_));
 sg13g2_mux2_1 _17715_ (.A0(_10169_),
    .A1(\top_ihp.oisc.regs[37][15] ),
    .S(net557),
    .X(_01450_));
 sg13g2_nand2_1 _17716_ (.Y(_11133_),
    .A(\top_ihp.oisc.regs[37][16] ),
    .B(net555));
 sg13g2_o21ai_1 _17717_ (.B1(_11133_),
    .Y(_01451_),
    .A1(_11094_),
    .A2(net556));
 sg13g2_nand2_1 _17718_ (.Y(_11134_),
    .A(\top_ihp.oisc.regs[37][17] ),
    .B(net555));
 sg13g2_o21ai_1 _17719_ (.B1(_11134_),
    .Y(_01452_),
    .A1(net236),
    .A2(net556));
 sg13g2_nand2_1 _17720_ (.Y(_11135_),
    .A(\top_ihp.oisc.regs[37][18] ),
    .B(net555));
 sg13g2_o21ai_1 _17721_ (.B1(_11135_),
    .Y(_01453_),
    .A1(_11098_),
    .A2(_11127_));
 sg13g2_mux2_1 _17722_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[37][19] ),
    .S(net557),
    .X(_01454_));
 sg13g2_nand2_1 _17723_ (.Y(_11136_),
    .A(\top_ihp.oisc.regs[37][1] ),
    .B(net555));
 sg13g2_o21ai_1 _17724_ (.B1(_11136_),
    .Y(_01455_),
    .A1(net120),
    .A2(net556));
 sg13g2_buf_1 _17725_ (.A(_11125_),
    .X(_11137_));
 sg13g2_nand2_1 _17726_ (.Y(_11138_),
    .A(\top_ihp.oisc.regs[37][20] ),
    .B(net554));
 sg13g2_o21ai_1 _17727_ (.B1(_11138_),
    .Y(_01456_),
    .A1(net48),
    .A2(net556));
 sg13g2_nand2_1 _17728_ (.Y(_11139_),
    .A(\top_ihp.oisc.regs[37][21] ),
    .B(_11137_));
 sg13g2_o21ai_1 _17729_ (.B1(_11139_),
    .Y(_01457_),
    .A1(net111),
    .A2(net556));
 sg13g2_buf_1 _17730_ (.A(_11125_),
    .X(_11140_));
 sg13g2_nand2_1 _17731_ (.Y(_11141_),
    .A(\top_ihp.oisc.regs[37][22] ),
    .B(net554));
 sg13g2_o21ai_1 _17732_ (.B1(_11141_),
    .Y(_01458_),
    .A1(net110),
    .A2(net553));
 sg13g2_nand2_1 _17733_ (.Y(_11142_),
    .A(\top_ihp.oisc.regs[37][23] ),
    .B(_11137_));
 sg13g2_o21ai_1 _17734_ (.B1(_11142_),
    .Y(_01459_),
    .A1(net109),
    .A2(_11140_));
 sg13g2_mux2_1 _17735_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[37][24] ),
    .S(net557),
    .X(_01460_));
 sg13g2_nand2_1 _17736_ (.Y(_11143_),
    .A(\top_ihp.oisc.regs[37][25] ),
    .B(net554));
 sg13g2_o21ai_1 _17737_ (.B1(_11143_),
    .Y(_01461_),
    .A1(net124),
    .A2(net553));
 sg13g2_nand2_1 _17738_ (.Y(_11144_),
    .A(\top_ihp.oisc.regs[37][26] ),
    .B(net554));
 sg13g2_o21ai_1 _17739_ (.B1(_11144_),
    .Y(_01462_),
    .A1(net235),
    .A2(net553));
 sg13g2_mux2_1 _17740_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[37][27] ),
    .S(net557),
    .X(_01463_));
 sg13g2_nand2_1 _17741_ (.Y(_11145_),
    .A(\top_ihp.oisc.regs[37][28] ),
    .B(net554));
 sg13g2_o21ai_1 _17742_ (.B1(_11145_),
    .Y(_01464_),
    .A1(net29),
    .A2(net553));
 sg13g2_nand2_1 _17743_ (.Y(_11146_),
    .A(\top_ihp.oisc.regs[37][29] ),
    .B(net554));
 sg13g2_o21ai_1 _17744_ (.B1(_11146_),
    .Y(_01465_),
    .A1(net108),
    .A2(_11140_));
 sg13g2_buf_1 _17745_ (.A(net122),
    .X(_11147_));
 sg13g2_nand2_1 _17746_ (.Y(_11148_),
    .A(\top_ihp.oisc.regs[37][2] ),
    .B(net554));
 sg13g2_o21ai_1 _17747_ (.B1(_11148_),
    .Y(_01466_),
    .A1(net47),
    .A2(net553));
 sg13g2_buf_8 _17748_ (.A(net53),
    .X(_11149_));
 sg13g2_nand2_1 _17749_ (.Y(_11150_),
    .A(\top_ihp.oisc.regs[37][30] ),
    .B(net554));
 sg13g2_o21ai_1 _17750_ (.B1(_11150_),
    .Y(_01467_),
    .A1(net28),
    .A2(net553));
 sg13g2_buf_1 _17751_ (.A(_10737_),
    .X(_11151_));
 sg13g2_nand2_1 _17752_ (.Y(_11152_),
    .A(\top_ihp.oisc.regs[37][31] ),
    .B(_11125_));
 sg13g2_o21ai_1 _17753_ (.B1(_11152_),
    .Y(_01468_),
    .A1(net106),
    .A2(net553));
 sg13g2_mux2_1 _17754_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[37][3] ),
    .S(_11126_),
    .X(_01469_));
 sg13g2_mux2_1 _17755_ (.A0(net56),
    .A1(\top_ihp.oisc.regs[37][4] ),
    .S(net557),
    .X(_01470_));
 sg13g2_mux2_1 _17756_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[37][5] ),
    .S(_11126_),
    .X(_01471_));
 sg13g2_mux2_1 _17757_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[37][6] ),
    .S(net555),
    .X(_01472_));
 sg13g2_nand2_1 _17758_ (.Y(_11153_),
    .A(\top_ihp.oisc.regs[37][7] ),
    .B(_11125_));
 sg13g2_o21ai_1 _17759_ (.B1(_11153_),
    .Y(_01473_),
    .A1(net234),
    .A2(net553));
 sg13g2_nand2_1 _17760_ (.Y(_11154_),
    .A(\top_ihp.oisc.regs[37][8] ),
    .B(_11125_));
 sg13g2_o21ai_1 _17761_ (.B1(_11154_),
    .Y(_01474_),
    .A1(_11122_),
    .A2(net557));
 sg13g2_mux2_1 _17762_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[37][9] ),
    .S(net555),
    .X(_01475_));
 sg13g2_buf_1 _17763_ (.A(net143),
    .X(_11155_));
 sg13g2_nand2_1 _17764_ (.Y(_11156_),
    .A(net740),
    .B(_11081_));
 sg13g2_buf_1 _17765_ (.A(_11156_),
    .X(_11157_));
 sg13g2_buf_2 _17766_ (.A(net656),
    .X(_11158_));
 sg13g2_mux2_1 _17767_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[38][0] ),
    .S(_11158_),
    .X(_01476_));
 sg13g2_mux2_1 _17768_ (.A0(net63),
    .A1(\top_ihp.oisc.regs[38][10] ),
    .S(net552),
    .X(_01477_));
 sg13g2_buf_1 _17769_ (.A(net656),
    .X(_11159_));
 sg13g2_buf_1 _17770_ (.A(_11156_),
    .X(_11160_));
 sg13g2_nand2_1 _17771_ (.Y(_11161_),
    .A(\top_ihp.oisc.regs[38][11] ),
    .B(net655));
 sg13g2_o21ai_1 _17772_ (.B1(_11161_),
    .Y(_01478_),
    .A1(_10991_),
    .A2(net551));
 sg13g2_nand2_1 _17773_ (.Y(_11162_),
    .A(\top_ihp.oisc.regs[38][12] ),
    .B(net655));
 sg13g2_o21ai_1 _17774_ (.B1(_11162_),
    .Y(_01479_),
    .A1(net51),
    .A2(net551));
 sg13g2_nand2_1 _17775_ (.Y(_11163_),
    .A(\top_ihp.oisc.regs[38][13] ),
    .B(net655));
 sg13g2_o21ai_1 _17776_ (.B1(_11163_),
    .Y(_01480_),
    .A1(net115),
    .A2(net551));
 sg13g2_nand2_1 _17777_ (.Y(_11164_),
    .A(\top_ihp.oisc.regs[38][14] ),
    .B(net655));
 sg13g2_o21ai_1 _17778_ (.B1(_11164_),
    .Y(_01481_),
    .A1(_11091_),
    .A2(net551));
 sg13g2_buf_1 _17779_ (.A(net399),
    .X(_11165_));
 sg13g2_nand2_1 _17780_ (.Y(_11166_),
    .A(\top_ihp.oisc.regs[38][15] ),
    .B(net655));
 sg13g2_o21ai_1 _17781_ (.B1(_11166_),
    .Y(_01482_),
    .A1(net233),
    .A2(net551));
 sg13g2_nand2_1 _17782_ (.Y(_11167_),
    .A(\top_ihp.oisc.regs[38][16] ),
    .B(_11160_));
 sg13g2_o21ai_1 _17783_ (.B1(_11167_),
    .Y(_01483_),
    .A1(net113),
    .A2(net551));
 sg13g2_nand2_1 _17784_ (.Y(_11168_),
    .A(\top_ihp.oisc.regs[38][17] ),
    .B(_11160_));
 sg13g2_o21ai_1 _17785_ (.B1(_11168_),
    .Y(_01484_),
    .A1(net236),
    .A2(_11159_));
 sg13g2_nand2_1 _17786_ (.Y(_11169_),
    .A(\top_ihp.oisc.regs[38][18] ),
    .B(net655));
 sg13g2_o21ai_1 _17787_ (.B1(_11169_),
    .Y(_01485_),
    .A1(net112),
    .A2(net551));
 sg13g2_buf_1 _17788_ (.A(_11157_),
    .X(_11170_));
 sg13g2_nand2_1 _17789_ (.Y(_11171_),
    .A(\top_ihp.oisc.regs[38][19] ),
    .B(_11170_));
 sg13g2_o21ai_1 _17790_ (.B1(_11171_),
    .Y(_01486_),
    .A1(net60),
    .A2(net551));
 sg13g2_buf_1 _17791_ (.A(net656),
    .X(_11172_));
 sg13g2_nand2_1 _17792_ (.Y(_11173_),
    .A(\top_ihp.oisc.regs[38][1] ),
    .B(net550));
 sg13g2_o21ai_1 _17793_ (.B1(_11173_),
    .Y(_01487_),
    .A1(net120),
    .A2(net549));
 sg13g2_nand2_1 _17794_ (.Y(_11174_),
    .A(\top_ihp.oisc.regs[38][20] ),
    .B(net550));
 sg13g2_o21ai_1 _17795_ (.B1(_11174_),
    .Y(_01488_),
    .A1(net48),
    .A2(net549));
 sg13g2_nand2_1 _17796_ (.Y(_11175_),
    .A(\top_ihp.oisc.regs[38][21] ),
    .B(net550));
 sg13g2_o21ai_1 _17797_ (.B1(_11175_),
    .Y(_01489_),
    .A1(net111),
    .A2(net549));
 sg13g2_nand2_1 _17798_ (.Y(_11176_),
    .A(\top_ihp.oisc.regs[38][22] ),
    .B(net550));
 sg13g2_o21ai_1 _17799_ (.B1(_11176_),
    .Y(_01490_),
    .A1(net110),
    .A2(_11172_));
 sg13g2_nand2_1 _17800_ (.Y(_11177_),
    .A(\top_ihp.oisc.regs[38][23] ),
    .B(net550));
 sg13g2_o21ai_1 _17801_ (.B1(_11177_),
    .Y(_01491_),
    .A1(net109),
    .A2(net549));
 sg13g2_mux2_1 _17802_ (.A0(net270),
    .A1(\top_ihp.oisc.regs[38][24] ),
    .S(net552),
    .X(_01492_));
 sg13g2_nand2_1 _17803_ (.Y(_11178_),
    .A(\top_ihp.oisc.regs[38][25] ),
    .B(_11170_));
 sg13g2_o21ai_1 _17804_ (.B1(_11178_),
    .Y(_01493_),
    .A1(net59),
    .A2(net549));
 sg13g2_nand2_1 _17805_ (.Y(_11179_),
    .A(\top_ihp.oisc.regs[38][26] ),
    .B(net550));
 sg13g2_o21ai_1 _17806_ (.B1(_11179_),
    .Y(_01494_),
    .A1(net235),
    .A2(net549));
 sg13g2_nand2_1 _17807_ (.Y(_11180_),
    .A(\top_ihp.oisc.regs[38][27] ),
    .B(net550));
 sg13g2_o21ai_1 _17808_ (.B1(_11180_),
    .Y(_01495_),
    .A1(net31),
    .A2(net549));
 sg13g2_nand2_1 _17809_ (.Y(_11181_),
    .A(\top_ihp.oisc.regs[38][28] ),
    .B(net550));
 sg13g2_o21ai_1 _17810_ (.B1(_11181_),
    .Y(_01496_),
    .A1(net29),
    .A2(net549));
 sg13g2_nand2_1 _17811_ (.Y(_11182_),
    .A(\top_ihp.oisc.regs[38][29] ),
    .B(net656));
 sg13g2_o21ai_1 _17812_ (.B1(_11182_),
    .Y(_01497_),
    .A1(net108),
    .A2(_11172_));
 sg13g2_nand2_1 _17813_ (.Y(_11183_),
    .A(\top_ihp.oisc.regs[38][2] ),
    .B(net656));
 sg13g2_o21ai_1 _17814_ (.B1(_11183_),
    .Y(_01498_),
    .A1(net47),
    .A2(net552));
 sg13g2_nand2_1 _17815_ (.Y(_11184_),
    .A(\top_ihp.oisc.regs[38][30] ),
    .B(net656));
 sg13g2_o21ai_1 _17816_ (.B1(_11184_),
    .Y(_01499_),
    .A1(_11149_),
    .A2(net552));
 sg13g2_inv_1 _17817_ (.Y(_11185_),
    .A(\top_ihp.oisc.regs[38][31] ));
 sg13g2_nor2_1 _17818_ (.A(net821),
    .B(_11157_),
    .Y(_11186_));
 sg13g2_a22oi_1 _17819_ (.Y(_01500_),
    .B1(_11186_),
    .B2(net129),
    .A2(_11159_),
    .A1(_11185_));
 sg13g2_mux2_1 _17820_ (.A0(net57),
    .A1(\top_ihp.oisc.regs[38][3] ),
    .S(_11158_),
    .X(_01501_));
 sg13g2_mux2_1 _17821_ (.A0(_10600_),
    .A1(\top_ihp.oisc.regs[38][4] ),
    .S(net552),
    .X(_01502_));
 sg13g2_mux2_1 _17822_ (.A0(net133),
    .A1(\top_ihp.oisc.regs[38][5] ),
    .S(net552),
    .X(_01503_));
 sg13g2_mux2_1 _17823_ (.A0(net55),
    .A1(\top_ihp.oisc.regs[38][6] ),
    .S(net655),
    .X(_01504_));
 sg13g2_nand2_1 _17824_ (.Y(_11187_),
    .A(\top_ihp.oisc.regs[38][7] ),
    .B(net656));
 sg13g2_o21ai_1 _17825_ (.B1(_11187_),
    .Y(_01505_),
    .A1(net234),
    .A2(net552));
 sg13g2_nand2_1 _17826_ (.Y(_11188_),
    .A(\top_ihp.oisc.regs[38][8] ),
    .B(net656));
 sg13g2_o21ai_1 _17827_ (.B1(_11188_),
    .Y(_01506_),
    .A1(net107),
    .A2(net552));
 sg13g2_mux2_1 _17828_ (.A0(net54),
    .A1(\top_ihp.oisc.regs[38][9] ),
    .S(net655),
    .X(_01507_));
 sg13g2_nand2_1 _17829_ (.Y(_11189_),
    .A(_10747_),
    .B(_11081_));
 sg13g2_buf_1 _17830_ (.A(_11189_),
    .X(_11190_));
 sg13g2_buf_2 _17831_ (.A(net654),
    .X(_11191_));
 sg13g2_mux2_1 _17832_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[39][0] ),
    .S(net548),
    .X(_01508_));
 sg13g2_buf_2 _17833_ (.A(net142),
    .X(_11192_));
 sg13g2_mux2_1 _17834_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[39][10] ),
    .S(net548),
    .X(_01509_));
 sg13g2_buf_1 _17835_ (.A(net654),
    .X(_11193_));
 sg13g2_buf_1 _17836_ (.A(_11190_),
    .X(_11194_));
 sg13g2_nand2_1 _17837_ (.Y(_11195_),
    .A(\top_ihp.oisc.regs[39][11] ),
    .B(net546));
 sg13g2_o21ai_1 _17838_ (.B1(_11195_),
    .Y(_01510_),
    .A1(net49),
    .A2(net547));
 sg13g2_nand2_1 _17839_ (.Y(_11196_),
    .A(\top_ihp.oisc.regs[39][12] ),
    .B(net546));
 sg13g2_o21ai_1 _17840_ (.B1(_11196_),
    .Y(_01511_),
    .A1(net51),
    .A2(net547));
 sg13g2_nand2_1 _17841_ (.Y(_11197_),
    .A(\top_ihp.oisc.regs[39][13] ),
    .B(net546));
 sg13g2_o21ai_1 _17842_ (.B1(_11197_),
    .Y(_01512_),
    .A1(net115),
    .A2(net547));
 sg13g2_nand2_1 _17843_ (.Y(_11198_),
    .A(\top_ihp.oisc.regs[39][14] ),
    .B(_11194_));
 sg13g2_o21ai_1 _17844_ (.B1(_11198_),
    .Y(_01513_),
    .A1(net114),
    .A2(_11193_));
 sg13g2_nand2_1 _17845_ (.Y(_11199_),
    .A(\top_ihp.oisc.regs[39][15] ),
    .B(net546));
 sg13g2_o21ai_1 _17846_ (.B1(_11199_),
    .Y(_01514_),
    .A1(net233),
    .A2(net547));
 sg13g2_nand2_1 _17847_ (.Y(_11200_),
    .A(\top_ihp.oisc.regs[39][16] ),
    .B(_11194_));
 sg13g2_o21ai_1 _17848_ (.B1(_11200_),
    .Y(_01515_),
    .A1(net113),
    .A2(_11193_));
 sg13g2_nand2_1 _17849_ (.Y(_11201_),
    .A(\top_ihp.oisc.regs[39][17] ),
    .B(net546));
 sg13g2_o21ai_1 _17850_ (.B1(_11201_),
    .Y(_01516_),
    .A1(net236),
    .A2(net547));
 sg13g2_nand2_1 _17851_ (.Y(_11202_),
    .A(\top_ihp.oisc.regs[39][18] ),
    .B(net546));
 sg13g2_o21ai_1 _17852_ (.B1(_11202_),
    .Y(_01517_),
    .A1(net112),
    .A2(net547));
 sg13g2_mux2_1 _17853_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[39][19] ),
    .S(net548),
    .X(_01518_));
 sg13g2_buf_1 _17854_ (.A(_10318_),
    .X(_11203_));
 sg13g2_buf_1 _17855_ (.A(net654),
    .X(_11204_));
 sg13g2_nand2_1 _17856_ (.Y(_11205_),
    .A(\top_ihp.oisc.regs[39][1] ),
    .B(net545));
 sg13g2_o21ai_1 _17857_ (.B1(_11205_),
    .Y(_01519_),
    .A1(net105),
    .A2(net547));
 sg13g2_nand2_1 _17858_ (.Y(_11206_),
    .A(\top_ihp.oisc.regs[39][20] ),
    .B(net545));
 sg13g2_o21ai_1 _17859_ (.B1(_11206_),
    .Y(_01520_),
    .A1(_11102_),
    .A2(net547));
 sg13g2_buf_1 _17860_ (.A(net654),
    .X(_11207_));
 sg13g2_nand2_1 _17861_ (.Y(_11208_),
    .A(\top_ihp.oisc.regs[39][21] ),
    .B(_11204_));
 sg13g2_o21ai_1 _17862_ (.B1(_11208_),
    .Y(_01521_),
    .A1(net111),
    .A2(net544));
 sg13g2_nand2_1 _17863_ (.Y(_11209_),
    .A(\top_ihp.oisc.regs[39][22] ),
    .B(net545));
 sg13g2_o21ai_1 _17864_ (.B1(_11209_),
    .Y(_01522_),
    .A1(net110),
    .A2(net544));
 sg13g2_nand2_1 _17865_ (.Y(_11210_),
    .A(\top_ihp.oisc.regs[39][23] ),
    .B(_11204_));
 sg13g2_o21ai_1 _17866_ (.B1(_11210_),
    .Y(_01523_),
    .A1(_11109_),
    .A2(_11207_));
 sg13g2_buf_2 _17867_ (.A(net403),
    .X(_11211_));
 sg13g2_mux2_1 _17868_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[39][24] ),
    .S(net548),
    .X(_01524_));
 sg13g2_nand2_1 _17869_ (.Y(_11212_),
    .A(\top_ihp.oisc.regs[39][25] ),
    .B(net545));
 sg13g2_o21ai_1 _17870_ (.B1(_11212_),
    .Y(_01525_),
    .A1(net124),
    .A2(net544));
 sg13g2_nand2_1 _17871_ (.Y(_11213_),
    .A(\top_ihp.oisc.regs[39][26] ),
    .B(net545));
 sg13g2_o21ai_1 _17872_ (.B1(_11213_),
    .Y(_01526_),
    .A1(net235),
    .A2(_11207_));
 sg13g2_mux2_1 _17873_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[39][27] ),
    .S(net548),
    .X(_01527_));
 sg13g2_nand2_1 _17874_ (.Y(_11214_),
    .A(\top_ihp.oisc.regs[39][28] ),
    .B(net545));
 sg13g2_o21ai_1 _17875_ (.B1(_11214_),
    .Y(_01528_),
    .A1(net29),
    .A2(net544));
 sg13g2_nand2_1 _17876_ (.Y(_11215_),
    .A(\top_ihp.oisc.regs[39][29] ),
    .B(net545));
 sg13g2_o21ai_1 _17877_ (.B1(_11215_),
    .Y(_01529_),
    .A1(net108),
    .A2(net544));
 sg13g2_nand2_1 _17878_ (.Y(_11216_),
    .A(\top_ihp.oisc.regs[39][2] ),
    .B(net545));
 sg13g2_o21ai_1 _17879_ (.B1(_11216_),
    .Y(_01530_),
    .A1(_11147_),
    .A2(net544));
 sg13g2_nand2_1 _17880_ (.Y(_11217_),
    .A(\top_ihp.oisc.regs[39][30] ),
    .B(net654));
 sg13g2_o21ai_1 _17881_ (.B1(_11217_),
    .Y(_01531_),
    .A1(net28),
    .A2(net544));
 sg13g2_nand2_1 _17882_ (.Y(_11218_),
    .A(\top_ihp.oisc.regs[39][31] ),
    .B(net654));
 sg13g2_o21ai_1 _17883_ (.B1(_11218_),
    .Y(_01532_),
    .A1(net106),
    .A2(net544));
 sg13g2_buf_1 _17884_ (.A(net135),
    .X(_11219_));
 sg13g2_mux2_1 _17885_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[39][3] ),
    .S(_11191_),
    .X(_01533_));
 sg13g2_buf_1 _17886_ (.A(net134),
    .X(_11220_));
 sg13g2_mux2_1 _17887_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[39][4] ),
    .S(_11191_),
    .X(_01534_));
 sg13g2_buf_1 _17888_ (.A(_10625_),
    .X(_11221_));
 sg13g2_mux2_1 _17889_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[39][5] ),
    .S(net548),
    .X(_01535_));
 sg13g2_buf_1 _17890_ (.A(net132),
    .X(_11222_));
 sg13g2_mux2_1 _17891_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[39][6] ),
    .S(net546),
    .X(_01536_));
 sg13g2_nand2_1 _17892_ (.Y(_11223_),
    .A(\top_ihp.oisc.regs[39][7] ),
    .B(net654));
 sg13g2_o21ai_1 _17893_ (.B1(_11223_),
    .Y(_01537_),
    .A1(_11120_),
    .A2(net548));
 sg13g2_nand2_1 _17894_ (.Y(_11224_),
    .A(\top_ihp.oisc.regs[39][8] ),
    .B(net654));
 sg13g2_o21ai_1 _17895_ (.B1(_11224_),
    .Y(_01538_),
    .A1(net107),
    .A2(net548));
 sg13g2_buf_1 _17896_ (.A(_10687_),
    .X(_11225_));
 sg13g2_mux2_1 _17897_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[39][9] ),
    .S(net546),
    .X(_01539_));
 sg13g2_and2_1 _17898_ (.A(_09915_),
    .B(_10749_),
    .X(_11226_));
 sg13g2_buf_1 _17899_ (.A(_11226_),
    .X(_11227_));
 sg13g2_buf_1 _17900_ (.A(_11227_),
    .X(_11228_));
 sg13g2_mux2_1 _17901_ (.A0(\top_ihp.oisc.regs[3][0] ),
    .A1(net119),
    .S(net387),
    .X(_01540_));
 sg13g2_mux2_1 _17902_ (.A0(\top_ihp.oisc.regs[3][10] ),
    .A1(net130),
    .S(_11228_),
    .X(_01541_));
 sg13g2_nor2_1 _17903_ (.A(\top_ihp.oisc.regs[3][11] ),
    .B(net543),
    .Y(_11229_));
 sg13g2_a21oi_1 _17904_ (.A1(_10917_),
    .A2(_11228_),
    .Y(_01542_),
    .B1(_11229_));
 sg13g2_nor2_1 _17905_ (.A(\top_ihp.oisc.regs[3][12] ),
    .B(net543),
    .Y(_11230_));
 sg13g2_a21oi_1 _17906_ (.A1(_10855_),
    .A2(net387),
    .Y(_01543_),
    .B1(_11230_));
 sg13g2_nand2_1 _17907_ (.Y(_11231_),
    .A(_09915_),
    .B(_10749_));
 sg13g2_buf_1 _17908_ (.A(_11231_),
    .X(_11232_));
 sg13g2_buf_1 _17909_ (.A(net542),
    .X(_11233_));
 sg13g2_buf_1 _17910_ (.A(_11232_),
    .X(_11234_));
 sg13g2_nand2_1 _17911_ (.Y(_11235_),
    .A(\top_ihp.oisc.regs[3][13] ),
    .B(net385));
 sg13g2_o21ai_1 _17912_ (.B1(_11235_),
    .Y(_01544_),
    .A1(_11089_),
    .A2(net386));
 sg13g2_nand2_1 _17913_ (.Y(_11236_),
    .A(\top_ihp.oisc.regs[3][14] ),
    .B(net385));
 sg13g2_o21ai_1 _17914_ (.B1(_11236_),
    .Y(_01545_),
    .A1(_11091_),
    .A2(net386));
 sg13g2_buf_1 _17915_ (.A(net542),
    .X(_11237_));
 sg13g2_nand2_1 _17916_ (.Y(_11238_),
    .A(\top_ihp.oisc.regs[3][15] ),
    .B(net384));
 sg13g2_o21ai_1 _17917_ (.B1(_11238_),
    .Y(_01546_),
    .A1(_11165_),
    .A2(net386));
 sg13g2_nand2_1 _17918_ (.Y(_11239_),
    .A(\top_ihp.oisc.regs[3][16] ),
    .B(net384));
 sg13g2_o21ai_1 _17919_ (.B1(_11239_),
    .Y(_01547_),
    .A1(_11094_),
    .A2(net386));
 sg13g2_nand2_1 _17920_ (.Y(_11240_),
    .A(\top_ihp.oisc.regs[3][17] ),
    .B(_11237_));
 sg13g2_o21ai_1 _17921_ (.B1(_11240_),
    .Y(_01548_),
    .A1(_11096_),
    .A2(net386));
 sg13g2_nand2_1 _17922_ (.Y(_11241_),
    .A(\top_ihp.oisc.regs[3][18] ),
    .B(net384));
 sg13g2_o21ai_1 _17923_ (.B1(_11241_),
    .Y(_01549_),
    .A1(_11098_),
    .A2(net386));
 sg13g2_mux2_1 _17924_ (.A0(\top_ihp.oisc.regs[3][19] ),
    .A1(_10931_),
    .S(net387),
    .X(_01550_));
 sg13g2_nor2_1 _17925_ (.A(\top_ihp.oisc.regs[3][1] ),
    .B(net543),
    .Y(_11242_));
 sg13g2_a21oi_1 _17926_ (.A1(_10932_),
    .A2(net387),
    .Y(_01551_),
    .B1(_11242_));
 sg13g2_nand2_1 _17927_ (.Y(_11243_),
    .A(\top_ihp.oisc.regs[3][20] ),
    .B(_11237_));
 sg13g2_o21ai_1 _17928_ (.B1(_11243_),
    .Y(_01552_),
    .A1(_11102_),
    .A2(_11233_));
 sg13g2_nand2_1 _17929_ (.Y(_11244_),
    .A(\top_ihp.oisc.regs[3][21] ),
    .B(net384));
 sg13g2_o21ai_1 _17930_ (.B1(_11244_),
    .Y(_01553_),
    .A1(_11104_),
    .A2(net386));
 sg13g2_nand2_1 _17931_ (.Y(_11245_),
    .A(\top_ihp.oisc.regs[3][22] ),
    .B(net384));
 sg13g2_o21ai_1 _17932_ (.B1(_11245_),
    .Y(_01554_),
    .A1(_11107_),
    .A2(net386));
 sg13g2_nand2_1 _17933_ (.Y(_11246_),
    .A(\top_ihp.oisc.regs[3][23] ),
    .B(net384));
 sg13g2_o21ai_1 _17934_ (.B1(_11246_),
    .Y(_01555_),
    .A1(_11109_),
    .A2(_11233_));
 sg13g2_mux2_1 _17935_ (.A0(\top_ihp.oisc.regs[3][24] ),
    .A1(_10726_),
    .S(net387),
    .X(_01556_));
 sg13g2_nand2_1 _17936_ (.Y(_11247_),
    .A(\top_ihp.oisc.regs[3][25] ),
    .B(net384));
 sg13g2_o21ai_1 _17937_ (.B1(_11247_),
    .Y(_01557_),
    .A1(_10773_),
    .A2(net385));
 sg13g2_nand2_1 _17938_ (.Y(_11248_),
    .A(\top_ihp.oisc.regs[3][26] ),
    .B(net384));
 sg13g2_o21ai_1 _17939_ (.B1(_11248_),
    .Y(_01558_),
    .A1(_11112_),
    .A2(_11234_));
 sg13g2_mux2_1 _17940_ (.A0(\top_ihp.oisc.regs[3][27] ),
    .A1(_10940_),
    .S(net387),
    .X(_01559_));
 sg13g2_nor2_1 _17941_ (.A(\top_ihp.oisc.regs[3][28] ),
    .B(net543),
    .Y(_11249_));
 sg13g2_a21oi_1 _17942_ (.A1(_10941_),
    .A2(net387),
    .Y(_01560_),
    .B1(_11249_));
 sg13g2_nand2_1 _17943_ (.Y(_11250_),
    .A(\top_ihp.oisc.regs[3][29] ),
    .B(net542));
 sg13g2_o21ai_1 _17944_ (.B1(_11250_),
    .Y(_01561_),
    .A1(_11115_),
    .A2(_11234_));
 sg13g2_nand2_1 _17945_ (.Y(_11251_),
    .A(\top_ihp.oisc.regs[3][2] ),
    .B(net542));
 sg13g2_o21ai_1 _17946_ (.B1(_11251_),
    .Y(_01562_),
    .A1(_11147_),
    .A2(net385));
 sg13g2_nand2_1 _17947_ (.Y(_11252_),
    .A(\top_ihp.oisc.regs[3][30] ),
    .B(net542));
 sg13g2_o21ai_1 _17948_ (.B1(_11252_),
    .Y(_01563_),
    .A1(_11149_),
    .A2(net385));
 sg13g2_nand2_1 _17949_ (.Y(_11253_),
    .A(\top_ihp.oisc.regs[3][31] ),
    .B(net542));
 sg13g2_o21ai_1 _17950_ (.B1(_11253_),
    .Y(_01564_),
    .A1(_11151_),
    .A2(net385));
 sg13g2_mux2_1 _17951_ (.A0(\top_ihp.oisc.regs[3][3] ),
    .A1(net128),
    .S(net387),
    .X(_01565_));
 sg13g2_mux2_1 _17952_ (.A0(\top_ihp.oisc.regs[3][4] ),
    .A1(net127),
    .S(net543),
    .X(_01566_));
 sg13g2_mux2_1 _17953_ (.A0(\top_ihp.oisc.regs[3][5] ),
    .A1(_10741_),
    .S(net543),
    .X(_01567_));
 sg13g2_mux2_1 _17954_ (.A0(\top_ihp.oisc.regs[3][6] ),
    .A1(_10742_),
    .S(net543),
    .X(_01568_));
 sg13g2_nand2_1 _17955_ (.Y(_11254_),
    .A(\top_ihp.oisc.regs[3][7] ),
    .B(net542));
 sg13g2_o21ai_1 _17956_ (.B1(_11254_),
    .Y(_01569_),
    .A1(_11120_),
    .A2(net385));
 sg13g2_nand2_1 _17957_ (.Y(_11255_),
    .A(\top_ihp.oisc.regs[3][8] ),
    .B(net542));
 sg13g2_o21ai_1 _17958_ (.B1(_11255_),
    .Y(_01570_),
    .A1(_11122_),
    .A2(net385));
 sg13g2_mux2_1 _17959_ (.A0(\top_ihp.oisc.regs[3][9] ),
    .A1(_10745_),
    .S(net543),
    .X(_01571_));
 sg13g2_buf_1 _17960_ (.A(_09887_),
    .X(_11256_));
 sg13g2_and2_1 _17961_ (.A(_10694_),
    .B(_10985_),
    .X(_11257_));
 sg13g2_buf_2 _17962_ (.A(_11257_),
    .X(_11258_));
 sg13g2_and2_1 _17963_ (.A(_09939_),
    .B(_11258_),
    .X(_11259_));
 sg13g2_buf_1 _17964_ (.A(_11259_),
    .X(_11260_));
 sg13g2_buf_1 _17965_ (.A(net383),
    .X(_11261_));
 sg13g2_mux2_1 _17966_ (.A0(\top_ihp.oisc.regs[40][0] ),
    .A1(net103),
    .S(net231),
    .X(_01572_));
 sg13g2_buf_1 _17967_ (.A(_10008_),
    .X(_11262_));
 sg13g2_mux2_1 _17968_ (.A0(\top_ihp.oisc.regs[40][10] ),
    .A1(net102),
    .S(net231),
    .X(_01573_));
 sg13g2_nor2_1 _17969_ (.A(\top_ihp.oisc.regs[40][11] ),
    .B(_11260_),
    .Y(_11263_));
 sg13g2_a21oi_1 _17970_ (.A1(net50),
    .A2(_11261_),
    .Y(_01574_),
    .B1(_11263_));
 sg13g2_nor2_1 _17971_ (.A(\top_ihp.oisc.regs[40][12] ),
    .B(net383),
    .Y(_11264_));
 sg13g2_a21oi_1 _17972_ (.A1(net52),
    .A2(net231),
    .Y(_01575_),
    .B1(_11264_));
 sg13g2_nand2_1 _17973_ (.Y(_11265_),
    .A(_09939_),
    .B(_11258_));
 sg13g2_buf_2 _17974_ (.A(_11265_),
    .X(_11266_));
 sg13g2_buf_2 _17975_ (.A(_11266_),
    .X(_11267_));
 sg13g2_buf_1 _17976_ (.A(_11266_),
    .X(_11268_));
 sg13g2_nand2_1 _17977_ (.Y(_11269_),
    .A(\top_ihp.oisc.regs[40][13] ),
    .B(_11268_));
 sg13g2_o21ai_1 _17978_ (.B1(_11269_),
    .Y(_01576_),
    .A1(net115),
    .A2(_11267_));
 sg13g2_nand2_1 _17979_ (.Y(_11270_),
    .A(\top_ihp.oisc.regs[40][14] ),
    .B(net229));
 sg13g2_o21ai_1 _17980_ (.B1(_11270_),
    .Y(_01577_),
    .A1(net114),
    .A2(net230));
 sg13g2_mux2_1 _17981_ (.A0(\top_ihp.oisc.regs[40][15] ),
    .A1(net663),
    .S(net231),
    .X(_01578_));
 sg13g2_nand2_1 _17982_ (.Y(_11271_),
    .A(\top_ihp.oisc.regs[40][16] ),
    .B(_11268_));
 sg13g2_o21ai_1 _17983_ (.B1(_11271_),
    .Y(_01579_),
    .A1(net113),
    .A2(net230));
 sg13g2_buf_2 _17984_ (.A(_11266_),
    .X(_11272_));
 sg13g2_nand2_1 _17985_ (.Y(_11273_),
    .A(\top_ihp.oisc.regs[40][17] ),
    .B(net228));
 sg13g2_o21ai_1 _17986_ (.B1(_11273_),
    .Y(_01580_),
    .A1(net236),
    .A2(_11267_));
 sg13g2_nand2_1 _17987_ (.Y(_11274_),
    .A(\top_ihp.oisc.regs[40][18] ),
    .B(_11272_));
 sg13g2_o21ai_1 _17988_ (.B1(_11274_),
    .Y(_01581_),
    .A1(net112),
    .A2(net230));
 sg13g2_buf_1 _17989_ (.A(_10271_),
    .X(_11275_));
 sg13g2_mux2_1 _17990_ (.A0(\top_ihp.oisc.regs[40][19] ),
    .A1(net227),
    .S(net231),
    .X(_01582_));
 sg13g2_nor2_1 _17991_ (.A(\top_ihp.oisc.regs[40][1] ),
    .B(net383),
    .Y(_11276_));
 sg13g2_a21oi_1 _17992_ (.A1(net118),
    .A2(_11261_),
    .Y(_01583_),
    .B1(_11276_));
 sg13g2_nand2_1 _17993_ (.Y(_11277_),
    .A(\top_ihp.oisc.regs[40][20] ),
    .B(net228));
 sg13g2_o21ai_1 _17994_ (.B1(_11277_),
    .Y(_01584_),
    .A1(net48),
    .A2(net230));
 sg13g2_nand2_1 _17995_ (.Y(_11278_),
    .A(\top_ihp.oisc.regs[40][21] ),
    .B(net228));
 sg13g2_o21ai_1 _17996_ (.B1(_11278_),
    .Y(_01585_),
    .A1(net111),
    .A2(net230));
 sg13g2_nand2_1 _17997_ (.Y(_11279_),
    .A(\top_ihp.oisc.regs[40][22] ),
    .B(net228));
 sg13g2_o21ai_1 _17998_ (.B1(_11279_),
    .Y(_01586_),
    .A1(net110),
    .A2(net230));
 sg13g2_nand2_1 _17999_ (.Y(_11280_),
    .A(\top_ihp.oisc.regs[40][23] ),
    .B(net228));
 sg13g2_o21ai_1 _18000_ (.B1(_11280_),
    .Y(_01587_),
    .A1(net109),
    .A2(net230));
 sg13g2_buf_1 _18001_ (.A(_10414_),
    .X(_11281_));
 sg13g2_mux2_1 _18002_ (.A0(\top_ihp.oisc.regs[40][24] ),
    .A1(net382),
    .S(net231),
    .X(_01588_));
 sg13g2_nand2_1 _18003_ (.Y(_11282_),
    .A(\top_ihp.oisc.regs[40][25] ),
    .B(net228));
 sg13g2_o21ai_1 _18004_ (.B1(_11282_),
    .Y(_01589_),
    .A1(net124),
    .A2(net230));
 sg13g2_nand2_1 _18005_ (.Y(_11283_),
    .A(\top_ihp.oisc.regs[40][26] ),
    .B(_11272_));
 sg13g2_o21ai_1 _18006_ (.B1(_11283_),
    .Y(_01590_),
    .A1(_11112_),
    .A2(net229));
 sg13g2_buf_1 _18007_ (.A(_10447_),
    .X(_11284_));
 sg13g2_mux2_1 _18008_ (.A0(\top_ihp.oisc.regs[40][27] ),
    .A1(net101),
    .S(net231),
    .X(_01591_));
 sg13g2_nor2_1 _18009_ (.A(\top_ihp.oisc.regs[40][28] ),
    .B(net383),
    .Y(_11285_));
 sg13g2_a21oi_1 _18010_ (.A1(net30),
    .A2(net231),
    .Y(_01592_),
    .B1(_11285_));
 sg13g2_nand2_1 _18011_ (.Y(_11286_),
    .A(\top_ihp.oisc.regs[40][29] ),
    .B(net228));
 sg13g2_o21ai_1 _18012_ (.B1(_11286_),
    .Y(_01593_),
    .A1(net108),
    .A2(net229));
 sg13g2_nand2_1 _18013_ (.Y(_11287_),
    .A(\top_ihp.oisc.regs[40][2] ),
    .B(net228));
 sg13g2_o21ai_1 _18014_ (.B1(_11287_),
    .Y(_01594_),
    .A1(net47),
    .A2(net229));
 sg13g2_nand2_1 _18015_ (.Y(_11288_),
    .A(\top_ihp.oisc.regs[40][30] ),
    .B(_11266_));
 sg13g2_o21ai_1 _18016_ (.B1(_11288_),
    .Y(_01595_),
    .A1(net28),
    .A2(net229));
 sg13g2_nand2_1 _18017_ (.Y(_11289_),
    .A(\top_ihp.oisc.regs[40][31] ),
    .B(_11266_));
 sg13g2_o21ai_1 _18018_ (.B1(_11289_),
    .Y(_01596_),
    .A1(net106),
    .A2(net229));
 sg13g2_buf_1 _18019_ (.A(_10566_),
    .X(_11290_));
 sg13g2_mux2_1 _18020_ (.A0(\top_ihp.oisc.regs[40][3] ),
    .A1(net100),
    .S(_11260_),
    .X(_01597_));
 sg13g2_buf_2 _18021_ (.A(_10598_),
    .X(_11291_));
 sg13g2_mux2_1 _18022_ (.A0(\top_ihp.oisc.regs[40][4] ),
    .A1(net99),
    .S(net383),
    .X(_01598_));
 sg13g2_buf_2 _18023_ (.A(_10624_),
    .X(_11292_));
 sg13g2_mux2_1 _18024_ (.A0(\top_ihp.oisc.regs[40][5] ),
    .A1(net226),
    .S(net383),
    .X(_01599_));
 sg13g2_buf_1 _18025_ (.A(_10647_),
    .X(_11293_));
 sg13g2_mux2_1 _18026_ (.A0(\top_ihp.oisc.regs[40][6] ),
    .A1(net98),
    .S(net383),
    .X(_01600_));
 sg13g2_nand2_1 _18027_ (.Y(_11294_),
    .A(\top_ihp.oisc.regs[40][7] ),
    .B(_11266_));
 sg13g2_o21ai_1 _18028_ (.B1(_11294_),
    .Y(_01601_),
    .A1(net234),
    .A2(net229));
 sg13g2_nand2_1 _18029_ (.Y(_11295_),
    .A(\top_ihp.oisc.regs[40][8] ),
    .B(_11266_));
 sg13g2_o21ai_1 _18030_ (.B1(_11295_),
    .Y(_01602_),
    .A1(net107),
    .A2(net229));
 sg13g2_buf_1 _18031_ (.A(_10686_),
    .X(_11296_));
 sg13g2_mux2_1 _18032_ (.A0(\top_ihp.oisc.regs[40][9] ),
    .A1(net97),
    .S(net383),
    .X(_01603_));
 sg13g2_nand2_1 _18033_ (.Y(_11297_),
    .A(_10822_),
    .B(_11258_));
 sg13g2_buf_1 _18034_ (.A(_11297_),
    .X(_11298_));
 sg13g2_buf_2 _18035_ (.A(net381),
    .X(_11299_));
 sg13g2_mux2_1 _18036_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[41][0] ),
    .S(net225),
    .X(_01604_));
 sg13g2_mux2_1 _18037_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[41][10] ),
    .S(net225),
    .X(_01605_));
 sg13g2_buf_2 _18038_ (.A(net381),
    .X(_11300_));
 sg13g2_buf_2 _18039_ (.A(net381),
    .X(_11301_));
 sg13g2_nand2_1 _18040_ (.Y(_11302_),
    .A(\top_ihp.oisc.regs[41][11] ),
    .B(net223));
 sg13g2_o21ai_1 _18041_ (.B1(_11302_),
    .Y(_01606_),
    .A1(_10041_),
    .A2(net224));
 sg13g2_buf_1 _18042_ (.A(net141),
    .X(_11303_));
 sg13g2_nand2_1 _18043_ (.Y(_11304_),
    .A(\top_ihp.oisc.regs[41][12] ),
    .B(net223));
 sg13g2_o21ai_1 _18044_ (.B1(_11304_),
    .Y(_01607_),
    .A1(net40),
    .A2(net224));
 sg13g2_nand2_1 _18045_ (.Y(_11305_),
    .A(\top_ihp.oisc.regs[41][13] ),
    .B(net223));
 sg13g2_o21ai_1 _18046_ (.B1(_11305_),
    .Y(_01608_),
    .A1(net115),
    .A2(net224));
 sg13g2_nand2_1 _18047_ (.Y(_11306_),
    .A(\top_ihp.oisc.regs[41][14] ),
    .B(_11301_));
 sg13g2_o21ai_1 _18048_ (.B1(_11306_),
    .Y(_01609_),
    .A1(net114),
    .A2(_11300_));
 sg13g2_nand2_1 _18049_ (.Y(_11307_),
    .A(\top_ihp.oisc.regs[41][15] ),
    .B(net223));
 sg13g2_o21ai_1 _18050_ (.B1(_11307_),
    .Y(_01610_),
    .A1(net233),
    .A2(net224));
 sg13g2_nand2_1 _18051_ (.Y(_11308_),
    .A(\top_ihp.oisc.regs[41][16] ),
    .B(net223));
 sg13g2_o21ai_1 _18052_ (.B1(_11308_),
    .Y(_01611_),
    .A1(net113),
    .A2(net224));
 sg13g2_nand2_1 _18053_ (.Y(_11309_),
    .A(\top_ihp.oisc.regs[41][17] ),
    .B(_11301_));
 sg13g2_o21ai_1 _18054_ (.B1(_11309_),
    .Y(_01612_),
    .A1(_11096_),
    .A2(net224));
 sg13g2_nand2_1 _18055_ (.Y(_11310_),
    .A(\top_ihp.oisc.regs[41][18] ),
    .B(net223));
 sg13g2_o21ai_1 _18056_ (.B1(_11310_),
    .Y(_01613_),
    .A1(net112),
    .A2(net224));
 sg13g2_mux2_1 _18057_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[41][19] ),
    .S(_11299_),
    .X(_01614_));
 sg13g2_buf_1 _18058_ (.A(net381),
    .X(_11311_));
 sg13g2_nand2_1 _18059_ (.Y(_11312_),
    .A(\top_ihp.oisc.regs[41][1] ),
    .B(net222));
 sg13g2_o21ai_1 _18060_ (.B1(_11312_),
    .Y(_01615_),
    .A1(net105),
    .A2(net224));
 sg13g2_nand2_1 _18061_ (.Y(_11313_),
    .A(\top_ihp.oisc.regs[41][20] ),
    .B(net222));
 sg13g2_o21ai_1 _18062_ (.B1(_11313_),
    .Y(_01616_),
    .A1(net48),
    .A2(_11300_));
 sg13g2_buf_1 _18063_ (.A(net381),
    .X(_11314_));
 sg13g2_nand2_1 _18064_ (.Y(_11315_),
    .A(\top_ihp.oisc.regs[41][21] ),
    .B(_11311_));
 sg13g2_o21ai_1 _18065_ (.B1(_11315_),
    .Y(_01617_),
    .A1(net111),
    .A2(_11314_));
 sg13g2_nand2_1 _18066_ (.Y(_11316_),
    .A(\top_ihp.oisc.regs[41][22] ),
    .B(_11311_));
 sg13g2_o21ai_1 _18067_ (.B1(_11316_),
    .Y(_01618_),
    .A1(net110),
    .A2(_11314_));
 sg13g2_nand2_1 _18068_ (.Y(_11317_),
    .A(\top_ihp.oisc.regs[41][23] ),
    .B(net222));
 sg13g2_o21ai_1 _18069_ (.B1(_11317_),
    .Y(_01619_),
    .A1(net109),
    .A2(net221));
 sg13g2_mux2_1 _18070_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[41][24] ),
    .S(net225),
    .X(_01620_));
 sg13g2_nand2_1 _18071_ (.Y(_11318_),
    .A(\top_ihp.oisc.regs[41][25] ),
    .B(net222));
 sg13g2_o21ai_1 _18072_ (.B1(_11318_),
    .Y(_01621_),
    .A1(net124),
    .A2(net221));
 sg13g2_nand2_1 _18073_ (.Y(_11319_),
    .A(\top_ihp.oisc.regs[41][26] ),
    .B(net222));
 sg13g2_o21ai_1 _18074_ (.B1(_11319_),
    .Y(_01622_),
    .A1(net235),
    .A2(net221));
 sg13g2_mux2_1 _18075_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[41][27] ),
    .S(net225),
    .X(_01623_));
 sg13g2_nand2_1 _18076_ (.Y(_11320_),
    .A(\top_ihp.oisc.regs[41][28] ),
    .B(net222));
 sg13g2_o21ai_1 _18077_ (.B1(_11320_),
    .Y(_01624_),
    .A1(_10974_),
    .A2(net221));
 sg13g2_nand2_1 _18078_ (.Y(_11321_),
    .A(\top_ihp.oisc.regs[41][29] ),
    .B(net222));
 sg13g2_o21ai_1 _18079_ (.B1(_11321_),
    .Y(_01625_),
    .A1(net108),
    .A2(net221));
 sg13g2_nand2_1 _18080_ (.Y(_11322_),
    .A(\top_ihp.oisc.regs[41][2] ),
    .B(net222));
 sg13g2_o21ai_1 _18081_ (.B1(_11322_),
    .Y(_01626_),
    .A1(net47),
    .A2(net221));
 sg13g2_nand2_1 _18082_ (.Y(_11323_),
    .A(\top_ihp.oisc.regs[41][30] ),
    .B(net381));
 sg13g2_o21ai_1 _18083_ (.B1(_11323_),
    .Y(_01627_),
    .A1(net28),
    .A2(net221));
 sg13g2_nand2_1 _18084_ (.Y(_11324_),
    .A(\top_ihp.oisc.regs[41][31] ),
    .B(net381));
 sg13g2_o21ai_1 _18085_ (.B1(_11324_),
    .Y(_01628_),
    .A1(net106),
    .A2(net221));
 sg13g2_mux2_1 _18086_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[41][3] ),
    .S(_11299_),
    .X(_01629_));
 sg13g2_mux2_1 _18087_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[41][4] ),
    .S(net225),
    .X(_01630_));
 sg13g2_mux2_1 _18088_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[41][5] ),
    .S(net225),
    .X(_01631_));
 sg13g2_mux2_1 _18089_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[41][6] ),
    .S(net223),
    .X(_01632_));
 sg13g2_nand2_1 _18090_ (.Y(_11325_),
    .A(\top_ihp.oisc.regs[41][7] ),
    .B(_11298_));
 sg13g2_o21ai_1 _18091_ (.B1(_11325_),
    .Y(_01633_),
    .A1(net234),
    .A2(net225));
 sg13g2_nand2_1 _18092_ (.Y(_11326_),
    .A(\top_ihp.oisc.regs[41][8] ),
    .B(net381));
 sg13g2_o21ai_1 _18093_ (.B1(_11326_),
    .Y(_01634_),
    .A1(net107),
    .A2(net225));
 sg13g2_mux2_1 _18094_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[41][9] ),
    .S(net223),
    .X(_01635_));
 sg13g2_nand2_1 _18095_ (.Y(_11327_),
    .A(net740),
    .B(_11258_));
 sg13g2_buf_1 _18096_ (.A(_11327_),
    .X(_11328_));
 sg13g2_buf_2 _18097_ (.A(net380),
    .X(_11329_));
 sg13g2_mux2_1 _18098_ (.A0(_11155_),
    .A1(\top_ihp.oisc.regs[42][0] ),
    .S(_11329_),
    .X(_01636_));
 sg13g2_mux2_1 _18099_ (.A0(_11192_),
    .A1(\top_ihp.oisc.regs[42][10] ),
    .S(net220),
    .X(_01637_));
 sg13g2_buf_1 _18100_ (.A(_11328_),
    .X(_11330_));
 sg13g2_buf_1 _18101_ (.A(_11327_),
    .X(_11331_));
 sg13g2_nand2_1 _18102_ (.Y(_11332_),
    .A(\top_ihp.oisc.regs[42][11] ),
    .B(net379));
 sg13g2_o21ai_1 _18103_ (.B1(_11332_),
    .Y(_01638_),
    .A1(net49),
    .A2(net219));
 sg13g2_nand2_1 _18104_ (.Y(_11333_),
    .A(\top_ihp.oisc.regs[42][12] ),
    .B(net379));
 sg13g2_o21ai_1 _18105_ (.B1(_11333_),
    .Y(_01639_),
    .A1(net40),
    .A2(net219));
 sg13g2_nand2_1 _18106_ (.Y(_11334_),
    .A(\top_ihp.oisc.regs[42][13] ),
    .B(net379));
 sg13g2_o21ai_1 _18107_ (.B1(_11334_),
    .Y(_01640_),
    .A1(net115),
    .A2(net219));
 sg13g2_nand2_1 _18108_ (.Y(_11335_),
    .A(\top_ihp.oisc.regs[42][14] ),
    .B(_11331_));
 sg13g2_o21ai_1 _18109_ (.B1(_11335_),
    .Y(_01641_),
    .A1(net114),
    .A2(_11330_));
 sg13g2_nand2_1 _18110_ (.Y(_11336_),
    .A(\top_ihp.oisc.regs[42][15] ),
    .B(net379));
 sg13g2_o21ai_1 _18111_ (.B1(_11336_),
    .Y(_01642_),
    .A1(net233),
    .A2(net219));
 sg13g2_nand2_1 _18112_ (.Y(_11337_),
    .A(\top_ihp.oisc.regs[42][16] ),
    .B(_11331_));
 sg13g2_o21ai_1 _18113_ (.B1(_11337_),
    .Y(_01643_),
    .A1(net113),
    .A2(net219));
 sg13g2_nand2_1 _18114_ (.Y(_11338_),
    .A(\top_ihp.oisc.regs[42][17] ),
    .B(net379));
 sg13g2_o21ai_1 _18115_ (.B1(_11338_),
    .Y(_01644_),
    .A1(net236),
    .A2(net219));
 sg13g2_nand2_1 _18116_ (.Y(_11339_),
    .A(\top_ihp.oisc.regs[42][18] ),
    .B(net379));
 sg13g2_o21ai_1 _18117_ (.B1(_11339_),
    .Y(_01645_),
    .A1(net112),
    .A2(net219));
 sg13g2_buf_1 _18118_ (.A(net380),
    .X(_11340_));
 sg13g2_nand2_1 _18119_ (.Y(_11341_),
    .A(\top_ihp.oisc.regs[42][19] ),
    .B(net218));
 sg13g2_o21ai_1 _18120_ (.B1(_11341_),
    .Y(_01646_),
    .A1(net60),
    .A2(net219));
 sg13g2_buf_1 _18121_ (.A(net380),
    .X(_11342_));
 sg13g2_nand2_1 _18122_ (.Y(_11343_),
    .A(\top_ihp.oisc.regs[42][1] ),
    .B(_11340_));
 sg13g2_o21ai_1 _18123_ (.B1(_11343_),
    .Y(_01647_),
    .A1(net105),
    .A2(net217));
 sg13g2_nand2_1 _18124_ (.Y(_11344_),
    .A(\top_ihp.oisc.regs[42][20] ),
    .B(net218));
 sg13g2_o21ai_1 _18125_ (.B1(_11344_),
    .Y(_01648_),
    .A1(net48),
    .A2(_11342_));
 sg13g2_nand2_1 _18126_ (.Y(_11345_),
    .A(\top_ihp.oisc.regs[42][21] ),
    .B(_11340_));
 sg13g2_o21ai_1 _18127_ (.B1(_11345_),
    .Y(_01649_),
    .A1(net111),
    .A2(_11342_));
 sg13g2_nand2_1 _18128_ (.Y(_11346_),
    .A(\top_ihp.oisc.regs[42][22] ),
    .B(net218));
 sg13g2_o21ai_1 _18129_ (.B1(_11346_),
    .Y(_01650_),
    .A1(net110),
    .A2(net217));
 sg13g2_nand2_1 _18130_ (.Y(_11347_),
    .A(\top_ihp.oisc.regs[42][23] ),
    .B(net218));
 sg13g2_o21ai_1 _18131_ (.B1(_11347_),
    .Y(_01651_),
    .A1(net109),
    .A2(net217));
 sg13g2_mux2_1 _18132_ (.A0(_11211_),
    .A1(\top_ihp.oisc.regs[42][24] ),
    .S(net220),
    .X(_01652_));
 sg13g2_nand2_1 _18133_ (.Y(_11348_),
    .A(\top_ihp.oisc.regs[42][25] ),
    .B(net218));
 sg13g2_o21ai_1 _18134_ (.B1(_11348_),
    .Y(_01653_),
    .A1(net59),
    .A2(net217));
 sg13g2_nand2_1 _18135_ (.Y(_11349_),
    .A(\top_ihp.oisc.regs[42][26] ),
    .B(net218));
 sg13g2_o21ai_1 _18136_ (.B1(_11349_),
    .Y(_01654_),
    .A1(net235),
    .A2(net217));
 sg13g2_nand2_1 _18137_ (.Y(_11350_),
    .A(\top_ihp.oisc.regs[42][27] ),
    .B(net218));
 sg13g2_o21ai_1 _18138_ (.B1(_11350_),
    .Y(_01655_),
    .A1(net31),
    .A2(net217));
 sg13g2_nand2_1 _18139_ (.Y(_11351_),
    .A(\top_ihp.oisc.regs[42][28] ),
    .B(net218));
 sg13g2_o21ai_1 _18140_ (.B1(_11351_),
    .Y(_01656_),
    .A1(net29),
    .A2(net217));
 sg13g2_nand2_1 _18141_ (.Y(_11352_),
    .A(\top_ihp.oisc.regs[42][29] ),
    .B(net380));
 sg13g2_o21ai_1 _18142_ (.B1(_11352_),
    .Y(_01657_),
    .A1(net108),
    .A2(net217));
 sg13g2_nand2_1 _18143_ (.Y(_11353_),
    .A(\top_ihp.oisc.regs[42][2] ),
    .B(net380));
 sg13g2_o21ai_1 _18144_ (.B1(_11353_),
    .Y(_01658_),
    .A1(net47),
    .A2(net220));
 sg13g2_nand2_1 _18145_ (.Y(_11354_),
    .A(\top_ihp.oisc.regs[42][30] ),
    .B(net380));
 sg13g2_o21ai_1 _18146_ (.B1(_11354_),
    .Y(_01659_),
    .A1(net28),
    .A2(net220));
 sg13g2_inv_1 _18147_ (.Y(_11355_),
    .A(\top_ihp.oisc.regs[42][31] ));
 sg13g2_nor2_1 _18148_ (.A(net821),
    .B(_11328_),
    .Y(_11356_));
 sg13g2_a22oi_1 _18149_ (.Y(_01660_),
    .B1(_11356_),
    .B2(net129),
    .A2(_11330_),
    .A1(_11355_));
 sg13g2_mux2_1 _18150_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[42][3] ),
    .S(_11329_),
    .X(_01661_));
 sg13g2_mux2_1 _18151_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[42][4] ),
    .S(net220),
    .X(_01662_));
 sg13g2_mux2_1 _18152_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[42][5] ),
    .S(net220),
    .X(_01663_));
 sg13g2_mux2_1 _18153_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[42][6] ),
    .S(net379),
    .X(_01664_));
 sg13g2_nand2_1 _18154_ (.Y(_11357_),
    .A(\top_ihp.oisc.regs[42][7] ),
    .B(net380));
 sg13g2_o21ai_1 _18155_ (.B1(_11357_),
    .Y(_01665_),
    .A1(net234),
    .A2(net220));
 sg13g2_nand2_1 _18156_ (.Y(_11358_),
    .A(\top_ihp.oisc.regs[42][8] ),
    .B(net380));
 sg13g2_o21ai_1 _18157_ (.B1(_11358_),
    .Y(_01666_),
    .A1(net107),
    .A2(net220));
 sg13g2_mux2_1 _18158_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[42][9] ),
    .S(net379),
    .X(_01667_));
 sg13g2_and2_1 _18159_ (.A(_10747_),
    .B(_11258_),
    .X(_11359_));
 sg13g2_buf_2 _18160_ (.A(_11359_),
    .X(_11360_));
 sg13g2_buf_1 _18161_ (.A(_11360_),
    .X(_11361_));
 sg13g2_mux2_1 _18162_ (.A0(\top_ihp.oisc.regs[43][0] ),
    .A1(net103),
    .S(net216),
    .X(_01668_));
 sg13g2_mux2_1 _18163_ (.A0(\top_ihp.oisc.regs[43][10] ),
    .A1(net102),
    .S(net216),
    .X(_01669_));
 sg13g2_nand2_1 _18164_ (.Y(_11362_),
    .A(_10747_),
    .B(_11258_));
 sg13g2_buf_1 _18165_ (.A(_11362_),
    .X(_11363_));
 sg13g2_buf_1 _18166_ (.A(_11363_),
    .X(_11364_));
 sg13g2_buf_1 _18167_ (.A(_11362_),
    .X(_11365_));
 sg13g2_nand2_1 _18168_ (.Y(_11366_),
    .A(\top_ihp.oisc.regs[43][11] ),
    .B(net377));
 sg13g2_o21ai_1 _18169_ (.B1(_11366_),
    .Y(_01670_),
    .A1(_10041_),
    .A2(net215));
 sg13g2_nor2_1 _18170_ (.A(\top_ihp.oisc.regs[43][12] ),
    .B(_11360_),
    .Y(_11367_));
 sg13g2_a21oi_1 _18171_ (.A1(net52),
    .A2(net216),
    .Y(_01671_),
    .B1(_11367_));
 sg13g2_buf_1 _18172_ (.A(_11363_),
    .X(_11368_));
 sg13g2_nand2_1 _18173_ (.Y(_11369_),
    .A(\top_ihp.oisc.regs[43][13] ),
    .B(net214));
 sg13g2_o21ai_1 _18174_ (.B1(_11369_),
    .Y(_01672_),
    .A1(net115),
    .A2(net215));
 sg13g2_nand2_1 _18175_ (.Y(_11370_),
    .A(\top_ihp.oisc.regs[43][14] ),
    .B(_11368_));
 sg13g2_o21ai_1 _18176_ (.B1(_11370_),
    .Y(_01673_),
    .A1(net114),
    .A2(_11364_));
 sg13g2_nand2_1 _18177_ (.Y(_11371_),
    .A(\top_ihp.oisc.regs[43][15] ),
    .B(net214));
 sg13g2_o21ai_1 _18178_ (.B1(_11371_),
    .Y(_01674_),
    .A1(net233),
    .A2(net215));
 sg13g2_nand2_1 _18179_ (.Y(_11372_),
    .A(\top_ihp.oisc.regs[43][16] ),
    .B(net214));
 sg13g2_o21ai_1 _18180_ (.B1(_11372_),
    .Y(_01675_),
    .A1(net113),
    .A2(net215));
 sg13g2_nand2_1 _18181_ (.Y(_11373_),
    .A(\top_ihp.oisc.regs[43][17] ),
    .B(net214));
 sg13g2_o21ai_1 _18182_ (.B1(_11373_),
    .Y(_01676_),
    .A1(net236),
    .A2(net215));
 sg13g2_nand2_1 _18183_ (.Y(_11374_),
    .A(\top_ihp.oisc.regs[43][18] ),
    .B(_11368_));
 sg13g2_o21ai_1 _18184_ (.B1(_11374_),
    .Y(_01677_),
    .A1(net112),
    .A2(_11364_));
 sg13g2_mux2_1 _18185_ (.A0(\top_ihp.oisc.regs[43][19] ),
    .A1(net227),
    .S(net216),
    .X(_01678_));
 sg13g2_nor2_1 _18186_ (.A(\top_ihp.oisc.regs[43][1] ),
    .B(_11360_),
    .Y(_11375_));
 sg13g2_a21oi_1 _18187_ (.A1(net118),
    .A2(_11361_),
    .Y(_01679_),
    .B1(_11375_));
 sg13g2_nand2_1 _18188_ (.Y(_11376_),
    .A(\top_ihp.oisc.regs[43][20] ),
    .B(net214));
 sg13g2_o21ai_1 _18189_ (.B1(_11376_),
    .Y(_01680_),
    .A1(net48),
    .A2(net215));
 sg13g2_nand2_1 _18190_ (.Y(_11377_),
    .A(\top_ihp.oisc.regs[43][21] ),
    .B(net214));
 sg13g2_o21ai_1 _18191_ (.B1(_11377_),
    .Y(_01681_),
    .A1(_11104_),
    .A2(net215));
 sg13g2_nand2_1 _18192_ (.Y(_11378_),
    .A(\top_ihp.oisc.regs[43][22] ),
    .B(net214));
 sg13g2_o21ai_1 _18193_ (.B1(_11378_),
    .Y(_01682_),
    .A1(net110),
    .A2(net215));
 sg13g2_nand2_1 _18194_ (.Y(_11379_),
    .A(\top_ihp.oisc.regs[43][23] ),
    .B(net214));
 sg13g2_o21ai_1 _18195_ (.B1(_11379_),
    .Y(_01683_),
    .A1(net109),
    .A2(_11365_));
 sg13g2_mux2_1 _18196_ (.A0(\top_ihp.oisc.regs[43][24] ),
    .A1(_11281_),
    .S(net216),
    .X(_01684_));
 sg13g2_buf_1 _18197_ (.A(_10426_),
    .X(_11380_));
 sg13g2_nand2_1 _18198_ (.Y(_11381_),
    .A(\top_ihp.oisc.regs[43][25] ),
    .B(net378));
 sg13g2_o21ai_1 _18199_ (.B1(_11381_),
    .Y(_01685_),
    .A1(net213),
    .A2(net377));
 sg13g2_nand2_1 _18200_ (.Y(_11382_),
    .A(\top_ihp.oisc.regs[43][26] ),
    .B(net378));
 sg13g2_o21ai_1 _18201_ (.B1(_11382_),
    .Y(_01686_),
    .A1(net235),
    .A2(_11365_));
 sg13g2_mux2_1 _18202_ (.A0(\top_ihp.oisc.regs[43][27] ),
    .A1(_11284_),
    .S(net216),
    .X(_01687_));
 sg13g2_nor2_1 _18203_ (.A(\top_ihp.oisc.regs[43][28] ),
    .B(_11360_),
    .Y(_11383_));
 sg13g2_a21oi_1 _18204_ (.A1(net30),
    .A2(net216),
    .Y(_01688_),
    .B1(_11383_));
 sg13g2_nand2_1 _18205_ (.Y(_11384_),
    .A(\top_ihp.oisc.regs[43][29] ),
    .B(net378));
 sg13g2_o21ai_1 _18206_ (.B1(_11384_),
    .Y(_01689_),
    .A1(net108),
    .A2(net377));
 sg13g2_nand2_1 _18207_ (.Y(_11385_),
    .A(\top_ihp.oisc.regs[43][2] ),
    .B(net378));
 sg13g2_o21ai_1 _18208_ (.B1(_11385_),
    .Y(_01690_),
    .A1(net47),
    .A2(net377));
 sg13g2_nand2_1 _18209_ (.Y(_02870_),
    .A(\top_ihp.oisc.regs[43][30] ),
    .B(net378));
 sg13g2_o21ai_1 _18210_ (.B1(_02870_),
    .Y(_01691_),
    .A1(net28),
    .A2(net377));
 sg13g2_nand2_1 _18211_ (.Y(_02871_),
    .A(\top_ihp.oisc.regs[43][31] ),
    .B(net378));
 sg13g2_o21ai_1 _18212_ (.B1(_02871_),
    .Y(_01692_),
    .A1(net106),
    .A2(net377));
 sg13g2_mux2_1 _18213_ (.A0(\top_ihp.oisc.regs[43][3] ),
    .A1(net100),
    .S(net216),
    .X(_01693_));
 sg13g2_mux2_1 _18214_ (.A0(\top_ihp.oisc.regs[43][4] ),
    .A1(net99),
    .S(_11361_),
    .X(_01694_));
 sg13g2_mux2_1 _18215_ (.A0(\top_ihp.oisc.regs[43][5] ),
    .A1(net226),
    .S(_11360_),
    .X(_01695_));
 sg13g2_mux2_1 _18216_ (.A0(\top_ihp.oisc.regs[43][6] ),
    .A1(_11293_),
    .S(_11360_),
    .X(_01696_));
 sg13g2_nand2_1 _18217_ (.Y(_02872_),
    .A(\top_ihp.oisc.regs[43][7] ),
    .B(net378));
 sg13g2_o21ai_1 _18218_ (.B1(_02872_),
    .Y(_01697_),
    .A1(net234),
    .A2(net377));
 sg13g2_nand2_1 _18219_ (.Y(_02873_),
    .A(\top_ihp.oisc.regs[43][8] ),
    .B(net378));
 sg13g2_o21ai_1 _18220_ (.B1(_02873_),
    .Y(_01698_),
    .A1(net107),
    .A2(net377));
 sg13g2_mux2_1 _18221_ (.A0(\top_ihp.oisc.regs[43][9] ),
    .A1(net97),
    .S(_11360_),
    .X(_01699_));
 sg13g2_nor2_1 _18222_ (.A(_10847_),
    .B(_10984_),
    .Y(_02874_));
 sg13g2_buf_2 _18223_ (.A(_02874_),
    .X(_02875_));
 sg13g2_and2_1 _18224_ (.A(_09939_),
    .B(_02875_),
    .X(_02876_));
 sg13g2_buf_1 _18225_ (.A(_02876_),
    .X(_02877_));
 sg13g2_buf_2 _18226_ (.A(net541),
    .X(_02878_));
 sg13g2_mux2_1 _18227_ (.A0(\top_ihp.oisc.regs[44][0] ),
    .A1(net103),
    .S(net376),
    .X(_01700_));
 sg13g2_mux2_1 _18228_ (.A0(\top_ihp.oisc.regs[44][10] ),
    .A1(net102),
    .S(net376),
    .X(_01701_));
 sg13g2_nor2_1 _18229_ (.A(\top_ihp.oisc.regs[44][11] ),
    .B(net541),
    .Y(_02879_));
 sg13g2_a21oi_1 _18230_ (.A1(_10041_),
    .A2(net376),
    .Y(_01702_),
    .B1(_02879_));
 sg13g2_nor2_1 _18231_ (.A(\top_ihp.oisc.regs[44][12] ),
    .B(_02877_),
    .Y(_02880_));
 sg13g2_a21oi_1 _18232_ (.A1(net52),
    .A2(_02878_),
    .Y(_01703_),
    .B1(_02880_));
 sg13g2_nand2_1 _18233_ (.Y(_02881_),
    .A(_09939_),
    .B(_02875_));
 sg13g2_buf_1 _18234_ (.A(_02881_),
    .X(_02882_));
 sg13g2_buf_1 _18235_ (.A(net540),
    .X(_02883_));
 sg13g2_buf_2 _18236_ (.A(net540),
    .X(_02884_));
 sg13g2_nand2_1 _18237_ (.Y(_02885_),
    .A(\top_ihp.oisc.regs[44][13] ),
    .B(_02884_));
 sg13g2_o21ai_1 _18238_ (.B1(_02885_),
    .Y(_01704_),
    .A1(net115),
    .A2(_02883_));
 sg13g2_nand2_1 _18239_ (.Y(_02886_),
    .A(\top_ihp.oisc.regs[44][14] ),
    .B(_02884_));
 sg13g2_o21ai_1 _18240_ (.B1(_02886_),
    .Y(_01705_),
    .A1(net114),
    .A2(_02883_));
 sg13g2_buf_1 _18241_ (.A(net540),
    .X(_02887_));
 sg13g2_nand2_1 _18242_ (.Y(_02888_),
    .A(\top_ihp.oisc.regs[44][15] ),
    .B(net373));
 sg13g2_o21ai_1 _18243_ (.B1(_02888_),
    .Y(_01706_),
    .A1(net233),
    .A2(net375));
 sg13g2_nand2_1 _18244_ (.Y(_02889_),
    .A(\top_ihp.oisc.regs[44][16] ),
    .B(_02887_));
 sg13g2_o21ai_1 _18245_ (.B1(_02889_),
    .Y(_01707_),
    .A1(net113),
    .A2(net375));
 sg13g2_nand2_1 _18246_ (.Y(_02890_),
    .A(\top_ihp.oisc.regs[44][17] ),
    .B(net373));
 sg13g2_o21ai_1 _18247_ (.B1(_02890_),
    .Y(_01708_),
    .A1(net236),
    .A2(net375));
 sg13g2_nand2_1 _18248_ (.Y(_02891_),
    .A(\top_ihp.oisc.regs[44][18] ),
    .B(_02887_));
 sg13g2_o21ai_1 _18249_ (.B1(_02891_),
    .Y(_01709_),
    .A1(net112),
    .A2(net375));
 sg13g2_mux2_1 _18250_ (.A0(\top_ihp.oisc.regs[44][19] ),
    .A1(_11275_),
    .S(net376),
    .X(_01710_));
 sg13g2_nor2_1 _18251_ (.A(\top_ihp.oisc.regs[44][1] ),
    .B(net541),
    .Y(_02892_));
 sg13g2_a21oi_1 _18252_ (.A1(net118),
    .A2(net376),
    .Y(_01711_),
    .B1(_02892_));
 sg13g2_nand2_1 _18253_ (.Y(_02893_),
    .A(\top_ihp.oisc.regs[44][20] ),
    .B(net373));
 sg13g2_o21ai_1 _18254_ (.B1(_02893_),
    .Y(_01712_),
    .A1(net48),
    .A2(net375));
 sg13g2_nand2_1 _18255_ (.Y(_02894_),
    .A(\top_ihp.oisc.regs[44][21] ),
    .B(net373));
 sg13g2_o21ai_1 _18256_ (.B1(_02894_),
    .Y(_01713_),
    .A1(net111),
    .A2(net375));
 sg13g2_nand2_1 _18257_ (.Y(_02895_),
    .A(\top_ihp.oisc.regs[44][22] ),
    .B(net373));
 sg13g2_o21ai_1 _18258_ (.B1(_02895_),
    .Y(_01714_),
    .A1(_11107_),
    .A2(net375));
 sg13g2_nand2_1 _18259_ (.Y(_02896_),
    .A(\top_ihp.oisc.regs[44][23] ),
    .B(net373));
 sg13g2_o21ai_1 _18260_ (.B1(_02896_),
    .Y(_01715_),
    .A1(net109),
    .A2(net375));
 sg13g2_mux2_1 _18261_ (.A0(\top_ihp.oisc.regs[44][24] ),
    .A1(net382),
    .S(net376),
    .X(_01716_));
 sg13g2_nand2_1 _18262_ (.Y(_02897_),
    .A(\top_ihp.oisc.regs[44][25] ),
    .B(net373));
 sg13g2_o21ai_1 _18263_ (.B1(_02897_),
    .Y(_01717_),
    .A1(_11380_),
    .A2(net374));
 sg13g2_nand2_1 _18264_ (.Y(_02898_),
    .A(\top_ihp.oisc.regs[44][26] ),
    .B(net373));
 sg13g2_o21ai_1 _18265_ (.B1(_02898_),
    .Y(_01718_),
    .A1(net235),
    .A2(net374));
 sg13g2_mux2_1 _18266_ (.A0(\top_ihp.oisc.regs[44][27] ),
    .A1(net101),
    .S(net376),
    .X(_01719_));
 sg13g2_nor2_1 _18267_ (.A(\top_ihp.oisc.regs[44][28] ),
    .B(net541),
    .Y(_02899_));
 sg13g2_a21oi_1 _18268_ (.A1(net116),
    .A2(net376),
    .Y(_01720_),
    .B1(_02899_));
 sg13g2_nand2_1 _18269_ (.Y(_02900_),
    .A(\top_ihp.oisc.regs[44][29] ),
    .B(net540));
 sg13g2_o21ai_1 _18270_ (.B1(_02900_),
    .Y(_01721_),
    .A1(_11115_),
    .A2(net374));
 sg13g2_nand2_1 _18271_ (.Y(_02901_),
    .A(\top_ihp.oisc.regs[44][2] ),
    .B(net540));
 sg13g2_o21ai_1 _18272_ (.B1(_02901_),
    .Y(_01722_),
    .A1(net47),
    .A2(net374));
 sg13g2_nand2_1 _18273_ (.Y(_02902_),
    .A(\top_ihp.oisc.regs[44][30] ),
    .B(net540));
 sg13g2_o21ai_1 _18274_ (.B1(_02902_),
    .Y(_01723_),
    .A1(net28),
    .A2(net374));
 sg13g2_nand2_1 _18275_ (.Y(_02903_),
    .A(\top_ihp.oisc.regs[44][31] ),
    .B(net540));
 sg13g2_o21ai_1 _18276_ (.B1(_02903_),
    .Y(_01724_),
    .A1(net106),
    .A2(net374));
 sg13g2_mux2_1 _18277_ (.A0(\top_ihp.oisc.regs[44][3] ),
    .A1(net100),
    .S(_02878_),
    .X(_01725_));
 sg13g2_mux2_1 _18278_ (.A0(\top_ihp.oisc.regs[44][4] ),
    .A1(net99),
    .S(net541),
    .X(_01726_));
 sg13g2_mux2_1 _18279_ (.A0(\top_ihp.oisc.regs[44][5] ),
    .A1(net226),
    .S(net541),
    .X(_01727_));
 sg13g2_mux2_1 _18280_ (.A0(\top_ihp.oisc.regs[44][6] ),
    .A1(net98),
    .S(net541),
    .X(_01728_));
 sg13g2_nand2_1 _18281_ (.Y(_02904_),
    .A(\top_ihp.oisc.regs[44][7] ),
    .B(_02882_));
 sg13g2_o21ai_1 _18282_ (.B1(_02904_),
    .Y(_01729_),
    .A1(net234),
    .A2(net374));
 sg13g2_nand2_1 _18283_ (.Y(_02905_),
    .A(\top_ihp.oisc.regs[44][8] ),
    .B(net540));
 sg13g2_o21ai_1 _18284_ (.B1(_02905_),
    .Y(_01730_),
    .A1(net107),
    .A2(net374));
 sg13g2_mux2_1 _18285_ (.A0(\top_ihp.oisc.regs[44][9] ),
    .A1(net97),
    .S(net541),
    .X(_01731_));
 sg13g2_nand2_1 _18286_ (.Y(_02906_),
    .A(_10822_),
    .B(_02875_));
 sg13g2_buf_2 _18287_ (.A(_02906_),
    .X(_02907_));
 sg13g2_buf_2 _18288_ (.A(_02907_),
    .X(_02908_));
 sg13g2_mux2_1 _18289_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[45][0] ),
    .S(_02908_),
    .X(_01732_));
 sg13g2_mux2_1 _18290_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[45][10] ),
    .S(net372),
    .X(_01733_));
 sg13g2_buf_1 _18291_ (.A(_02907_),
    .X(_02909_));
 sg13g2_buf_2 _18292_ (.A(_02907_),
    .X(_02910_));
 sg13g2_nand2_1 _18293_ (.Y(_02911_),
    .A(\top_ihp.oisc.regs[45][11] ),
    .B(net370));
 sg13g2_o21ai_1 _18294_ (.B1(_02911_),
    .Y(_01734_),
    .A1(_10991_),
    .A2(net371));
 sg13g2_nand2_1 _18295_ (.Y(_02912_),
    .A(\top_ihp.oisc.regs[45][12] ),
    .B(net370));
 sg13g2_o21ai_1 _18296_ (.B1(_02912_),
    .Y(_01735_),
    .A1(net40),
    .A2(net371));
 sg13g2_buf_1 _18297_ (.A(net261),
    .X(_02913_));
 sg13g2_nand2_1 _18298_ (.Y(_02914_),
    .A(\top_ihp.oisc.regs[45][13] ),
    .B(net370));
 sg13g2_o21ai_1 _18299_ (.B1(_02914_),
    .Y(_01736_),
    .A1(net96),
    .A2(net371));
 sg13g2_buf_1 _18300_ (.A(net260),
    .X(_02915_));
 sg13g2_nand2_1 _18301_ (.Y(_02916_),
    .A(\top_ihp.oisc.regs[45][14] ),
    .B(_02910_));
 sg13g2_o21ai_1 _18302_ (.B1(_02916_),
    .Y(_01737_),
    .A1(net95),
    .A2(net371));
 sg13g2_mux2_1 _18303_ (.A0(net663),
    .A1(\top_ihp.oisc.regs[45][15] ),
    .S(net372),
    .X(_01738_));
 sg13g2_buf_1 _18304_ (.A(net276),
    .X(_02917_));
 sg13g2_nand2_1 _18305_ (.Y(_02918_),
    .A(\top_ihp.oisc.regs[45][16] ),
    .B(net370));
 sg13g2_o21ai_1 _18306_ (.B1(_02918_),
    .Y(_01739_),
    .A1(net94),
    .A2(net371));
 sg13g2_buf_1 _18307_ (.A(_10800_),
    .X(_02919_));
 sg13g2_nand2_1 _18308_ (.Y(_02920_),
    .A(\top_ihp.oisc.regs[45][17] ),
    .B(net370));
 sg13g2_o21ai_1 _18309_ (.B1(_02920_),
    .Y(_01740_),
    .A1(net212),
    .A2(_02909_));
 sg13g2_buf_1 _18310_ (.A(net259),
    .X(_02921_));
 sg13g2_nand2_1 _18311_ (.Y(_02922_),
    .A(\top_ihp.oisc.regs[45][18] ),
    .B(_02910_));
 sg13g2_o21ai_1 _18312_ (.B1(_02922_),
    .Y(_01741_),
    .A1(net93),
    .A2(_02909_));
 sg13g2_mux2_1 _18313_ (.A0(net263),
    .A1(\top_ihp.oisc.regs[45][19] ),
    .S(net372),
    .X(_01742_));
 sg13g2_nand2_1 _18314_ (.Y(_02923_),
    .A(\top_ihp.oisc.regs[45][1] ),
    .B(net370));
 sg13g2_o21ai_1 _18315_ (.B1(_02923_),
    .Y(_01743_),
    .A1(_11203_),
    .A2(net371));
 sg13g2_buf_1 _18316_ (.A(net121),
    .X(_02924_));
 sg13g2_buf_1 _18317_ (.A(_02907_),
    .X(_02925_));
 sg13g2_nand2_1 _18318_ (.Y(_02926_),
    .A(\top_ihp.oisc.regs[45][20] ),
    .B(_02925_));
 sg13g2_o21ai_1 _18319_ (.B1(_02926_),
    .Y(_01744_),
    .A1(net39),
    .A2(net371));
 sg13g2_buf_1 _18320_ (.A(net273),
    .X(_02927_));
 sg13g2_nand2_1 _18321_ (.Y(_02928_),
    .A(\top_ihp.oisc.regs[45][21] ),
    .B(net369));
 sg13g2_o21ai_1 _18322_ (.B1(_02928_),
    .Y(_01745_),
    .A1(net92),
    .A2(net371));
 sg13g2_buf_2 _18323_ (.A(_10807_),
    .X(_02929_));
 sg13g2_buf_1 _18324_ (.A(_02907_),
    .X(_02930_));
 sg13g2_nand2_1 _18325_ (.Y(_02931_),
    .A(\top_ihp.oisc.regs[45][22] ),
    .B(_02925_));
 sg13g2_o21ai_1 _18326_ (.B1(_02931_),
    .Y(_01746_),
    .A1(net91),
    .A2(net368));
 sg13g2_buf_1 _18327_ (.A(_10808_),
    .X(_02932_));
 sg13g2_nand2_1 _18328_ (.Y(_02933_),
    .A(\top_ihp.oisc.regs[45][23] ),
    .B(net369));
 sg13g2_o21ai_1 _18329_ (.B1(_02933_),
    .Y(_01747_),
    .A1(net90),
    .A2(net368));
 sg13g2_mux2_1 _18330_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[45][24] ),
    .S(net372),
    .X(_01748_));
 sg13g2_nand2_1 _18331_ (.Y(_02934_),
    .A(\top_ihp.oisc.regs[45][25] ),
    .B(net369));
 sg13g2_o21ai_1 _18332_ (.B1(_02934_),
    .Y(_01749_),
    .A1(net213),
    .A2(net368));
 sg13g2_buf_2 _18333_ (.A(net397),
    .X(_02935_));
 sg13g2_nand2_1 _18334_ (.Y(_02936_),
    .A(\top_ihp.oisc.regs[45][26] ),
    .B(net369));
 sg13g2_o21ai_1 _18335_ (.B1(_02936_),
    .Y(_01750_),
    .A1(net211),
    .A2(_02930_));
 sg13g2_mux2_1 _18336_ (.A0(net123),
    .A1(\top_ihp.oisc.regs[45][27] ),
    .S(net372),
    .X(_01751_));
 sg13g2_buf_1 _18337_ (.A(_10459_),
    .X(_02937_));
 sg13g2_nand2_1 _18338_ (.Y(_02938_),
    .A(\top_ihp.oisc.regs[45][28] ),
    .B(net369));
 sg13g2_o21ai_1 _18339_ (.B1(_02938_),
    .Y(_01752_),
    .A1(net27),
    .A2(net368));
 sg13g2_buf_1 _18340_ (.A(net256),
    .X(_02939_));
 sg13g2_nand2_1 _18341_ (.Y(_02940_),
    .A(\top_ihp.oisc.regs[45][29] ),
    .B(net369));
 sg13g2_o21ai_1 _18342_ (.B1(_02940_),
    .Y(_01753_),
    .A1(net89),
    .A2(_02930_));
 sg13g2_nand2_1 _18343_ (.Y(_02941_),
    .A(\top_ihp.oisc.regs[45][2] ),
    .B(net369));
 sg13g2_o21ai_1 _18344_ (.B1(_02941_),
    .Y(_01754_),
    .A1(net47),
    .A2(net368));
 sg13g2_nand2_1 _18345_ (.Y(_02942_),
    .A(\top_ihp.oisc.regs[45][30] ),
    .B(net369));
 sg13g2_o21ai_1 _18346_ (.B1(_02942_),
    .Y(_01755_),
    .A1(net28),
    .A2(net368));
 sg13g2_nand2_1 _18347_ (.Y(_02943_),
    .A(\top_ihp.oisc.regs[45][31] ),
    .B(_02907_));
 sg13g2_o21ai_1 _18348_ (.B1(_02943_),
    .Y(_01756_),
    .A1(net106),
    .A2(net368));
 sg13g2_mux2_1 _18349_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[45][3] ),
    .S(_02908_),
    .X(_01757_));
 sg13g2_mux2_1 _18350_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[45][4] ),
    .S(net372),
    .X(_01758_));
 sg13g2_mux2_1 _18351_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[45][5] ),
    .S(net372),
    .X(_01759_));
 sg13g2_mux2_1 _18352_ (.A0(_11222_),
    .A1(\top_ihp.oisc.regs[45][6] ),
    .S(net370),
    .X(_01760_));
 sg13g2_buf_2 _18353_ (.A(net396),
    .X(_02944_));
 sg13g2_nand2_1 _18354_ (.Y(_02945_),
    .A(\top_ihp.oisc.regs[45][7] ),
    .B(_02907_));
 sg13g2_o21ai_1 _18355_ (.B1(_02945_),
    .Y(_01761_),
    .A1(net210),
    .A2(net368));
 sg13g2_buf_2 _18356_ (.A(net255),
    .X(_02946_));
 sg13g2_nand2_1 _18357_ (.Y(_02947_),
    .A(\top_ihp.oisc.regs[45][8] ),
    .B(_02907_));
 sg13g2_o21ai_1 _18358_ (.B1(_02947_),
    .Y(_01762_),
    .A1(net88),
    .A2(net372));
 sg13g2_mux2_1 _18359_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[45][9] ),
    .S(net370),
    .X(_01763_));
 sg13g2_and2_1 _18360_ (.A(net740),
    .B(_02875_),
    .X(_02948_));
 sg13g2_buf_1 _18361_ (.A(_02948_),
    .X(_02949_));
 sg13g2_buf_2 _18362_ (.A(_02949_),
    .X(_02950_));
 sg13g2_mux2_1 _18363_ (.A0(\top_ihp.oisc.regs[46][0] ),
    .A1(net103),
    .S(_02950_),
    .X(_01764_));
 sg13g2_mux2_1 _18364_ (.A0(\top_ihp.oisc.regs[46][10] ),
    .A1(net102),
    .S(net367),
    .X(_01765_));
 sg13g2_nand2_1 _18365_ (.Y(_02951_),
    .A(net740),
    .B(_02875_));
 sg13g2_buf_2 _18366_ (.A(_02951_),
    .X(_02952_));
 sg13g2_buf_1 _18367_ (.A(_02952_),
    .X(_02953_));
 sg13g2_buf_1 _18368_ (.A(_02952_),
    .X(_02954_));
 sg13g2_nand2_1 _18369_ (.Y(_02955_),
    .A(\top_ihp.oisc.regs[46][11] ),
    .B(net365));
 sg13g2_o21ai_1 _18370_ (.B1(_02955_),
    .Y(_01766_),
    .A1(net49),
    .A2(net366));
 sg13g2_nor2_1 _18371_ (.A(\top_ihp.oisc.regs[46][12] ),
    .B(_02949_),
    .Y(_02956_));
 sg13g2_a21oi_1 _18372_ (.A1(net52),
    .A2(net367),
    .Y(_01767_),
    .B1(_02956_));
 sg13g2_nand2_1 _18373_ (.Y(_02957_),
    .A(\top_ihp.oisc.regs[46][13] ),
    .B(net365));
 sg13g2_o21ai_1 _18374_ (.B1(_02957_),
    .Y(_01768_),
    .A1(net96),
    .A2(net366));
 sg13g2_nand2_1 _18375_ (.Y(_02958_),
    .A(\top_ihp.oisc.regs[46][14] ),
    .B(net365));
 sg13g2_o21ai_1 _18376_ (.B1(_02958_),
    .Y(_01769_),
    .A1(net95),
    .A2(net366));
 sg13g2_nand2_1 _18377_ (.Y(_02959_),
    .A(\top_ihp.oisc.regs[46][15] ),
    .B(net365));
 sg13g2_o21ai_1 _18378_ (.B1(_02959_),
    .Y(_01770_),
    .A1(net233),
    .A2(net366));
 sg13g2_nand2_1 _18379_ (.Y(_02960_),
    .A(\top_ihp.oisc.regs[46][16] ),
    .B(net365));
 sg13g2_o21ai_1 _18380_ (.B1(_02960_),
    .Y(_01771_),
    .A1(net94),
    .A2(_02953_));
 sg13g2_nand2_1 _18381_ (.Y(_02961_),
    .A(\top_ihp.oisc.regs[46][17] ),
    .B(_02954_));
 sg13g2_o21ai_1 _18382_ (.B1(_02961_),
    .Y(_01772_),
    .A1(net212),
    .A2(_02953_));
 sg13g2_nand2_1 _18383_ (.Y(_02962_),
    .A(\top_ihp.oisc.regs[46][18] ),
    .B(net365));
 sg13g2_o21ai_1 _18384_ (.B1(_02962_),
    .Y(_01773_),
    .A1(net93),
    .A2(net366));
 sg13g2_nand2_1 _18385_ (.Y(_02963_),
    .A(\top_ihp.oisc.regs[46][19] ),
    .B(_02954_));
 sg13g2_o21ai_1 _18386_ (.B1(_02963_),
    .Y(_01774_),
    .A1(net60),
    .A2(net366));
 sg13g2_nor2_1 _18387_ (.A(\top_ihp.oisc.regs[46][1] ),
    .B(_02949_),
    .Y(_02964_));
 sg13g2_a21oi_1 _18388_ (.A1(net118),
    .A2(net367),
    .Y(_01775_),
    .B1(_02964_));
 sg13g2_buf_1 _18389_ (.A(_02952_),
    .X(_02965_));
 sg13g2_nand2_1 _18390_ (.Y(_02966_),
    .A(\top_ihp.oisc.regs[46][20] ),
    .B(net364));
 sg13g2_o21ai_1 _18391_ (.B1(_02966_),
    .Y(_01776_),
    .A1(net39),
    .A2(net366));
 sg13g2_buf_1 _18392_ (.A(_02952_),
    .X(_02967_));
 sg13g2_nand2_1 _18393_ (.Y(_02968_),
    .A(\top_ihp.oisc.regs[46][21] ),
    .B(_02965_));
 sg13g2_o21ai_1 _18394_ (.B1(_02968_),
    .Y(_01777_),
    .A1(net92),
    .A2(net363));
 sg13g2_nand2_1 _18395_ (.Y(_02969_),
    .A(\top_ihp.oisc.regs[46][22] ),
    .B(net364));
 sg13g2_o21ai_1 _18396_ (.B1(_02969_),
    .Y(_01778_),
    .A1(_02929_),
    .A2(net363));
 sg13g2_nand2_1 _18397_ (.Y(_02970_),
    .A(\top_ihp.oisc.regs[46][23] ),
    .B(net364));
 sg13g2_o21ai_1 _18398_ (.B1(_02970_),
    .Y(_01779_),
    .A1(net90),
    .A2(net363));
 sg13g2_mux2_1 _18399_ (.A0(\top_ihp.oisc.regs[46][24] ),
    .A1(net382),
    .S(net367),
    .X(_01780_));
 sg13g2_nand2_1 _18400_ (.Y(_02971_),
    .A(\top_ihp.oisc.regs[46][25] ),
    .B(net364));
 sg13g2_o21ai_1 _18401_ (.B1(_02971_),
    .Y(_01781_),
    .A1(_10428_),
    .A2(net363));
 sg13g2_nand2_1 _18402_ (.Y(_02972_),
    .A(\top_ihp.oisc.regs[46][26] ),
    .B(net364));
 sg13g2_o21ai_1 _18403_ (.B1(_02972_),
    .Y(_01782_),
    .A1(net211),
    .A2(_02967_));
 sg13g2_nand2_1 _18404_ (.Y(_02973_),
    .A(\top_ihp.oisc.regs[46][27] ),
    .B(net364));
 sg13g2_o21ai_1 _18405_ (.B1(_02973_),
    .Y(_01783_),
    .A1(net31),
    .A2(net363));
 sg13g2_nand2_1 _18406_ (.Y(_02974_),
    .A(\top_ihp.oisc.regs[46][28] ),
    .B(_02965_));
 sg13g2_o21ai_1 _18407_ (.B1(_02974_),
    .Y(_01784_),
    .A1(net27),
    .A2(net363));
 sg13g2_nand2_1 _18408_ (.Y(_02975_),
    .A(\top_ihp.oisc.regs[46][29] ),
    .B(net364));
 sg13g2_o21ai_1 _18409_ (.B1(_02975_),
    .Y(_01785_),
    .A1(net89),
    .A2(_02967_));
 sg13g2_buf_1 _18410_ (.A(net122),
    .X(_02976_));
 sg13g2_nand2_1 _18411_ (.Y(_02977_),
    .A(\top_ihp.oisc.regs[46][2] ),
    .B(net364));
 sg13g2_o21ai_1 _18412_ (.B1(_02977_),
    .Y(_01786_),
    .A1(net38),
    .A2(net363));
 sg13g2_buf_1 _18413_ (.A(net53),
    .X(_02978_));
 sg13g2_nand2_1 _18414_ (.Y(_02979_),
    .A(\top_ihp.oisc.regs[46][30] ),
    .B(_02952_));
 sg13g2_o21ai_1 _18415_ (.B1(_02979_),
    .Y(_01787_),
    .A1(net26),
    .A2(net363));
 sg13g2_inv_1 _18416_ (.Y(_02980_),
    .A(\top_ihp.oisc.regs[46][31] ));
 sg13g2_nor2_1 _18417_ (.A(net821),
    .B(_02952_),
    .Y(_02981_));
 sg13g2_a22oi_1 _18418_ (.Y(_01788_),
    .B1(_02981_),
    .B2(net129),
    .A2(net366),
    .A1(_02980_));
 sg13g2_mux2_1 _18419_ (.A0(\top_ihp.oisc.regs[46][3] ),
    .A1(net100),
    .S(net367),
    .X(_01789_));
 sg13g2_mux2_1 _18420_ (.A0(\top_ihp.oisc.regs[46][4] ),
    .A1(net99),
    .S(net367),
    .X(_01790_));
 sg13g2_mux2_1 _18421_ (.A0(\top_ihp.oisc.regs[46][5] ),
    .A1(net226),
    .S(net367),
    .X(_01791_));
 sg13g2_mux2_1 _18422_ (.A0(\top_ihp.oisc.regs[46][6] ),
    .A1(net98),
    .S(net367),
    .X(_01792_));
 sg13g2_nand2_1 _18423_ (.Y(_02982_),
    .A(\top_ihp.oisc.regs[46][7] ),
    .B(_02952_));
 sg13g2_o21ai_1 _18424_ (.B1(_02982_),
    .Y(_01793_),
    .A1(net210),
    .A2(net365));
 sg13g2_nand2_1 _18425_ (.Y(_02983_),
    .A(\top_ihp.oisc.regs[46][8] ),
    .B(_02952_));
 sg13g2_o21ai_1 _18426_ (.B1(_02983_),
    .Y(_01794_),
    .A1(net88),
    .A2(net365));
 sg13g2_mux2_1 _18427_ (.A0(\top_ihp.oisc.regs[46][9] ),
    .A1(_11296_),
    .S(_02950_),
    .X(_01795_));
 sg13g2_nand2_1 _18428_ (.Y(_02984_),
    .A(_10747_),
    .B(_02875_));
 sg13g2_buf_2 _18429_ (.A(_02984_),
    .X(_02985_));
 sg13g2_buf_2 _18430_ (.A(_02985_),
    .X(_02986_));
 sg13g2_mux2_1 _18431_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[47][0] ),
    .S(net362),
    .X(_01796_));
 sg13g2_mux2_1 _18432_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[47][10] ),
    .S(net362),
    .X(_01797_));
 sg13g2_buf_2 _18433_ (.A(_02985_),
    .X(_02987_));
 sg13g2_buf_1 _18434_ (.A(_02985_),
    .X(_02988_));
 sg13g2_nand2_1 _18435_ (.Y(_02989_),
    .A(\top_ihp.oisc.regs[47][11] ),
    .B(net360));
 sg13g2_o21ai_1 _18436_ (.B1(_02989_),
    .Y(_01798_),
    .A1(net49),
    .A2(net361));
 sg13g2_nand2_1 _18437_ (.Y(_02990_),
    .A(\top_ihp.oisc.regs[47][12] ),
    .B(net360));
 sg13g2_o21ai_1 _18438_ (.B1(_02990_),
    .Y(_01799_),
    .A1(net40),
    .A2(net361));
 sg13g2_nand2_1 _18439_ (.Y(_02991_),
    .A(\top_ihp.oisc.regs[47][13] ),
    .B(_02988_));
 sg13g2_o21ai_1 _18440_ (.B1(_02991_),
    .Y(_01800_),
    .A1(net96),
    .A2(net361));
 sg13g2_nand2_1 _18441_ (.Y(_02992_),
    .A(\top_ihp.oisc.regs[47][14] ),
    .B(net360));
 sg13g2_o21ai_1 _18442_ (.B1(_02992_),
    .Y(_01801_),
    .A1(net95),
    .A2(_02987_));
 sg13g2_mux2_1 _18443_ (.A0(net663),
    .A1(\top_ihp.oisc.regs[47][15] ),
    .S(net362),
    .X(_01802_));
 sg13g2_nand2_1 _18444_ (.Y(_02993_),
    .A(\top_ihp.oisc.regs[47][16] ),
    .B(_02988_));
 sg13g2_o21ai_1 _18445_ (.B1(_02993_),
    .Y(_01803_),
    .A1(net94),
    .A2(_02987_));
 sg13g2_nand2_1 _18446_ (.Y(_02994_),
    .A(\top_ihp.oisc.regs[47][17] ),
    .B(net360));
 sg13g2_o21ai_1 _18447_ (.B1(_02994_),
    .Y(_01804_),
    .A1(net212),
    .A2(net361));
 sg13g2_nand2_1 _18448_ (.Y(_02995_),
    .A(\top_ihp.oisc.regs[47][18] ),
    .B(net360));
 sg13g2_o21ai_1 _18449_ (.B1(_02995_),
    .Y(_01805_),
    .A1(net93),
    .A2(net361));
 sg13g2_mux2_1 _18450_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[47][19] ),
    .S(net362),
    .X(_01806_));
 sg13g2_nand2_1 _18451_ (.Y(_02996_),
    .A(\top_ihp.oisc.regs[47][1] ),
    .B(net360));
 sg13g2_o21ai_1 _18452_ (.B1(_02996_),
    .Y(_01807_),
    .A1(net105),
    .A2(net361));
 sg13g2_buf_1 _18453_ (.A(_02985_),
    .X(_02997_));
 sg13g2_nand2_1 _18454_ (.Y(_02998_),
    .A(\top_ihp.oisc.regs[47][20] ),
    .B(_02997_));
 sg13g2_o21ai_1 _18455_ (.B1(_02998_),
    .Y(_01808_),
    .A1(net39),
    .A2(net361));
 sg13g2_nand2_1 _18456_ (.Y(_02999_),
    .A(\top_ihp.oisc.regs[47][21] ),
    .B(_02997_));
 sg13g2_o21ai_1 _18457_ (.B1(_02999_),
    .Y(_01809_),
    .A1(net92),
    .A2(net361));
 sg13g2_buf_2 _18458_ (.A(_02985_),
    .X(_03000_));
 sg13g2_nand2_1 _18459_ (.Y(_03001_),
    .A(\top_ihp.oisc.regs[47][22] ),
    .B(net359));
 sg13g2_o21ai_1 _18460_ (.B1(_03001_),
    .Y(_01810_),
    .A1(net91),
    .A2(net358));
 sg13g2_nand2_1 _18461_ (.Y(_03002_),
    .A(\top_ihp.oisc.regs[47][23] ),
    .B(net359));
 sg13g2_o21ai_1 _18462_ (.B1(_03002_),
    .Y(_01811_),
    .A1(net90),
    .A2(_03000_));
 sg13g2_mux2_1 _18463_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[47][24] ),
    .S(net362),
    .X(_01812_));
 sg13g2_nand2_1 _18464_ (.Y(_03003_),
    .A(\top_ihp.oisc.regs[47][25] ),
    .B(net359));
 sg13g2_o21ai_1 _18465_ (.B1(_03003_),
    .Y(_01813_),
    .A1(net213),
    .A2(net358));
 sg13g2_nand2_1 _18466_ (.Y(_03004_),
    .A(\top_ihp.oisc.regs[47][26] ),
    .B(net359));
 sg13g2_o21ai_1 _18467_ (.B1(_03004_),
    .Y(_01814_),
    .A1(net211),
    .A2(net358));
 sg13g2_mux2_1 _18468_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[47][27] ),
    .S(net362),
    .X(_01815_));
 sg13g2_nand2_1 _18469_ (.Y(_03005_),
    .A(\top_ihp.oisc.regs[47][28] ),
    .B(net359));
 sg13g2_o21ai_1 _18470_ (.B1(_03005_),
    .Y(_01816_),
    .A1(net27),
    .A2(net358));
 sg13g2_nand2_1 _18471_ (.Y(_03006_),
    .A(\top_ihp.oisc.regs[47][29] ),
    .B(net359));
 sg13g2_o21ai_1 _18472_ (.B1(_03006_),
    .Y(_01817_),
    .A1(net89),
    .A2(net358));
 sg13g2_nand2_1 _18473_ (.Y(_03007_),
    .A(\top_ihp.oisc.regs[47][2] ),
    .B(net359));
 sg13g2_o21ai_1 _18474_ (.B1(_03007_),
    .Y(_01818_),
    .A1(net38),
    .A2(net358));
 sg13g2_nand2_1 _18475_ (.Y(_03008_),
    .A(\top_ihp.oisc.regs[47][30] ),
    .B(net359));
 sg13g2_o21ai_1 _18476_ (.B1(_03008_),
    .Y(_01819_),
    .A1(net26),
    .A2(net358));
 sg13g2_nand2_1 _18477_ (.Y(_03009_),
    .A(\top_ihp.oisc.regs[47][31] ),
    .B(_02985_));
 sg13g2_o21ai_1 _18478_ (.B1(_03009_),
    .Y(_01820_),
    .A1(net106),
    .A2(_03000_));
 sg13g2_mux2_1 _18479_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[47][3] ),
    .S(_02986_),
    .X(_01821_));
 sg13g2_mux2_1 _18480_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[47][4] ),
    .S(net362),
    .X(_01822_));
 sg13g2_mux2_1 _18481_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[47][5] ),
    .S(_02986_),
    .X(_01823_));
 sg13g2_mux2_1 _18482_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[47][6] ),
    .S(net360),
    .X(_01824_));
 sg13g2_nand2_1 _18483_ (.Y(_03010_),
    .A(\top_ihp.oisc.regs[47][7] ),
    .B(_02985_));
 sg13g2_o21ai_1 _18484_ (.B1(_03010_),
    .Y(_01825_),
    .A1(net210),
    .A2(net358));
 sg13g2_nand2_1 _18485_ (.Y(_03011_),
    .A(\top_ihp.oisc.regs[47][8] ),
    .B(_02985_));
 sg13g2_o21ai_1 _18486_ (.B1(_03011_),
    .Y(_01826_),
    .A1(net88),
    .A2(net362));
 sg13g2_mux2_1 _18487_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[47][9] ),
    .S(net360),
    .X(_01827_));
 sg13g2_nor2b_1 _18488_ (.A(_09921_),
    .B_N(_09926_),
    .Y(_03012_));
 sg13g2_buf_1 _18489_ (.A(_03012_),
    .X(_03013_));
 sg13g2_and2_1 _18490_ (.A(_09939_),
    .B(_03013_),
    .X(_03014_));
 sg13g2_buf_1 _18491_ (.A(_03014_),
    .X(_03015_));
 sg13g2_nand2_1 _18492_ (.Y(_03016_),
    .A(net692),
    .B(_03015_));
 sg13g2_buf_1 _18493_ (.A(_03016_),
    .X(_03017_));
 sg13g2_buf_2 _18494_ (.A(net539),
    .X(_03018_));
 sg13g2_mux2_1 _18495_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[48][0] ),
    .S(net357),
    .X(_01828_));
 sg13g2_mux2_1 _18496_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[48][10] ),
    .S(net357),
    .X(_01829_));
 sg13g2_buf_1 _18497_ (.A(_10050_),
    .X(_03019_));
 sg13g2_buf_1 _18498_ (.A(net539),
    .X(_03020_));
 sg13g2_buf_1 _18499_ (.A(net539),
    .X(_03021_));
 sg13g2_nand2_1 _18500_ (.Y(_03022_),
    .A(\top_ihp.oisc.regs[48][11] ),
    .B(net355));
 sg13g2_o21ai_1 _18501_ (.B1(_03022_),
    .Y(_01830_),
    .A1(net37),
    .A2(net356));
 sg13g2_nand2_1 _18502_ (.Y(_03023_),
    .A(\top_ihp.oisc.regs[48][12] ),
    .B(net355));
 sg13g2_o21ai_1 _18503_ (.B1(_03023_),
    .Y(_01831_),
    .A1(net40),
    .A2(net356));
 sg13g2_nand2_1 _18504_ (.Y(_03024_),
    .A(\top_ihp.oisc.regs[48][13] ),
    .B(net355));
 sg13g2_o21ai_1 _18505_ (.B1(_03024_),
    .Y(_01832_),
    .A1(net96),
    .A2(_03020_));
 sg13g2_nand2_1 _18506_ (.Y(_03025_),
    .A(\top_ihp.oisc.regs[48][14] ),
    .B(_03021_));
 sg13g2_o21ai_1 _18507_ (.B1(_03025_),
    .Y(_01833_),
    .A1(net95),
    .A2(net356));
 sg13g2_nand2_1 _18508_ (.Y(_03026_),
    .A(\top_ihp.oisc.regs[48][15] ),
    .B(net355));
 sg13g2_o21ai_1 _18509_ (.B1(_03026_),
    .Y(_01834_),
    .A1(net233),
    .A2(net356));
 sg13g2_nand2_1 _18510_ (.Y(_03027_),
    .A(\top_ihp.oisc.regs[48][16] ),
    .B(_03021_));
 sg13g2_o21ai_1 _18511_ (.B1(_03027_),
    .Y(_01835_),
    .A1(net94),
    .A2(net356));
 sg13g2_nand2_1 _18512_ (.Y(_03028_),
    .A(\top_ihp.oisc.regs[48][17] ),
    .B(net355));
 sg13g2_o21ai_1 _18513_ (.B1(_03028_),
    .Y(_01836_),
    .A1(net212),
    .A2(_03020_));
 sg13g2_nand2_1 _18514_ (.Y(_03029_),
    .A(\top_ihp.oisc.regs[48][18] ),
    .B(net355));
 sg13g2_o21ai_1 _18515_ (.B1(_03029_),
    .Y(_01837_),
    .A1(net93),
    .A2(net356));
 sg13g2_mux2_1 _18516_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[48][19] ),
    .S(net357),
    .X(_01838_));
 sg13g2_buf_1 _18517_ (.A(net539),
    .X(_03030_));
 sg13g2_nand2_1 _18518_ (.Y(_03031_),
    .A(\top_ihp.oisc.regs[48][1] ),
    .B(_03030_));
 sg13g2_o21ai_1 _18519_ (.B1(_03031_),
    .Y(_01839_),
    .A1(net105),
    .A2(net356));
 sg13g2_nand2_1 _18520_ (.Y(_03032_),
    .A(\top_ihp.oisc.regs[48][20] ),
    .B(_03030_));
 sg13g2_o21ai_1 _18521_ (.B1(_03032_),
    .Y(_01840_),
    .A1(_02924_),
    .A2(net356));
 sg13g2_buf_1 _18522_ (.A(net539),
    .X(_03033_));
 sg13g2_nand2_1 _18523_ (.Y(_03034_),
    .A(\top_ihp.oisc.regs[48][21] ),
    .B(net354));
 sg13g2_o21ai_1 _18524_ (.B1(_03034_),
    .Y(_01841_),
    .A1(net92),
    .A2(_03033_));
 sg13g2_nand2_1 _18525_ (.Y(_03035_),
    .A(\top_ihp.oisc.regs[48][22] ),
    .B(net354));
 sg13g2_o21ai_1 _18526_ (.B1(_03035_),
    .Y(_01842_),
    .A1(net91),
    .A2(net353));
 sg13g2_nand2_1 _18527_ (.Y(_03036_),
    .A(\top_ihp.oisc.regs[48][23] ),
    .B(net354));
 sg13g2_o21ai_1 _18528_ (.B1(_03036_),
    .Y(_01843_),
    .A1(net90),
    .A2(net353));
 sg13g2_mux2_1 _18529_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[48][24] ),
    .S(net357),
    .X(_01844_));
 sg13g2_nand2_1 _18530_ (.Y(_03037_),
    .A(\top_ihp.oisc.regs[48][25] ),
    .B(net354));
 sg13g2_o21ai_1 _18531_ (.B1(_03037_),
    .Y(_01845_),
    .A1(net213),
    .A2(net353));
 sg13g2_nand2_1 _18532_ (.Y(_03038_),
    .A(\top_ihp.oisc.regs[48][26] ),
    .B(net354));
 sg13g2_o21ai_1 _18533_ (.B1(_03038_),
    .Y(_01846_),
    .A1(net211),
    .A2(net353));
 sg13g2_mux2_1 _18534_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[48][27] ),
    .S(_03018_),
    .X(_01847_));
 sg13g2_nand2_1 _18535_ (.Y(_03039_),
    .A(\top_ihp.oisc.regs[48][28] ),
    .B(net354));
 sg13g2_o21ai_1 _18536_ (.B1(_03039_),
    .Y(_01848_),
    .A1(_02937_),
    .A2(net353));
 sg13g2_nand2_1 _18537_ (.Y(_03040_),
    .A(\top_ihp.oisc.regs[48][29] ),
    .B(net354));
 sg13g2_o21ai_1 _18538_ (.B1(_03040_),
    .Y(_01849_),
    .A1(net89),
    .A2(net353));
 sg13g2_nand2_1 _18539_ (.Y(_03041_),
    .A(\top_ihp.oisc.regs[48][2] ),
    .B(net354));
 sg13g2_o21ai_1 _18540_ (.B1(_03041_),
    .Y(_01850_),
    .A1(net38),
    .A2(net353));
 sg13g2_nand2_1 _18541_ (.Y(_03042_),
    .A(\top_ihp.oisc.regs[48][30] ),
    .B(net539));
 sg13g2_o21ai_1 _18542_ (.B1(_03042_),
    .Y(_01851_),
    .A1(_02978_),
    .A2(net353));
 sg13g2_nand2_1 _18543_ (.Y(_03043_),
    .A(\top_ihp.oisc.regs[48][31] ),
    .B(net539));
 sg13g2_o21ai_1 _18544_ (.B1(_03043_),
    .Y(_01852_),
    .A1(_11151_),
    .A2(_03033_));
 sg13g2_mux2_1 _18545_ (.A0(_11219_),
    .A1(\top_ihp.oisc.regs[48][3] ),
    .S(net357),
    .X(_01853_));
 sg13g2_mux2_1 _18546_ (.A0(_11220_),
    .A1(\top_ihp.oisc.regs[48][4] ),
    .S(_03018_),
    .X(_01854_));
 sg13g2_mux2_1 _18547_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[48][5] ),
    .S(net357),
    .X(_01855_));
 sg13g2_mux2_1 _18548_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[48][6] ),
    .S(net355),
    .X(_01856_));
 sg13g2_nand2_1 _18549_ (.Y(_03044_),
    .A(\top_ihp.oisc.regs[48][7] ),
    .B(_03017_));
 sg13g2_o21ai_1 _18550_ (.B1(_03044_),
    .Y(_01857_),
    .A1(_02944_),
    .A2(net357));
 sg13g2_nand2_1 _18551_ (.Y(_03045_),
    .A(\top_ihp.oisc.regs[48][8] ),
    .B(net539));
 sg13g2_o21ai_1 _18552_ (.B1(_03045_),
    .Y(_01858_),
    .A1(net88),
    .A2(net357));
 sg13g2_mux2_1 _18553_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[48][9] ),
    .S(net355),
    .X(_01859_));
 sg13g2_nand2_1 _18554_ (.Y(_03046_),
    .A(_10822_),
    .B(_03013_));
 sg13g2_buf_2 _18555_ (.A(_03046_),
    .X(_03047_));
 sg13g2_nor2_1 _18556_ (.A(_10912_),
    .B(_03047_),
    .Y(_03048_));
 sg13g2_buf_2 _18557_ (.A(_03048_),
    .X(_03049_));
 sg13g2_buf_2 _18558_ (.A(net653),
    .X(_03050_));
 sg13g2_mux2_1 _18559_ (.A0(\top_ihp.oisc.regs[49][0] ),
    .A1(net103),
    .S(net538),
    .X(_01860_));
 sg13g2_mux2_1 _18560_ (.A0(\top_ihp.oisc.regs[49][10] ),
    .A1(net102),
    .S(net538),
    .X(_01861_));
 sg13g2_nor2_1 _18561_ (.A(\top_ihp.oisc.regs[49][11] ),
    .B(net653),
    .Y(_03051_));
 sg13g2_a21oi_1 _18562_ (.A1(net50),
    .A2(net538),
    .Y(_01862_),
    .B1(_03051_));
 sg13g2_nor2_1 _18563_ (.A(\top_ihp.oisc.regs[49][12] ),
    .B(net653),
    .Y(_03052_));
 sg13g2_a21oi_1 _18564_ (.A1(net52),
    .A2(net538),
    .Y(_01863_),
    .B1(_03052_));
 sg13g2_nand2b_1 _18565_ (.Y(_03053_),
    .B(net692),
    .A_N(_03047_));
 sg13g2_buf_2 _18566_ (.A(_03053_),
    .X(_03054_));
 sg13g2_buf_2 _18567_ (.A(_03054_),
    .X(_03055_));
 sg13g2_buf_2 _18568_ (.A(_03054_),
    .X(_03056_));
 sg13g2_nand2_1 _18569_ (.Y(_03057_),
    .A(\top_ihp.oisc.regs[49][13] ),
    .B(net351));
 sg13g2_o21ai_1 _18570_ (.B1(_03057_),
    .Y(_01864_),
    .A1(net96),
    .A2(net352));
 sg13g2_nand2_1 _18571_ (.Y(_03058_),
    .A(\top_ihp.oisc.regs[49][14] ),
    .B(_03056_));
 sg13g2_o21ai_1 _18572_ (.B1(_03058_),
    .Y(_01865_),
    .A1(net95),
    .A2(_03055_));
 sg13g2_mux2_1 _18573_ (.A0(\top_ihp.oisc.regs[49][15] ),
    .A1(net663),
    .S(net538),
    .X(_01866_));
 sg13g2_nand2_1 _18574_ (.Y(_03059_),
    .A(\top_ihp.oisc.regs[49][16] ),
    .B(_03056_));
 sg13g2_o21ai_1 _18575_ (.B1(_03059_),
    .Y(_01867_),
    .A1(net94),
    .A2(_03055_));
 sg13g2_buf_2 _18576_ (.A(_03054_),
    .X(_03060_));
 sg13g2_nand2_1 _18577_ (.Y(_03061_),
    .A(\top_ihp.oisc.regs[49][17] ),
    .B(_03060_));
 sg13g2_o21ai_1 _18578_ (.B1(_03061_),
    .Y(_01868_),
    .A1(net212),
    .A2(net352));
 sg13g2_nand2_1 _18579_ (.Y(_03062_),
    .A(\top_ihp.oisc.regs[49][18] ),
    .B(net350));
 sg13g2_o21ai_1 _18580_ (.B1(_03062_),
    .Y(_01869_),
    .A1(net93),
    .A2(net352));
 sg13g2_mux2_1 _18581_ (.A0(\top_ihp.oisc.regs[49][19] ),
    .A1(net227),
    .S(_03050_),
    .X(_01870_));
 sg13g2_nor2_1 _18582_ (.A(\top_ihp.oisc.regs[49][1] ),
    .B(net653),
    .Y(_03063_));
 sg13g2_a21oi_1 _18583_ (.A1(net118),
    .A2(net538),
    .Y(_01871_),
    .B1(_03063_));
 sg13g2_nand2_1 _18584_ (.Y(_03064_),
    .A(\top_ihp.oisc.regs[49][20] ),
    .B(net350));
 sg13g2_o21ai_1 _18585_ (.B1(_03064_),
    .Y(_01872_),
    .A1(net39),
    .A2(net352));
 sg13g2_nand2_1 _18586_ (.Y(_03065_),
    .A(\top_ihp.oisc.regs[49][21] ),
    .B(net350));
 sg13g2_o21ai_1 _18587_ (.B1(_03065_),
    .Y(_01873_),
    .A1(net92),
    .A2(net352));
 sg13g2_nand2_1 _18588_ (.Y(_03066_),
    .A(\top_ihp.oisc.regs[49][22] ),
    .B(net350));
 sg13g2_o21ai_1 _18589_ (.B1(_03066_),
    .Y(_01874_),
    .A1(net91),
    .A2(net352));
 sg13g2_nand2_1 _18590_ (.Y(_03067_),
    .A(\top_ihp.oisc.regs[49][23] ),
    .B(net350));
 sg13g2_o21ai_1 _18591_ (.B1(_03067_),
    .Y(_01875_),
    .A1(net90),
    .A2(net352));
 sg13g2_mux2_1 _18592_ (.A0(\top_ihp.oisc.regs[49][24] ),
    .A1(net382),
    .S(net538),
    .X(_01876_));
 sg13g2_nand2_1 _18593_ (.Y(_03068_),
    .A(\top_ihp.oisc.regs[49][25] ),
    .B(net350));
 sg13g2_o21ai_1 _18594_ (.B1(_03068_),
    .Y(_01877_),
    .A1(_11380_),
    .A2(net352));
 sg13g2_nand2_1 _18595_ (.Y(_03069_),
    .A(\top_ihp.oisc.regs[49][26] ),
    .B(net350));
 sg13g2_o21ai_1 _18596_ (.B1(_03069_),
    .Y(_01878_),
    .A1(net211),
    .A2(net351));
 sg13g2_mux2_1 _18597_ (.A0(\top_ihp.oisc.regs[49][27] ),
    .A1(_11284_),
    .S(_03050_),
    .X(_01879_));
 sg13g2_nor2_1 _18598_ (.A(\top_ihp.oisc.regs[49][28] ),
    .B(net653),
    .Y(_03070_));
 sg13g2_a21oi_1 _18599_ (.A1(net116),
    .A2(net538),
    .Y(_01880_),
    .B1(_03070_));
 sg13g2_nand2_1 _18600_ (.Y(_03071_),
    .A(\top_ihp.oisc.regs[49][29] ),
    .B(net350));
 sg13g2_o21ai_1 _18601_ (.B1(_03071_),
    .Y(_01881_),
    .A1(net89),
    .A2(net351));
 sg13g2_nand2_1 _18602_ (.Y(_03072_),
    .A(\top_ihp.oisc.regs[49][2] ),
    .B(_03060_));
 sg13g2_o21ai_1 _18603_ (.B1(_03072_),
    .Y(_01882_),
    .A1(_02976_),
    .A2(net351));
 sg13g2_nand2_1 _18604_ (.Y(_03073_),
    .A(\top_ihp.oisc.regs[49][30] ),
    .B(_03054_));
 sg13g2_o21ai_1 _18605_ (.B1(_03073_),
    .Y(_01883_),
    .A1(net26),
    .A2(net351));
 sg13g2_buf_1 _18606_ (.A(_10737_),
    .X(_03074_));
 sg13g2_nand2_1 _18607_ (.Y(_03075_),
    .A(\top_ihp.oisc.regs[49][31] ),
    .B(_03054_));
 sg13g2_o21ai_1 _18608_ (.B1(_03075_),
    .Y(_01884_),
    .A1(net87),
    .A2(net351));
 sg13g2_mux2_1 _18609_ (.A0(\top_ihp.oisc.regs[49][3] ),
    .A1(net100),
    .S(_03049_),
    .X(_01885_));
 sg13g2_mux2_1 _18610_ (.A0(\top_ihp.oisc.regs[49][4] ),
    .A1(_11291_),
    .S(_03049_),
    .X(_01886_));
 sg13g2_mux2_1 _18611_ (.A0(\top_ihp.oisc.regs[49][5] ),
    .A1(_11292_),
    .S(net653),
    .X(_01887_));
 sg13g2_mux2_1 _18612_ (.A0(\top_ihp.oisc.regs[49][6] ),
    .A1(_11293_),
    .S(net653),
    .X(_01888_));
 sg13g2_nand2_1 _18613_ (.Y(_03076_),
    .A(\top_ihp.oisc.regs[49][7] ),
    .B(_03054_));
 sg13g2_o21ai_1 _18614_ (.B1(_03076_),
    .Y(_01889_),
    .A1(net210),
    .A2(net351));
 sg13g2_nand2_1 _18615_ (.Y(_03077_),
    .A(\top_ihp.oisc.regs[49][8] ),
    .B(_03054_));
 sg13g2_o21ai_1 _18616_ (.B1(_03077_),
    .Y(_01890_),
    .A1(net88),
    .A2(net351));
 sg13g2_mux2_1 _18617_ (.A0(\top_ihp.oisc.regs[49][9] ),
    .A1(net97),
    .S(net653),
    .X(_01891_));
 sg13g2_nor3_1 _18618_ (.A(_09910_),
    .B(_11077_),
    .C(_11078_),
    .Y(_03078_));
 sg13g2_buf_2 _18619_ (.A(_03078_),
    .X(_03079_));
 sg13g2_nand2_1 _18620_ (.Y(_03080_),
    .A(_09941_),
    .B(net729));
 sg13g2_buf_1 _18621_ (.A(_03080_),
    .X(_03081_));
 sg13g2_buf_1 _18622_ (.A(net652),
    .X(_03082_));
 sg13g2_mux2_1 _18623_ (.A0(_11155_),
    .A1(\top_ihp.oisc.regs[4][0] ),
    .S(net537),
    .X(_01892_));
 sg13g2_mux2_1 _18624_ (.A0(_11192_),
    .A1(\top_ihp.oisc.regs[4][10] ),
    .S(net537),
    .X(_01893_));
 sg13g2_buf_1 _18625_ (.A(net652),
    .X(_03083_));
 sg13g2_buf_1 _18626_ (.A(_03080_),
    .X(_03084_));
 sg13g2_nand2_1 _18627_ (.Y(_03085_),
    .A(\top_ihp.oisc.regs[4][11] ),
    .B(net651));
 sg13g2_o21ai_1 _18628_ (.B1(_03085_),
    .Y(_01894_),
    .A1(net37),
    .A2(net536));
 sg13g2_nand2_1 _18629_ (.Y(_03086_),
    .A(\top_ihp.oisc.regs[4][12] ),
    .B(net651));
 sg13g2_o21ai_1 _18630_ (.B1(_03086_),
    .Y(_01895_),
    .A1(_11303_),
    .A2(net536));
 sg13g2_nand2_1 _18631_ (.Y(_03087_),
    .A(\top_ihp.oisc.regs[4][13] ),
    .B(net651));
 sg13g2_o21ai_1 _18632_ (.B1(_03087_),
    .Y(_01896_),
    .A1(_02913_),
    .A2(net536));
 sg13g2_nand2_1 _18633_ (.Y(_03088_),
    .A(\top_ihp.oisc.regs[4][14] ),
    .B(net651));
 sg13g2_o21ai_1 _18634_ (.B1(_03088_),
    .Y(_01897_),
    .A1(_02915_),
    .A2(net536));
 sg13g2_nand2_1 _18635_ (.Y(_03089_),
    .A(\top_ihp.oisc.regs[4][15] ),
    .B(net651));
 sg13g2_o21ai_1 _18636_ (.B1(_03089_),
    .Y(_01898_),
    .A1(_11165_),
    .A2(net536));
 sg13g2_nand2_1 _18637_ (.Y(_03090_),
    .A(\top_ihp.oisc.regs[4][16] ),
    .B(net651));
 sg13g2_o21ai_1 _18638_ (.B1(_03090_),
    .Y(_01899_),
    .A1(_02917_),
    .A2(net536));
 sg13g2_nand2_1 _18639_ (.Y(_03091_),
    .A(\top_ihp.oisc.regs[4][17] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18640_ (.B1(_03091_),
    .Y(_01900_),
    .A1(_02919_),
    .A2(_03083_));
 sg13g2_nand2_1 _18641_ (.Y(_03092_),
    .A(\top_ihp.oisc.regs[4][18] ),
    .B(_03084_));
 sg13g2_o21ai_1 _18642_ (.B1(_03092_),
    .Y(_01901_),
    .A1(_02921_),
    .A2(_03083_));
 sg13g2_buf_1 _18643_ (.A(net652),
    .X(_03093_));
 sg13g2_nand2_1 _18644_ (.Y(_03094_),
    .A(\top_ihp.oisc.regs[4][19] ),
    .B(net535));
 sg13g2_o21ai_1 _18645_ (.B1(_03094_),
    .Y(_01902_),
    .A1(_10274_),
    .A2(net536));
 sg13g2_buf_1 _18646_ (.A(net652),
    .X(_03095_));
 sg13g2_nand2_1 _18647_ (.Y(_03096_),
    .A(\top_ihp.oisc.regs[4][1] ),
    .B(net535));
 sg13g2_o21ai_1 _18648_ (.B1(_03096_),
    .Y(_01903_),
    .A1(_11203_),
    .A2(net534));
 sg13g2_nand2_1 _18649_ (.Y(_03097_),
    .A(\top_ihp.oisc.regs[4][20] ),
    .B(net535));
 sg13g2_o21ai_1 _18650_ (.B1(_03097_),
    .Y(_01904_),
    .A1(_02924_),
    .A2(net534));
 sg13g2_nand2_1 _18651_ (.Y(_03098_),
    .A(\top_ihp.oisc.regs[4][21] ),
    .B(net535));
 sg13g2_o21ai_1 _18652_ (.B1(_03098_),
    .Y(_01905_),
    .A1(_02927_),
    .A2(net534));
 sg13g2_nand2_1 _18653_ (.Y(_03099_),
    .A(\top_ihp.oisc.regs[4][22] ),
    .B(_03093_));
 sg13g2_o21ai_1 _18654_ (.B1(_03099_),
    .Y(_01906_),
    .A1(_02929_),
    .A2(net534));
 sg13g2_nand2_1 _18655_ (.Y(_03100_),
    .A(\top_ihp.oisc.regs[4][23] ),
    .B(net535));
 sg13g2_o21ai_1 _18656_ (.B1(_03100_),
    .Y(_01907_),
    .A1(net90),
    .A2(_03095_));
 sg13g2_mux2_1 _18657_ (.A0(_11211_),
    .A1(\top_ihp.oisc.regs[4][24] ),
    .S(net537),
    .X(_01908_));
 sg13g2_nand2_1 _18658_ (.Y(_03101_),
    .A(\top_ihp.oisc.regs[4][25] ),
    .B(net535));
 sg13g2_o21ai_1 _18659_ (.B1(_03101_),
    .Y(_01909_),
    .A1(_10428_),
    .A2(_03095_));
 sg13g2_nand2_1 _18660_ (.Y(_03102_),
    .A(\top_ihp.oisc.regs[4][26] ),
    .B(_03093_));
 sg13g2_o21ai_1 _18661_ (.B1(_03102_),
    .Y(_01910_),
    .A1(_02935_),
    .A2(net534));
 sg13g2_nand2_1 _18662_ (.Y(_03103_),
    .A(\top_ihp.oisc.regs[4][27] ),
    .B(net535));
 sg13g2_o21ai_1 _18663_ (.B1(_03103_),
    .Y(_01911_),
    .A1(_10450_),
    .A2(net534));
 sg13g2_nand2_1 _18664_ (.Y(_03104_),
    .A(\top_ihp.oisc.regs[4][28] ),
    .B(net535));
 sg13g2_o21ai_1 _18665_ (.B1(_03104_),
    .Y(_01912_),
    .A1(_02937_),
    .A2(net534));
 sg13g2_nand2_1 _18666_ (.Y(_03105_),
    .A(\top_ihp.oisc.regs[4][29] ),
    .B(_03081_));
 sg13g2_o21ai_1 _18667_ (.B1(_03105_),
    .Y(_01913_),
    .A1(_02939_),
    .A2(net534));
 sg13g2_nand2_1 _18668_ (.Y(_03106_),
    .A(\top_ihp.oisc.regs[4][2] ),
    .B(_03081_));
 sg13g2_o21ai_1 _18669_ (.B1(_03106_),
    .Y(_01914_),
    .A1(_02976_),
    .A2(net537));
 sg13g2_nand2_1 _18670_ (.Y(_03107_),
    .A(\top_ihp.oisc.regs[4][30] ),
    .B(net652));
 sg13g2_o21ai_1 _18671_ (.B1(_03107_),
    .Y(_01915_),
    .A1(_02978_),
    .A2(net537));
 sg13g2_inv_1 _18672_ (.Y(_03108_),
    .A(\top_ihp.oisc.regs[4][31] ));
 sg13g2_nor2_1 _18673_ (.A(_10536_),
    .B(net652),
    .Y(_03109_));
 sg13g2_a22oi_1 _18674_ (.Y(_01916_),
    .B1(_03109_),
    .B2(_10738_),
    .A2(net536),
    .A1(_03108_));
 sg13g2_mux2_1 _18675_ (.A0(_11219_),
    .A1(\top_ihp.oisc.regs[4][3] ),
    .S(net537),
    .X(_01917_));
 sg13g2_mux2_1 _18676_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[4][4] ),
    .S(net537),
    .X(_01918_));
 sg13g2_mux2_1 _18677_ (.A0(_11221_),
    .A1(\top_ihp.oisc.regs[4][5] ),
    .S(net537),
    .X(_01919_));
 sg13g2_mux2_1 _18678_ (.A0(_11222_),
    .A1(\top_ihp.oisc.regs[4][6] ),
    .S(net651),
    .X(_01920_));
 sg13g2_nand2_1 _18679_ (.Y(_03110_),
    .A(\top_ihp.oisc.regs[4][7] ),
    .B(net652));
 sg13g2_o21ai_1 _18680_ (.B1(_03110_),
    .Y(_01921_),
    .A1(_02944_),
    .A2(_03082_));
 sg13g2_nand2_1 _18681_ (.Y(_03111_),
    .A(\top_ihp.oisc.regs[4][8] ),
    .B(net652));
 sg13g2_o21ai_1 _18682_ (.B1(_03111_),
    .Y(_01922_),
    .A1(_02946_),
    .A2(_03082_));
 sg13g2_mux2_1 _18683_ (.A0(_11225_),
    .A1(\top_ihp.oisc.regs[4][9] ),
    .S(net651),
    .X(_01923_));
 sg13g2_nand2_1 _18684_ (.Y(_03112_),
    .A(net740),
    .B(_03013_));
 sg13g2_nor2_1 _18685_ (.A(_10912_),
    .B(_03112_),
    .Y(_03113_));
 sg13g2_buf_1 _18686_ (.A(_03113_),
    .X(_03114_));
 sg13g2_buf_2 _18687_ (.A(net650),
    .X(_03115_));
 sg13g2_mux2_1 _18688_ (.A0(\top_ihp.oisc.regs[50][0] ),
    .A1(net103),
    .S(_03115_),
    .X(_01924_));
 sg13g2_mux2_1 _18689_ (.A0(\top_ihp.oisc.regs[50][10] ),
    .A1(net102),
    .S(net533),
    .X(_01925_));
 sg13g2_nor2_1 _18690_ (.A(\top_ihp.oisc.regs[50][11] ),
    .B(net650),
    .Y(_03116_));
 sg13g2_a21oi_1 _18691_ (.A1(net50),
    .A2(net533),
    .Y(_01926_),
    .B1(_03116_));
 sg13g2_nor2_1 _18692_ (.A(\top_ihp.oisc.regs[50][12] ),
    .B(net650),
    .Y(_03117_));
 sg13g2_a21oi_1 _18693_ (.A1(net52),
    .A2(net533),
    .Y(_01927_),
    .B1(_03117_));
 sg13g2_and2_1 _18694_ (.A(net740),
    .B(_03013_),
    .X(_03118_));
 sg13g2_buf_1 _18695_ (.A(_03118_),
    .X(_03119_));
 sg13g2_nand2_1 _18696_ (.Y(_03120_),
    .A(net692),
    .B(_03119_));
 sg13g2_buf_1 _18697_ (.A(_03120_),
    .X(_03121_));
 sg13g2_buf_1 _18698_ (.A(net532),
    .X(_03122_));
 sg13g2_buf_1 _18699_ (.A(_03120_),
    .X(_03123_));
 sg13g2_nand2_1 _18700_ (.Y(_03124_),
    .A(\top_ihp.oisc.regs[50][13] ),
    .B(_03123_));
 sg13g2_o21ai_1 _18701_ (.B1(_03124_),
    .Y(_01928_),
    .A1(net96),
    .A2(net349));
 sg13g2_buf_1 _18702_ (.A(net532),
    .X(_03125_));
 sg13g2_nand2_1 _18703_ (.Y(_03126_),
    .A(\top_ihp.oisc.regs[50][14] ),
    .B(_03125_));
 sg13g2_o21ai_1 _18704_ (.B1(_03126_),
    .Y(_01929_),
    .A1(net95),
    .A2(_03122_));
 sg13g2_buf_1 _18705_ (.A(net399),
    .X(_03127_));
 sg13g2_nand2_1 _18706_ (.Y(_03128_),
    .A(\top_ihp.oisc.regs[50][15] ),
    .B(net348));
 sg13g2_o21ai_1 _18707_ (.B1(_03128_),
    .Y(_01930_),
    .A1(net209),
    .A2(net349));
 sg13g2_nand2_1 _18708_ (.Y(_03129_),
    .A(\top_ihp.oisc.regs[50][16] ),
    .B(net348));
 sg13g2_o21ai_1 _18709_ (.B1(_03129_),
    .Y(_01931_),
    .A1(net94),
    .A2(_03122_));
 sg13g2_nand2_1 _18710_ (.Y(_03130_),
    .A(\top_ihp.oisc.regs[50][17] ),
    .B(net348));
 sg13g2_o21ai_1 _18711_ (.B1(_03130_),
    .Y(_01932_),
    .A1(net212),
    .A2(net349));
 sg13g2_nand2_1 _18712_ (.Y(_03131_),
    .A(\top_ihp.oisc.regs[50][18] ),
    .B(_03125_));
 sg13g2_o21ai_1 _18713_ (.B1(_03131_),
    .Y(_01933_),
    .A1(_02921_),
    .A2(net349));
 sg13g2_nand2_1 _18714_ (.Y(_03132_),
    .A(\top_ihp.oisc.regs[50][19] ),
    .B(net348));
 sg13g2_o21ai_1 _18715_ (.B1(_03132_),
    .Y(_01934_),
    .A1(net60),
    .A2(net349));
 sg13g2_nor2_1 _18716_ (.A(\top_ihp.oisc.regs[50][1] ),
    .B(_03114_),
    .Y(_03133_));
 sg13g2_a21oi_1 _18717_ (.A1(net118),
    .A2(net533),
    .Y(_01935_),
    .B1(_03133_));
 sg13g2_nand2_1 _18718_ (.Y(_03134_),
    .A(\top_ihp.oisc.regs[50][20] ),
    .B(net348));
 sg13g2_o21ai_1 _18719_ (.B1(_03134_),
    .Y(_01936_),
    .A1(net39),
    .A2(net349));
 sg13g2_nand2_1 _18720_ (.Y(_03135_),
    .A(\top_ihp.oisc.regs[50][21] ),
    .B(net348));
 sg13g2_o21ai_1 _18721_ (.B1(_03135_),
    .Y(_01937_),
    .A1(_02927_),
    .A2(net349));
 sg13g2_nand2_1 _18722_ (.Y(_03136_),
    .A(\top_ihp.oisc.regs[50][22] ),
    .B(net348));
 sg13g2_o21ai_1 _18723_ (.B1(_03136_),
    .Y(_01938_),
    .A1(net91),
    .A2(net531));
 sg13g2_nand2_1 _18724_ (.Y(_03137_),
    .A(\top_ihp.oisc.regs[50][23] ),
    .B(net348));
 sg13g2_o21ai_1 _18725_ (.B1(_03137_),
    .Y(_01939_),
    .A1(_02932_),
    .A2(_03123_));
 sg13g2_mux2_1 _18726_ (.A0(\top_ihp.oisc.regs[50][24] ),
    .A1(net382),
    .S(net533),
    .X(_01940_));
 sg13g2_nor2_1 _18727_ (.A(\top_ihp.oisc.regs[50][25] ),
    .B(net650),
    .Y(_03138_));
 sg13g2_a21oi_1 _18728_ (.A1(net59),
    .A2(net533),
    .Y(_01941_),
    .B1(_03138_));
 sg13g2_nand2_1 _18729_ (.Y(_03139_),
    .A(\top_ihp.oisc.regs[50][26] ),
    .B(net532));
 sg13g2_o21ai_1 _18730_ (.B1(_03139_),
    .Y(_01942_),
    .A1(net211),
    .A2(net531));
 sg13g2_nand2_1 _18731_ (.Y(_03140_),
    .A(\top_ihp.oisc.regs[50][27] ),
    .B(net532));
 sg13g2_o21ai_1 _18732_ (.B1(_03140_),
    .Y(_01943_),
    .A1(net31),
    .A2(net531));
 sg13g2_nor2_1 _18733_ (.A(\top_ihp.oisc.regs[50][28] ),
    .B(net650),
    .Y(_03141_));
 sg13g2_a21oi_1 _18734_ (.A1(net30),
    .A2(net533),
    .Y(_01944_),
    .B1(_03141_));
 sg13g2_nand2_1 _18735_ (.Y(_03142_),
    .A(\top_ihp.oisc.regs[50][29] ),
    .B(net532));
 sg13g2_o21ai_1 _18736_ (.B1(_03142_),
    .Y(_01945_),
    .A1(net89),
    .A2(net531));
 sg13g2_nand2_1 _18737_ (.Y(_03143_),
    .A(\top_ihp.oisc.regs[50][2] ),
    .B(net532));
 sg13g2_o21ai_1 _18738_ (.B1(_03143_),
    .Y(_01946_),
    .A1(net38),
    .A2(net531));
 sg13g2_nand2_1 _18739_ (.Y(_03144_),
    .A(\top_ihp.oisc.regs[50][30] ),
    .B(net532));
 sg13g2_o21ai_1 _18740_ (.B1(_03144_),
    .Y(_01947_),
    .A1(net26),
    .A2(net531));
 sg13g2_inv_1 _18741_ (.Y(_03145_),
    .A(\top_ihp.oisc.regs[50][31] ));
 sg13g2_nor2_1 _18742_ (.A(net821),
    .B(net532),
    .Y(_03146_));
 sg13g2_a22oi_1 _18743_ (.Y(_01948_),
    .B1(_03146_),
    .B2(net129),
    .A2(net349),
    .A1(_03145_));
 sg13g2_mux2_1 _18744_ (.A0(\top_ihp.oisc.regs[50][3] ),
    .A1(net100),
    .S(_03115_),
    .X(_01949_));
 sg13g2_mux2_1 _18745_ (.A0(\top_ihp.oisc.regs[50][4] ),
    .A1(net99),
    .S(net533),
    .X(_01950_));
 sg13g2_mux2_1 _18746_ (.A0(\top_ihp.oisc.regs[50][5] ),
    .A1(net226),
    .S(net650),
    .X(_01951_));
 sg13g2_mux2_1 _18747_ (.A0(\top_ihp.oisc.regs[50][6] ),
    .A1(net98),
    .S(net650),
    .X(_01952_));
 sg13g2_nand2_1 _18748_ (.Y(_03147_),
    .A(\top_ihp.oisc.regs[50][7] ),
    .B(_03121_));
 sg13g2_o21ai_1 _18749_ (.B1(_03147_),
    .Y(_01953_),
    .A1(net210),
    .A2(net531));
 sg13g2_nand2_1 _18750_ (.Y(_03148_),
    .A(\top_ihp.oisc.regs[50][8] ),
    .B(_03121_));
 sg13g2_o21ai_1 _18751_ (.B1(_03148_),
    .Y(_01954_),
    .A1(net88),
    .A2(net531));
 sg13g2_mux2_1 _18752_ (.A0(\top_ihp.oisc.regs[50][9] ),
    .A1(_11296_),
    .S(net650),
    .X(_01955_));
 sg13g2_and2_1 _18753_ (.A(_10747_),
    .B(_03013_),
    .X(_03149_));
 sg13g2_buf_2 _18754_ (.A(_03149_),
    .X(_03150_));
 sg13g2_and2_1 _18755_ (.A(net692),
    .B(_03150_),
    .X(_03151_));
 sg13g2_buf_2 _18756_ (.A(_03151_),
    .X(_03152_));
 sg13g2_buf_2 _18757_ (.A(net530),
    .X(_03153_));
 sg13g2_mux2_1 _18758_ (.A0(\top_ihp.oisc.regs[51][0] ),
    .A1(net103),
    .S(_03153_),
    .X(_01956_));
 sg13g2_mux2_1 _18759_ (.A0(\top_ihp.oisc.regs[51][10] ),
    .A1(net102),
    .S(net347),
    .X(_01957_));
 sg13g2_nor2_1 _18760_ (.A(\top_ihp.oisc.regs[51][11] ),
    .B(net530),
    .Y(_03154_));
 sg13g2_a21oi_1 _18761_ (.A1(net50),
    .A2(net347),
    .Y(_01958_),
    .B1(_03154_));
 sg13g2_nor2_1 _18762_ (.A(\top_ihp.oisc.regs[51][12] ),
    .B(_03152_),
    .Y(_03155_));
 sg13g2_a21oi_1 _18763_ (.A1(net52),
    .A2(_03153_),
    .Y(_01959_),
    .B1(_03155_));
 sg13g2_nand2_1 _18764_ (.Y(_03156_),
    .A(net692),
    .B(_03150_));
 sg13g2_buf_2 _18765_ (.A(_03156_),
    .X(_03157_));
 sg13g2_buf_1 _18766_ (.A(_03157_),
    .X(_03158_));
 sg13g2_buf_2 _18767_ (.A(_03157_),
    .X(_03159_));
 sg13g2_nand2_1 _18768_ (.Y(_03160_),
    .A(\top_ihp.oisc.regs[51][13] ),
    .B(_03159_));
 sg13g2_o21ai_1 _18769_ (.B1(_03160_),
    .Y(_01960_),
    .A1(_02913_),
    .A2(net346));
 sg13g2_nand2_1 _18770_ (.Y(_03161_),
    .A(\top_ihp.oisc.regs[51][14] ),
    .B(_03159_));
 sg13g2_o21ai_1 _18771_ (.B1(_03161_),
    .Y(_01961_),
    .A1(net95),
    .A2(net346));
 sg13g2_mux2_1 _18772_ (.A0(\top_ihp.oisc.regs[51][15] ),
    .A1(net663),
    .S(net347),
    .X(_01962_));
 sg13g2_nand2_1 _18773_ (.Y(_03162_),
    .A(\top_ihp.oisc.regs[51][16] ),
    .B(net345));
 sg13g2_o21ai_1 _18774_ (.B1(_03162_),
    .Y(_01963_),
    .A1(net94),
    .A2(net346));
 sg13g2_buf_1 _18775_ (.A(_03157_),
    .X(_03163_));
 sg13g2_nand2_1 _18776_ (.Y(_03164_),
    .A(\top_ihp.oisc.regs[51][17] ),
    .B(_03163_));
 sg13g2_o21ai_1 _18777_ (.B1(_03164_),
    .Y(_01964_),
    .A1(net212),
    .A2(_03158_));
 sg13g2_nand2_1 _18778_ (.Y(_03165_),
    .A(\top_ihp.oisc.regs[51][18] ),
    .B(_03163_));
 sg13g2_o21ai_1 _18779_ (.B1(_03165_),
    .Y(_01965_),
    .A1(net93),
    .A2(_03158_));
 sg13g2_mux2_1 _18780_ (.A0(\top_ihp.oisc.regs[51][19] ),
    .A1(net227),
    .S(net347),
    .X(_01966_));
 sg13g2_nor2_1 _18781_ (.A(\top_ihp.oisc.regs[51][1] ),
    .B(net530),
    .Y(_03166_));
 sg13g2_a21oi_1 _18782_ (.A1(net118),
    .A2(net347),
    .Y(_01967_),
    .B1(_03166_));
 sg13g2_nand2_1 _18783_ (.Y(_03167_),
    .A(\top_ihp.oisc.regs[51][20] ),
    .B(net344));
 sg13g2_o21ai_1 _18784_ (.B1(_03167_),
    .Y(_01968_),
    .A1(net39),
    .A2(net346));
 sg13g2_nand2_1 _18785_ (.Y(_03168_),
    .A(\top_ihp.oisc.regs[51][21] ),
    .B(net344));
 sg13g2_o21ai_1 _18786_ (.B1(_03168_),
    .Y(_01969_),
    .A1(net92),
    .A2(net346));
 sg13g2_nand2_1 _18787_ (.Y(_03169_),
    .A(\top_ihp.oisc.regs[51][22] ),
    .B(net344));
 sg13g2_o21ai_1 _18788_ (.B1(_03169_),
    .Y(_01970_),
    .A1(net91),
    .A2(net346));
 sg13g2_nand2_1 _18789_ (.Y(_03170_),
    .A(\top_ihp.oisc.regs[51][23] ),
    .B(net344));
 sg13g2_o21ai_1 _18790_ (.B1(_03170_),
    .Y(_01971_),
    .A1(_02932_),
    .A2(net346));
 sg13g2_mux2_1 _18791_ (.A0(\top_ihp.oisc.regs[51][24] ),
    .A1(net382),
    .S(net347),
    .X(_01972_));
 sg13g2_nand2_1 _18792_ (.Y(_03171_),
    .A(\top_ihp.oisc.regs[51][25] ),
    .B(net344));
 sg13g2_o21ai_1 _18793_ (.B1(_03171_),
    .Y(_01973_),
    .A1(net213),
    .A2(net346));
 sg13g2_nand2_1 _18794_ (.Y(_03172_),
    .A(\top_ihp.oisc.regs[51][26] ),
    .B(net344));
 sg13g2_o21ai_1 _18795_ (.B1(_03172_),
    .Y(_01974_),
    .A1(net211),
    .A2(net345));
 sg13g2_mux2_1 _18796_ (.A0(\top_ihp.oisc.regs[51][27] ),
    .A1(net101),
    .S(net347),
    .X(_01975_));
 sg13g2_nor2_1 _18797_ (.A(\top_ihp.oisc.regs[51][28] ),
    .B(net530),
    .Y(_03173_));
 sg13g2_a21oi_1 _18798_ (.A1(net116),
    .A2(net347),
    .Y(_01976_),
    .B1(_03173_));
 sg13g2_nand2_1 _18799_ (.Y(_03174_),
    .A(\top_ihp.oisc.regs[51][29] ),
    .B(net344));
 sg13g2_o21ai_1 _18800_ (.B1(_03174_),
    .Y(_01977_),
    .A1(_02939_),
    .A2(net345));
 sg13g2_nand2_1 _18801_ (.Y(_03175_),
    .A(\top_ihp.oisc.regs[51][2] ),
    .B(net344));
 sg13g2_o21ai_1 _18802_ (.B1(_03175_),
    .Y(_01978_),
    .A1(net38),
    .A2(net345));
 sg13g2_nand2_1 _18803_ (.Y(_03176_),
    .A(\top_ihp.oisc.regs[51][30] ),
    .B(_03157_));
 sg13g2_o21ai_1 _18804_ (.B1(_03176_),
    .Y(_01979_),
    .A1(net26),
    .A2(net345));
 sg13g2_nand2_1 _18805_ (.Y(_03177_),
    .A(\top_ihp.oisc.regs[51][31] ),
    .B(_03157_));
 sg13g2_o21ai_1 _18806_ (.B1(_03177_),
    .Y(_01980_),
    .A1(net87),
    .A2(net345));
 sg13g2_mux2_1 _18807_ (.A0(\top_ihp.oisc.regs[51][3] ),
    .A1(_11290_),
    .S(net530),
    .X(_01981_));
 sg13g2_mux2_1 _18808_ (.A0(\top_ihp.oisc.regs[51][4] ),
    .A1(net99),
    .S(net530),
    .X(_01982_));
 sg13g2_mux2_1 _18809_ (.A0(\top_ihp.oisc.regs[51][5] ),
    .A1(net226),
    .S(_03152_),
    .X(_01983_));
 sg13g2_mux2_1 _18810_ (.A0(\top_ihp.oisc.regs[51][6] ),
    .A1(net98),
    .S(net530),
    .X(_01984_));
 sg13g2_nand2_1 _18811_ (.Y(_03178_),
    .A(\top_ihp.oisc.regs[51][7] ),
    .B(_03157_));
 sg13g2_o21ai_1 _18812_ (.B1(_03178_),
    .Y(_01985_),
    .A1(net210),
    .A2(net345));
 sg13g2_nand2_1 _18813_ (.Y(_03179_),
    .A(\top_ihp.oisc.regs[51][8] ),
    .B(_03157_));
 sg13g2_o21ai_1 _18814_ (.B1(_03179_),
    .Y(_01986_),
    .A1(_02946_),
    .A2(net345));
 sg13g2_mux2_1 _18815_ (.A0(\top_ihp.oisc.regs[51][9] ),
    .A1(net97),
    .S(net530),
    .X(_01987_));
 sg13g2_nand2_1 _18816_ (.Y(_03180_),
    .A(net729),
    .B(_03015_));
 sg13g2_buf_1 _18817_ (.A(_03180_),
    .X(_03181_));
 sg13g2_buf_2 _18818_ (.A(net649),
    .X(_03182_));
 sg13g2_mux2_1 _18819_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[52][0] ),
    .S(_03182_),
    .X(_01988_));
 sg13g2_mux2_1 _18820_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[52][10] ),
    .S(net529),
    .X(_01989_));
 sg13g2_buf_1 _18821_ (.A(net649),
    .X(_03183_));
 sg13g2_buf_2 _18822_ (.A(net649),
    .X(_03184_));
 sg13g2_nand2_1 _18823_ (.Y(_03185_),
    .A(\top_ihp.oisc.regs[52][11] ),
    .B(net527));
 sg13g2_o21ai_1 _18824_ (.B1(_03185_),
    .Y(_01990_),
    .A1(net37),
    .A2(net528));
 sg13g2_nand2_1 _18825_ (.Y(_03186_),
    .A(\top_ihp.oisc.regs[52][12] ),
    .B(net527));
 sg13g2_o21ai_1 _18826_ (.B1(_03186_),
    .Y(_01991_),
    .A1(net40),
    .A2(net528));
 sg13g2_nand2_1 _18827_ (.Y(_03187_),
    .A(\top_ihp.oisc.regs[52][13] ),
    .B(net527));
 sg13g2_o21ai_1 _18828_ (.B1(_03187_),
    .Y(_01992_),
    .A1(net96),
    .A2(net528));
 sg13g2_nand2_1 _18829_ (.Y(_03188_),
    .A(\top_ihp.oisc.regs[52][14] ),
    .B(net527));
 sg13g2_o21ai_1 _18830_ (.B1(_03188_),
    .Y(_01993_),
    .A1(_02915_),
    .A2(net528));
 sg13g2_nand2_1 _18831_ (.Y(_03189_),
    .A(\top_ihp.oisc.regs[52][15] ),
    .B(net527));
 sg13g2_o21ai_1 _18832_ (.B1(_03189_),
    .Y(_01994_),
    .A1(net209),
    .A2(net528));
 sg13g2_nand2_1 _18833_ (.Y(_03190_),
    .A(\top_ihp.oisc.regs[52][16] ),
    .B(_03184_));
 sg13g2_o21ai_1 _18834_ (.B1(_03190_),
    .Y(_01995_),
    .A1(_02917_),
    .A2(net528));
 sg13g2_nand2_1 _18835_ (.Y(_03191_),
    .A(\top_ihp.oisc.regs[52][17] ),
    .B(net527));
 sg13g2_o21ai_1 _18836_ (.B1(_03191_),
    .Y(_01996_),
    .A1(_02919_),
    .A2(_03183_));
 sg13g2_nand2_1 _18837_ (.Y(_03192_),
    .A(\top_ihp.oisc.regs[52][18] ),
    .B(net527));
 sg13g2_o21ai_1 _18838_ (.B1(_03192_),
    .Y(_01997_),
    .A1(net93),
    .A2(_03183_));
 sg13g2_mux2_1 _18839_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[52][19] ),
    .S(_03182_),
    .X(_01998_));
 sg13g2_buf_1 _18840_ (.A(net649),
    .X(_03193_));
 sg13g2_nand2_1 _18841_ (.Y(_03194_),
    .A(\top_ihp.oisc.regs[52][1] ),
    .B(_03193_));
 sg13g2_o21ai_1 _18842_ (.B1(_03194_),
    .Y(_01999_),
    .A1(net105),
    .A2(net528));
 sg13g2_nand2_1 _18843_ (.Y(_03195_),
    .A(\top_ihp.oisc.regs[52][20] ),
    .B(net526));
 sg13g2_o21ai_1 _18844_ (.B1(_03195_),
    .Y(_02000_),
    .A1(net39),
    .A2(net528));
 sg13g2_buf_1 _18845_ (.A(net649),
    .X(_03196_));
 sg13g2_nand2_1 _18846_ (.Y(_03197_),
    .A(\top_ihp.oisc.regs[52][21] ),
    .B(_03193_));
 sg13g2_o21ai_1 _18847_ (.B1(_03197_),
    .Y(_02001_),
    .A1(net92),
    .A2(net525));
 sg13g2_nand2_1 _18848_ (.Y(_03198_),
    .A(\top_ihp.oisc.regs[52][22] ),
    .B(net526));
 sg13g2_o21ai_1 _18849_ (.B1(_03198_),
    .Y(_02002_),
    .A1(net91),
    .A2(net525));
 sg13g2_nand2_1 _18850_ (.Y(_03199_),
    .A(\top_ihp.oisc.regs[52][23] ),
    .B(net526));
 sg13g2_o21ai_1 _18851_ (.B1(_03199_),
    .Y(_02003_),
    .A1(net90),
    .A2(net525));
 sg13g2_mux2_1 _18852_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[52][24] ),
    .S(net529),
    .X(_02004_));
 sg13g2_nand2_1 _18853_ (.Y(_03200_),
    .A(\top_ihp.oisc.regs[52][25] ),
    .B(net526));
 sg13g2_o21ai_1 _18854_ (.B1(_03200_),
    .Y(_02005_),
    .A1(net213),
    .A2(_03196_));
 sg13g2_nand2_1 _18855_ (.Y(_03201_),
    .A(\top_ihp.oisc.regs[52][26] ),
    .B(net526));
 sg13g2_o21ai_1 _18856_ (.B1(_03201_),
    .Y(_02006_),
    .A1(net211),
    .A2(net525));
 sg13g2_mux2_1 _18857_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[52][27] ),
    .S(net529),
    .X(_02007_));
 sg13g2_nand2_1 _18858_ (.Y(_03202_),
    .A(\top_ihp.oisc.regs[52][28] ),
    .B(net526));
 sg13g2_o21ai_1 _18859_ (.B1(_03202_),
    .Y(_02008_),
    .A1(net27),
    .A2(net525));
 sg13g2_nand2_1 _18860_ (.Y(_03203_),
    .A(\top_ihp.oisc.regs[52][29] ),
    .B(net526));
 sg13g2_o21ai_1 _18861_ (.B1(_03203_),
    .Y(_02009_),
    .A1(net89),
    .A2(net525));
 sg13g2_nand2_1 _18862_ (.Y(_03204_),
    .A(\top_ihp.oisc.regs[52][2] ),
    .B(net526));
 sg13g2_o21ai_1 _18863_ (.B1(_03204_),
    .Y(_02010_),
    .A1(net38),
    .A2(net525));
 sg13g2_nand2_1 _18864_ (.Y(_03205_),
    .A(\top_ihp.oisc.regs[52][30] ),
    .B(net649));
 sg13g2_o21ai_1 _18865_ (.B1(_03205_),
    .Y(_02011_),
    .A1(net26),
    .A2(net525));
 sg13g2_nand2_1 _18866_ (.Y(_03206_),
    .A(\top_ihp.oisc.regs[52][31] ),
    .B(net649));
 sg13g2_o21ai_1 _18867_ (.B1(_03206_),
    .Y(_02012_),
    .A1(net87),
    .A2(_03196_));
 sg13g2_mux2_1 _18868_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[52][3] ),
    .S(net529),
    .X(_02013_));
 sg13g2_mux2_1 _18869_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[52][4] ),
    .S(net529),
    .X(_02014_));
 sg13g2_mux2_1 _18870_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[52][5] ),
    .S(net529),
    .X(_02015_));
 sg13g2_mux2_1 _18871_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[52][6] ),
    .S(net527),
    .X(_02016_));
 sg13g2_nand2_1 _18872_ (.Y(_03207_),
    .A(\top_ihp.oisc.regs[52][7] ),
    .B(net649));
 sg13g2_o21ai_1 _18873_ (.B1(_03207_),
    .Y(_02017_),
    .A1(net210),
    .A2(net529));
 sg13g2_nand2_1 _18874_ (.Y(_03208_),
    .A(\top_ihp.oisc.regs[52][8] ),
    .B(_03181_));
 sg13g2_o21ai_1 _18875_ (.B1(_03208_),
    .Y(_02018_),
    .A1(net88),
    .A2(net529));
 sg13g2_mux2_1 _18876_ (.A0(_11225_),
    .A1(\top_ihp.oisc.regs[52][9] ),
    .S(_03184_),
    .X(_02019_));
 sg13g2_nor2_1 _18877_ (.A(_11080_),
    .B(_03047_),
    .Y(_03209_));
 sg13g2_buf_1 _18878_ (.A(_03209_),
    .X(_03210_));
 sg13g2_buf_2 _18879_ (.A(_03210_),
    .X(_03211_));
 sg13g2_mux2_1 _18880_ (.A0(\top_ihp.oisc.regs[53][0] ),
    .A1(net103),
    .S(_03211_),
    .X(_02020_));
 sg13g2_mux2_1 _18881_ (.A0(\top_ihp.oisc.regs[53][10] ),
    .A1(_11262_),
    .S(net524),
    .X(_02021_));
 sg13g2_nor2_1 _18882_ (.A(\top_ihp.oisc.regs[53][11] ),
    .B(net648),
    .Y(_03212_));
 sg13g2_a21oi_1 _18883_ (.A1(net50),
    .A2(net524),
    .Y(_02022_),
    .B1(_03212_));
 sg13g2_nor2_1 _18884_ (.A(\top_ihp.oisc.regs[53][12] ),
    .B(net648),
    .Y(_03213_));
 sg13g2_a21oi_1 _18885_ (.A1(net52),
    .A2(net524),
    .Y(_02023_),
    .B1(_03213_));
 sg13g2_or2_1 _18886_ (.X(_03214_),
    .B(_03047_),
    .A(_11080_));
 sg13g2_buf_1 _18887_ (.A(_03214_),
    .X(_03215_));
 sg13g2_buf_1 _18888_ (.A(net647),
    .X(_03216_));
 sg13g2_buf_1 _18889_ (.A(net647),
    .X(_03217_));
 sg13g2_nand2_1 _18890_ (.Y(_03218_),
    .A(\top_ihp.oisc.regs[53][13] ),
    .B(_03217_));
 sg13g2_o21ai_1 _18891_ (.B1(_03218_),
    .Y(_02024_),
    .A1(net96),
    .A2(net523));
 sg13g2_nand2_1 _18892_ (.Y(_03219_),
    .A(\top_ihp.oisc.regs[53][14] ),
    .B(_03217_));
 sg13g2_o21ai_1 _18893_ (.B1(_03219_),
    .Y(_02025_),
    .A1(net95),
    .A2(net523));
 sg13g2_buf_1 _18894_ (.A(_03215_),
    .X(_03220_));
 sg13g2_nand2_1 _18895_ (.Y(_03221_),
    .A(\top_ihp.oisc.regs[53][15] ),
    .B(net521));
 sg13g2_o21ai_1 _18896_ (.B1(_03221_),
    .Y(_02026_),
    .A1(net209),
    .A2(net523));
 sg13g2_nand2_1 _18897_ (.Y(_03222_),
    .A(\top_ihp.oisc.regs[53][16] ),
    .B(net521));
 sg13g2_o21ai_1 _18898_ (.B1(_03222_),
    .Y(_02027_),
    .A1(net94),
    .A2(net523));
 sg13g2_nand2_1 _18899_ (.Y(_03223_),
    .A(\top_ihp.oisc.regs[53][17] ),
    .B(_03220_));
 sg13g2_o21ai_1 _18900_ (.B1(_03223_),
    .Y(_02028_),
    .A1(net212),
    .A2(_03216_));
 sg13g2_nand2_1 _18901_ (.Y(_03224_),
    .A(\top_ihp.oisc.regs[53][18] ),
    .B(_03220_));
 sg13g2_o21ai_1 _18902_ (.B1(_03224_),
    .Y(_02029_),
    .A1(net93),
    .A2(_03216_));
 sg13g2_mux2_1 _18903_ (.A0(\top_ihp.oisc.regs[53][19] ),
    .A1(net227),
    .S(net524),
    .X(_02030_));
 sg13g2_nor2_1 _18904_ (.A(\top_ihp.oisc.regs[53][1] ),
    .B(net648),
    .Y(_03225_));
 sg13g2_a21oi_1 _18905_ (.A1(_10932_),
    .A2(net524),
    .Y(_02031_),
    .B1(_03225_));
 sg13g2_nand2_1 _18906_ (.Y(_03226_),
    .A(\top_ihp.oisc.regs[53][20] ),
    .B(net521));
 sg13g2_o21ai_1 _18907_ (.B1(_03226_),
    .Y(_02032_),
    .A1(net39),
    .A2(net523));
 sg13g2_nand2_1 _18908_ (.Y(_03227_),
    .A(\top_ihp.oisc.regs[53][21] ),
    .B(net521));
 sg13g2_o21ai_1 _18909_ (.B1(_03227_),
    .Y(_02033_),
    .A1(net92),
    .A2(net523));
 sg13g2_nand2_1 _18910_ (.Y(_03228_),
    .A(\top_ihp.oisc.regs[53][22] ),
    .B(net521));
 sg13g2_o21ai_1 _18911_ (.B1(_03228_),
    .Y(_02034_),
    .A1(net91),
    .A2(net523));
 sg13g2_nand2_1 _18912_ (.Y(_03229_),
    .A(\top_ihp.oisc.regs[53][23] ),
    .B(net521));
 sg13g2_o21ai_1 _18913_ (.B1(_03229_),
    .Y(_02035_),
    .A1(net90),
    .A2(net523));
 sg13g2_mux2_1 _18914_ (.A0(\top_ihp.oisc.regs[53][24] ),
    .A1(_11281_),
    .S(net524),
    .X(_02036_));
 sg13g2_nand2_1 _18915_ (.Y(_03230_),
    .A(\top_ihp.oisc.regs[53][25] ),
    .B(net521));
 sg13g2_o21ai_1 _18916_ (.B1(_03230_),
    .Y(_02037_),
    .A1(net213),
    .A2(net522));
 sg13g2_nand2_1 _18917_ (.Y(_03231_),
    .A(\top_ihp.oisc.regs[53][26] ),
    .B(net521));
 sg13g2_o21ai_1 _18918_ (.B1(_03231_),
    .Y(_02038_),
    .A1(_02935_),
    .A2(net522));
 sg13g2_mux2_1 _18919_ (.A0(\top_ihp.oisc.regs[53][27] ),
    .A1(net101),
    .S(net524),
    .X(_02039_));
 sg13g2_nor2_1 _18920_ (.A(\top_ihp.oisc.regs[53][28] ),
    .B(net648),
    .Y(_03232_));
 sg13g2_a21oi_1 _18921_ (.A1(net116),
    .A2(net524),
    .Y(_02040_),
    .B1(_03232_));
 sg13g2_nand2_1 _18922_ (.Y(_03233_),
    .A(\top_ihp.oisc.regs[53][29] ),
    .B(net647));
 sg13g2_o21ai_1 _18923_ (.B1(_03233_),
    .Y(_02041_),
    .A1(net89),
    .A2(net522));
 sg13g2_nand2_1 _18924_ (.Y(_03234_),
    .A(\top_ihp.oisc.regs[53][2] ),
    .B(net647));
 sg13g2_o21ai_1 _18925_ (.B1(_03234_),
    .Y(_02042_),
    .A1(net38),
    .A2(net522));
 sg13g2_nand2_1 _18926_ (.Y(_03235_),
    .A(\top_ihp.oisc.regs[53][30] ),
    .B(net647));
 sg13g2_o21ai_1 _18927_ (.B1(_03235_),
    .Y(_02043_),
    .A1(net26),
    .A2(net522));
 sg13g2_nand2_1 _18928_ (.Y(_03236_),
    .A(\top_ihp.oisc.regs[53][31] ),
    .B(net647));
 sg13g2_o21ai_1 _18929_ (.B1(_03236_),
    .Y(_02044_),
    .A1(net87),
    .A2(net522));
 sg13g2_mux2_1 _18930_ (.A0(\top_ihp.oisc.regs[53][3] ),
    .A1(_11290_),
    .S(_03211_),
    .X(_02045_));
 sg13g2_mux2_1 _18931_ (.A0(\top_ihp.oisc.regs[53][4] ),
    .A1(_11291_),
    .S(net648),
    .X(_02046_));
 sg13g2_mux2_1 _18932_ (.A0(\top_ihp.oisc.regs[53][5] ),
    .A1(net226),
    .S(net648),
    .X(_02047_));
 sg13g2_mux2_1 _18933_ (.A0(\top_ihp.oisc.regs[53][6] ),
    .A1(net98),
    .S(net648),
    .X(_02048_));
 sg13g2_nand2_1 _18934_ (.Y(_03237_),
    .A(\top_ihp.oisc.regs[53][7] ),
    .B(net647));
 sg13g2_o21ai_1 _18935_ (.B1(_03237_),
    .Y(_02049_),
    .A1(net210),
    .A2(net522));
 sg13g2_nand2_1 _18936_ (.Y(_03238_),
    .A(\top_ihp.oisc.regs[53][8] ),
    .B(net647));
 sg13g2_o21ai_1 _18937_ (.B1(_03238_),
    .Y(_02050_),
    .A1(net88),
    .A2(net522));
 sg13g2_mux2_1 _18938_ (.A0(\top_ihp.oisc.regs[53][9] ),
    .A1(net97),
    .S(net648),
    .X(_02051_));
 sg13g2_nor2_1 _18939_ (.A(_11080_),
    .B(_03112_),
    .Y(_03239_));
 sg13g2_buf_1 _18940_ (.A(_03239_),
    .X(_03240_));
 sg13g2_buf_2 _18941_ (.A(net690),
    .X(_03241_));
 sg13g2_mux2_1 _18942_ (.A0(\top_ihp.oisc.regs[54][0] ),
    .A1(_11256_),
    .S(net646),
    .X(_02052_));
 sg13g2_mux2_1 _18943_ (.A0(\top_ihp.oisc.regs[54][10] ),
    .A1(net102),
    .S(net646),
    .X(_02053_));
 sg13g2_nor2_1 _18944_ (.A(\top_ihp.oisc.regs[54][11] ),
    .B(net690),
    .Y(_03242_));
 sg13g2_a21oi_1 _18945_ (.A1(net50),
    .A2(_03241_),
    .Y(_02054_),
    .B1(_03242_));
 sg13g2_nor2_1 _18946_ (.A(\top_ihp.oisc.regs[54][12] ),
    .B(_03240_),
    .Y(_03243_));
 sg13g2_a21oi_1 _18947_ (.A1(net61),
    .A2(net646),
    .Y(_02055_),
    .B1(_03243_));
 sg13g2_buf_1 _18948_ (.A(net261),
    .X(_03244_));
 sg13g2_nand2_1 _18949_ (.Y(_03245_),
    .A(net729),
    .B(_03119_));
 sg13g2_buf_1 _18950_ (.A(_03245_),
    .X(_03246_));
 sg13g2_buf_2 _18951_ (.A(net645),
    .X(_03247_));
 sg13g2_buf_1 _18952_ (.A(_03245_),
    .X(_03248_));
 sg13g2_nand2_1 _18953_ (.Y(_03249_),
    .A(\top_ihp.oisc.regs[54][13] ),
    .B(_03248_));
 sg13g2_o21ai_1 _18954_ (.B1(_03249_),
    .Y(_02056_),
    .A1(net86),
    .A2(net520));
 sg13g2_buf_1 _18955_ (.A(net260),
    .X(_03250_));
 sg13g2_buf_2 _18956_ (.A(net645),
    .X(_03251_));
 sg13g2_nand2_1 _18957_ (.Y(_03252_),
    .A(\top_ihp.oisc.regs[54][14] ),
    .B(net519));
 sg13g2_o21ai_1 _18958_ (.B1(_03252_),
    .Y(_02057_),
    .A1(net85),
    .A2(net520));
 sg13g2_nand2_1 _18959_ (.Y(_03253_),
    .A(\top_ihp.oisc.regs[54][15] ),
    .B(net519));
 sg13g2_o21ai_1 _18960_ (.B1(_03253_),
    .Y(_02058_),
    .A1(net209),
    .A2(net520));
 sg13g2_buf_1 _18961_ (.A(net276),
    .X(_03254_));
 sg13g2_nand2_1 _18962_ (.Y(_03255_),
    .A(\top_ihp.oisc.regs[54][16] ),
    .B(_03251_));
 sg13g2_o21ai_1 _18963_ (.B1(_03255_),
    .Y(_02059_),
    .A1(net84),
    .A2(net520));
 sg13g2_buf_1 _18964_ (.A(net398),
    .X(_03256_));
 sg13g2_nand2_1 _18965_ (.Y(_03257_),
    .A(\top_ihp.oisc.regs[54][17] ),
    .B(net519));
 sg13g2_o21ai_1 _18966_ (.B1(_03257_),
    .Y(_02060_),
    .A1(_03256_),
    .A2(net520));
 sg13g2_buf_1 _18967_ (.A(net259),
    .X(_03258_));
 sg13g2_nand2_1 _18968_ (.Y(_03259_),
    .A(\top_ihp.oisc.regs[54][18] ),
    .B(net519));
 sg13g2_o21ai_1 _18969_ (.B1(_03259_),
    .Y(_02061_),
    .A1(net83),
    .A2(net520));
 sg13g2_nand2_1 _18970_ (.Y(_03260_),
    .A(\top_ihp.oisc.regs[54][19] ),
    .B(_03251_));
 sg13g2_o21ai_1 _18971_ (.B1(_03260_),
    .Y(_02062_),
    .A1(_10273_),
    .A2(_03247_));
 sg13g2_nor2_1 _18972_ (.A(\top_ihp.oisc.regs[54][1] ),
    .B(net690),
    .Y(_03261_));
 sg13g2_a21oi_1 _18973_ (.A1(net139),
    .A2(net646),
    .Y(_02063_),
    .B1(_03261_));
 sg13g2_buf_1 _18974_ (.A(net121),
    .X(_03262_));
 sg13g2_nand2_1 _18975_ (.Y(_03263_),
    .A(\top_ihp.oisc.regs[54][20] ),
    .B(net519));
 sg13g2_o21ai_1 _18976_ (.B1(_03263_),
    .Y(_02064_),
    .A1(net36),
    .A2(net520));
 sg13g2_buf_1 _18977_ (.A(_10361_),
    .X(_03264_));
 sg13g2_nand2_1 _18978_ (.Y(_03265_),
    .A(\top_ihp.oisc.regs[54][21] ),
    .B(net519));
 sg13g2_o21ai_1 _18979_ (.B1(_03265_),
    .Y(_02065_),
    .A1(_03264_),
    .A2(_03247_));
 sg13g2_buf_2 _18980_ (.A(net258),
    .X(_03266_));
 sg13g2_nand2_1 _18981_ (.Y(_03267_),
    .A(\top_ihp.oisc.regs[54][22] ),
    .B(net519));
 sg13g2_o21ai_1 _18982_ (.B1(_03267_),
    .Y(_02066_),
    .A1(net81),
    .A2(net644));
 sg13g2_buf_2 _18983_ (.A(_10392_),
    .X(_03268_));
 sg13g2_nand2_1 _18984_ (.Y(_03269_),
    .A(\top_ihp.oisc.regs[54][23] ),
    .B(net519));
 sg13g2_o21ai_1 _18985_ (.B1(_03269_),
    .Y(_02067_),
    .A1(net207),
    .A2(net644));
 sg13g2_mux2_1 _18986_ (.A0(\top_ihp.oisc.regs[54][24] ),
    .A1(net382),
    .S(net646),
    .X(_02068_));
 sg13g2_nor2_1 _18987_ (.A(\top_ihp.oisc.regs[54][25] ),
    .B(net690),
    .Y(_03270_));
 sg13g2_a21oi_1 _18988_ (.A1(net59),
    .A2(net646),
    .Y(_02069_),
    .B1(_03270_));
 sg13g2_buf_1 _18989_ (.A(net397),
    .X(_03271_));
 sg13g2_nand2_1 _18990_ (.Y(_03272_),
    .A(\top_ihp.oisc.regs[54][26] ),
    .B(net645));
 sg13g2_o21ai_1 _18991_ (.B1(_03272_),
    .Y(_02070_),
    .A1(net206),
    .A2(net644));
 sg13g2_nand2_1 _18992_ (.Y(_03273_),
    .A(\top_ihp.oisc.regs[54][27] ),
    .B(net645));
 sg13g2_o21ai_1 _18993_ (.B1(_03273_),
    .Y(_02071_),
    .A1(net31),
    .A2(net644));
 sg13g2_nor2_1 _18994_ (.A(\top_ihp.oisc.regs[54][28] ),
    .B(net690),
    .Y(_03274_));
 sg13g2_a21oi_1 _18995_ (.A1(net30),
    .A2(net646),
    .Y(_02072_),
    .B1(_03274_));
 sg13g2_buf_1 _18996_ (.A(net256),
    .X(_03275_));
 sg13g2_nand2_1 _18997_ (.Y(_03276_),
    .A(\top_ihp.oisc.regs[54][29] ),
    .B(net645));
 sg13g2_o21ai_1 _18998_ (.B1(_03276_),
    .Y(_02073_),
    .A1(_03275_),
    .A2(net644));
 sg13g2_nand2_1 _18999_ (.Y(_03277_),
    .A(\top_ihp.oisc.regs[54][2] ),
    .B(net645));
 sg13g2_o21ai_1 _19000_ (.B1(_03277_),
    .Y(_02074_),
    .A1(net38),
    .A2(net644));
 sg13g2_nand2_1 _19001_ (.Y(_03278_),
    .A(\top_ihp.oisc.regs[54][30] ),
    .B(_03246_));
 sg13g2_o21ai_1 _19002_ (.B1(_03278_),
    .Y(_02075_),
    .A1(net26),
    .A2(net644));
 sg13g2_inv_1 _19003_ (.Y(_03279_),
    .A(\top_ihp.oisc.regs[54][31] ));
 sg13g2_nor2_1 _19004_ (.A(_10535_),
    .B(net645),
    .Y(_03280_));
 sg13g2_a22oi_1 _19005_ (.Y(_02076_),
    .B1(_03280_),
    .B2(net129),
    .A2(net520),
    .A1(_03279_));
 sg13g2_mux2_1 _19006_ (.A0(\top_ihp.oisc.regs[54][3] ),
    .A1(net100),
    .S(_03241_),
    .X(_02077_));
 sg13g2_mux2_1 _19007_ (.A0(\top_ihp.oisc.regs[54][4] ),
    .A1(net99),
    .S(net646),
    .X(_02078_));
 sg13g2_mux2_1 _19008_ (.A0(\top_ihp.oisc.regs[54][5] ),
    .A1(net226),
    .S(net690),
    .X(_02079_));
 sg13g2_mux2_1 _19009_ (.A0(\top_ihp.oisc.regs[54][6] ),
    .A1(net98),
    .S(net690),
    .X(_02080_));
 sg13g2_buf_1 _19010_ (.A(_10661_),
    .X(_03281_));
 sg13g2_nand2_1 _19011_ (.Y(_03282_),
    .A(\top_ihp.oisc.regs[54][7] ),
    .B(net645));
 sg13g2_o21ai_1 _19012_ (.B1(_03282_),
    .Y(_02081_),
    .A1(net343),
    .A2(net644));
 sg13g2_buf_2 _19013_ (.A(_10673_),
    .X(_03283_));
 sg13g2_nand2_1 _19014_ (.Y(_03284_),
    .A(\top_ihp.oisc.regs[54][8] ),
    .B(_03246_));
 sg13g2_o21ai_1 _19015_ (.B1(_03284_),
    .Y(_02082_),
    .A1(net205),
    .A2(_03248_));
 sg13g2_mux2_1 _19016_ (.A0(\top_ihp.oisc.regs[54][9] ),
    .A1(net97),
    .S(net690),
    .X(_02083_));
 sg13g2_and2_1 _19017_ (.A(net729),
    .B(_03150_),
    .X(_03285_));
 sg13g2_buf_1 _19018_ (.A(_03285_),
    .X(_03286_));
 sg13g2_buf_2 _19019_ (.A(_03286_),
    .X(_03287_));
 sg13g2_mux2_1 _19020_ (.A0(\top_ihp.oisc.regs[55][0] ),
    .A1(_11256_),
    .S(_03287_),
    .X(_02084_));
 sg13g2_mux2_1 _19021_ (.A0(\top_ihp.oisc.regs[55][10] ),
    .A1(_11262_),
    .S(net518),
    .X(_02085_));
 sg13g2_nand2_1 _19022_ (.Y(_03288_),
    .A(net729),
    .B(_03150_));
 sg13g2_buf_1 _19023_ (.A(_03288_),
    .X(_03289_));
 sg13g2_buf_1 _19024_ (.A(_03289_),
    .X(_03290_));
 sg13g2_buf_1 _19025_ (.A(_03289_),
    .X(_03291_));
 sg13g2_nand2_1 _19026_ (.Y(_03292_),
    .A(\top_ihp.oisc.regs[55][11] ),
    .B(_03291_));
 sg13g2_o21ai_1 _19027_ (.B1(_03292_),
    .Y(_02086_),
    .A1(net37),
    .A2(_03290_));
 sg13g2_nand2_1 _19028_ (.Y(_03293_),
    .A(\top_ihp.oisc.regs[55][12] ),
    .B(_03291_));
 sg13g2_o21ai_1 _19029_ (.B1(_03293_),
    .Y(_02087_),
    .A1(_11303_),
    .A2(_03290_));
 sg13g2_nand2_1 _19030_ (.Y(_03294_),
    .A(\top_ihp.oisc.regs[55][13] ),
    .B(net516));
 sg13g2_o21ai_1 _19031_ (.B1(_03294_),
    .Y(_02088_),
    .A1(net86),
    .A2(net517));
 sg13g2_nand2_1 _19032_ (.Y(_03295_),
    .A(\top_ihp.oisc.regs[55][14] ),
    .B(net516));
 sg13g2_o21ai_1 _19033_ (.B1(_03295_),
    .Y(_02089_),
    .A1(net85),
    .A2(net517));
 sg13g2_mux2_1 _19034_ (.A0(\top_ihp.oisc.regs[55][15] ),
    .A1(net663),
    .S(net518),
    .X(_02090_));
 sg13g2_nand2_1 _19035_ (.Y(_03296_),
    .A(\top_ihp.oisc.regs[55][16] ),
    .B(net516));
 sg13g2_o21ai_1 _19036_ (.B1(_03296_),
    .Y(_02091_),
    .A1(net84),
    .A2(net517));
 sg13g2_nand2_1 _19037_ (.Y(_03297_),
    .A(\top_ihp.oisc.regs[55][17] ),
    .B(net516));
 sg13g2_o21ai_1 _19038_ (.B1(_03297_),
    .Y(_02092_),
    .A1(net208),
    .A2(net517));
 sg13g2_nand2_1 _19039_ (.Y(_03298_),
    .A(\top_ihp.oisc.regs[55][18] ),
    .B(net516));
 sg13g2_o21ai_1 _19040_ (.B1(_03298_),
    .Y(_02093_),
    .A1(net83),
    .A2(net517));
 sg13g2_mux2_1 _19041_ (.A0(\top_ihp.oisc.regs[55][19] ),
    .A1(net227),
    .S(net518),
    .X(_02094_));
 sg13g2_nand2_1 _19042_ (.Y(_03299_),
    .A(\top_ihp.oisc.regs[55][1] ),
    .B(net516));
 sg13g2_o21ai_1 _19043_ (.B1(_03299_),
    .Y(_02095_),
    .A1(net105),
    .A2(net517));
 sg13g2_nand2_1 _19044_ (.Y(_03300_),
    .A(\top_ihp.oisc.regs[55][20] ),
    .B(net516));
 sg13g2_o21ai_1 _19045_ (.B1(_03300_),
    .Y(_02096_),
    .A1(net36),
    .A2(net517));
 sg13g2_nand2_1 _19046_ (.Y(_03301_),
    .A(\top_ihp.oisc.regs[55][21] ),
    .B(net516));
 sg13g2_o21ai_1 _19047_ (.B1(_03301_),
    .Y(_02097_),
    .A1(net82),
    .A2(net517));
 sg13g2_buf_1 _19048_ (.A(_03289_),
    .X(_03302_));
 sg13g2_buf_1 _19049_ (.A(_03289_),
    .X(_03303_));
 sg13g2_nand2_1 _19050_ (.Y(_03304_),
    .A(\top_ihp.oisc.regs[55][22] ),
    .B(net514));
 sg13g2_o21ai_1 _19051_ (.B1(_03304_),
    .Y(_02098_),
    .A1(net81),
    .A2(net515));
 sg13g2_nand2_1 _19052_ (.Y(_03305_),
    .A(\top_ihp.oisc.regs[55][23] ),
    .B(net514));
 sg13g2_o21ai_1 _19053_ (.B1(_03305_),
    .Y(_02099_),
    .A1(net207),
    .A2(net515));
 sg13g2_mux2_1 _19054_ (.A0(\top_ihp.oisc.regs[55][24] ),
    .A1(net382),
    .S(net518),
    .X(_02100_));
 sg13g2_nand2_1 _19055_ (.Y(_03306_),
    .A(\top_ihp.oisc.regs[55][25] ),
    .B(net514));
 sg13g2_o21ai_1 _19056_ (.B1(_03306_),
    .Y(_02101_),
    .A1(net213),
    .A2(net515));
 sg13g2_nand2_1 _19057_ (.Y(_03307_),
    .A(\top_ihp.oisc.regs[55][26] ),
    .B(net514));
 sg13g2_o21ai_1 _19058_ (.B1(_03307_),
    .Y(_02102_),
    .A1(net206),
    .A2(net515));
 sg13g2_mux2_1 _19059_ (.A0(\top_ihp.oisc.regs[55][27] ),
    .A1(net101),
    .S(net518),
    .X(_02103_));
 sg13g2_nor2_1 _19060_ (.A(\top_ihp.oisc.regs[55][28] ),
    .B(_03286_),
    .Y(_03308_));
 sg13g2_a21oi_1 _19061_ (.A1(net116),
    .A2(net518),
    .Y(_02104_),
    .B1(_03308_));
 sg13g2_nand2_1 _19062_ (.Y(_03309_),
    .A(\top_ihp.oisc.regs[55][29] ),
    .B(net514));
 sg13g2_o21ai_1 _19063_ (.B1(_03309_),
    .Y(_02105_),
    .A1(net80),
    .A2(net515));
 sg13g2_buf_2 _19064_ (.A(_10499_),
    .X(_03310_));
 sg13g2_nand2_1 _19065_ (.Y(_03311_),
    .A(\top_ihp.oisc.regs[55][2] ),
    .B(net514));
 sg13g2_o21ai_1 _19066_ (.B1(_03311_),
    .Y(_02106_),
    .A1(net79),
    .A2(net515));
 sg13g2_buf_1 _19067_ (.A(_10508_),
    .X(_03312_));
 sg13g2_nand2_1 _19068_ (.Y(_03313_),
    .A(\top_ihp.oisc.regs[55][30] ),
    .B(net514));
 sg13g2_o21ai_1 _19069_ (.B1(_03313_),
    .Y(_02107_),
    .A1(net35),
    .A2(net515));
 sg13g2_nand2_1 _19070_ (.Y(_03314_),
    .A(\top_ihp.oisc.regs[55][31] ),
    .B(net514));
 sg13g2_o21ai_1 _19071_ (.B1(_03314_),
    .Y(_02108_),
    .A1(_03074_),
    .A2(net515));
 sg13g2_mux2_1 _19072_ (.A0(\top_ihp.oisc.regs[55][3] ),
    .A1(net100),
    .S(net518),
    .X(_02109_));
 sg13g2_mux2_1 _19073_ (.A0(\top_ihp.oisc.regs[55][4] ),
    .A1(net99),
    .S(net518),
    .X(_02110_));
 sg13g2_mux2_1 _19074_ (.A0(\top_ihp.oisc.regs[55][5] ),
    .A1(_11292_),
    .S(_03287_),
    .X(_02111_));
 sg13g2_mux2_1 _19075_ (.A0(\top_ihp.oisc.regs[55][6] ),
    .A1(net98),
    .S(_03286_),
    .X(_02112_));
 sg13g2_nand2_1 _19076_ (.Y(_03315_),
    .A(\top_ihp.oisc.regs[55][7] ),
    .B(_03303_));
 sg13g2_o21ai_1 _19077_ (.B1(_03315_),
    .Y(_02113_),
    .A1(net343),
    .A2(_03302_));
 sg13g2_nand2_1 _19078_ (.Y(_03316_),
    .A(\top_ihp.oisc.regs[55][8] ),
    .B(_03303_));
 sg13g2_o21ai_1 _19079_ (.B1(_03316_),
    .Y(_02114_),
    .A1(net205),
    .A2(_03302_));
 sg13g2_mux2_1 _19080_ (.A0(\top_ihp.oisc.regs[55][9] ),
    .A1(net97),
    .S(_03286_),
    .X(_02115_));
 sg13g2_nand2_1 _19081_ (.Y(_03317_),
    .A(_10694_),
    .B(_03015_));
 sg13g2_buf_1 _19082_ (.A(_03317_),
    .X(_03318_));
 sg13g2_buf_2 _19083_ (.A(net643),
    .X(_03319_));
 sg13g2_mux2_1 _19084_ (.A0(net46),
    .A1(\top_ihp.oisc.regs[56][0] ),
    .S(net513),
    .X(_02116_));
 sg13g2_mux2_1 _19085_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[56][10] ),
    .S(net513),
    .X(_02117_));
 sg13g2_buf_1 _19086_ (.A(net643),
    .X(_03320_));
 sg13g2_buf_2 _19087_ (.A(net643),
    .X(_03321_));
 sg13g2_nand2_1 _19088_ (.Y(_03322_),
    .A(\top_ihp.oisc.regs[56][11] ),
    .B(net511));
 sg13g2_o21ai_1 _19089_ (.B1(_03322_),
    .Y(_02118_),
    .A1(net37),
    .A2(net512));
 sg13g2_nand2_1 _19090_ (.Y(_03323_),
    .A(\top_ihp.oisc.regs[56][12] ),
    .B(net511));
 sg13g2_o21ai_1 _19091_ (.B1(_03323_),
    .Y(_02119_),
    .A1(net40),
    .A2(net512));
 sg13g2_nand2_1 _19092_ (.Y(_03324_),
    .A(\top_ihp.oisc.regs[56][13] ),
    .B(net511));
 sg13g2_o21ai_1 _19093_ (.B1(_03324_),
    .Y(_02120_),
    .A1(net86),
    .A2(net512));
 sg13g2_nand2_1 _19094_ (.Y(_03325_),
    .A(\top_ihp.oisc.regs[56][14] ),
    .B(_03321_));
 sg13g2_o21ai_1 _19095_ (.B1(_03325_),
    .Y(_02121_),
    .A1(_03250_),
    .A2(net512));
 sg13g2_nand2_1 _19096_ (.Y(_03326_),
    .A(\top_ihp.oisc.regs[56][15] ),
    .B(net511));
 sg13g2_o21ai_1 _19097_ (.B1(_03326_),
    .Y(_02122_),
    .A1(_03127_),
    .A2(net512));
 sg13g2_nand2_1 _19098_ (.Y(_03327_),
    .A(\top_ihp.oisc.regs[56][16] ),
    .B(_03321_));
 sg13g2_o21ai_1 _19099_ (.B1(_03327_),
    .Y(_02123_),
    .A1(_03254_),
    .A2(net512));
 sg13g2_nand2_1 _19100_ (.Y(_03328_),
    .A(\top_ihp.oisc.regs[56][17] ),
    .B(net511));
 sg13g2_o21ai_1 _19101_ (.B1(_03328_),
    .Y(_02124_),
    .A1(net208),
    .A2(_03320_));
 sg13g2_nand2_1 _19102_ (.Y(_03329_),
    .A(\top_ihp.oisc.regs[56][18] ),
    .B(net511));
 sg13g2_o21ai_1 _19103_ (.B1(_03329_),
    .Y(_02125_),
    .A1(_03258_),
    .A2(net512));
 sg13g2_mux2_1 _19104_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[56][19] ),
    .S(net513),
    .X(_02126_));
 sg13g2_buf_1 _19105_ (.A(net643),
    .X(_03330_));
 sg13g2_nand2_1 _19106_ (.Y(_03331_),
    .A(\top_ihp.oisc.regs[56][1] ),
    .B(net510));
 sg13g2_o21ai_1 _19107_ (.B1(_03331_),
    .Y(_02127_),
    .A1(net105),
    .A2(net512));
 sg13g2_nand2_1 _19108_ (.Y(_03332_),
    .A(\top_ihp.oisc.regs[56][20] ),
    .B(_03330_));
 sg13g2_o21ai_1 _19109_ (.B1(_03332_),
    .Y(_02128_),
    .A1(net36),
    .A2(_03320_));
 sg13g2_buf_1 _19110_ (.A(net643),
    .X(_03333_));
 sg13g2_nand2_1 _19111_ (.Y(_03334_),
    .A(\top_ihp.oisc.regs[56][21] ),
    .B(_03330_));
 sg13g2_o21ai_1 _19112_ (.B1(_03334_),
    .Y(_02129_),
    .A1(net82),
    .A2(net509));
 sg13g2_nand2_1 _19113_ (.Y(_03335_),
    .A(\top_ihp.oisc.regs[56][22] ),
    .B(net510));
 sg13g2_o21ai_1 _19114_ (.B1(_03335_),
    .Y(_02130_),
    .A1(net81),
    .A2(net509));
 sg13g2_nand2_1 _19115_ (.Y(_03336_),
    .A(\top_ihp.oisc.regs[56][23] ),
    .B(net510));
 sg13g2_o21ai_1 _19116_ (.B1(_03336_),
    .Y(_02131_),
    .A1(net207),
    .A2(net509));
 sg13g2_mux2_1 _19117_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[56][24] ),
    .S(net513),
    .X(_02132_));
 sg13g2_nand2_1 _19118_ (.Y(_03337_),
    .A(\top_ihp.oisc.regs[56][25] ),
    .B(net510));
 sg13g2_o21ai_1 _19119_ (.B1(_03337_),
    .Y(_02133_),
    .A1(net262),
    .A2(_03333_));
 sg13g2_nand2_1 _19120_ (.Y(_03338_),
    .A(\top_ihp.oisc.regs[56][26] ),
    .B(net510));
 sg13g2_o21ai_1 _19121_ (.B1(_03338_),
    .Y(_02134_),
    .A1(net206),
    .A2(net509));
 sg13g2_mux2_1 _19122_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[56][27] ),
    .S(net513),
    .X(_02135_));
 sg13g2_nand2_1 _19123_ (.Y(_03339_),
    .A(\top_ihp.oisc.regs[56][28] ),
    .B(net510));
 sg13g2_o21ai_1 _19124_ (.B1(_03339_),
    .Y(_02136_),
    .A1(net27),
    .A2(net509));
 sg13g2_nand2_1 _19125_ (.Y(_03340_),
    .A(\top_ihp.oisc.regs[56][29] ),
    .B(net510));
 sg13g2_o21ai_1 _19126_ (.B1(_03340_),
    .Y(_02137_),
    .A1(net80),
    .A2(net509));
 sg13g2_nand2_1 _19127_ (.Y(_03341_),
    .A(\top_ihp.oisc.regs[56][2] ),
    .B(net510));
 sg13g2_o21ai_1 _19128_ (.B1(_03341_),
    .Y(_02138_),
    .A1(net79),
    .A2(net509));
 sg13g2_nand2_1 _19129_ (.Y(_03342_),
    .A(\top_ihp.oisc.regs[56][30] ),
    .B(net643));
 sg13g2_o21ai_1 _19130_ (.B1(_03342_),
    .Y(_02139_),
    .A1(_03312_),
    .A2(_03333_));
 sg13g2_nand2_1 _19131_ (.Y(_03343_),
    .A(\top_ihp.oisc.regs[56][31] ),
    .B(net643));
 sg13g2_o21ai_1 _19132_ (.B1(_03343_),
    .Y(_02140_),
    .A1(net87),
    .A2(net509));
 sg13g2_mux2_1 _19133_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[56][3] ),
    .S(_03319_),
    .X(_02141_));
 sg13g2_mux2_1 _19134_ (.A0(_11220_),
    .A1(\top_ihp.oisc.regs[56][4] ),
    .S(_03319_),
    .X(_02142_));
 sg13g2_mux2_1 _19135_ (.A0(net104),
    .A1(\top_ihp.oisc.regs[56][5] ),
    .S(net513),
    .X(_02143_));
 sg13g2_mux2_1 _19136_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[56][6] ),
    .S(net511),
    .X(_02144_));
 sg13g2_nand2_1 _19137_ (.Y(_03344_),
    .A(\top_ihp.oisc.regs[56][7] ),
    .B(net643));
 sg13g2_o21ai_1 _19138_ (.B1(_03344_),
    .Y(_02145_),
    .A1(net343),
    .A2(net513));
 sg13g2_nand2_1 _19139_ (.Y(_03345_),
    .A(\top_ihp.oisc.regs[56][8] ),
    .B(_03318_));
 sg13g2_o21ai_1 _19140_ (.B1(_03345_),
    .Y(_02146_),
    .A1(net205),
    .A2(net513));
 sg13g2_mux2_1 _19141_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[56][9] ),
    .S(net511),
    .X(_02147_));
 sg13g2_nor2_1 _19142_ (.A(_10706_),
    .B(_03047_),
    .Y(_03346_));
 sg13g2_buf_1 _19143_ (.A(_03346_),
    .X(_03347_));
 sg13g2_buf_2 _19144_ (.A(net642),
    .X(_03348_));
 sg13g2_mux2_1 _19145_ (.A0(\top_ihp.oisc.regs[57][0] ),
    .A1(net143),
    .S(net508),
    .X(_02148_));
 sg13g2_mux2_1 _19146_ (.A0(\top_ihp.oisc.regs[57][10] ),
    .A1(net142),
    .S(net508),
    .X(_02149_));
 sg13g2_nor2_1 _19147_ (.A(\top_ihp.oisc.regs[57][11] ),
    .B(net642),
    .Y(_03349_));
 sg13g2_a21oi_1 _19148_ (.A1(net50),
    .A2(net508),
    .Y(_02150_),
    .B1(_03349_));
 sg13g2_nor2_1 _19149_ (.A(\top_ihp.oisc.regs[57][12] ),
    .B(_03347_),
    .Y(_03350_));
 sg13g2_a21oi_1 _19150_ (.A1(net61),
    .A2(_03348_),
    .Y(_02151_),
    .B1(_03350_));
 sg13g2_or2_1 _19151_ (.X(_03351_),
    .B(_03047_),
    .A(_10706_));
 sg13g2_buf_1 _19152_ (.A(_03351_),
    .X(_03352_));
 sg13g2_buf_2 _19153_ (.A(net641),
    .X(_03353_));
 sg13g2_buf_2 _19154_ (.A(net641),
    .X(_03354_));
 sg13g2_nand2_1 _19155_ (.Y(_03355_),
    .A(\top_ihp.oisc.regs[57][13] ),
    .B(_03354_));
 sg13g2_o21ai_1 _19156_ (.B1(_03355_),
    .Y(_02152_),
    .A1(_03244_),
    .A2(net507));
 sg13g2_nand2_1 _19157_ (.Y(_03356_),
    .A(\top_ihp.oisc.regs[57][14] ),
    .B(_03354_));
 sg13g2_o21ai_1 _19158_ (.B1(_03356_),
    .Y(_02153_),
    .A1(net85),
    .A2(_03353_));
 sg13g2_buf_2 _19159_ (.A(net641),
    .X(_03357_));
 sg13g2_nand2_1 _19160_ (.Y(_03358_),
    .A(\top_ihp.oisc.regs[57][15] ),
    .B(net505));
 sg13g2_o21ai_1 _19161_ (.B1(_03358_),
    .Y(_02154_),
    .A1(net209),
    .A2(net507));
 sg13g2_nand2_1 _19162_ (.Y(_03359_),
    .A(\top_ihp.oisc.regs[57][16] ),
    .B(_03357_));
 sg13g2_o21ai_1 _19163_ (.B1(_03359_),
    .Y(_02155_),
    .A1(net84),
    .A2(net507));
 sg13g2_nand2_1 _19164_ (.Y(_03360_),
    .A(\top_ihp.oisc.regs[57][17] ),
    .B(net505));
 sg13g2_o21ai_1 _19165_ (.B1(_03360_),
    .Y(_02156_),
    .A1(net208),
    .A2(net507));
 sg13g2_nand2_1 _19166_ (.Y(_03361_),
    .A(\top_ihp.oisc.regs[57][18] ),
    .B(_03357_));
 sg13g2_o21ai_1 _19167_ (.B1(_03361_),
    .Y(_02157_),
    .A1(net83),
    .A2(_03353_));
 sg13g2_mux2_1 _19168_ (.A0(\top_ihp.oisc.regs[57][19] ),
    .A1(net227),
    .S(net508),
    .X(_02158_));
 sg13g2_nor2_1 _19169_ (.A(\top_ihp.oisc.regs[57][1] ),
    .B(net642),
    .Y(_03362_));
 sg13g2_a21oi_1 _19170_ (.A1(net139),
    .A2(net508),
    .Y(_02159_),
    .B1(_03362_));
 sg13g2_nand2_1 _19171_ (.Y(_03363_),
    .A(\top_ihp.oisc.regs[57][20] ),
    .B(net505));
 sg13g2_o21ai_1 _19172_ (.B1(_03363_),
    .Y(_02160_),
    .A1(net36),
    .A2(net507));
 sg13g2_nand2_1 _19173_ (.Y(_03364_),
    .A(\top_ihp.oisc.regs[57][21] ),
    .B(net505));
 sg13g2_o21ai_1 _19174_ (.B1(_03364_),
    .Y(_02161_),
    .A1(net82),
    .A2(net507));
 sg13g2_nand2_1 _19175_ (.Y(_03365_),
    .A(\top_ihp.oisc.regs[57][22] ),
    .B(net505));
 sg13g2_o21ai_1 _19176_ (.B1(_03365_),
    .Y(_02162_),
    .A1(net81),
    .A2(net507));
 sg13g2_nand2_1 _19177_ (.Y(_03366_),
    .A(\top_ihp.oisc.regs[57][23] ),
    .B(net505));
 sg13g2_o21ai_1 _19178_ (.B1(_03366_),
    .Y(_02163_),
    .A1(net207),
    .A2(net507));
 sg13g2_mux2_1 _19179_ (.A0(\top_ihp.oisc.regs[57][24] ),
    .A1(net403),
    .S(net508),
    .X(_02164_));
 sg13g2_nand2_1 _19180_ (.Y(_03367_),
    .A(\top_ihp.oisc.regs[57][25] ),
    .B(net505));
 sg13g2_o21ai_1 _19181_ (.B1(_03367_),
    .Y(_02165_),
    .A1(net262),
    .A2(net506));
 sg13g2_nand2_1 _19182_ (.Y(_03368_),
    .A(\top_ihp.oisc.regs[57][26] ),
    .B(net505));
 sg13g2_o21ai_1 _19183_ (.B1(_03368_),
    .Y(_02166_),
    .A1(net206),
    .A2(net506));
 sg13g2_mux2_1 _19184_ (.A0(\top_ihp.oisc.regs[57][27] ),
    .A1(net101),
    .S(net508),
    .X(_02167_));
 sg13g2_nor2_1 _19185_ (.A(\top_ihp.oisc.regs[57][28] ),
    .B(net642),
    .Y(_03369_));
 sg13g2_a21oi_1 _19186_ (.A1(net116),
    .A2(net508),
    .Y(_02168_),
    .B1(_03369_));
 sg13g2_nand2_1 _19187_ (.Y(_03370_),
    .A(\top_ihp.oisc.regs[57][29] ),
    .B(net641));
 sg13g2_o21ai_1 _19188_ (.B1(_03370_),
    .Y(_02169_),
    .A1(net80),
    .A2(net506));
 sg13g2_nand2_1 _19189_ (.Y(_03371_),
    .A(\top_ihp.oisc.regs[57][2] ),
    .B(_03352_));
 sg13g2_o21ai_1 _19190_ (.B1(_03371_),
    .Y(_02170_),
    .A1(net79),
    .A2(net506));
 sg13g2_nand2_1 _19191_ (.Y(_03372_),
    .A(\top_ihp.oisc.regs[57][30] ),
    .B(net641));
 sg13g2_o21ai_1 _19192_ (.B1(_03372_),
    .Y(_02171_),
    .A1(net35),
    .A2(net506));
 sg13g2_nand2_1 _19193_ (.Y(_03373_),
    .A(\top_ihp.oisc.regs[57][31] ),
    .B(net641));
 sg13g2_o21ai_1 _19194_ (.B1(_03373_),
    .Y(_02172_),
    .A1(net87),
    .A2(net506));
 sg13g2_mux2_1 _19195_ (.A0(\top_ihp.oisc.regs[57][3] ),
    .A1(net135),
    .S(_03348_),
    .X(_02173_));
 sg13g2_mux2_1 _19196_ (.A0(\top_ihp.oisc.regs[57][4] ),
    .A1(net134),
    .S(net642),
    .X(_02174_));
 sg13g2_mux2_1 _19197_ (.A0(\top_ihp.oisc.regs[57][5] ),
    .A1(net267),
    .S(net642),
    .X(_02175_));
 sg13g2_mux2_1 _19198_ (.A0(\top_ihp.oisc.regs[57][6] ),
    .A1(net132),
    .S(net642),
    .X(_02176_));
 sg13g2_nand2_1 _19199_ (.Y(_03374_),
    .A(\top_ihp.oisc.regs[57][7] ),
    .B(net641));
 sg13g2_o21ai_1 _19200_ (.B1(_03374_),
    .Y(_02177_),
    .A1(net343),
    .A2(net506));
 sg13g2_nand2_1 _19201_ (.Y(_03375_),
    .A(\top_ihp.oisc.regs[57][8] ),
    .B(net641));
 sg13g2_o21ai_1 _19202_ (.B1(_03375_),
    .Y(_02178_),
    .A1(net205),
    .A2(net506));
 sg13g2_mux2_1 _19203_ (.A0(\top_ihp.oisc.regs[57][9] ),
    .A1(net131),
    .S(net642),
    .X(_02179_));
 sg13g2_nor2_1 _19204_ (.A(_10706_),
    .B(_03112_),
    .Y(_03376_));
 sg13g2_buf_2 _19205_ (.A(_03376_),
    .X(_03377_));
 sg13g2_mux2_1 _19206_ (.A0(\top_ihp.oisc.regs[58][0] ),
    .A1(net143),
    .S(_03377_),
    .X(_02180_));
 sg13g2_mux2_1 _19207_ (.A0(\top_ihp.oisc.regs[58][10] ),
    .A1(net142),
    .S(net640),
    .X(_02181_));
 sg13g2_nor2_1 _19208_ (.A(\top_ihp.oisc.regs[58][11] ),
    .B(_03376_),
    .Y(_03378_));
 sg13g2_a21oi_1 _19209_ (.A1(net50),
    .A2(net640),
    .Y(_02182_),
    .B1(_03378_));
 sg13g2_nand2_1 _19210_ (.Y(_03379_),
    .A(_10694_),
    .B(_03119_));
 sg13g2_buf_2 _19211_ (.A(_03379_),
    .X(_03380_));
 sg13g2_buf_1 _19212_ (.A(_03380_),
    .X(_03381_));
 sg13g2_buf_2 _19213_ (.A(_03380_),
    .X(_03382_));
 sg13g2_nand2_1 _19214_ (.Y(_03383_),
    .A(\top_ihp.oisc.regs[58][12] ),
    .B(net503));
 sg13g2_o21ai_1 _19215_ (.B1(_03383_),
    .Y(_02183_),
    .A1(net40),
    .A2(net504));
 sg13g2_nand2_1 _19216_ (.Y(_03384_),
    .A(\top_ihp.oisc.regs[58][13] ),
    .B(_03382_));
 sg13g2_o21ai_1 _19217_ (.B1(_03384_),
    .Y(_02184_),
    .A1(net86),
    .A2(_03381_));
 sg13g2_nand2_1 _19218_ (.Y(_03385_),
    .A(\top_ihp.oisc.regs[58][14] ),
    .B(net503));
 sg13g2_o21ai_1 _19219_ (.B1(_03385_),
    .Y(_02185_),
    .A1(net85),
    .A2(net504));
 sg13g2_nand2_1 _19220_ (.Y(_03386_),
    .A(\top_ihp.oisc.regs[58][15] ),
    .B(net503));
 sg13g2_o21ai_1 _19221_ (.B1(_03386_),
    .Y(_02186_),
    .A1(net209),
    .A2(net504));
 sg13g2_nand2_1 _19222_ (.Y(_03387_),
    .A(\top_ihp.oisc.regs[58][16] ),
    .B(net503));
 sg13g2_o21ai_1 _19223_ (.B1(_03387_),
    .Y(_02187_),
    .A1(net84),
    .A2(net504));
 sg13g2_nand2_1 _19224_ (.Y(_03388_),
    .A(\top_ihp.oisc.regs[58][17] ),
    .B(_03382_));
 sg13g2_o21ai_1 _19225_ (.B1(_03388_),
    .Y(_02188_),
    .A1(net208),
    .A2(_03381_));
 sg13g2_nand2_1 _19226_ (.Y(_03389_),
    .A(\top_ihp.oisc.regs[58][18] ),
    .B(net503));
 sg13g2_o21ai_1 _19227_ (.B1(_03389_),
    .Y(_02189_),
    .A1(net83),
    .A2(net504));
 sg13g2_nand2_1 _19228_ (.Y(_03390_),
    .A(\top_ihp.oisc.regs[58][19] ),
    .B(net503));
 sg13g2_o21ai_1 _19229_ (.B1(_03390_),
    .Y(_02190_),
    .A1(_10273_),
    .A2(net504));
 sg13g2_nor2_1 _19230_ (.A(\top_ihp.oisc.regs[58][1] ),
    .B(_03376_),
    .Y(_03391_));
 sg13g2_a21oi_1 _19231_ (.A1(net139),
    .A2(net640),
    .Y(_02191_),
    .B1(_03391_));
 sg13g2_buf_2 _19232_ (.A(_03380_),
    .X(_03392_));
 sg13g2_nand2_1 _19233_ (.Y(_03393_),
    .A(\top_ihp.oisc.regs[58][20] ),
    .B(_03392_));
 sg13g2_o21ai_1 _19234_ (.B1(_03393_),
    .Y(_02192_),
    .A1(net36),
    .A2(net504));
 sg13g2_buf_1 _19235_ (.A(_03380_),
    .X(_03394_));
 sg13g2_nand2_1 _19236_ (.Y(_03395_),
    .A(\top_ihp.oisc.regs[58][21] ),
    .B(net502));
 sg13g2_o21ai_1 _19237_ (.B1(_03395_),
    .Y(_02193_),
    .A1(net82),
    .A2(_03394_));
 sg13g2_nand2_1 _19238_ (.Y(_03396_),
    .A(\top_ihp.oisc.regs[58][22] ),
    .B(net502));
 sg13g2_o21ai_1 _19239_ (.B1(_03396_),
    .Y(_02194_),
    .A1(net81),
    .A2(net501));
 sg13g2_nand2_1 _19240_ (.Y(_03397_),
    .A(\top_ihp.oisc.regs[58][23] ),
    .B(net502));
 sg13g2_o21ai_1 _19241_ (.B1(_03397_),
    .Y(_02195_),
    .A1(net207),
    .A2(net501));
 sg13g2_mux2_1 _19242_ (.A0(\top_ihp.oisc.regs[58][24] ),
    .A1(net403),
    .S(net640),
    .X(_02196_));
 sg13g2_nand2_1 _19243_ (.Y(_03398_),
    .A(\top_ihp.oisc.regs[58][25] ),
    .B(net502));
 sg13g2_o21ai_1 _19244_ (.B1(_03398_),
    .Y(_02197_),
    .A1(_10428_),
    .A2(net501));
 sg13g2_nand2_1 _19245_ (.Y(_03399_),
    .A(\top_ihp.oisc.regs[58][26] ),
    .B(net502));
 sg13g2_o21ai_1 _19246_ (.B1(_03399_),
    .Y(_02198_),
    .A1(net206),
    .A2(net501));
 sg13g2_nand2_1 _19247_ (.Y(_03400_),
    .A(\top_ihp.oisc.regs[58][27] ),
    .B(net502));
 sg13g2_o21ai_1 _19248_ (.B1(_03400_),
    .Y(_02199_),
    .A1(_10449_),
    .A2(net501));
 sg13g2_nand2_1 _19249_ (.Y(_03401_),
    .A(\top_ihp.oisc.regs[58][28] ),
    .B(_03392_));
 sg13g2_o21ai_1 _19250_ (.B1(_03401_),
    .Y(_02200_),
    .A1(net27),
    .A2(net501));
 sg13g2_nand2_1 _19251_ (.Y(_03402_),
    .A(\top_ihp.oisc.regs[58][29] ),
    .B(net502));
 sg13g2_o21ai_1 _19252_ (.B1(_03402_),
    .Y(_02201_),
    .A1(net80),
    .A2(net501));
 sg13g2_nand2_1 _19253_ (.Y(_03403_),
    .A(\top_ihp.oisc.regs[58][2] ),
    .B(net502));
 sg13g2_o21ai_1 _19254_ (.B1(_03403_),
    .Y(_02202_),
    .A1(net79),
    .A2(_03394_));
 sg13g2_nand2_1 _19255_ (.Y(_03404_),
    .A(\top_ihp.oisc.regs[58][30] ),
    .B(_03380_));
 sg13g2_o21ai_1 _19256_ (.B1(_03404_),
    .Y(_02203_),
    .A1(net35),
    .A2(net501));
 sg13g2_inv_1 _19257_ (.Y(_03405_),
    .A(\top_ihp.oisc.regs[58][31] ));
 sg13g2_nor2_1 _19258_ (.A(_10535_),
    .B(_03380_),
    .Y(_03406_));
 sg13g2_a22oi_1 _19259_ (.Y(_02204_),
    .B1(_03406_),
    .B2(net268),
    .A2(net504),
    .A1(_03405_));
 sg13g2_mux2_1 _19260_ (.A0(\top_ihp.oisc.regs[58][3] ),
    .A1(net135),
    .S(_03377_),
    .X(_02205_));
 sg13g2_mux2_1 _19261_ (.A0(\top_ihp.oisc.regs[58][4] ),
    .A1(net134),
    .S(net640),
    .X(_02206_));
 sg13g2_mux2_1 _19262_ (.A0(\top_ihp.oisc.regs[58][5] ),
    .A1(net267),
    .S(net640),
    .X(_02207_));
 sg13g2_mux2_1 _19263_ (.A0(\top_ihp.oisc.regs[58][6] ),
    .A1(net132),
    .S(net640),
    .X(_02208_));
 sg13g2_nand2_1 _19264_ (.Y(_03407_),
    .A(\top_ihp.oisc.regs[58][7] ),
    .B(_03380_));
 sg13g2_o21ai_1 _19265_ (.B1(_03407_),
    .Y(_02209_),
    .A1(_03281_),
    .A2(net503));
 sg13g2_nand2_1 _19266_ (.Y(_03408_),
    .A(\top_ihp.oisc.regs[58][8] ),
    .B(_03380_));
 sg13g2_o21ai_1 _19267_ (.B1(_03408_),
    .Y(_02210_),
    .A1(net205),
    .A2(net503));
 sg13g2_mux2_1 _19268_ (.A0(\top_ihp.oisc.regs[58][9] ),
    .A1(net131),
    .S(net640),
    .X(_02211_));
 sg13g2_nand2_1 _19269_ (.Y(_03409_),
    .A(_10694_),
    .B(_03150_));
 sg13g2_buf_2 _19270_ (.A(_03409_),
    .X(_03410_));
 sg13g2_buf_2 _19271_ (.A(_03410_),
    .X(_03411_));
 sg13g2_mux2_1 _19272_ (.A0(net119),
    .A1(\top_ihp.oisc.regs[59][0] ),
    .S(net500),
    .X(_02212_));
 sg13g2_mux2_1 _19273_ (.A0(net45),
    .A1(\top_ihp.oisc.regs[59][10] ),
    .S(net500),
    .X(_02213_));
 sg13g2_buf_1 _19274_ (.A(_03410_),
    .X(_03412_));
 sg13g2_buf_1 _19275_ (.A(_03410_),
    .X(_03413_));
 sg13g2_nand2_1 _19276_ (.Y(_03414_),
    .A(\top_ihp.oisc.regs[59][11] ),
    .B(net498));
 sg13g2_o21ai_1 _19277_ (.B1(_03414_),
    .Y(_02214_),
    .A1(net37),
    .A2(net499));
 sg13g2_nand2_1 _19278_ (.Y(_03415_),
    .A(\top_ihp.oisc.regs[59][12] ),
    .B(net498));
 sg13g2_o21ai_1 _19279_ (.B1(_03415_),
    .Y(_02215_),
    .A1(net141),
    .A2(net499));
 sg13g2_nand2_1 _19280_ (.Y(_03416_),
    .A(\top_ihp.oisc.regs[59][13] ),
    .B(net498));
 sg13g2_o21ai_1 _19281_ (.B1(_03416_),
    .Y(_02216_),
    .A1(net86),
    .A2(net499));
 sg13g2_nand2_1 _19282_ (.Y(_03417_),
    .A(\top_ihp.oisc.regs[59][14] ),
    .B(_03413_));
 sg13g2_o21ai_1 _19283_ (.B1(_03417_),
    .Y(_02217_),
    .A1(net85),
    .A2(net499));
 sg13g2_mux2_1 _19284_ (.A0(net663),
    .A1(\top_ihp.oisc.regs[59][15] ),
    .S(net500),
    .X(_02218_));
 sg13g2_nand2_1 _19285_ (.Y(_03418_),
    .A(\top_ihp.oisc.regs[59][16] ),
    .B(_03413_));
 sg13g2_o21ai_1 _19286_ (.B1(_03418_),
    .Y(_02219_),
    .A1(net84),
    .A2(_03412_));
 sg13g2_nand2_1 _19287_ (.Y(_03419_),
    .A(\top_ihp.oisc.regs[59][17] ),
    .B(net498));
 sg13g2_o21ai_1 _19288_ (.B1(_03419_),
    .Y(_02220_),
    .A1(net208),
    .A2(net499));
 sg13g2_nand2_1 _19289_ (.Y(_03420_),
    .A(\top_ihp.oisc.regs[59][18] ),
    .B(net498));
 sg13g2_o21ai_1 _19290_ (.B1(_03420_),
    .Y(_02221_),
    .A1(net83),
    .A2(net499));
 sg13g2_mux2_1 _19291_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[59][19] ),
    .S(net500),
    .X(_02222_));
 sg13g2_nand2_1 _19292_ (.Y(_03421_),
    .A(\top_ihp.oisc.regs[59][1] ),
    .B(net498));
 sg13g2_o21ai_1 _19293_ (.B1(_03421_),
    .Y(_02223_),
    .A1(net274),
    .A2(net499));
 sg13g2_buf_1 _19294_ (.A(_03410_),
    .X(_03422_));
 sg13g2_nand2_1 _19295_ (.Y(_03423_),
    .A(\top_ihp.oisc.regs[59][20] ),
    .B(_03422_));
 sg13g2_o21ai_1 _19296_ (.B1(_03423_),
    .Y(_02224_),
    .A1(net36),
    .A2(_03412_));
 sg13g2_nand2_1 _19297_ (.Y(_03424_),
    .A(\top_ihp.oisc.regs[59][21] ),
    .B(net497));
 sg13g2_o21ai_1 _19298_ (.B1(_03424_),
    .Y(_02225_),
    .A1(net82),
    .A2(net499));
 sg13g2_buf_1 _19299_ (.A(_03410_),
    .X(_03425_));
 sg13g2_nand2_1 _19300_ (.Y(_03426_),
    .A(\top_ihp.oisc.regs[59][22] ),
    .B(net497));
 sg13g2_o21ai_1 _19301_ (.B1(_03426_),
    .Y(_02226_),
    .A1(net81),
    .A2(net496));
 sg13g2_nand2_1 _19302_ (.Y(_03427_),
    .A(\top_ihp.oisc.regs[59][23] ),
    .B(net497));
 sg13g2_o21ai_1 _19303_ (.B1(_03427_),
    .Y(_02227_),
    .A1(net207),
    .A2(net496));
 sg13g2_mux2_1 _19304_ (.A0(net232),
    .A1(\top_ihp.oisc.regs[59][24] ),
    .S(net500),
    .X(_02228_));
 sg13g2_nand2_1 _19305_ (.Y(_03428_),
    .A(\top_ihp.oisc.regs[59][25] ),
    .B(net497));
 sg13g2_o21ai_1 _19306_ (.B1(_03428_),
    .Y(_02229_),
    .A1(net262),
    .A2(net496));
 sg13g2_nand2_1 _19307_ (.Y(_03429_),
    .A(\top_ihp.oisc.regs[59][26] ),
    .B(net497));
 sg13g2_o21ai_1 _19308_ (.B1(_03429_),
    .Y(_02230_),
    .A1(net206),
    .A2(net496));
 sg13g2_mux2_1 _19309_ (.A0(_10940_),
    .A1(\top_ihp.oisc.regs[59][27] ),
    .S(net500),
    .X(_02231_));
 sg13g2_nand2_1 _19310_ (.Y(_03430_),
    .A(\top_ihp.oisc.regs[59][28] ),
    .B(_03422_));
 sg13g2_o21ai_1 _19311_ (.B1(_03430_),
    .Y(_02232_),
    .A1(net27),
    .A2(_03425_));
 sg13g2_nand2_1 _19312_ (.Y(_03431_),
    .A(\top_ihp.oisc.regs[59][29] ),
    .B(net497));
 sg13g2_o21ai_1 _19313_ (.B1(_03431_),
    .Y(_02233_),
    .A1(net80),
    .A2(net496));
 sg13g2_nand2_1 _19314_ (.Y(_03432_),
    .A(\top_ihp.oisc.regs[59][2] ),
    .B(net497));
 sg13g2_o21ai_1 _19315_ (.B1(_03432_),
    .Y(_02234_),
    .A1(_03310_),
    .A2(net496));
 sg13g2_nand2_1 _19316_ (.Y(_03433_),
    .A(\top_ihp.oisc.regs[59][30] ),
    .B(net497));
 sg13g2_o21ai_1 _19317_ (.B1(_03433_),
    .Y(_02235_),
    .A1(net35),
    .A2(net496));
 sg13g2_nand2_1 _19318_ (.Y(_03434_),
    .A(\top_ihp.oisc.regs[59][31] ),
    .B(_03410_));
 sg13g2_o21ai_1 _19319_ (.B1(_03434_),
    .Y(_02236_),
    .A1(net87),
    .A2(net496));
 sg13g2_mux2_1 _19320_ (.A0(net44),
    .A1(\top_ihp.oisc.regs[59][3] ),
    .S(_03411_),
    .X(_02237_));
 sg13g2_mux2_1 _19321_ (.A0(net43),
    .A1(\top_ihp.oisc.regs[59][4] ),
    .S(net500),
    .X(_02238_));
 sg13g2_mux2_1 _19322_ (.A0(_11221_),
    .A1(\top_ihp.oisc.regs[59][5] ),
    .S(_03411_),
    .X(_02239_));
 sg13g2_mux2_1 _19323_ (.A0(net42),
    .A1(\top_ihp.oisc.regs[59][6] ),
    .S(net498),
    .X(_02240_));
 sg13g2_nand2_1 _19324_ (.Y(_03435_),
    .A(\top_ihp.oisc.regs[59][7] ),
    .B(_03410_));
 sg13g2_o21ai_1 _19325_ (.B1(_03435_),
    .Y(_02241_),
    .A1(net343),
    .A2(_03425_));
 sg13g2_nand2_1 _19326_ (.Y(_03436_),
    .A(\top_ihp.oisc.regs[59][8] ),
    .B(_03410_));
 sg13g2_o21ai_1 _19327_ (.B1(_03436_),
    .Y(_02242_),
    .A1(_03283_),
    .A2(net500));
 sg13g2_mux2_1 _19328_ (.A0(net41),
    .A1(\top_ihp.oisc.regs[59][9] ),
    .S(net498),
    .X(_02243_));
 sg13g2_nor2_1 _19329_ (.A(_10913_),
    .B(_11080_),
    .Y(_03437_));
 sg13g2_buf_1 _19330_ (.A(_03437_),
    .X(_03438_));
 sg13g2_buf_1 _19331_ (.A(_03438_),
    .X(_03439_));
 sg13g2_mux2_1 _19332_ (.A0(\top_ihp.oisc.regs[5][0] ),
    .A1(net143),
    .S(net639),
    .X(_02244_));
 sg13g2_mux2_1 _19333_ (.A0(\top_ihp.oisc.regs[5][10] ),
    .A1(net142),
    .S(net639),
    .X(_02245_));
 sg13g2_nor2_1 _19334_ (.A(\top_ihp.oisc.regs[5][11] ),
    .B(net689),
    .Y(_03440_));
 sg13g2_a21oi_1 _19335_ (.A1(net62),
    .A2(net639),
    .Y(_02246_),
    .B1(_03440_));
 sg13g2_nor2_1 _19336_ (.A(\top_ihp.oisc.regs[5][12] ),
    .B(net689),
    .Y(_03441_));
 sg13g2_a21oi_1 _19337_ (.A1(net61),
    .A2(net639),
    .Y(_02247_),
    .B1(_03441_));
 sg13g2_nand2_1 _19338_ (.Y(_03442_),
    .A(_10824_),
    .B(net729));
 sg13g2_buf_1 _19339_ (.A(_03442_),
    .X(_03443_));
 sg13g2_buf_1 _19340_ (.A(net638),
    .X(_03444_));
 sg13g2_buf_1 _19341_ (.A(_03443_),
    .X(_03445_));
 sg13g2_nand2_1 _19342_ (.Y(_03446_),
    .A(\top_ihp.oisc.regs[5][13] ),
    .B(net494));
 sg13g2_o21ai_1 _19343_ (.B1(_03446_),
    .Y(_02248_),
    .A1(_03244_),
    .A2(_03444_));
 sg13g2_nand2_1 _19344_ (.Y(_03447_),
    .A(\top_ihp.oisc.regs[5][14] ),
    .B(net494));
 sg13g2_o21ai_1 _19345_ (.B1(_03447_),
    .Y(_02249_),
    .A1(_03250_),
    .A2(net495));
 sg13g2_buf_1 _19346_ (.A(net638),
    .X(_03448_));
 sg13g2_nand2_1 _19347_ (.Y(_03449_),
    .A(\top_ihp.oisc.regs[5][15] ),
    .B(net493));
 sg13g2_o21ai_1 _19348_ (.B1(_03449_),
    .Y(_02250_),
    .A1(_03127_),
    .A2(net495));
 sg13g2_nand2_1 _19349_ (.Y(_03450_),
    .A(\top_ihp.oisc.regs[5][16] ),
    .B(_03448_));
 sg13g2_o21ai_1 _19350_ (.B1(_03450_),
    .Y(_02251_),
    .A1(_03254_),
    .A2(_03444_));
 sg13g2_nand2_1 _19351_ (.Y(_03451_),
    .A(\top_ihp.oisc.regs[5][17] ),
    .B(net493));
 sg13g2_o21ai_1 _19352_ (.B1(_03451_),
    .Y(_02252_),
    .A1(_03256_),
    .A2(net495));
 sg13g2_nand2_1 _19353_ (.Y(_03452_),
    .A(\top_ihp.oisc.regs[5][18] ),
    .B(net493));
 sg13g2_o21ai_1 _19354_ (.B1(_03452_),
    .Y(_02253_),
    .A1(_03258_),
    .A2(net495));
 sg13g2_mux2_1 _19355_ (.A0(\top_ihp.oisc.regs[5][19] ),
    .A1(_11275_),
    .S(net639),
    .X(_02254_));
 sg13g2_nor2_1 _19356_ (.A(\top_ihp.oisc.regs[5][1] ),
    .B(net689),
    .Y(_03453_));
 sg13g2_a21oi_1 _19357_ (.A1(net139),
    .A2(_03439_),
    .Y(_02255_),
    .B1(_03453_));
 sg13g2_nand2_1 _19358_ (.Y(_03454_),
    .A(\top_ihp.oisc.regs[5][20] ),
    .B(net493));
 sg13g2_o21ai_1 _19359_ (.B1(_03454_),
    .Y(_02256_),
    .A1(_03262_),
    .A2(net495));
 sg13g2_nand2_1 _19360_ (.Y(_03455_),
    .A(\top_ihp.oisc.regs[5][21] ),
    .B(net493));
 sg13g2_o21ai_1 _19361_ (.B1(_03455_),
    .Y(_02257_),
    .A1(_03264_),
    .A2(net495));
 sg13g2_nand2_1 _19362_ (.Y(_03456_),
    .A(\top_ihp.oisc.regs[5][22] ),
    .B(net493));
 sg13g2_o21ai_1 _19363_ (.B1(_03456_),
    .Y(_02258_),
    .A1(_03266_),
    .A2(net495));
 sg13g2_nand2_1 _19364_ (.Y(_03457_),
    .A(\top_ihp.oisc.regs[5][23] ),
    .B(_03448_));
 sg13g2_o21ai_1 _19365_ (.B1(_03457_),
    .Y(_02259_),
    .A1(_03268_),
    .A2(net495));
 sg13g2_mux2_1 _19366_ (.A0(\top_ihp.oisc.regs[5][24] ),
    .A1(net403),
    .S(net639),
    .X(_02260_));
 sg13g2_nand2_1 _19367_ (.Y(_03458_),
    .A(\top_ihp.oisc.regs[5][25] ),
    .B(net493));
 sg13g2_o21ai_1 _19368_ (.B1(_03458_),
    .Y(_02261_),
    .A1(_10772_),
    .A2(net494));
 sg13g2_nand2_1 _19369_ (.Y(_03459_),
    .A(\top_ihp.oisc.regs[5][26] ),
    .B(net493));
 sg13g2_o21ai_1 _19370_ (.B1(_03459_),
    .Y(_02262_),
    .A1(_03271_),
    .A2(_03445_));
 sg13g2_mux2_1 _19371_ (.A0(\top_ihp.oisc.regs[5][27] ),
    .A1(net101),
    .S(net639),
    .X(_02263_));
 sg13g2_nor2_1 _19372_ (.A(\top_ihp.oisc.regs[5][28] ),
    .B(net689),
    .Y(_03460_));
 sg13g2_a21oi_1 _19373_ (.A1(_10941_),
    .A2(_03439_),
    .Y(_02264_),
    .B1(_03460_));
 sg13g2_nand2_1 _19374_ (.Y(_03461_),
    .A(\top_ihp.oisc.regs[5][29] ),
    .B(net638));
 sg13g2_o21ai_1 _19375_ (.B1(_03461_),
    .Y(_02265_),
    .A1(_03275_),
    .A2(_03445_));
 sg13g2_nand2_1 _19376_ (.Y(_03462_),
    .A(\top_ihp.oisc.regs[5][2] ),
    .B(net638));
 sg13g2_o21ai_1 _19377_ (.B1(_03462_),
    .Y(_02266_),
    .A1(_03310_),
    .A2(net494));
 sg13g2_nand2_1 _19378_ (.Y(_03463_),
    .A(\top_ihp.oisc.regs[5][30] ),
    .B(net638));
 sg13g2_o21ai_1 _19379_ (.B1(_03463_),
    .Y(_02267_),
    .A1(_03312_),
    .A2(net494));
 sg13g2_nand2_1 _19380_ (.Y(_03464_),
    .A(\top_ihp.oisc.regs[5][31] ),
    .B(net638));
 sg13g2_o21ai_1 _19381_ (.B1(_03464_),
    .Y(_02268_),
    .A1(_03074_),
    .A2(net494));
 sg13g2_mux2_1 _19382_ (.A0(\top_ihp.oisc.regs[5][3] ),
    .A1(net135),
    .S(net639),
    .X(_02269_));
 sg13g2_mux2_1 _19383_ (.A0(\top_ihp.oisc.regs[5][4] ),
    .A1(net134),
    .S(net689),
    .X(_02270_));
 sg13g2_mux2_1 _19384_ (.A0(\top_ihp.oisc.regs[5][5] ),
    .A1(net267),
    .S(net689),
    .X(_02271_));
 sg13g2_mux2_1 _19385_ (.A0(\top_ihp.oisc.regs[5][6] ),
    .A1(net132),
    .S(net689),
    .X(_02272_));
 sg13g2_nand2_1 _19386_ (.Y(_03465_),
    .A(\top_ihp.oisc.regs[5][7] ),
    .B(net638));
 sg13g2_o21ai_1 _19387_ (.B1(_03465_),
    .Y(_02273_),
    .A1(_03281_),
    .A2(net494));
 sg13g2_nand2_1 _19388_ (.Y(_03466_),
    .A(\top_ihp.oisc.regs[5][8] ),
    .B(net638));
 sg13g2_o21ai_1 _19389_ (.B1(_03466_),
    .Y(_02274_),
    .A1(_03283_),
    .A2(net494));
 sg13g2_mux2_1 _19390_ (.A0(\top_ihp.oisc.regs[5][9] ),
    .A1(net131),
    .S(net689),
    .X(_02275_));
 sg13g2_nand2_1 _19391_ (.Y(_03467_),
    .A(_10787_),
    .B(_03015_));
 sg13g2_buf_1 _19392_ (.A(_03467_),
    .X(_03468_));
 sg13g2_buf_2 _19393_ (.A(net637),
    .X(_03469_));
 sg13g2_mux2_1 _19394_ (.A0(net119),
    .A1(\top_ihp.oisc.regs[60][0] ),
    .S(_03469_),
    .X(_02276_));
 sg13g2_mux2_1 _19395_ (.A0(net130),
    .A1(\top_ihp.oisc.regs[60][10] ),
    .S(net492),
    .X(_02277_));
 sg13g2_buf_1 _19396_ (.A(net637),
    .X(_03470_));
 sg13g2_buf_1 _19397_ (.A(_03468_),
    .X(_03471_));
 sg13g2_nand2_1 _19398_ (.Y(_03472_),
    .A(\top_ihp.oisc.regs[60][11] ),
    .B(net490));
 sg13g2_o21ai_1 _19399_ (.B1(_03472_),
    .Y(_02278_),
    .A1(net37),
    .A2(net491));
 sg13g2_nand2_1 _19400_ (.Y(_03473_),
    .A(\top_ihp.oisc.regs[60][12] ),
    .B(net490));
 sg13g2_o21ai_1 _19401_ (.B1(_03473_),
    .Y(_02279_),
    .A1(net141),
    .A2(net491));
 sg13g2_nand2_1 _19402_ (.Y(_03474_),
    .A(\top_ihp.oisc.regs[60][13] ),
    .B(_03471_));
 sg13g2_o21ai_1 _19403_ (.B1(_03474_),
    .Y(_02280_),
    .A1(net86),
    .A2(net491));
 sg13g2_nand2_1 _19404_ (.Y(_03475_),
    .A(\top_ihp.oisc.regs[60][14] ),
    .B(net490));
 sg13g2_o21ai_1 _19405_ (.B1(_03475_),
    .Y(_02281_),
    .A1(net85),
    .A2(_03470_));
 sg13g2_nand2_1 _19406_ (.Y(_03476_),
    .A(\top_ihp.oisc.regs[60][15] ),
    .B(net490));
 sg13g2_o21ai_1 _19407_ (.B1(_03476_),
    .Y(_02282_),
    .A1(net209),
    .A2(net491));
 sg13g2_nand2_1 _19408_ (.Y(_03477_),
    .A(\top_ihp.oisc.regs[60][16] ),
    .B(net490));
 sg13g2_o21ai_1 _19409_ (.B1(_03477_),
    .Y(_02283_),
    .A1(net84),
    .A2(_03470_));
 sg13g2_nand2_1 _19410_ (.Y(_03478_),
    .A(\top_ihp.oisc.regs[60][17] ),
    .B(net490));
 sg13g2_o21ai_1 _19411_ (.B1(_03478_),
    .Y(_02284_),
    .A1(net208),
    .A2(net491));
 sg13g2_nand2_1 _19412_ (.Y(_03479_),
    .A(\top_ihp.oisc.regs[60][18] ),
    .B(_03471_));
 sg13g2_o21ai_1 _19413_ (.B1(_03479_),
    .Y(_02285_),
    .A1(net83),
    .A2(net491));
 sg13g2_mux2_1 _19414_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[60][19] ),
    .S(net492),
    .X(_02286_));
 sg13g2_buf_2 _19415_ (.A(net637),
    .X(_03480_));
 sg13g2_nand2_1 _19416_ (.Y(_03481_),
    .A(\top_ihp.oisc.regs[60][1] ),
    .B(net489));
 sg13g2_o21ai_1 _19417_ (.B1(_03481_),
    .Y(_02287_),
    .A1(net274),
    .A2(net491));
 sg13g2_nand2_1 _19418_ (.Y(_03482_),
    .A(\top_ihp.oisc.regs[60][20] ),
    .B(_03480_));
 sg13g2_o21ai_1 _19419_ (.B1(_03482_),
    .Y(_02288_),
    .A1(net36),
    .A2(net491));
 sg13g2_buf_1 _19420_ (.A(net637),
    .X(_03483_));
 sg13g2_nand2_1 _19421_ (.Y(_03484_),
    .A(\top_ihp.oisc.regs[60][21] ),
    .B(_03480_));
 sg13g2_o21ai_1 _19422_ (.B1(_03484_),
    .Y(_02289_),
    .A1(net82),
    .A2(_03483_));
 sg13g2_nand2_1 _19423_ (.Y(_03485_),
    .A(\top_ihp.oisc.regs[60][22] ),
    .B(net489));
 sg13g2_o21ai_1 _19424_ (.B1(_03485_),
    .Y(_02290_),
    .A1(net81),
    .A2(net488));
 sg13g2_nand2_1 _19425_ (.Y(_03486_),
    .A(\top_ihp.oisc.regs[60][23] ),
    .B(net489));
 sg13g2_o21ai_1 _19426_ (.B1(_03486_),
    .Y(_02291_),
    .A1(net207),
    .A2(net488));
 sg13g2_mux2_1 _19427_ (.A0(net400),
    .A1(\top_ihp.oisc.regs[60][24] ),
    .S(net492),
    .X(_02292_));
 sg13g2_nand2_1 _19428_ (.Y(_03487_),
    .A(\top_ihp.oisc.regs[60][25] ),
    .B(net489));
 sg13g2_o21ai_1 _19429_ (.B1(_03487_),
    .Y(_02293_),
    .A1(net262),
    .A2(net488));
 sg13g2_nand2_1 _19430_ (.Y(_03488_),
    .A(\top_ihp.oisc.regs[60][26] ),
    .B(net489));
 sg13g2_o21ai_1 _19431_ (.B1(_03488_),
    .Y(_02294_),
    .A1(net206),
    .A2(net488));
 sg13g2_mux2_1 _19432_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[60][27] ),
    .S(net492),
    .X(_02295_));
 sg13g2_nand2_1 _19433_ (.Y(_03489_),
    .A(\top_ihp.oisc.regs[60][28] ),
    .B(net489));
 sg13g2_o21ai_1 _19434_ (.B1(_03489_),
    .Y(_02296_),
    .A1(net27),
    .A2(net488));
 sg13g2_nand2_1 _19435_ (.Y(_03490_),
    .A(\top_ihp.oisc.regs[60][29] ),
    .B(net489));
 sg13g2_o21ai_1 _19436_ (.B1(_03490_),
    .Y(_02297_),
    .A1(net80),
    .A2(net488));
 sg13g2_nand2_1 _19437_ (.Y(_03491_),
    .A(\top_ihp.oisc.regs[60][2] ),
    .B(net489));
 sg13g2_o21ai_1 _19438_ (.B1(_03491_),
    .Y(_02298_),
    .A1(net79),
    .A2(net488));
 sg13g2_nand2_1 _19439_ (.Y(_03492_),
    .A(\top_ihp.oisc.regs[60][30] ),
    .B(net637));
 sg13g2_o21ai_1 _19440_ (.B1(_03492_),
    .Y(_02299_),
    .A1(net35),
    .A2(net488));
 sg13g2_nand2_1 _19441_ (.Y(_03493_),
    .A(\top_ihp.oisc.regs[60][31] ),
    .B(net637));
 sg13g2_o21ai_1 _19442_ (.B1(_03493_),
    .Y(_02300_),
    .A1(net87),
    .A2(_03483_));
 sg13g2_mux2_1 _19443_ (.A0(net128),
    .A1(\top_ihp.oisc.regs[60][3] ),
    .S(net492),
    .X(_02301_));
 sg13g2_mux2_1 _19444_ (.A0(net127),
    .A1(\top_ihp.oisc.regs[60][4] ),
    .S(net492),
    .X(_02302_));
 sg13g2_mux2_1 _19445_ (.A0(net264),
    .A1(\top_ihp.oisc.regs[60][5] ),
    .S(net492),
    .X(_02303_));
 sg13g2_mux2_1 _19446_ (.A0(net126),
    .A1(\top_ihp.oisc.regs[60][6] ),
    .S(net490),
    .X(_02304_));
 sg13g2_nand2_1 _19447_ (.Y(_03494_),
    .A(\top_ihp.oisc.regs[60][7] ),
    .B(net637));
 sg13g2_o21ai_1 _19448_ (.B1(_03494_),
    .Y(_02305_),
    .A1(net343),
    .A2(net492));
 sg13g2_nand2_1 _19449_ (.Y(_03495_),
    .A(\top_ihp.oisc.regs[60][8] ),
    .B(net637));
 sg13g2_o21ai_1 _19450_ (.B1(_03495_),
    .Y(_02306_),
    .A1(net205),
    .A2(_03469_));
 sg13g2_mux2_1 _19451_ (.A0(net125),
    .A1(\top_ihp.oisc.regs[60][9] ),
    .S(net490),
    .X(_02307_));
 sg13g2_nor2_1 _19452_ (.A(_10847_),
    .B(_03047_),
    .Y(_03496_));
 sg13g2_buf_1 _19453_ (.A(_03496_),
    .X(_03497_));
 sg13g2_buf_2 _19454_ (.A(net636),
    .X(_03498_));
 sg13g2_mux2_1 _19455_ (.A0(\top_ihp.oisc.regs[61][0] ),
    .A1(net143),
    .S(net487),
    .X(_02308_));
 sg13g2_mux2_1 _19456_ (.A0(\top_ihp.oisc.regs[61][10] ),
    .A1(net142),
    .S(net487),
    .X(_02309_));
 sg13g2_nor2_1 _19457_ (.A(\top_ihp.oisc.regs[61][11] ),
    .B(net636),
    .Y(_03499_));
 sg13g2_a21oi_1 _19458_ (.A1(_10041_),
    .A2(net487),
    .Y(_02310_),
    .B1(_03499_));
 sg13g2_nor2_1 _19459_ (.A(\top_ihp.oisc.regs[61][12] ),
    .B(net636),
    .Y(_03500_));
 sg13g2_a21oi_1 _19460_ (.A1(net61),
    .A2(_03498_),
    .Y(_02311_),
    .B1(_03500_));
 sg13g2_or2_1 _19461_ (.X(_03501_),
    .B(_03047_),
    .A(_10847_));
 sg13g2_buf_1 _19462_ (.A(_03501_),
    .X(_03502_));
 sg13g2_buf_2 _19463_ (.A(net635),
    .X(_03503_));
 sg13g2_buf_2 _19464_ (.A(net635),
    .X(_03504_));
 sg13g2_nand2_1 _19465_ (.Y(_03505_),
    .A(\top_ihp.oisc.regs[61][13] ),
    .B(_03504_));
 sg13g2_o21ai_1 _19466_ (.B1(_03505_),
    .Y(_02312_),
    .A1(net86),
    .A2(net486));
 sg13g2_nand2_1 _19467_ (.Y(_03506_),
    .A(\top_ihp.oisc.regs[61][14] ),
    .B(net485));
 sg13g2_o21ai_1 _19468_ (.B1(_03506_),
    .Y(_02313_),
    .A1(net85),
    .A2(_03503_));
 sg13g2_buf_2 _19469_ (.A(net635),
    .X(_03507_));
 sg13g2_nand2_1 _19470_ (.Y(_03508_),
    .A(\top_ihp.oisc.regs[61][15] ),
    .B(net484));
 sg13g2_o21ai_1 _19471_ (.B1(_03508_),
    .Y(_02314_),
    .A1(net209),
    .A2(net486));
 sg13g2_nand2_1 _19472_ (.Y(_03509_),
    .A(\top_ihp.oisc.regs[61][16] ),
    .B(net484));
 sg13g2_o21ai_1 _19473_ (.B1(_03509_),
    .Y(_02315_),
    .A1(net84),
    .A2(net486));
 sg13g2_nand2_1 _19474_ (.Y(_03510_),
    .A(\top_ihp.oisc.regs[61][17] ),
    .B(_03507_));
 sg13g2_o21ai_1 _19475_ (.B1(_03510_),
    .Y(_02316_),
    .A1(net208),
    .A2(_03503_));
 sg13g2_nand2_1 _19476_ (.Y(_03511_),
    .A(\top_ihp.oisc.regs[61][18] ),
    .B(_03507_));
 sg13g2_o21ai_1 _19477_ (.B1(_03511_),
    .Y(_02317_),
    .A1(net83),
    .A2(net486));
 sg13g2_mux2_1 _19478_ (.A0(\top_ihp.oisc.regs[61][19] ),
    .A1(net227),
    .S(net487),
    .X(_02318_));
 sg13g2_nor2_1 _19479_ (.A(\top_ihp.oisc.regs[61][1] ),
    .B(net636),
    .Y(_03512_));
 sg13g2_a21oi_1 _19480_ (.A1(net139),
    .A2(net487),
    .Y(_02319_),
    .B1(_03512_));
 sg13g2_nand2_1 _19481_ (.Y(_03513_),
    .A(\top_ihp.oisc.regs[61][20] ),
    .B(net484));
 sg13g2_o21ai_1 _19482_ (.B1(_03513_),
    .Y(_02320_),
    .A1(net36),
    .A2(net486));
 sg13g2_nand2_1 _19483_ (.Y(_03514_),
    .A(\top_ihp.oisc.regs[61][21] ),
    .B(net484));
 sg13g2_o21ai_1 _19484_ (.B1(_03514_),
    .Y(_02321_),
    .A1(net82),
    .A2(net486));
 sg13g2_nand2_1 _19485_ (.Y(_03515_),
    .A(\top_ihp.oisc.regs[61][22] ),
    .B(net484));
 sg13g2_o21ai_1 _19486_ (.B1(_03515_),
    .Y(_02322_),
    .A1(net81),
    .A2(net486));
 sg13g2_nand2_1 _19487_ (.Y(_03516_),
    .A(\top_ihp.oisc.regs[61][23] ),
    .B(net484));
 sg13g2_o21ai_1 _19488_ (.B1(_03516_),
    .Y(_02323_),
    .A1(_03268_),
    .A2(net486));
 sg13g2_mux2_1 _19489_ (.A0(\top_ihp.oisc.regs[61][24] ),
    .A1(net403),
    .S(net487),
    .X(_02324_));
 sg13g2_nand2_1 _19490_ (.Y(_03517_),
    .A(\top_ihp.oisc.regs[61][25] ),
    .B(net484));
 sg13g2_o21ai_1 _19491_ (.B1(_03517_),
    .Y(_02325_),
    .A1(net262),
    .A2(net485));
 sg13g2_nand2_1 _19492_ (.Y(_03518_),
    .A(\top_ihp.oisc.regs[61][26] ),
    .B(net484));
 sg13g2_o21ai_1 _19493_ (.B1(_03518_),
    .Y(_02326_),
    .A1(_03271_),
    .A2(_03504_));
 sg13g2_mux2_1 _19494_ (.A0(\top_ihp.oisc.regs[61][27] ),
    .A1(net101),
    .S(_03498_),
    .X(_02327_));
 sg13g2_nor2_1 _19495_ (.A(\top_ihp.oisc.regs[61][28] ),
    .B(net636),
    .Y(_03519_));
 sg13g2_a21oi_1 _19496_ (.A1(net116),
    .A2(net487),
    .Y(_02328_),
    .B1(_03519_));
 sg13g2_nand2_1 _19497_ (.Y(_03520_),
    .A(\top_ihp.oisc.regs[61][29] ),
    .B(net635));
 sg13g2_o21ai_1 _19498_ (.B1(_03520_),
    .Y(_02329_),
    .A1(net80),
    .A2(net485));
 sg13g2_nand2_1 _19499_ (.Y(_03521_),
    .A(\top_ihp.oisc.regs[61][2] ),
    .B(net635));
 sg13g2_o21ai_1 _19500_ (.B1(_03521_),
    .Y(_02330_),
    .A1(net79),
    .A2(net485));
 sg13g2_nand2_1 _19501_ (.Y(_03522_),
    .A(\top_ihp.oisc.regs[61][30] ),
    .B(net635));
 sg13g2_o21ai_1 _19502_ (.B1(_03522_),
    .Y(_02331_),
    .A1(net35),
    .A2(net485));
 sg13g2_nand2_1 _19503_ (.Y(_03523_),
    .A(\top_ihp.oisc.regs[61][31] ),
    .B(_03502_));
 sg13g2_o21ai_1 _19504_ (.B1(_03523_),
    .Y(_02332_),
    .A1(net265),
    .A2(net485));
 sg13g2_mux2_1 _19505_ (.A0(\top_ihp.oisc.regs[61][3] ),
    .A1(net135),
    .S(net487),
    .X(_02333_));
 sg13g2_mux2_1 _19506_ (.A0(\top_ihp.oisc.regs[61][4] ),
    .A1(net134),
    .S(net636),
    .X(_02334_));
 sg13g2_mux2_1 _19507_ (.A0(\top_ihp.oisc.regs[61][5] ),
    .A1(net267),
    .S(_03497_),
    .X(_02335_));
 sg13g2_mux2_1 _19508_ (.A0(\top_ihp.oisc.regs[61][6] ),
    .A1(net132),
    .S(net636),
    .X(_02336_));
 sg13g2_nand2_1 _19509_ (.Y(_03524_),
    .A(\top_ihp.oisc.regs[61][7] ),
    .B(net635));
 sg13g2_o21ai_1 _19510_ (.B1(_03524_),
    .Y(_02337_),
    .A1(net343),
    .A2(net485));
 sg13g2_nand2_1 _19511_ (.Y(_03525_),
    .A(\top_ihp.oisc.regs[61][8] ),
    .B(net635));
 sg13g2_o21ai_1 _19512_ (.B1(_03525_),
    .Y(_02338_),
    .A1(net205),
    .A2(net485));
 sg13g2_mux2_1 _19513_ (.A0(\top_ihp.oisc.regs[61][9] ),
    .A1(net131),
    .S(net636),
    .X(_02339_));
 sg13g2_nor2_1 _19514_ (.A(_10847_),
    .B(_03112_),
    .Y(_03526_));
 sg13g2_buf_1 _19515_ (.A(_03526_),
    .X(_03527_));
 sg13g2_buf_2 _19516_ (.A(net688),
    .X(_03528_));
 sg13g2_mux2_1 _19517_ (.A0(\top_ihp.oisc.regs[62][0] ),
    .A1(net143),
    .S(net634),
    .X(_02340_));
 sg13g2_mux2_1 _19518_ (.A0(\top_ihp.oisc.regs[62][10] ),
    .A1(net142),
    .S(net634),
    .X(_02341_));
 sg13g2_nor2_1 _19519_ (.A(\top_ihp.oisc.regs[62][11] ),
    .B(net688),
    .Y(_03529_));
 sg13g2_a21oi_1 _19520_ (.A1(net62),
    .A2(net634),
    .Y(_02342_),
    .B1(_03529_));
 sg13g2_nor2_1 _19521_ (.A(\top_ihp.oisc.regs[62][12] ),
    .B(_03527_),
    .Y(_03530_));
 sg13g2_a21oi_1 _19522_ (.A1(net61),
    .A2(net634),
    .Y(_02343_),
    .B1(_03530_));
 sg13g2_nand2_1 _19523_ (.Y(_03531_),
    .A(_10787_),
    .B(_03119_));
 sg13g2_buf_1 _19524_ (.A(_03531_),
    .X(_03532_));
 sg13g2_buf_1 _19525_ (.A(_03532_),
    .X(_03533_));
 sg13g2_buf_1 _19526_ (.A(_03531_),
    .X(_03534_));
 sg13g2_nand2_1 _19527_ (.Y(_03535_),
    .A(\top_ihp.oisc.regs[62][13] ),
    .B(_03534_));
 sg13g2_o21ai_1 _19528_ (.B1(_03535_),
    .Y(_02344_),
    .A1(net86),
    .A2(net483));
 sg13g2_buf_2 _19529_ (.A(net633),
    .X(_03536_));
 sg13g2_nand2_1 _19530_ (.Y(_03537_),
    .A(\top_ihp.oisc.regs[62][14] ),
    .B(net482));
 sg13g2_o21ai_1 _19531_ (.B1(_03537_),
    .Y(_02345_),
    .A1(net85),
    .A2(net483));
 sg13g2_nand2_1 _19532_ (.Y(_03538_),
    .A(\top_ihp.oisc.regs[62][15] ),
    .B(net482));
 sg13g2_o21ai_1 _19533_ (.B1(_03538_),
    .Y(_02346_),
    .A1(net399),
    .A2(net483));
 sg13g2_nand2_1 _19534_ (.Y(_03539_),
    .A(\top_ihp.oisc.regs[62][16] ),
    .B(net482));
 sg13g2_o21ai_1 _19535_ (.B1(_03539_),
    .Y(_02347_),
    .A1(net84),
    .A2(net483));
 sg13g2_nand2_1 _19536_ (.Y(_03540_),
    .A(\top_ihp.oisc.regs[62][17] ),
    .B(net482));
 sg13g2_o21ai_1 _19537_ (.B1(_03540_),
    .Y(_02348_),
    .A1(net208),
    .A2(net483));
 sg13g2_nand2_1 _19538_ (.Y(_03541_),
    .A(\top_ihp.oisc.regs[62][18] ),
    .B(net482));
 sg13g2_o21ai_1 _19539_ (.B1(_03541_),
    .Y(_02349_),
    .A1(net83),
    .A2(net483));
 sg13g2_nand2_1 _19540_ (.Y(_03542_),
    .A(\top_ihp.oisc.regs[62][19] ),
    .B(_03536_));
 sg13g2_o21ai_1 _19541_ (.B1(_03542_),
    .Y(_02350_),
    .A1(_10273_),
    .A2(net483));
 sg13g2_nor2_1 _19542_ (.A(\top_ihp.oisc.regs[62][1] ),
    .B(net688),
    .Y(_03543_));
 sg13g2_a21oi_1 _19543_ (.A1(net139),
    .A2(net634),
    .Y(_02351_),
    .B1(_03543_));
 sg13g2_nand2_1 _19544_ (.Y(_03544_),
    .A(\top_ihp.oisc.regs[62][20] ),
    .B(net482));
 sg13g2_o21ai_1 _19545_ (.B1(_03544_),
    .Y(_02352_),
    .A1(_03262_),
    .A2(_03533_));
 sg13g2_nand2_1 _19546_ (.Y(_03545_),
    .A(\top_ihp.oisc.regs[62][21] ),
    .B(_03536_));
 sg13g2_o21ai_1 _19547_ (.B1(_03545_),
    .Y(_02353_),
    .A1(net82),
    .A2(_03533_));
 sg13g2_nand2_1 _19548_ (.Y(_03546_),
    .A(\top_ihp.oisc.regs[62][22] ),
    .B(net482));
 sg13g2_o21ai_1 _19549_ (.B1(_03546_),
    .Y(_02354_),
    .A1(_03266_),
    .A2(_03534_));
 sg13g2_nand2_1 _19550_ (.Y(_03547_),
    .A(\top_ihp.oisc.regs[62][23] ),
    .B(net482));
 sg13g2_o21ai_1 _19551_ (.B1(_03547_),
    .Y(_02355_),
    .A1(net207),
    .A2(net632));
 sg13g2_mux2_1 _19552_ (.A0(\top_ihp.oisc.regs[62][24] ),
    .A1(net403),
    .S(net634),
    .X(_02356_));
 sg13g2_nor2_1 _19553_ (.A(\top_ihp.oisc.regs[62][25] ),
    .B(net688),
    .Y(_03548_));
 sg13g2_a21oi_1 _19554_ (.A1(net59),
    .A2(net634),
    .Y(_02357_),
    .B1(_03548_));
 sg13g2_nand2_1 _19555_ (.Y(_03549_),
    .A(\top_ihp.oisc.regs[62][26] ),
    .B(net633));
 sg13g2_o21ai_1 _19556_ (.B1(_03549_),
    .Y(_02358_),
    .A1(net206),
    .A2(net632));
 sg13g2_nand2_1 _19557_ (.Y(_03550_),
    .A(\top_ihp.oisc.regs[62][27] ),
    .B(net633));
 sg13g2_o21ai_1 _19558_ (.B1(_03550_),
    .Y(_02359_),
    .A1(_10449_),
    .A2(net632));
 sg13g2_nor2_1 _19559_ (.A(\top_ihp.oisc.regs[62][28] ),
    .B(net688),
    .Y(_03551_));
 sg13g2_a21oi_1 _19560_ (.A1(net30),
    .A2(net634),
    .Y(_02360_),
    .B1(_03551_));
 sg13g2_nand2_1 _19561_ (.Y(_03552_),
    .A(\top_ihp.oisc.regs[62][29] ),
    .B(net633));
 sg13g2_o21ai_1 _19562_ (.B1(_03552_),
    .Y(_02361_),
    .A1(net80),
    .A2(net632));
 sg13g2_nand2_1 _19563_ (.Y(_03553_),
    .A(\top_ihp.oisc.regs[62][2] ),
    .B(net633));
 sg13g2_o21ai_1 _19564_ (.B1(_03553_),
    .Y(_02362_),
    .A1(net79),
    .A2(net632));
 sg13g2_nand2_1 _19565_ (.Y(_03554_),
    .A(\top_ihp.oisc.regs[62][30] ),
    .B(net633));
 sg13g2_o21ai_1 _19566_ (.B1(_03554_),
    .Y(_02363_),
    .A1(net35),
    .A2(net632));
 sg13g2_inv_1 _19567_ (.Y(_03555_),
    .A(\top_ihp.oisc.regs[62][31] ));
 sg13g2_nor2_1 _19568_ (.A(_10535_),
    .B(_03532_),
    .Y(_03556_));
 sg13g2_a22oi_1 _19569_ (.Y(_02364_),
    .B1(_03556_),
    .B2(net268),
    .A2(net483),
    .A1(_03555_));
 sg13g2_mux2_1 _19570_ (.A0(\top_ihp.oisc.regs[62][3] ),
    .A1(net135),
    .S(_03528_),
    .X(_02365_));
 sg13g2_mux2_1 _19571_ (.A0(\top_ihp.oisc.regs[62][4] ),
    .A1(_10599_),
    .S(_03528_),
    .X(_02366_));
 sg13g2_mux2_1 _19572_ (.A0(\top_ihp.oisc.regs[62][5] ),
    .A1(net267),
    .S(net688),
    .X(_02367_));
 sg13g2_mux2_1 _19573_ (.A0(\top_ihp.oisc.regs[62][6] ),
    .A1(net132),
    .S(net688),
    .X(_02368_));
 sg13g2_nand2_1 _19574_ (.Y(_03557_),
    .A(\top_ihp.oisc.regs[62][7] ),
    .B(net633));
 sg13g2_o21ai_1 _19575_ (.B1(_03557_),
    .Y(_02369_),
    .A1(net343),
    .A2(net632));
 sg13g2_nand2_1 _19576_ (.Y(_03558_),
    .A(\top_ihp.oisc.regs[62][8] ),
    .B(net633));
 sg13g2_o21ai_1 _19577_ (.B1(_03558_),
    .Y(_02370_),
    .A1(net205),
    .A2(net632));
 sg13g2_mux2_1 _19578_ (.A0(\top_ihp.oisc.regs[62][9] ),
    .A1(net131),
    .S(net688),
    .X(_02371_));
 sg13g2_nand2_1 _19579_ (.Y(_03559_),
    .A(_10787_),
    .B(_03150_));
 sg13g2_buf_2 _19580_ (.A(_03559_),
    .X(_03560_));
 sg13g2_buf_2 _19581_ (.A(_03560_),
    .X(_03561_));
 sg13g2_mux2_1 _19582_ (.A0(net119),
    .A1(\top_ihp.oisc.regs[63][0] ),
    .S(net481),
    .X(_02372_));
 sg13g2_mux2_1 _19583_ (.A0(_10704_),
    .A1(\top_ihp.oisc.regs[63][10] ),
    .S(net481),
    .X(_02373_));
 sg13g2_buf_1 _19584_ (.A(_03560_),
    .X(_03562_));
 sg13g2_buf_1 _19585_ (.A(_03560_),
    .X(_03563_));
 sg13g2_nand2_1 _19586_ (.Y(_03564_),
    .A(\top_ihp.oisc.regs[63][11] ),
    .B(net479));
 sg13g2_o21ai_1 _19587_ (.B1(_03564_),
    .Y(_02374_),
    .A1(net37),
    .A2(net480));
 sg13g2_nand2_1 _19588_ (.Y(_03565_),
    .A(\top_ihp.oisc.regs[63][12] ),
    .B(net479));
 sg13g2_o21ai_1 _19589_ (.B1(_03565_),
    .Y(_02375_),
    .A1(net141),
    .A2(net480));
 sg13g2_nand2_1 _19590_ (.Y(_03566_),
    .A(\top_ihp.oisc.regs[63][13] ),
    .B(_03563_));
 sg13g2_o21ai_1 _19591_ (.B1(_03566_),
    .Y(_02376_),
    .A1(net261),
    .A2(net480));
 sg13g2_nand2_1 _19592_ (.Y(_03567_),
    .A(\top_ihp.oisc.regs[63][14] ),
    .B(net479));
 sg13g2_o21ai_1 _19593_ (.B1(_03567_),
    .Y(_02377_),
    .A1(net260),
    .A2(net480));
 sg13g2_mux2_1 _19594_ (.A0(_10169_),
    .A1(\top_ihp.oisc.regs[63][15] ),
    .S(_03561_),
    .X(_02378_));
 sg13g2_nand2_1 _19595_ (.Y(_03568_),
    .A(\top_ihp.oisc.regs[63][16] ),
    .B(net479));
 sg13g2_o21ai_1 _19596_ (.B1(_03568_),
    .Y(_02379_),
    .A1(net276),
    .A2(_03562_));
 sg13g2_nand2_1 _19597_ (.Y(_03569_),
    .A(\top_ihp.oisc.regs[63][17] ),
    .B(_03563_));
 sg13g2_o21ai_1 _19598_ (.B1(_03569_),
    .Y(_02380_),
    .A1(_10800_),
    .A2(net480));
 sg13g2_nand2_1 _19599_ (.Y(_03570_),
    .A(\top_ihp.oisc.regs[63][18] ),
    .B(net479));
 sg13g2_o21ai_1 _19600_ (.B1(_03570_),
    .Y(_02381_),
    .A1(net259),
    .A2(_03562_));
 sg13g2_mux2_1 _19601_ (.A0(net254),
    .A1(\top_ihp.oisc.regs[63][19] ),
    .S(_03561_),
    .X(_02382_));
 sg13g2_nand2_1 _19602_ (.Y(_03571_),
    .A(\top_ihp.oisc.regs[63][1] ),
    .B(net479));
 sg13g2_o21ai_1 _19603_ (.B1(_03571_),
    .Y(_02383_),
    .A1(net274),
    .A2(net480));
 sg13g2_buf_1 _19604_ (.A(_03560_),
    .X(_03572_));
 sg13g2_nand2_1 _19605_ (.Y(_03573_),
    .A(\top_ihp.oisc.regs[63][20] ),
    .B(net478));
 sg13g2_o21ai_1 _19606_ (.B1(_03573_),
    .Y(_02384_),
    .A1(net121),
    .A2(net480));
 sg13g2_nand2_1 _19607_ (.Y(_03574_),
    .A(\top_ihp.oisc.regs[63][21] ),
    .B(net478));
 sg13g2_o21ai_1 _19608_ (.B1(_03574_),
    .Y(_02385_),
    .A1(net273),
    .A2(net480));
 sg13g2_buf_1 _19609_ (.A(_03560_),
    .X(_03575_));
 sg13g2_nand2_1 _19610_ (.Y(_03576_),
    .A(\top_ihp.oisc.regs[63][22] ),
    .B(net478));
 sg13g2_o21ai_1 _19611_ (.B1(_03576_),
    .Y(_02386_),
    .A1(net258),
    .A2(_03575_));
 sg13g2_nand2_1 _19612_ (.Y(_03577_),
    .A(\top_ihp.oisc.regs[63][23] ),
    .B(net478));
 sg13g2_o21ai_1 _19613_ (.B1(_03577_),
    .Y(_02387_),
    .A1(net257),
    .A2(net477));
 sg13g2_mux2_1 _19614_ (.A0(net400),
    .A1(\top_ihp.oisc.regs[63][24] ),
    .S(net481),
    .X(_02388_));
 sg13g2_nand2_1 _19615_ (.Y(_03578_),
    .A(\top_ihp.oisc.regs[63][25] ),
    .B(_03572_));
 sg13g2_o21ai_1 _19616_ (.B1(_03578_),
    .Y(_02389_),
    .A1(net262),
    .A2(net477));
 sg13g2_nand2_1 _19617_ (.Y(_03579_),
    .A(\top_ihp.oisc.regs[63][26] ),
    .B(net478));
 sg13g2_o21ai_1 _19618_ (.B1(_03579_),
    .Y(_02390_),
    .A1(_10810_),
    .A2(net477));
 sg13g2_mux2_1 _19619_ (.A0(net117),
    .A1(\top_ihp.oisc.regs[63][27] ),
    .S(net481),
    .X(_02391_));
 sg13g2_nand2_1 _19620_ (.Y(_03580_),
    .A(\top_ihp.oisc.regs[63][28] ),
    .B(net478));
 sg13g2_o21ai_1 _19621_ (.B1(_03580_),
    .Y(_02392_),
    .A1(_10459_),
    .A2(net477));
 sg13g2_nand2_1 _19622_ (.Y(_03581_),
    .A(\top_ihp.oisc.regs[63][29] ),
    .B(net478));
 sg13g2_o21ai_1 _19623_ (.B1(_03581_),
    .Y(_02393_),
    .A1(_10812_),
    .A2(net477));
 sg13g2_nand2_1 _19624_ (.Y(_03582_),
    .A(\top_ihp.oisc.regs[63][2] ),
    .B(_03572_));
 sg13g2_o21ai_1 _19625_ (.B1(_03582_),
    .Y(_02394_),
    .A1(net79),
    .A2(_03575_));
 sg13g2_nand2_1 _19626_ (.Y(_03583_),
    .A(\top_ihp.oisc.regs[63][30] ),
    .B(net478));
 sg13g2_o21ai_1 _19627_ (.B1(_03583_),
    .Y(_02395_),
    .A1(net35),
    .A2(net477));
 sg13g2_nand2_1 _19628_ (.Y(_03584_),
    .A(\top_ihp.oisc.regs[63][31] ),
    .B(_03560_));
 sg13g2_o21ai_1 _19629_ (.B1(_03584_),
    .Y(_02396_),
    .A1(net265),
    .A2(net477));
 sg13g2_mux2_1 _19630_ (.A0(_10739_),
    .A1(\top_ihp.oisc.regs[63][3] ),
    .S(net481),
    .X(_02397_));
 sg13g2_mux2_1 _19631_ (.A0(_10740_),
    .A1(\top_ihp.oisc.regs[63][4] ),
    .S(net481),
    .X(_02398_));
 sg13g2_mux2_1 _19632_ (.A0(net264),
    .A1(\top_ihp.oisc.regs[63][5] ),
    .S(net481),
    .X(_02399_));
 sg13g2_mux2_1 _19633_ (.A0(net126),
    .A1(\top_ihp.oisc.regs[63][6] ),
    .S(net479),
    .X(_02400_));
 sg13g2_nand2_1 _19634_ (.Y(_03585_),
    .A(\top_ihp.oisc.regs[63][7] ),
    .B(_03560_));
 sg13g2_o21ai_1 _19635_ (.B1(_03585_),
    .Y(_02401_),
    .A1(net396),
    .A2(net477));
 sg13g2_nand2_1 _19636_ (.Y(_03586_),
    .A(\top_ihp.oisc.regs[63][8] ),
    .B(_03560_));
 sg13g2_o21ai_1 _19637_ (.B1(_03586_),
    .Y(_02402_),
    .A1(net255),
    .A2(net481));
 sg13g2_mux2_1 _19638_ (.A0(net125),
    .A1(\top_ihp.oisc.regs[63][9] ),
    .S(net479),
    .X(_02403_));
 sg13g2_nor2_1 _19639_ (.A(_10707_),
    .B(_11080_),
    .Y(_03587_));
 sg13g2_buf_4 _19640_ (.X(_03588_),
    .A(_03587_));
 sg13g2_mux2_1 _19641_ (.A0(\top_ihp.oisc.regs[6][0] ),
    .A1(net143),
    .S(_03588_),
    .X(_02404_));
 sg13g2_mux2_1 _19642_ (.A0(\top_ihp.oisc.regs[6][10] ),
    .A1(net142),
    .S(_03588_),
    .X(_02405_));
 sg13g2_nand2_1 _19643_ (.Y(_03589_),
    .A(_10698_),
    .B(net729));
 sg13g2_buf_1 _19644_ (.A(_03589_),
    .X(_03590_));
 sg13g2_buf_1 _19645_ (.A(_03590_),
    .X(_03591_));
 sg13g2_buf_1 _19646_ (.A(net476),
    .X(_03592_));
 sg13g2_buf_1 _19647_ (.A(_03590_),
    .X(_03593_));
 sg13g2_nand2_1 _19648_ (.Y(_03594_),
    .A(\top_ihp.oisc.regs[6][11] ),
    .B(net475));
 sg13g2_o21ai_1 _19649_ (.B1(_03594_),
    .Y(_02406_),
    .A1(_03019_),
    .A2(net342));
 sg13g2_nand2_1 _19650_ (.Y(_03595_),
    .A(\top_ihp.oisc.regs[6][12] ),
    .B(net475));
 sg13g2_o21ai_1 _19651_ (.B1(_03595_),
    .Y(_02407_),
    .A1(net141),
    .A2(net342));
 sg13g2_nand2_1 _19652_ (.Y(_03596_),
    .A(\top_ihp.oisc.regs[6][13] ),
    .B(net475));
 sg13g2_o21ai_1 _19653_ (.B1(_03596_),
    .Y(_02408_),
    .A1(net261),
    .A2(_03592_));
 sg13g2_nand2_1 _19654_ (.Y(_03597_),
    .A(\top_ihp.oisc.regs[6][14] ),
    .B(net475));
 sg13g2_o21ai_1 _19655_ (.B1(_03597_),
    .Y(_02409_),
    .A1(net260),
    .A2(net342));
 sg13g2_nand2_1 _19656_ (.Y(_03598_),
    .A(\top_ihp.oisc.regs[6][15] ),
    .B(net475));
 sg13g2_o21ai_1 _19657_ (.B1(_03598_),
    .Y(_02410_),
    .A1(net399),
    .A2(_03592_));
 sg13g2_nand2_1 _19658_ (.Y(_03599_),
    .A(\top_ihp.oisc.regs[6][16] ),
    .B(net475));
 sg13g2_o21ai_1 _19659_ (.B1(_03599_),
    .Y(_02411_),
    .A1(net276),
    .A2(net342));
 sg13g2_buf_1 _19660_ (.A(_03590_),
    .X(_03600_));
 sg13g2_nand2_1 _19661_ (.Y(_03601_),
    .A(\top_ihp.oisc.regs[6][17] ),
    .B(net474));
 sg13g2_o21ai_1 _19662_ (.B1(_03601_),
    .Y(_02412_),
    .A1(net398),
    .A2(net342));
 sg13g2_nand2_1 _19663_ (.Y(_03602_),
    .A(\top_ihp.oisc.regs[6][18] ),
    .B(net474));
 sg13g2_o21ai_1 _19664_ (.B1(_03602_),
    .Y(_02413_),
    .A1(net259),
    .A2(net342));
 sg13g2_nand2_1 _19665_ (.Y(_03603_),
    .A(\top_ihp.oisc.regs[6][19] ),
    .B(net474));
 sg13g2_o21ai_1 _19666_ (.B1(_03603_),
    .Y(_02414_),
    .A1(_10273_),
    .A2(net342));
 sg13g2_buf_1 _19667_ (.A(net476),
    .X(_03604_));
 sg13g2_nand2_1 _19668_ (.Y(_03605_),
    .A(\top_ihp.oisc.regs[6][1] ),
    .B(net474));
 sg13g2_o21ai_1 _19669_ (.B1(_03605_),
    .Y(_02415_),
    .A1(net274),
    .A2(net341));
 sg13g2_nand2_1 _19670_ (.Y(_03606_),
    .A(\top_ihp.oisc.regs[6][20] ),
    .B(net474));
 sg13g2_o21ai_1 _19671_ (.B1(_03606_),
    .Y(_02416_),
    .A1(net121),
    .A2(_03604_));
 sg13g2_nand2_1 _19672_ (.Y(_03607_),
    .A(\top_ihp.oisc.regs[6][21] ),
    .B(net474));
 sg13g2_o21ai_1 _19673_ (.B1(_03607_),
    .Y(_02417_),
    .A1(net273),
    .A2(net341));
 sg13g2_nand2_1 _19674_ (.Y(_03608_),
    .A(\top_ihp.oisc.regs[6][22] ),
    .B(net474));
 sg13g2_o21ai_1 _19675_ (.B1(_03608_),
    .Y(_02418_),
    .A1(net258),
    .A2(net341));
 sg13g2_nand2_1 _19676_ (.Y(_03609_),
    .A(\top_ihp.oisc.regs[6][23] ),
    .B(_03600_));
 sg13g2_o21ai_1 _19677_ (.B1(_03609_),
    .Y(_02419_),
    .A1(net257),
    .A2(_03604_));
 sg13g2_mux2_1 _19678_ (.A0(\top_ihp.oisc.regs[6][24] ),
    .A1(net403),
    .S(_03588_),
    .X(_02420_));
 sg13g2_nand2_1 _19679_ (.Y(_03610_),
    .A(\top_ihp.oisc.regs[6][25] ),
    .B(net474));
 sg13g2_o21ai_1 _19680_ (.B1(_03610_),
    .Y(_02421_),
    .A1(_10428_),
    .A2(net341));
 sg13g2_nand2_1 _19681_ (.Y(_03611_),
    .A(\top_ihp.oisc.regs[6][26] ),
    .B(_03600_));
 sg13g2_o21ai_1 _19682_ (.B1(_03611_),
    .Y(_02422_),
    .A1(net397),
    .A2(net341));
 sg13g2_nand2_1 _19683_ (.Y(_03612_),
    .A(\top_ihp.oisc.regs[6][27] ),
    .B(_03591_));
 sg13g2_o21ai_1 _19684_ (.B1(_03612_),
    .Y(_02423_),
    .A1(_10449_),
    .A2(net341));
 sg13g2_nand2_1 _19685_ (.Y(_03613_),
    .A(\top_ihp.oisc.regs[6][28] ),
    .B(net476));
 sg13g2_o21ai_1 _19686_ (.B1(_03613_),
    .Y(_02424_),
    .A1(_10459_),
    .A2(net341));
 sg13g2_nand2_1 _19687_ (.Y(_03614_),
    .A(\top_ihp.oisc.regs[6][29] ),
    .B(net476));
 sg13g2_o21ai_1 _19688_ (.B1(_03614_),
    .Y(_02425_),
    .A1(net256),
    .A2(net341));
 sg13g2_nand2_1 _19689_ (.Y(_03615_),
    .A(\top_ihp.oisc.regs[6][2] ),
    .B(net476));
 sg13g2_o21ai_1 _19690_ (.B1(_03615_),
    .Y(_02426_),
    .A1(net122),
    .A2(net475));
 sg13g2_nand2_1 _19691_ (.Y(_03616_),
    .A(\top_ihp.oisc.regs[6][30] ),
    .B(net476));
 sg13g2_o21ai_1 _19692_ (.B1(_03616_),
    .Y(_02427_),
    .A1(net53),
    .A2(net475));
 sg13g2_inv_1 _19693_ (.Y(_03617_),
    .A(\top_ihp.oisc.regs[6][31] ));
 sg13g2_nor2_1 _19694_ (.A(_10535_),
    .B(net476),
    .Y(_03618_));
 sg13g2_a22oi_1 _19695_ (.Y(_02428_),
    .B1(_03618_),
    .B2(_10533_),
    .A2(net342),
    .A1(_03617_));
 sg13g2_mux2_1 _19696_ (.A0(\top_ihp.oisc.regs[6][3] ),
    .A1(net135),
    .S(_03588_),
    .X(_02429_));
 sg13g2_mux2_1 _19697_ (.A0(\top_ihp.oisc.regs[6][4] ),
    .A1(net134),
    .S(_03588_),
    .X(_02430_));
 sg13g2_mux2_1 _19698_ (.A0(\top_ihp.oisc.regs[6][5] ),
    .A1(net267),
    .S(_03588_),
    .X(_02431_));
 sg13g2_mux2_1 _19699_ (.A0(\top_ihp.oisc.regs[6][6] ),
    .A1(net132),
    .S(_03588_),
    .X(_02432_));
 sg13g2_nand2_1 _19700_ (.Y(_03619_),
    .A(\top_ihp.oisc.regs[6][7] ),
    .B(_03591_));
 sg13g2_o21ai_1 _19701_ (.B1(_03619_),
    .Y(_02433_),
    .A1(net396),
    .A2(_03593_));
 sg13g2_nand2_1 _19702_ (.Y(_03620_),
    .A(\top_ihp.oisc.regs[6][8] ),
    .B(net476));
 sg13g2_o21ai_1 _19703_ (.B1(_03620_),
    .Y(_02434_),
    .A1(net255),
    .A2(_03593_));
 sg13g2_mux2_1 _19704_ (.A0(\top_ihp.oisc.regs[6][9] ),
    .A1(net131),
    .S(_03588_),
    .X(_02435_));
 sg13g2_and2_1 _19705_ (.A(_10749_),
    .B(net729),
    .X(_03621_));
 sg13g2_buf_1 _19706_ (.A(_03621_),
    .X(_03622_));
 sg13g2_buf_1 _19707_ (.A(net631),
    .X(_03623_));
 sg13g2_mux2_1 _19708_ (.A0(\top_ihp.oisc.regs[7][0] ),
    .A1(_09888_),
    .S(net473),
    .X(_02436_));
 sg13g2_mux2_1 _19709_ (.A0(\top_ihp.oisc.regs[7][10] ),
    .A1(_10009_),
    .S(net473),
    .X(_02437_));
 sg13g2_nor2_1 _19710_ (.A(\top_ihp.oisc.regs[7][11] ),
    .B(net631),
    .Y(_03624_));
 sg13g2_a21oi_1 _19711_ (.A1(_10051_),
    .A2(_03623_),
    .Y(_02438_),
    .B1(_03624_));
 sg13g2_nor2_1 _19712_ (.A(\top_ihp.oisc.regs[7][12] ),
    .B(net631),
    .Y(_03625_));
 sg13g2_a21oi_1 _19713_ (.A1(_10090_),
    .A2(net473),
    .Y(_02439_),
    .B1(_03625_));
 sg13g2_nand2_1 _19714_ (.Y(_03626_),
    .A(_10749_),
    .B(_03079_));
 sg13g2_buf_1 _19715_ (.A(_03626_),
    .X(_03627_));
 sg13g2_buf_1 _19716_ (.A(net630),
    .X(_03628_));
 sg13g2_buf_1 _19717_ (.A(net630),
    .X(_03629_));
 sg13g2_nand2_1 _19718_ (.Y(_03630_),
    .A(\top_ihp.oisc.regs[7][13] ),
    .B(net471));
 sg13g2_o21ai_1 _19719_ (.B1(_03630_),
    .Y(_02440_),
    .A1(net261),
    .A2(net472));
 sg13g2_nand2_1 _19720_ (.Y(_03631_),
    .A(\top_ihp.oisc.regs[7][14] ),
    .B(net471));
 sg13g2_o21ai_1 _19721_ (.B1(_03631_),
    .Y(_02441_),
    .A1(net260),
    .A2(net472));
 sg13g2_buf_1 _19722_ (.A(_03627_),
    .X(_03632_));
 sg13g2_nand2_1 _19723_ (.Y(_03633_),
    .A(\top_ihp.oisc.regs[7][15] ),
    .B(_03632_));
 sg13g2_o21ai_1 _19724_ (.B1(_03633_),
    .Y(_02442_),
    .A1(_10798_),
    .A2(net472));
 sg13g2_nand2_1 _19725_ (.Y(_03634_),
    .A(\top_ihp.oisc.regs[7][16] ),
    .B(net470));
 sg13g2_o21ai_1 _19726_ (.B1(_03634_),
    .Y(_02443_),
    .A1(net276),
    .A2(net472));
 sg13g2_nand2_1 _19727_ (.Y(_03635_),
    .A(\top_ihp.oisc.regs[7][17] ),
    .B(net470));
 sg13g2_o21ai_1 _19728_ (.B1(_03635_),
    .Y(_02444_),
    .A1(net398),
    .A2(net472));
 sg13g2_nand2_1 _19729_ (.Y(_03636_),
    .A(\top_ihp.oisc.regs[7][18] ),
    .B(net470));
 sg13g2_o21ai_1 _19730_ (.B1(_03636_),
    .Y(_02445_),
    .A1(net259),
    .A2(net472));
 sg13g2_mux2_1 _19731_ (.A0(\top_ihp.oisc.regs[7][19] ),
    .A1(_10271_),
    .S(net473),
    .X(_02446_));
 sg13g2_nor2_1 _19732_ (.A(\top_ihp.oisc.regs[7][1] ),
    .B(_03622_),
    .Y(_03637_));
 sg13g2_a21oi_1 _19733_ (.A1(_10319_),
    .A2(net473),
    .Y(_02447_),
    .B1(_03637_));
 sg13g2_nand2_1 _19734_ (.Y(_03638_),
    .A(\top_ihp.oisc.regs[7][20] ),
    .B(net470));
 sg13g2_o21ai_1 _19735_ (.B1(_03638_),
    .Y(_02448_),
    .A1(net121),
    .A2(net472));
 sg13g2_nand2_1 _19736_ (.Y(_03639_),
    .A(\top_ihp.oisc.regs[7][21] ),
    .B(net470));
 sg13g2_o21ai_1 _19737_ (.B1(_03639_),
    .Y(_02449_),
    .A1(net273),
    .A2(net472));
 sg13g2_nand2_1 _19738_ (.Y(_03640_),
    .A(\top_ihp.oisc.regs[7][22] ),
    .B(_03632_));
 sg13g2_o21ai_1 _19739_ (.B1(_03640_),
    .Y(_02450_),
    .A1(net258),
    .A2(_03628_));
 sg13g2_nand2_1 _19740_ (.Y(_03641_),
    .A(\top_ihp.oisc.regs[7][23] ),
    .B(net470));
 sg13g2_o21ai_1 _19741_ (.B1(_03641_),
    .Y(_02451_),
    .A1(net257),
    .A2(_03628_));
 sg13g2_mux2_1 _19742_ (.A0(\top_ihp.oisc.regs[7][24] ),
    .A1(_10415_),
    .S(net473),
    .X(_02452_));
 sg13g2_nand2_1 _19743_ (.Y(_03642_),
    .A(\top_ihp.oisc.regs[7][25] ),
    .B(net470));
 sg13g2_o21ai_1 _19744_ (.B1(_03642_),
    .Y(_02453_),
    .A1(_10772_),
    .A2(net471));
 sg13g2_nand2_1 _19745_ (.Y(_03643_),
    .A(\top_ihp.oisc.regs[7][26] ),
    .B(net470));
 sg13g2_o21ai_1 _19746_ (.B1(_03643_),
    .Y(_02454_),
    .A1(net397),
    .A2(net471));
 sg13g2_mux2_1 _19747_ (.A0(\top_ihp.oisc.regs[7][27] ),
    .A1(_10447_),
    .S(_03623_),
    .X(_02455_));
 sg13g2_nor2_1 _19748_ (.A(\top_ihp.oisc.regs[7][28] ),
    .B(net631),
    .Y(_03644_));
 sg13g2_a21oi_1 _19749_ (.A1(_10456_),
    .A2(net473),
    .Y(_02456_),
    .B1(_03644_));
 sg13g2_nand2_1 _19750_ (.Y(_03645_),
    .A(\top_ihp.oisc.regs[7][29] ),
    .B(net630));
 sg13g2_o21ai_1 _19751_ (.B1(_03645_),
    .Y(_02457_),
    .A1(net256),
    .A2(net471));
 sg13g2_nand2_1 _19752_ (.Y(_03646_),
    .A(\top_ihp.oisc.regs[7][2] ),
    .B(net630));
 sg13g2_o21ai_1 _19753_ (.B1(_03646_),
    .Y(_02458_),
    .A1(net122),
    .A2(net471));
 sg13g2_nand2_1 _19754_ (.Y(_03647_),
    .A(\top_ihp.oisc.regs[7][30] ),
    .B(net630));
 sg13g2_o21ai_1 _19755_ (.B1(_03647_),
    .Y(_02459_),
    .A1(net53),
    .A2(net471));
 sg13g2_nand2_1 _19756_ (.Y(_03648_),
    .A(\top_ihp.oisc.regs[7][31] ),
    .B(net630));
 sg13g2_o21ai_1 _19757_ (.B1(_03648_),
    .Y(_02460_),
    .A1(net265),
    .A2(net471));
 sg13g2_mux2_1 _19758_ (.A0(\top_ihp.oisc.regs[7][3] ),
    .A1(_10567_),
    .S(net473),
    .X(_02461_));
 sg13g2_mux2_1 _19759_ (.A0(\top_ihp.oisc.regs[7][4] ),
    .A1(_10599_),
    .S(net631),
    .X(_02462_));
 sg13g2_mux2_1 _19760_ (.A0(\top_ihp.oisc.regs[7][5] ),
    .A1(_10625_),
    .S(net631),
    .X(_02463_));
 sg13g2_mux2_1 _19761_ (.A0(\top_ihp.oisc.regs[7][6] ),
    .A1(_10648_),
    .S(net631),
    .X(_02464_));
 sg13g2_nand2_1 _19762_ (.Y(_03649_),
    .A(\top_ihp.oisc.regs[7][7] ),
    .B(net630));
 sg13g2_o21ai_1 _19763_ (.B1(_03649_),
    .Y(_02465_),
    .A1(net396),
    .A2(_03629_));
 sg13g2_nand2_1 _19764_ (.Y(_03650_),
    .A(\top_ihp.oisc.regs[7][8] ),
    .B(net630));
 sg13g2_o21ai_1 _19765_ (.B1(_03650_),
    .Y(_02466_),
    .A1(net255),
    .A2(_03629_));
 sg13g2_mux2_1 _19766_ (.A0(\top_ihp.oisc.regs[7][9] ),
    .A1(_10687_),
    .S(net631),
    .X(_02467_));
 sg13g2_nand2_1 _19767_ (.Y(_03651_),
    .A(_09941_),
    .B(_10694_));
 sg13g2_buf_1 _19768_ (.A(_03651_),
    .X(_03652_));
 sg13g2_buf_1 _19769_ (.A(net629),
    .X(_03653_));
 sg13g2_mux2_1 _19770_ (.A0(_10845_),
    .A1(\top_ihp.oisc.regs[8][0] ),
    .S(net469),
    .X(_02468_));
 sg13g2_mux2_1 _19771_ (.A0(_10704_),
    .A1(\top_ihp.oisc.regs[8][10] ),
    .S(net469),
    .X(_02469_));
 sg13g2_buf_2 _19772_ (.A(net629),
    .X(_03654_));
 sg13g2_buf_1 _19773_ (.A(_03651_),
    .X(_03655_));
 sg13g2_nand2_1 _19774_ (.Y(_03656_),
    .A(\top_ihp.oisc.regs[8][11] ),
    .B(net628));
 sg13g2_o21ai_1 _19775_ (.B1(_03656_),
    .Y(_02470_),
    .A1(_03019_),
    .A2(net468));
 sg13g2_nand2_1 _19776_ (.Y(_03657_),
    .A(\top_ihp.oisc.regs[8][12] ),
    .B(net628));
 sg13g2_o21ai_1 _19777_ (.B1(_03657_),
    .Y(_02471_),
    .A1(net141),
    .A2(net468));
 sg13g2_nand2_1 _19778_ (.Y(_03658_),
    .A(\top_ihp.oisc.regs[8][13] ),
    .B(net628));
 sg13g2_o21ai_1 _19779_ (.B1(_03658_),
    .Y(_02472_),
    .A1(_10796_),
    .A2(net468));
 sg13g2_nand2_1 _19780_ (.Y(_03659_),
    .A(\top_ihp.oisc.regs[8][14] ),
    .B(net628));
 sg13g2_o21ai_1 _19781_ (.B1(_03659_),
    .Y(_02473_),
    .A1(_10797_),
    .A2(_03654_));
 sg13g2_nand2_1 _19782_ (.Y(_03660_),
    .A(\top_ihp.oisc.regs[8][15] ),
    .B(net628));
 sg13g2_o21ai_1 _19783_ (.B1(_03660_),
    .Y(_02474_),
    .A1(net399),
    .A2(net468));
 sg13g2_nand2_1 _19784_ (.Y(_03661_),
    .A(\top_ihp.oisc.regs[8][16] ),
    .B(_03655_));
 sg13g2_o21ai_1 _19785_ (.B1(_03661_),
    .Y(_02475_),
    .A1(net276),
    .A2(net468));
 sg13g2_nand2_1 _19786_ (.Y(_03662_),
    .A(\top_ihp.oisc.regs[8][17] ),
    .B(net628));
 sg13g2_o21ai_1 _19787_ (.B1(_03662_),
    .Y(_02476_),
    .A1(net398),
    .A2(_03654_));
 sg13g2_nand2_1 _19788_ (.Y(_03663_),
    .A(\top_ihp.oisc.regs[8][18] ),
    .B(_03655_));
 sg13g2_o21ai_1 _19789_ (.B1(_03663_),
    .Y(_02477_),
    .A1(_10801_),
    .A2(net468));
 sg13g2_buf_1 _19790_ (.A(net629),
    .X(_03664_));
 sg13g2_nand2_1 _19791_ (.Y(_03665_),
    .A(\top_ihp.oisc.regs[8][19] ),
    .B(net467));
 sg13g2_o21ai_1 _19792_ (.B1(_03665_),
    .Y(_02478_),
    .A1(_10273_),
    .A2(net468));
 sg13g2_buf_1 _19793_ (.A(net629),
    .X(_03666_));
 sg13g2_nand2_1 _19794_ (.Y(_03667_),
    .A(\top_ihp.oisc.regs[8][1] ),
    .B(net467));
 sg13g2_o21ai_1 _19795_ (.B1(_03667_),
    .Y(_02479_),
    .A1(net274),
    .A2(net466));
 sg13g2_nand2_1 _19796_ (.Y(_03668_),
    .A(\top_ihp.oisc.regs[8][20] ),
    .B(net467));
 sg13g2_o21ai_1 _19797_ (.B1(_03668_),
    .Y(_02480_),
    .A1(_10804_),
    .A2(net466));
 sg13g2_nand2_1 _19798_ (.Y(_03669_),
    .A(\top_ihp.oisc.regs[8][21] ),
    .B(net467));
 sg13g2_o21ai_1 _19799_ (.B1(_03669_),
    .Y(_02481_),
    .A1(net273),
    .A2(net466));
 sg13g2_nand2_1 _19800_ (.Y(_03670_),
    .A(\top_ihp.oisc.regs[8][22] ),
    .B(net467));
 sg13g2_o21ai_1 _19801_ (.B1(_03670_),
    .Y(_02482_),
    .A1(net258),
    .A2(net466));
 sg13g2_nand2_1 _19802_ (.Y(_03671_),
    .A(\top_ihp.oisc.regs[8][23] ),
    .B(_03664_));
 sg13g2_o21ai_1 _19803_ (.B1(_03671_),
    .Y(_02483_),
    .A1(net257),
    .A2(net466));
 sg13g2_mux2_1 _19804_ (.A0(_10726_),
    .A1(\top_ihp.oisc.regs[8][24] ),
    .S(net469),
    .X(_02484_));
 sg13g2_nand2_1 _19805_ (.Y(_03672_),
    .A(\top_ihp.oisc.regs[8][25] ),
    .B(net467));
 sg13g2_o21ai_1 _19806_ (.B1(_03672_),
    .Y(_02485_),
    .A1(_10428_),
    .A2(net466));
 sg13g2_nand2_1 _19807_ (.Y(_03673_),
    .A(\top_ihp.oisc.regs[8][26] ),
    .B(net467));
 sg13g2_o21ai_1 _19808_ (.B1(_03673_),
    .Y(_02486_),
    .A1(_10810_),
    .A2(net466));
 sg13g2_nand2_1 _19809_ (.Y(_03674_),
    .A(\top_ihp.oisc.regs[8][27] ),
    .B(net467));
 sg13g2_o21ai_1 _19810_ (.B1(_03674_),
    .Y(_02487_),
    .A1(_10449_),
    .A2(net466));
 sg13g2_nand2_1 _19811_ (.Y(_03675_),
    .A(\top_ihp.oisc.regs[8][28] ),
    .B(_03664_));
 sg13g2_o21ai_1 _19812_ (.B1(_03675_),
    .Y(_02488_),
    .A1(_10459_),
    .A2(_03666_));
 sg13g2_nand2_1 _19813_ (.Y(_03676_),
    .A(\top_ihp.oisc.regs[8][29] ),
    .B(net629));
 sg13g2_o21ai_1 _19814_ (.B1(_03676_),
    .Y(_02489_),
    .A1(_10812_),
    .A2(_03666_));
 sg13g2_nand2_1 _19815_ (.Y(_03677_),
    .A(\top_ihp.oisc.regs[8][2] ),
    .B(net629));
 sg13g2_o21ai_1 _19816_ (.B1(_03677_),
    .Y(_02490_),
    .A1(net122),
    .A2(net469));
 sg13g2_nand2_1 _19817_ (.Y(_03678_),
    .A(\top_ihp.oisc.regs[8][30] ),
    .B(net629));
 sg13g2_o21ai_1 _19818_ (.B1(_03678_),
    .Y(_02491_),
    .A1(net53),
    .A2(net469));
 sg13g2_inv_1 _19819_ (.Y(_03679_),
    .A(\top_ihp.oisc.regs[8][31] ));
 sg13g2_nor2_1 _19820_ (.A(_10535_),
    .B(net629),
    .Y(_03680_));
 sg13g2_a22oi_1 _19821_ (.Y(_02492_),
    .B1(_03680_),
    .B2(_10533_),
    .A2(net468),
    .A1(_03679_));
 sg13g2_mux2_1 _19822_ (.A0(net128),
    .A1(\top_ihp.oisc.regs[8][3] ),
    .S(net469),
    .X(_02493_));
 sg13g2_mux2_1 _19823_ (.A0(net127),
    .A1(\top_ihp.oisc.regs[8][4] ),
    .S(net469),
    .X(_02494_));
 sg13g2_mux2_1 _19824_ (.A0(_10741_),
    .A1(\top_ihp.oisc.regs[8][5] ),
    .S(net469),
    .X(_02495_));
 sg13g2_mux2_1 _19825_ (.A0(_10742_),
    .A1(\top_ihp.oisc.regs[8][6] ),
    .S(net628),
    .X(_02496_));
 sg13g2_nand2_1 _19826_ (.Y(_03681_),
    .A(\top_ihp.oisc.regs[8][7] ),
    .B(_03652_));
 sg13g2_o21ai_1 _19827_ (.B1(_03681_),
    .Y(_02497_),
    .A1(net396),
    .A2(_03653_));
 sg13g2_nand2_1 _19828_ (.Y(_03682_),
    .A(\top_ihp.oisc.regs[8][8] ),
    .B(_03652_));
 sg13g2_o21ai_1 _19829_ (.B1(_03682_),
    .Y(_02498_),
    .A1(net255),
    .A2(_03653_));
 sg13g2_mux2_1 _19830_ (.A0(_10745_),
    .A1(\top_ihp.oisc.regs[8][9] ),
    .S(net628),
    .X(_02499_));
 sg13g2_nor2_1 _19831_ (.A(_10706_),
    .B(_10913_),
    .Y(_03683_));
 sg13g2_buf_1 _19832_ (.A(_03683_),
    .X(_03684_));
 sg13g2_buf_1 _19833_ (.A(_03684_),
    .X(_03685_));
 sg13g2_mux2_1 _19834_ (.A0(\top_ihp.oisc.regs[9][0] ),
    .A1(_09888_),
    .S(net465),
    .X(_02500_));
 sg13g2_mux2_1 _19835_ (.A0(\top_ihp.oisc.regs[9][10] ),
    .A1(_10009_),
    .S(net465),
    .X(_02501_));
 sg13g2_nor2_1 _19836_ (.A(\top_ihp.oisc.regs[9][11] ),
    .B(net627),
    .Y(_03686_));
 sg13g2_a21oi_1 _19837_ (.A1(_10051_),
    .A2(_03685_),
    .Y(_02502_),
    .B1(_03686_));
 sg13g2_nor2_1 _19838_ (.A(\top_ihp.oisc.regs[9][12] ),
    .B(net627),
    .Y(_03687_));
 sg13g2_a21oi_1 _19839_ (.A1(_10090_),
    .A2(net465),
    .Y(_02503_),
    .B1(_03687_));
 sg13g2_nand2_1 _19840_ (.Y(_03688_),
    .A(_10694_),
    .B(_10824_));
 sg13g2_buf_1 _19841_ (.A(_03688_),
    .X(_03689_));
 sg13g2_buf_1 _19842_ (.A(net626),
    .X(_03690_));
 sg13g2_buf_1 _19843_ (.A(net626),
    .X(_03691_));
 sg13g2_nand2_1 _19844_ (.Y(_03692_),
    .A(\top_ihp.oisc.regs[9][13] ),
    .B(net463));
 sg13g2_o21ai_1 _19845_ (.B1(_03692_),
    .Y(_02504_),
    .A1(_10796_),
    .A2(net464));
 sg13g2_nand2_1 _19846_ (.Y(_03693_),
    .A(\top_ihp.oisc.regs[9][14] ),
    .B(net463));
 sg13g2_o21ai_1 _19847_ (.B1(_03693_),
    .Y(_02505_),
    .A1(_10797_),
    .A2(net464));
 sg13g2_buf_1 _19848_ (.A(_03689_),
    .X(_03694_));
 sg13g2_nand2_1 _19849_ (.Y(_03695_),
    .A(\top_ihp.oisc.regs[9][15] ),
    .B(net462));
 sg13g2_o21ai_1 _19850_ (.B1(_03695_),
    .Y(_02506_),
    .A1(_10798_),
    .A2(net464));
 sg13g2_nand2_1 _19851_ (.Y(_03696_),
    .A(\top_ihp.oisc.regs[9][16] ),
    .B(net462));
 sg13g2_o21ai_1 _19852_ (.B1(_03696_),
    .Y(_02507_),
    .A1(_10205_),
    .A2(net464));
 sg13g2_nand2_1 _19853_ (.Y(_03697_),
    .A(\top_ihp.oisc.regs[9][17] ),
    .B(net462));
 sg13g2_o21ai_1 _19854_ (.B1(_03697_),
    .Y(_02508_),
    .A1(net398),
    .A2(net464));
 sg13g2_nand2_1 _19855_ (.Y(_03698_),
    .A(\top_ihp.oisc.regs[9][18] ),
    .B(net462));
 sg13g2_o21ai_1 _19856_ (.B1(_03698_),
    .Y(_02509_),
    .A1(_10801_),
    .A2(net464));
 sg13g2_mux2_1 _19857_ (.A0(\top_ihp.oisc.regs[9][19] ),
    .A1(_10271_),
    .S(net465),
    .X(_02510_));
 sg13g2_nor2_1 _19858_ (.A(\top_ihp.oisc.regs[9][1] ),
    .B(net627),
    .Y(_03699_));
 sg13g2_a21oi_1 _19859_ (.A1(_10319_),
    .A2(net465),
    .Y(_02511_),
    .B1(_03699_));
 sg13g2_nand2_1 _19860_ (.Y(_03700_),
    .A(\top_ihp.oisc.regs[9][20] ),
    .B(net462));
 sg13g2_o21ai_1 _19861_ (.B1(_03700_),
    .Y(_02512_),
    .A1(net121),
    .A2(net464));
 sg13g2_nand2_1 _19862_ (.Y(_03701_),
    .A(\top_ihp.oisc.regs[9][21] ),
    .B(net462));
 sg13g2_o21ai_1 _19863_ (.B1(_03701_),
    .Y(_02513_),
    .A1(net273),
    .A2(net464));
 sg13g2_nand2_1 _19864_ (.Y(_03702_),
    .A(\top_ihp.oisc.regs[9][22] ),
    .B(_03694_));
 sg13g2_o21ai_1 _19865_ (.B1(_03702_),
    .Y(_02514_),
    .A1(net258),
    .A2(_03690_));
 sg13g2_nand2_1 _19866_ (.Y(_03703_),
    .A(\top_ihp.oisc.regs[9][23] ),
    .B(net462));
 sg13g2_o21ai_1 _19867_ (.B1(_03703_),
    .Y(_02515_),
    .A1(net257),
    .A2(_03690_));
 sg13g2_mux2_1 _19868_ (.A0(\top_ihp.oisc.regs[9][24] ),
    .A1(_10415_),
    .S(net465),
    .X(_02516_));
 sg13g2_nand2_1 _19869_ (.Y(_03704_),
    .A(\top_ihp.oisc.regs[9][25] ),
    .B(net462));
 sg13g2_o21ai_1 _19870_ (.B1(_03704_),
    .Y(_02517_),
    .A1(net262),
    .A2(net463));
 sg13g2_nand2_1 _19871_ (.Y(_03705_),
    .A(\top_ihp.oisc.regs[9][26] ),
    .B(_03694_));
 sg13g2_o21ai_1 _19872_ (.B1(_03705_),
    .Y(_02518_),
    .A1(net397),
    .A2(net463));
 sg13g2_mux2_1 _19873_ (.A0(\top_ihp.oisc.regs[9][27] ),
    .A1(_10447_),
    .S(net465),
    .X(_02519_));
 sg13g2_nor2_1 _19874_ (.A(\top_ihp.oisc.regs[9][28] ),
    .B(net627),
    .Y(_03706_));
 sg13g2_a21oi_1 _19875_ (.A1(_10456_),
    .A2(_03685_),
    .Y(_02520_),
    .B1(_03706_));
 sg13g2_nand2_1 _19876_ (.Y(_03707_),
    .A(\top_ihp.oisc.regs[9][29] ),
    .B(net626));
 sg13g2_o21ai_1 _19877_ (.B1(_03707_),
    .Y(_02521_),
    .A1(net256),
    .A2(net463));
 sg13g2_nand2_1 _19878_ (.Y(_03708_),
    .A(\top_ihp.oisc.regs[9][2] ),
    .B(net626));
 sg13g2_o21ai_1 _19879_ (.B1(_03708_),
    .Y(_02522_),
    .A1(_10779_),
    .A2(net463));
 sg13g2_nand2_1 _19880_ (.Y(_03709_),
    .A(\top_ihp.oisc.regs[9][30] ),
    .B(net626));
 sg13g2_o21ai_1 _19881_ (.B1(_03709_),
    .Y(_02523_),
    .A1(_10813_),
    .A2(net463));
 sg13g2_nand2_1 _19882_ (.Y(_03710_),
    .A(\top_ihp.oisc.regs[9][31] ),
    .B(net626));
 sg13g2_o21ai_1 _19883_ (.B1(_03710_),
    .Y(_02524_),
    .A1(net265),
    .A2(net463));
 sg13g2_mux2_1 _19884_ (.A0(\top_ihp.oisc.regs[9][3] ),
    .A1(_10567_),
    .S(net465),
    .X(_02525_));
 sg13g2_mux2_1 _19885_ (.A0(\top_ihp.oisc.regs[9][4] ),
    .A1(net134),
    .S(net627),
    .X(_02526_));
 sg13g2_mux2_1 _19886_ (.A0(\top_ihp.oisc.regs[9][5] ),
    .A1(net267),
    .S(net627),
    .X(_02527_));
 sg13g2_mux2_1 _19887_ (.A0(\top_ihp.oisc.regs[9][6] ),
    .A1(_10648_),
    .S(net627),
    .X(_02528_));
 sg13g2_nand2_1 _19888_ (.Y(_03711_),
    .A(\top_ihp.oisc.regs[9][7] ),
    .B(net626));
 sg13g2_o21ai_1 _19889_ (.B1(_03711_),
    .Y(_02529_),
    .A1(_10818_),
    .A2(_03691_));
 sg13g2_nand2_1 _19890_ (.Y(_03712_),
    .A(\top_ihp.oisc.regs[9][8] ),
    .B(net626));
 sg13g2_o21ai_1 _19891_ (.B1(_03712_),
    .Y(_02530_),
    .A1(_10819_),
    .A2(_03691_));
 sg13g2_mux2_1 _19892_ (.A0(\top_ihp.oisc.regs[9][9] ),
    .A1(net131),
    .S(net627),
    .X(_02531_));
 sg13g2_nor2_1 _19893_ (.A(_08615_),
    .B(net793),
    .Y(_03713_));
 sg13g2_buf_2 _19894_ (.A(_03713_),
    .X(_03714_));
 sg13g2_buf_2 _19895_ (.A(net748),
    .X(_03715_));
 sg13g2_buf_1 _19896_ (.A(net739),
    .X(_03716_));
 sg13g2_buf_1 _19897_ (.A(net728),
    .X(_03717_));
 sg13g2_nor3_1 _19898_ (.A(net1032),
    .B(_09001_),
    .C(net719),
    .Y(_03718_));
 sg13g2_and4_1 _19899_ (.A(_08944_),
    .B(_08957_),
    .C(_08975_),
    .D(_08976_),
    .X(_03719_));
 sg13g2_buf_2 _19900_ (.A(_03719_),
    .X(_03720_));
 sg13g2_a21oi_1 _19901_ (.A1(_08201_),
    .A2(_03720_),
    .Y(_03721_),
    .B1(_08415_));
 sg13g2_nor2_1 _19902_ (.A(net890),
    .B(_03721_),
    .Y(_03722_));
 sg13g2_o21ai_1 _19903_ (.B1(_03720_),
    .Y(_03723_),
    .A1(net934),
    .A2(_09001_));
 sg13g2_buf_1 _19904_ (.A(_03723_),
    .X(_03724_));
 sg13g2_o21ai_1 _19905_ (.B1(_09007_),
    .Y(_03725_),
    .A1(net1032),
    .A2(_03724_));
 sg13g2_a22oi_1 _19906_ (.Y(_03726_),
    .B1(_03725_),
    .B2(_13699_),
    .A2(_03722_),
    .A1(net959));
 sg13g2_nand2b_1 _19907_ (.Y(_02532_),
    .B(_03726_),
    .A_N(_03718_));
 sg13g2_buf_1 _19908_ (.A(net934),
    .X(_03727_));
 sg13g2_buf_1 _19909_ (.A(net1000),
    .X(_03728_));
 sg13g2_buf_1 _19910_ (.A(_00078_),
    .X(_03729_));
 sg13g2_nand3_1 _19911_ (.B(_03729_),
    .C(_03724_),
    .A(net948),
    .Y(_03730_));
 sg13g2_nor2_1 _19912_ (.A(net890),
    .B(_03730_),
    .Y(_03731_));
 sg13g2_a21oi_1 _19913_ (.A1(_03727_),
    .A2(net890),
    .Y(_03732_),
    .B1(_03731_));
 sg13g2_buf_1 _19914_ (.A(net728),
    .X(_03733_));
 sg13g2_nor2_1 _19915_ (.A(net959),
    .B(net718),
    .Y(_03734_));
 sg13g2_a22oi_1 _19916_ (.Y(_02533_),
    .B1(_03734_),
    .B2(_03730_),
    .A2(_03732_),
    .A1(net959));
 sg13g2_nor2_1 _19917_ (.A(_08615_),
    .B(_03720_),
    .Y(_03735_));
 sg13g2_buf_2 _19918_ (.A(_03735_),
    .X(_03736_));
 sg13g2_buf_1 _19919_ (.A(_03736_),
    .X(_03737_));
 sg13g2_nand2_1 _19920_ (.Y(_03738_),
    .A(_03729_),
    .B(net747));
 sg13g2_nand2_1 _19921_ (.Y(_03739_),
    .A(net1037),
    .B(_03725_));
 sg13g2_o21ai_1 _19922_ (.B1(_03739_),
    .Y(_02534_),
    .A1(_03725_),
    .A2(_03738_));
 sg13g2_nand3_1 _19923_ (.B(net960),
    .C(net890),
    .A(net959),
    .Y(_03740_));
 sg13g2_nand2_1 _19924_ (.Y(_03741_),
    .A(_09671_),
    .B(_09004_));
 sg13g2_nand3_1 _19925_ (.B(_03729_),
    .C(_03724_),
    .A(net1037),
    .Y(_03742_));
 sg13g2_a21o_1 _19926_ (.A2(_03742_),
    .A1(_03741_),
    .B1(net1032),
    .X(_03743_));
 sg13g2_nand4_1 _19927_ (.B(_03729_),
    .C(net892),
    .A(net1037),
    .Y(_03744_),
    .D(_03724_));
 sg13g2_nand3_1 _19928_ (.B(_03743_),
    .C(_03744_),
    .A(_03740_),
    .Y(_02535_));
 sg13g2_nand2_1 _19929_ (.Y(_03745_),
    .A(net958),
    .B(_09004_));
 sg13g2_nand3_1 _19930_ (.B(_03729_),
    .C(_03724_),
    .A(net1008),
    .Y(_03746_));
 sg13g2_a21oi_1 _19931_ (.A1(_03745_),
    .A2(_03746_),
    .Y(_03747_),
    .B1(net959));
 sg13g2_nand4_1 _19932_ (.B(_03729_),
    .C(net892),
    .A(_09671_),
    .Y(_03748_),
    .D(_03724_));
 sg13g2_o21ai_1 _19933_ (.B1(_03748_),
    .Y(_03749_),
    .A1(net949),
    .A2(_09007_));
 sg13g2_or2_1 _19934_ (.X(_02536_),
    .B(_03749_),
    .A(_03747_));
 sg13g2_nand2_1 _19935_ (.Y(_03750_),
    .A(_09001_),
    .B(_03720_));
 sg13g2_nor2_1 _19936_ (.A(_09002_),
    .B(net892),
    .Y(_03751_));
 sg13g2_o21ai_1 _19937_ (.B1(_09779_),
    .Y(_03752_),
    .A1(_03722_),
    .A2(_03751_));
 sg13g2_o21ai_1 _19938_ (.B1(_03752_),
    .Y(_02537_),
    .A1(_09779_),
    .A2(_03750_));
 sg13g2_buf_1 _19939_ (.A(\top_ihp.oisc.wb_dat_o[0] ),
    .X(_03753_));
 sg13g2_nand2_1 _19940_ (.Y(_03754_),
    .A(_08201_),
    .B(net1008));
 sg13g2_buf_1 _19941_ (.A(_03754_),
    .X(_03755_));
 sg13g2_buf_1 _19942_ (.A(net900),
    .X(_03756_));
 sg13g2_mux2_1 _19943_ (.A0(_10845_),
    .A1(net1034),
    .S(net870),
    .X(_02538_));
 sg13g2_buf_2 _19944_ (.A(\top_ihp.oisc.wb_dat_o[10] ),
    .X(_03757_));
 sg13g2_mux2_1 _19945_ (.A0(net130),
    .A1(_03757_),
    .S(net870),
    .X(_02539_));
 sg13g2_buf_2 _19946_ (.A(\top_ihp.oisc.wb_dat_o[11] ),
    .X(_03758_));
 sg13g2_mux2_1 _19947_ (.A0(net1030),
    .A1(_03758_),
    .S(net870),
    .X(_02540_));
 sg13g2_buf_1 _19948_ (.A(net900),
    .X(_03759_));
 sg13g2_buf_2 _19949_ (.A(\top_ihp.oisc.wb_dat_o[12] ),
    .X(_03760_));
 sg13g2_buf_1 _19950_ (.A(net900),
    .X(_03761_));
 sg13g2_nand2_1 _19951_ (.Y(_03762_),
    .A(_03760_),
    .B(net868));
 sg13g2_o21ai_1 _19952_ (.B1(_03762_),
    .Y(_02541_),
    .A1(_10089_),
    .A2(net869));
 sg13g2_buf_2 _19953_ (.A(\top_ihp.oisc.wb_dat_o[13] ),
    .X(_03763_));
 sg13g2_mux2_1 _19954_ (.A0(net1055),
    .A1(_03763_),
    .S(net870),
    .X(_02542_));
 sg13g2_inv_1 _19955_ (.Y(_03764_),
    .A(net1051));
 sg13g2_buf_2 _19956_ (.A(\top_ihp.oisc.wb_dat_o[14] ),
    .X(_03765_));
 sg13g2_nand2_1 _19957_ (.Y(_03766_),
    .A(_03765_),
    .B(_03761_));
 sg13g2_o21ai_1 _19958_ (.B1(_03766_),
    .Y(_02543_),
    .A1(_03764_),
    .A2(_03759_));
 sg13g2_buf_1 _19959_ (.A(\top_ihp.oisc.wb_dat_o[15] ),
    .X(_03767_));
 sg13g2_mux2_1 _19960_ (.A0(_08287_),
    .A1(_03767_),
    .S(net870),
    .X(_02544_));
 sg13g2_buf_2 _19961_ (.A(\top_ihp.oisc.wb_dat_o[16] ),
    .X(_03768_));
 sg13g2_nand2_1 _19962_ (.Y(_03769_),
    .A(_03768_),
    .B(net868));
 sg13g2_o21ai_1 _19963_ (.B1(_03769_),
    .Y(_02545_),
    .A1(_08291_),
    .A2(net869));
 sg13g2_buf_1 _19964_ (.A(\top_ihp.oisc.wb_dat_o[17] ),
    .X(_03770_));
 sg13g2_mux2_1 _19965_ (.A0(net1052),
    .A1(_03770_),
    .S(net870),
    .X(_02546_));
 sg13g2_inv_1 _19966_ (.Y(_03771_),
    .A(net1059));
 sg13g2_buf_2 _19967_ (.A(\top_ihp.oisc.wb_dat_o[18] ),
    .X(_03772_));
 sg13g2_nand2_1 _19968_ (.Y(_03773_),
    .A(_03772_),
    .B(net868));
 sg13g2_o21ai_1 _19969_ (.B1(_03773_),
    .Y(_02547_),
    .A1(_03771_),
    .A2(net869));
 sg13g2_buf_2 _19970_ (.A(\top_ihp.oisc.wb_dat_o[19] ),
    .X(_03774_));
 sg13g2_nand2_1 _19971_ (.Y(_03775_),
    .A(_03774_),
    .B(net868));
 sg13g2_o21ai_1 _19972_ (.B1(_03775_),
    .Y(_02548_),
    .A1(_08224_),
    .A2(net869));
 sg13g2_buf_2 _19973_ (.A(\top_ihp.oisc.wb_dat_o[1] ),
    .X(_03776_));
 sg13g2_nand2_1 _19974_ (.Y(_03777_),
    .A(_03776_),
    .B(net868));
 sg13g2_o21ai_1 _19975_ (.B1(_03777_),
    .Y(_02549_),
    .A1(net274),
    .A2(net869));
 sg13g2_buf_1 _19976_ (.A(\top_ihp.oisc.wb_dat_o[20] ),
    .X(_03778_));
 sg13g2_buf_1 _19977_ (.A(_03755_),
    .X(_03779_));
 sg13g2_mux2_1 _19978_ (.A0(net1056),
    .A1(_03778_),
    .S(net867),
    .X(_02550_));
 sg13g2_buf_2 _19979_ (.A(\top_ihp.oisc.wb_dat_o[21] ),
    .X(_03780_));
 sg13g2_nand2_1 _19980_ (.Y(_03781_),
    .A(_03780_),
    .B(net868));
 sg13g2_o21ai_1 _19981_ (.B1(_03781_),
    .Y(_02551_),
    .A1(_08236_),
    .A2(net869));
 sg13g2_buf_2 _19982_ (.A(\top_ihp.oisc.wb_dat_o[22] ),
    .X(_03782_));
 sg13g2_nand2_1 _19983_ (.Y(_03783_),
    .A(_03782_),
    .B(net868));
 sg13g2_o21ai_1 _19984_ (.B1(_03783_),
    .Y(_02552_),
    .A1(_08508_),
    .A2(net869));
 sg13g2_buf_2 _19985_ (.A(\top_ihp.oisc.wb_dat_o[23] ),
    .X(_03784_));
 sg13g2_nand2_1 _19986_ (.Y(_03785_),
    .A(_03784_),
    .B(net900));
 sg13g2_o21ai_1 _19987_ (.B1(_03785_),
    .Y(_02553_),
    .A1(net257),
    .A2(_03759_));
 sg13g2_buf_1 _19988_ (.A(\top_ihp.oisc.wb_dat_o[24] ),
    .X(_03786_));
 sg13g2_mux2_1 _19989_ (.A0(net400),
    .A1(_03786_),
    .S(net867),
    .X(_02554_));
 sg13g2_buf_1 _19990_ (.A(\top_ihp.oisc.wb_dat_o[25] ),
    .X(_03787_));
 sg13g2_mux2_1 _19991_ (.A0(_08384_),
    .A1(_03787_),
    .S(net867),
    .X(_02555_));
 sg13g2_buf_1 _19992_ (.A(\top_ihp.oisc.wb_dat_o[26] ),
    .X(_03788_));
 sg13g2_mux2_1 _19993_ (.A0(net1031),
    .A1(_03788_),
    .S(net867),
    .X(_02556_));
 sg13g2_buf_1 _19994_ (.A(\top_ihp.oisc.wb_dat_o[27] ),
    .X(_03789_));
 sg13g2_mux2_1 _19995_ (.A0(net1046),
    .A1(_03789_),
    .S(net867),
    .X(_02557_));
 sg13g2_buf_2 _19996_ (.A(\top_ihp.oisc.wb_dat_o[28] ),
    .X(_03790_));
 sg13g2_nand2_1 _19997_ (.Y(_03791_),
    .A(_03790_),
    .B(_03755_));
 sg13g2_o21ai_1 _19998_ (.B1(_03791_),
    .Y(_02558_),
    .A1(_10516_),
    .A2(net869));
 sg13g2_buf_1 _19999_ (.A(\top_ihp.oisc.wb_dat_o[29] ),
    .X(_03792_));
 sg13g2_mux2_1 _20000_ (.A0(net1045),
    .A1(_03792_),
    .S(_03779_),
    .X(_02559_));
 sg13g2_buf_2 _20001_ (.A(\top_ihp.oisc.wb_dat_o[2] ),
    .X(_03793_));
 sg13g2_nand2_1 _20002_ (.Y(_03794_),
    .A(_03793_),
    .B(net900));
 sg13g2_o21ai_1 _20003_ (.B1(_03794_),
    .Y(_02560_),
    .A1(_10779_),
    .A2(_03756_));
 sg13g2_buf_2 _20004_ (.A(\top_ihp.oisc.wb_dat_o[30] ),
    .X(_03795_));
 sg13g2_nand2_1 _20005_ (.Y(_03796_),
    .A(_03795_),
    .B(net900));
 sg13g2_o21ai_1 _20006_ (.B1(_03796_),
    .Y(_02561_),
    .A1(_10813_),
    .A2(net870));
 sg13g2_buf_1 _20007_ (.A(\top_ihp.oisc.wb_dat_o[31] ),
    .X(_03797_));
 sg13g2_mux2_1 _20008_ (.A0(_09673_),
    .A1(_03797_),
    .S(net867),
    .X(_02562_));
 sg13g2_buf_2 _20009_ (.A(\top_ihp.oisc.wb_dat_o[3] ),
    .X(_03798_));
 sg13g2_mux2_1 _20010_ (.A0(_10739_),
    .A1(_03798_),
    .S(_03779_),
    .X(_02563_));
 sg13g2_buf_2 _20011_ (.A(\top_ihp.oisc.wb_dat_o[4] ),
    .X(_03799_));
 sg13g2_mux2_1 _20012_ (.A0(net127),
    .A1(_03799_),
    .S(net867),
    .X(_02564_));
 sg13g2_buf_2 _20013_ (.A(\top_ihp.oisc.wb_dat_o[5] ),
    .X(_03800_));
 sg13g2_mux2_1 _20014_ (.A0(net264),
    .A1(_03800_),
    .S(net867),
    .X(_02565_));
 sg13g2_buf_2 _20015_ (.A(\top_ihp.oisc.wb_dat_o[6] ),
    .X(_03801_));
 sg13g2_mux2_1 _20016_ (.A0(net126),
    .A1(_03801_),
    .S(net868),
    .X(_02566_));
 sg13g2_buf_2 _20017_ (.A(\top_ihp.oisc.wb_dat_o[7] ),
    .X(_03802_));
 sg13g2_nand2_1 _20018_ (.Y(_03803_),
    .A(_03802_),
    .B(net900));
 sg13g2_o21ai_1 _20019_ (.B1(_03803_),
    .Y(_02567_),
    .A1(net396),
    .A2(_03756_));
 sg13g2_buf_2 _20020_ (.A(\top_ihp.oisc.wb_dat_o[8] ),
    .X(_03804_));
 sg13g2_nand2_1 _20021_ (.Y(_03805_),
    .A(_03804_),
    .B(net900));
 sg13g2_o21ai_1 _20022_ (.B1(_03805_),
    .Y(_02568_),
    .A1(net255),
    .A2(net870));
 sg13g2_buf_1 _20023_ (.A(\top_ihp.oisc.wb_dat_o[9] ),
    .X(_03806_));
 sg13g2_mux2_1 _20024_ (.A0(net125),
    .A1(_03806_),
    .S(_03761_),
    .X(_02569_));
 sg13g2_xor2_1 _20025_ (.B(_10484_),
    .A(_08330_),
    .X(_03807_));
 sg13g2_a21o_1 _20026_ (.A2(_03807_),
    .A1(_08417_),
    .B1(net1028),
    .X(_03808_));
 sg13g2_nor3_1 _20027_ (.A(net1050),
    .B(_08423_),
    .C(_03807_),
    .Y(_03809_));
 sg13g2_a21oi_2 _20028_ (.B1(_03809_),
    .Y(_03810_),
    .A2(_03808_),
    .A1(net1050));
 sg13g2_o21ai_1 _20029_ (.B1(_08413_),
    .Y(_03811_),
    .A1(_08317_),
    .A2(_08321_));
 sg13g2_o21ai_1 _20030_ (.B1(_03811_),
    .Y(_03812_),
    .A1(_08613_),
    .A2(_09685_));
 sg13g2_buf_1 _20031_ (.A(_03812_),
    .X(_03813_));
 sg13g2_nor2_1 _20032_ (.A(_03810_),
    .B(_03813_),
    .Y(_03814_));
 sg13g2_a21o_1 _20033_ (.A2(_10591_),
    .A1(_08417_),
    .B1(_08419_),
    .X(_03815_));
 sg13g2_nor3_1 _20034_ (.A(net1049),
    .B(_08423_),
    .C(_10591_),
    .Y(_03816_));
 sg13g2_a21o_1 _20035_ (.A2(_03815_),
    .A1(net1049),
    .B1(_03816_),
    .X(_03817_));
 sg13g2_buf_1 _20036_ (.A(_03817_),
    .X(_03818_));
 sg13g2_a22oi_1 _20037_ (.Y(_03819_),
    .B1(net832),
    .B2(_10553_),
    .A2(_08326_),
    .A1(net984));
 sg13g2_buf_2 _20038_ (.A(_03819_),
    .X(_03820_));
 sg13g2_nor2_1 _20039_ (.A(_03818_),
    .B(_03820_),
    .Y(_03821_));
 sg13g2_nand2_1 _20040_ (.Y(_03822_),
    .A(_03814_),
    .B(_03821_));
 sg13g2_buf_1 _20041_ (.A(_03822_),
    .X(_03823_));
 sg13g2_buf_1 _20042_ (.A(net717),
    .X(_03824_));
 sg13g2_buf_1 _20043_ (.A(\top_ihp.wb_coproc.opb[4] ),
    .X(_03825_));
 sg13g2_inv_1 _20044_ (.Y(_03826_),
    .A(net1033));
 sg13g2_buf_1 _20045_ (.A(_03826_),
    .X(_03827_));
 sg13g2_buf_1 _20046_ (.A(\top_ihp.wb_coproc.opb[3] ),
    .X(_03828_));
 sg13g2_buf_1 _20047_ (.A(_03828_),
    .X(_03829_));
 sg13g2_buf_1 _20048_ (.A(net998),
    .X(_03830_));
 sg13g2_buf_1 _20049_ (.A(\top_ihp.wb_coproc.opb[1] ),
    .X(_03831_));
 sg13g2_buf_1 _20050_ (.A(_03831_),
    .X(_03832_));
 sg13g2_buf_1 _20051_ (.A(net997),
    .X(_03833_));
 sg13g2_mux2_1 _20052_ (.A0(_00190_),
    .A1(_00192_),
    .S(net945),
    .X(_03834_));
 sg13g2_buf_1 _20053_ (.A(net997),
    .X(_03835_));
 sg13g2_mux2_1 _20054_ (.A0(_00189_),
    .A1(_00191_),
    .S(net944),
    .X(_03836_));
 sg13g2_buf_1 _20055_ (.A(\top_ihp.wb_coproc.opb[0] ),
    .X(_03837_));
 sg13g2_inv_1 _20056_ (.Y(_03838_),
    .A(_03837_));
 sg13g2_buf_1 _20057_ (.A(_03838_),
    .X(_03839_));
 sg13g2_buf_1 _20058_ (.A(net943),
    .X(_03840_));
 sg13g2_mux2_1 _20059_ (.A0(_03834_),
    .A1(_03836_),
    .S(net899),
    .X(_03841_));
 sg13g2_buf_1 _20060_ (.A(_03831_),
    .X(_03842_));
 sg13g2_mux2_1 _20061_ (.A0(_00194_),
    .A1(_00196_),
    .S(net996),
    .X(_03843_));
 sg13g2_mux2_1 _20062_ (.A0(_00193_),
    .A1(_00195_),
    .S(net944),
    .X(_03844_));
 sg13g2_mux2_1 _20063_ (.A0(_03843_),
    .A1(_03844_),
    .S(net899),
    .X(_03845_));
 sg13g2_buf_1 _20064_ (.A(\top_ihp.wb_coproc.opb[2] ),
    .X(_03846_));
 sg13g2_buf_1 _20065_ (.A(_03846_),
    .X(_03847_));
 sg13g2_buf_1 _20066_ (.A(net995),
    .X(_03848_));
 sg13g2_mux2_1 _20067_ (.A0(_03841_),
    .A1(_03845_),
    .S(net942),
    .X(_03849_));
 sg13g2_buf_1 _20068_ (.A(_03828_),
    .X(_03850_));
 sg13g2_buf_1 _20069_ (.A(net945),
    .X(_03851_));
 sg13g2_mux2_1 _20070_ (.A0(_00186_),
    .A1(_00188_),
    .S(net898),
    .X(_03852_));
 sg13g2_mux2_1 _20071_ (.A0(_00185_),
    .A1(_00187_),
    .S(net944),
    .X(_03853_));
 sg13g2_mux2_1 _20072_ (.A0(_03852_),
    .A1(_03853_),
    .S(net899),
    .X(_03854_));
 sg13g2_buf_1 _20073_ (.A(_03847_),
    .X(_03855_));
 sg13g2_buf_1 _20074_ (.A(\top_ihp.wb_coproc.opa[0] ),
    .X(_03856_));
 sg13g2_buf_1 _20075_ (.A(\top_ihp.wb_coproc.opa[1] ),
    .X(_03857_));
 sg13g2_inv_1 _20076_ (.Y(_03858_),
    .A(_00183_));
 sg13g2_inv_1 _20077_ (.Y(_03859_),
    .A(_00184_));
 sg13g2_buf_1 _20078_ (.A(_03837_),
    .X(_03860_));
 sg13g2_mux4_1 _20079_ (.S0(net993),
    .A0(_03856_),
    .A1(_03857_),
    .A2(_03858_),
    .A3(_03859_),
    .S1(net898),
    .X(_03861_));
 sg13g2_nor2_1 _20080_ (.A(net941),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_a21oi_1 _20081_ (.A1(net942),
    .A2(_03854_),
    .Y(_03863_),
    .B1(_03862_));
 sg13g2_nor2_1 _20082_ (.A(net994),
    .B(_03863_),
    .Y(_03864_));
 sg13g2_a21oi_1 _20083_ (.A1(net946),
    .A2(_03849_),
    .Y(_03865_),
    .B1(_03864_));
 sg13g2_mux2_1 _20084_ (.A0(_00206_),
    .A1(_00208_),
    .S(net997),
    .X(_03866_));
 sg13g2_mux2_1 _20085_ (.A0(_00205_),
    .A1(_00207_),
    .S(net996),
    .X(_03867_));
 sg13g2_mux2_1 _20086_ (.A0(_03866_),
    .A1(_03867_),
    .S(net943),
    .X(_03868_));
 sg13g2_buf_1 _20087_ (.A(_03837_),
    .X(_03869_));
 sg13g2_buf_1 _20088_ (.A(\top_ihp.wb_coproc.opa[30] ),
    .X(_03870_));
 sg13g2_nand2_1 _20089_ (.Y(_03871_),
    .A(net997),
    .B(_03870_));
 sg13g2_o21ai_1 _20090_ (.B1(_03871_),
    .Y(_03872_),
    .A1(net997),
    .A2(_00209_));
 sg13g2_nor2_1 _20091_ (.A(net992),
    .B(_03872_),
    .Y(_03873_));
 sg13g2_buf_1 _20092_ (.A(\top_ihp.wb_coproc.opa[31] ),
    .X(_03874_));
 sg13g2_nand2_1 _20093_ (.Y(_03875_),
    .A(net996),
    .B(_03874_));
 sg13g2_or2_1 _20094_ (.X(_03876_),
    .B(_00210_),
    .A(net996));
 sg13g2_nand3_1 _20095_ (.B(_03875_),
    .C(_03876_),
    .A(_03869_),
    .Y(_03877_));
 sg13g2_nand2b_1 _20096_ (.Y(_03878_),
    .B(_03877_),
    .A_N(_03873_));
 sg13g2_buf_1 _20097_ (.A(_03846_),
    .X(_03879_));
 sg13g2_mux2_1 _20098_ (.A0(_03868_),
    .A1(_03878_),
    .S(net991),
    .X(_03880_));
 sg13g2_mux2_1 _20099_ (.A0(_00198_),
    .A1(_00200_),
    .S(net996),
    .X(_03881_));
 sg13g2_mux2_1 _20100_ (.A0(_00197_),
    .A1(_00199_),
    .S(net945),
    .X(_03882_));
 sg13g2_mux2_1 _20101_ (.A0(_03881_),
    .A1(_03882_),
    .S(net943),
    .X(_03883_));
 sg13g2_mux2_1 _20102_ (.A0(_00202_),
    .A1(_00204_),
    .S(_03832_),
    .X(_03884_));
 sg13g2_mux2_1 _20103_ (.A0(_00201_),
    .A1(_00203_),
    .S(net997),
    .X(_03885_));
 sg13g2_mux2_1 _20104_ (.A0(_03884_),
    .A1(_03885_),
    .S(net943),
    .X(_03886_));
 sg13g2_mux2_1 _20105_ (.A0(_03883_),
    .A1(_03886_),
    .S(net991),
    .X(_03887_));
 sg13g2_inv_1 _20106_ (.Y(_03888_),
    .A(_03828_));
 sg13g2_buf_1 _20107_ (.A(_03888_),
    .X(_03889_));
 sg13g2_mux2_1 _20108_ (.A0(_03880_),
    .A1(_03887_),
    .S(net940),
    .X(_03890_));
 sg13g2_nor2_1 _20109_ (.A(net947),
    .B(_03890_),
    .Y(_03891_));
 sg13g2_a21oi_1 _20110_ (.A1(net947),
    .A2(_03865_),
    .Y(_03892_),
    .B1(_03891_));
 sg13g2_a21o_1 _20111_ (.A2(_03808_),
    .A1(net1050),
    .B1(_03809_),
    .X(_03893_));
 sg13g2_nor2_1 _20112_ (.A(_03893_),
    .B(_03813_),
    .Y(_03894_));
 sg13g2_a21oi_2 _20113_ (.B1(_03816_),
    .Y(_03895_),
    .A2(_03815_),
    .A1(net1049));
 sg13g2_nor2_1 _20114_ (.A(_03895_),
    .B(_03820_),
    .Y(_03896_));
 sg13g2_nand2_1 _20115_ (.Y(_03897_),
    .A(_03894_),
    .B(_03896_));
 sg13g2_buf_2 _20116_ (.A(_03897_),
    .X(_03898_));
 sg13g2_buf_1 _20117_ (.A(_03898_),
    .X(_03899_));
 sg13g2_and2_1 _20118_ (.A(_03896_),
    .B(_03814_),
    .X(_03900_));
 sg13g2_buf_1 _20119_ (.A(_03900_),
    .X(_03901_));
 sg13g2_buf_1 _20120_ (.A(_03901_),
    .X(_03902_));
 sg13g2_inv_1 _20121_ (.Y(_03903_),
    .A(_03813_));
 sg13g2_and3_1 _20122_ (.X(_03904_),
    .A(_03893_),
    .B(_03903_),
    .C(_03820_));
 sg13g2_buf_1 _20123_ (.A(_03904_),
    .X(_03905_));
 sg13g2_nand2_1 _20124_ (.Y(_03906_),
    .A(_03818_),
    .B(_03905_));
 sg13g2_buf_1 _20125_ (.A(_03906_),
    .X(_03907_));
 sg13g2_buf_1 _20126_ (.A(_03907_),
    .X(_03908_));
 sg13g2_nand3_1 _20127_ (.B(_03856_),
    .C(net625),
    .A(net993),
    .Y(_03909_));
 sg13g2_o21ai_1 _20128_ (.B1(_03909_),
    .Y(_03910_),
    .A1(_03856_),
    .A2(net715));
 sg13g2_nand2_1 _20129_ (.Y(_03911_),
    .A(_03896_),
    .B(_03814_));
 sg13g2_nand2_1 _20130_ (.Y(_03912_),
    .A(_03898_),
    .B(_03911_));
 sg13g2_buf_1 _20131_ (.A(_03912_),
    .X(_03913_));
 sg13g2_buf_1 _20132_ (.A(_03913_),
    .X(_03914_));
 sg13g2_a21oi_1 _20133_ (.A1(_03856_),
    .A2(net624),
    .Y(_03915_),
    .B1(net993));
 sg13g2_a21o_1 _20134_ (.A2(_03910_),
    .A1(net716),
    .B1(_03915_),
    .X(_03916_));
 sg13g2_o21ai_1 _20135_ (.B1(_03916_),
    .Y(_03917_),
    .A1(_03824_),
    .A2(_03892_));
 sg13g2_nand3b_1 _20136_ (.B(_08213_),
    .C(_08604_),
    .Y(_03918_),
    .A_N(_08598_));
 sg13g2_buf_2 _20137_ (.A(_03918_),
    .X(_03919_));
 sg13g2_buf_1 _20138_ (.A(_03919_),
    .X(_03920_));
 sg13g2_mux2_1 _20139_ (.A0(_03917_),
    .A1(\top_ihp.wb_coproc.dat_o[0] ),
    .S(net204),
    .X(_02570_));
 sg13g2_mux2_1 _20140_ (.A0(_00204_),
    .A1(_00206_),
    .S(net996),
    .X(_03921_));
 sg13g2_mux2_1 _20141_ (.A0(_00203_),
    .A1(_00205_),
    .S(_03832_),
    .X(_03922_));
 sg13g2_mux2_1 _20142_ (.A0(_03921_),
    .A1(_03922_),
    .S(_03840_),
    .X(_03923_));
 sg13g2_mux2_1 _20143_ (.A0(_00200_),
    .A1(_00202_),
    .S(_03833_),
    .X(_03924_));
 sg13g2_mux2_1 _20144_ (.A0(_00199_),
    .A1(_00201_),
    .S(net996),
    .X(_03925_));
 sg13g2_mux2_1 _20145_ (.A0(_03924_),
    .A1(_03925_),
    .S(net943),
    .X(_03926_));
 sg13g2_nor2b_1 _20146_ (.A(_03879_),
    .B_N(_03926_),
    .Y(_03927_));
 sg13g2_a21oi_1 _20147_ (.A1(net941),
    .A2(_03923_),
    .Y(_03928_),
    .B1(_03927_));
 sg13g2_buf_1 _20148_ (.A(net940),
    .X(_03929_));
 sg13g2_nor2_1 _20149_ (.A(net897),
    .B(net1033),
    .Y(_03930_));
 sg13g2_nor2b_1 _20150_ (.A(net997),
    .B_N(_00207_),
    .Y(_03931_));
 sg13g2_a21oi_1 _20151_ (.A1(_03842_),
    .A2(_00209_),
    .Y(_03932_),
    .B1(_03931_));
 sg13g2_nand2_1 _20152_ (.Y(_03933_),
    .A(net943),
    .B(_03932_));
 sg13g2_nor2_1 _20153_ (.A(net997),
    .B(_00208_),
    .Y(_03934_));
 sg13g2_nor2b_1 _20154_ (.A(_00210_),
    .B_N(_03833_),
    .Y(_03935_));
 sg13g2_o21ai_1 _20155_ (.B1(net992),
    .Y(_03936_),
    .A1(_03934_),
    .A2(_03935_));
 sg13g2_and2_1 _20156_ (.A(_03933_),
    .B(_03936_),
    .X(_03937_));
 sg13g2_mux2_1 _20157_ (.A0(_03870_),
    .A1(_03874_),
    .S(_03837_),
    .X(_03938_));
 sg13g2_nand2b_1 _20158_ (.Y(_03939_),
    .B(_03938_),
    .A_N(_03851_));
 sg13g2_mux2_1 _20159_ (.A0(_03937_),
    .A1(_03939_),
    .S(net995),
    .X(_03940_));
 sg13g2_mux2_1 _20160_ (.A0(_00192_),
    .A1(_00194_),
    .S(net944),
    .X(_03941_));
 sg13g2_mux2_1 _20161_ (.A0(_00191_),
    .A1(_00193_),
    .S(net945),
    .X(_03942_));
 sg13g2_mux2_1 _20162_ (.A0(_03941_),
    .A1(_03942_),
    .S(net899),
    .X(_03943_));
 sg13g2_mux2_1 _20163_ (.A0(_00196_),
    .A1(_00198_),
    .S(net945),
    .X(_03944_));
 sg13g2_mux2_1 _20164_ (.A0(_00195_),
    .A1(_00197_),
    .S(net996),
    .X(_03945_));
 sg13g2_mux2_1 _20165_ (.A0(_03944_),
    .A1(_03945_),
    .S(net943),
    .X(_03946_));
 sg13g2_mux2_1 _20166_ (.A0(_03943_),
    .A1(_03946_),
    .S(net991),
    .X(_03947_));
 sg13g2_mux2_1 _20167_ (.A0(_03940_),
    .A1(_03947_),
    .S(_03826_),
    .X(_03948_));
 sg13g2_nor2_1 _20168_ (.A(net946),
    .B(_03948_),
    .Y(_03949_));
 sg13g2_a21oi_1 _20169_ (.A1(_03928_),
    .A2(_03930_),
    .Y(_03950_),
    .B1(_03949_));
 sg13g2_buf_1 _20170_ (.A(\top_ihp.wb_coproc.opa[10] ),
    .X(_03951_));
 sg13g2_nand3_1 _20171_ (.B(_03951_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[10] ),
    .Y(_03952_));
 sg13g2_o21ai_1 _20172_ (.B1(_03952_),
    .Y(_03953_),
    .A1(_03951_),
    .A2(net715));
 sg13g2_a21oi_1 _20173_ (.A1(_03951_),
    .A2(net624),
    .Y(_03954_),
    .B1(\top_ihp.wb_coproc.opb[10] ));
 sg13g2_a21o_1 _20174_ (.A2(_03953_),
    .A1(net716),
    .B1(_03954_),
    .X(_03955_));
 sg13g2_o21ai_1 _20175_ (.B1(_03955_),
    .Y(_03956_),
    .A1(net687),
    .A2(_03950_));
 sg13g2_mux2_1 _20176_ (.A0(_03956_),
    .A1(\top_ihp.wb_coproc.dat_o[10] ),
    .S(net204),
    .X(_02571_));
 sg13g2_mux2_1 _20177_ (.A0(_03844_),
    .A1(_03941_),
    .S(_03840_),
    .X(_03957_));
 sg13g2_mux2_1 _20178_ (.A0(_03882_),
    .A1(_03944_),
    .S(net899),
    .X(_03958_));
 sg13g2_mux2_1 _20179_ (.A0(_03957_),
    .A1(_03958_),
    .S(net941),
    .X(_03959_));
 sg13g2_buf_1 _20180_ (.A(\top_ihp.wb_coproc.opa[29] ),
    .X(_03960_));
 sg13g2_a21oi_1 _20181_ (.A1(_03842_),
    .A2(_03960_),
    .Y(_03961_),
    .B1(_03934_));
 sg13g2_nor2_1 _20182_ (.A(_03837_),
    .B(_03961_),
    .Y(_03962_));
 sg13g2_a21oi_1 _20183_ (.A1(net992),
    .A2(_03872_),
    .Y(_03963_),
    .B1(_03962_));
 sg13g2_inv_1 _20184_ (.Y(_03964_),
    .A(_03874_));
 sg13g2_nor3_2 _20185_ (.A(net992),
    .B(_03835_),
    .C(_03964_),
    .Y(_03965_));
 sg13g2_nand2_1 _20186_ (.Y(_03966_),
    .A(_03846_),
    .B(_03965_));
 sg13g2_o21ai_1 _20187_ (.B1(_03966_),
    .Y(_03967_),
    .A1(net995),
    .A2(_03963_));
 sg13g2_nand2_1 _20188_ (.Y(_03968_),
    .A(net1033),
    .B(_03967_));
 sg13g2_o21ai_1 _20189_ (.B1(_03968_),
    .Y(_03969_),
    .A1(net1033),
    .A2(_03959_));
 sg13g2_mux2_1 _20190_ (.A0(_03867_),
    .A1(_03921_),
    .S(net943),
    .X(_03970_));
 sg13g2_mux2_1 _20191_ (.A0(_03885_),
    .A1(_03924_),
    .S(_03839_),
    .X(_03971_));
 sg13g2_nor2b_1 _20192_ (.A(net991),
    .B_N(_03971_),
    .Y(_03972_));
 sg13g2_a21oi_1 _20193_ (.A1(net941),
    .A2(_03970_),
    .Y(_03973_),
    .B1(_03972_));
 sg13g2_a22oi_1 _20194_ (.Y(_03974_),
    .B1(_03973_),
    .B2(_03930_),
    .A2(_03969_),
    .A1(net897));
 sg13g2_buf_1 _20195_ (.A(\top_ihp.wb_coproc.opa[11] ),
    .X(_03975_));
 sg13g2_nand3_1 _20196_ (.B(_03975_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[11] ),
    .Y(_03976_));
 sg13g2_o21ai_1 _20197_ (.B1(_03976_),
    .Y(_03977_),
    .A1(_03975_),
    .A2(net715));
 sg13g2_a21oi_1 _20198_ (.A1(_03975_),
    .A2(net624),
    .Y(_03978_),
    .B1(\top_ihp.wb_coproc.opb[11] ));
 sg13g2_a21o_1 _20199_ (.A2(_03977_),
    .A1(net716),
    .B1(_03978_),
    .X(_03979_));
 sg13g2_o21ai_1 _20200_ (.B1(_03979_),
    .Y(_03980_),
    .A1(net687),
    .A2(_03974_));
 sg13g2_mux2_1 _20201_ (.A0(_03980_),
    .A1(\top_ihp.wb_coproc.dat_o[11] ),
    .S(net204),
    .X(_02572_));
 sg13g2_nor2b_1 _20202_ (.A(_03873_),
    .B_N(_03877_),
    .Y(_03981_));
 sg13g2_buf_1 _20203_ (.A(_03879_),
    .X(_03982_));
 sg13g2_nand2_1 _20204_ (.Y(_03983_),
    .A(net1033),
    .B(_00181_));
 sg13g2_nor2_1 _20205_ (.A(net939),
    .B(_03983_),
    .Y(_03984_));
 sg13g2_mux2_1 _20206_ (.A0(_03845_),
    .A1(_03883_),
    .S(net991),
    .X(_03985_));
 sg13g2_nor2b_1 _20207_ (.A(_03847_),
    .B_N(_03886_),
    .Y(_03986_));
 sg13g2_a21oi_1 _20208_ (.A1(net991),
    .A2(_03868_),
    .Y(_03987_),
    .B1(_03986_));
 sg13g2_nand2_1 _20209_ (.Y(_03988_),
    .A(net994),
    .B(_03987_));
 sg13g2_o21ai_1 _20210_ (.B1(_03988_),
    .Y(_03989_),
    .A1(net994),
    .A2(_03985_));
 sg13g2_a22oi_1 _20211_ (.Y(_03990_),
    .B1(_03989_),
    .B2(_03827_),
    .A2(_03984_),
    .A1(_03981_));
 sg13g2_buf_1 _20212_ (.A(\top_ihp.wb_coproc.opa[12] ),
    .X(_03991_));
 sg13g2_nand3_1 _20213_ (.B(_03991_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[12] ),
    .Y(_03992_));
 sg13g2_o21ai_1 _20214_ (.B1(_03992_),
    .Y(_03993_),
    .A1(_03991_),
    .A2(net715));
 sg13g2_a21oi_1 _20215_ (.A1(_03991_),
    .A2(net624),
    .Y(_03994_),
    .B1(\top_ihp.wb_coproc.opb[12] ));
 sg13g2_a21o_1 _20216_ (.A2(_03993_),
    .A1(net716),
    .B1(_03994_),
    .X(_03995_));
 sg13g2_o21ai_1 _20217_ (.B1(_03995_),
    .Y(_03996_),
    .A1(net687),
    .A2(_03990_));
 sg13g2_mux2_1 _20218_ (.A0(_03996_),
    .A1(\top_ihp.wb_coproc.dat_o[12] ),
    .S(net204),
    .X(_02573_));
 sg13g2_nand2b_1 _20219_ (.Y(_03997_),
    .B(_03960_),
    .A_N(net945));
 sg13g2_a21oi_1 _20220_ (.A1(_03875_),
    .A2(_03997_),
    .Y(_03998_),
    .B1(_03860_));
 sg13g2_nand3b_1 _20221_ (.B(_03870_),
    .C(net992),
    .Y(_03999_),
    .A_N(_03835_));
 sg13g2_nand2b_1 _20222_ (.Y(_04000_),
    .B(_03999_),
    .A_N(_03998_));
 sg13g2_and2_1 _20223_ (.A(_00182_),
    .B(_04000_),
    .X(_04001_));
 sg13g2_inv_1 _20224_ (.Y(_04002_),
    .A(_04001_));
 sg13g2_mux2_1 _20225_ (.A0(_03884_),
    .A1(_03922_),
    .S(_03869_),
    .X(_04003_));
 sg13g2_nor2_1 _20226_ (.A(_03837_),
    .B(_03866_),
    .Y(_04004_));
 sg13g2_a21oi_1 _20227_ (.A1(net992),
    .A2(_03932_),
    .Y(_04005_),
    .B1(_04004_));
 sg13g2_mux2_1 _20228_ (.A0(_04003_),
    .A1(_04005_),
    .S(net995),
    .X(_04006_));
 sg13g2_nor2_1 _20229_ (.A(net940),
    .B(_04006_),
    .Y(_04007_));
 sg13g2_mux2_1 _20230_ (.A0(_03843_),
    .A1(_03945_),
    .S(net992),
    .X(_04008_));
 sg13g2_mux2_1 _20231_ (.A0(_03881_),
    .A1(_03925_),
    .S(net992),
    .X(_04009_));
 sg13g2_mux2_1 _20232_ (.A0(_04008_),
    .A1(_04009_),
    .S(net995),
    .X(_04010_));
 sg13g2_nor2_1 _20233_ (.A(_03828_),
    .B(_04010_),
    .Y(_04011_));
 sg13g2_o21ai_1 _20234_ (.B1(_03826_),
    .Y(_04012_),
    .A1(_04007_),
    .A2(_04011_));
 sg13g2_o21ai_1 _20235_ (.B1(_04012_),
    .Y(_04013_),
    .A1(_03983_),
    .A2(_04002_));
 sg13g2_nor2b_1 _20236_ (.A(_03823_),
    .B_N(_04013_),
    .Y(_04014_));
 sg13g2_buf_1 _20237_ (.A(_03898_),
    .X(_04015_));
 sg13g2_buf_1 _20238_ (.A(\top_ihp.wb_coproc.opa[13] ),
    .X(_04016_));
 sg13g2_buf_1 _20239_ (.A(_03901_),
    .X(_04017_));
 sg13g2_buf_1 _20240_ (.A(_03907_),
    .X(_04018_));
 sg13g2_nand3_1 _20241_ (.B(_04016_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[13] ),
    .Y(_04019_));
 sg13g2_o21ai_1 _20242_ (.B1(_04019_),
    .Y(_04020_),
    .A1(_04016_),
    .A2(net713));
 sg13g2_buf_1 _20243_ (.A(_03913_),
    .X(_04021_));
 sg13g2_a21oi_1 _20244_ (.A1(_04016_),
    .A2(net622),
    .Y(_04022_),
    .B1(\top_ihp.wb_coproc.opb[13] ));
 sg13g2_a21oi_1 _20245_ (.A1(net714),
    .A2(_04020_),
    .Y(_04023_),
    .B1(_04022_));
 sg13g2_or2_1 _20246_ (.X(_04024_),
    .B(_04023_),
    .A(_04014_));
 sg13g2_mux2_1 _20247_ (.A0(_04024_),
    .A1(\top_ihp.wb_coproc.dat_o[13] ),
    .S(net204),
    .X(_02574_));
 sg13g2_nor2b_1 _20248_ (.A(_03851_),
    .B_N(_03938_),
    .Y(_04025_));
 sg13g2_buf_1 _20249_ (.A(net1033),
    .X(_04026_));
 sg13g2_mux2_1 _20250_ (.A0(_03923_),
    .A1(_03937_),
    .S(net941),
    .X(_04027_));
 sg13g2_mux2_1 _20251_ (.A0(_03946_),
    .A1(_03926_),
    .S(net991),
    .X(_04028_));
 sg13g2_mux2_1 _20252_ (.A0(_04027_),
    .A1(_04028_),
    .S(_03889_),
    .X(_04029_));
 sg13g2_nor2_1 _20253_ (.A(net990),
    .B(_04029_),
    .Y(_04030_));
 sg13g2_a21oi_1 _20254_ (.A1(_04025_),
    .A2(_03984_),
    .Y(_04031_),
    .B1(_04030_));
 sg13g2_buf_1 _20255_ (.A(\top_ihp.wb_coproc.opa[14] ),
    .X(_04032_));
 sg13g2_nand3_1 _20256_ (.B(_04032_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[14] ),
    .Y(_04033_));
 sg13g2_o21ai_1 _20257_ (.B1(_04033_),
    .Y(_04034_),
    .A1(_04032_),
    .A2(net715));
 sg13g2_a21oi_1 _20258_ (.A1(_04032_),
    .A2(net624),
    .Y(_04035_),
    .B1(\top_ihp.wb_coproc.opb[14] ));
 sg13g2_a21o_1 _20259_ (.A2(_04034_),
    .A1(net716),
    .B1(_04035_),
    .X(_04036_));
 sg13g2_o21ai_1 _20260_ (.B1(_04036_),
    .Y(_04037_),
    .A1(net687),
    .A2(_04031_));
 sg13g2_mux2_1 _20261_ (.A0(_04037_),
    .A1(\top_ihp.wb_coproc.dat_o[14] ),
    .S(_03920_),
    .X(_02575_));
 sg13g2_mux2_1 _20262_ (.A0(_03958_),
    .A1(_03971_),
    .S(_03848_),
    .X(_04038_));
 sg13g2_nor2b_1 _20263_ (.A(net995),
    .B_N(_03970_),
    .Y(_04039_));
 sg13g2_a21oi_1 _20264_ (.A1(_03855_),
    .A2(_03963_),
    .Y(_04040_),
    .B1(_04039_));
 sg13g2_nand2_1 _20265_ (.Y(_04041_),
    .A(_03850_),
    .B(_04040_));
 sg13g2_o21ai_1 _20266_ (.B1(_04041_),
    .Y(_04042_),
    .A1(net994),
    .A2(_04038_));
 sg13g2_a22oi_1 _20267_ (.Y(_04043_),
    .B1(_04042_),
    .B2(_03827_),
    .A2(_03984_),
    .A1(_03965_));
 sg13g2_buf_1 _20268_ (.A(\top_ihp.wb_coproc.opa[15] ),
    .X(_04044_));
 sg13g2_nand3_1 _20269_ (.B(_04044_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[15] ),
    .Y(_04045_));
 sg13g2_o21ai_1 _20270_ (.B1(_04045_),
    .Y(_04046_),
    .A1(_04044_),
    .A2(net715));
 sg13g2_a21oi_1 _20271_ (.A1(_04044_),
    .A2(net624),
    .Y(_04047_),
    .B1(\top_ihp.wb_coproc.opb[15] ));
 sg13g2_a21o_1 _20272_ (.A2(_04046_),
    .A1(net716),
    .B1(_04047_),
    .X(_04048_));
 sg13g2_o21ai_1 _20273_ (.B1(_04048_),
    .Y(_04049_),
    .A1(net687),
    .A2(_04043_));
 sg13g2_mux2_1 _20274_ (.A0(_04049_),
    .A1(\top_ihp.wb_coproc.dat_o[15] ),
    .S(net204),
    .X(_02576_));
 sg13g2_nand2b_1 _20275_ (.Y(_04050_),
    .B(_00180_),
    .A_N(_03890_));
 sg13g2_buf_1 _20276_ (.A(\top_ihp.wb_coproc.opa[16] ),
    .X(_04051_));
 sg13g2_nand3_1 _20277_ (.B(_04051_),
    .C(_03908_),
    .A(\top_ihp.wb_coproc.opb[16] ),
    .Y(_04052_));
 sg13g2_o21ai_1 _20278_ (.B1(_04052_),
    .Y(_04053_),
    .A1(_04051_),
    .A2(_03902_));
 sg13g2_a21oi_1 _20279_ (.A1(_04051_),
    .A2(net624),
    .Y(_04054_),
    .B1(\top_ihp.wb_coproc.opb[16] ));
 sg13g2_a21o_1 _20280_ (.A2(_04053_),
    .A1(_03899_),
    .B1(_04054_),
    .X(_04055_));
 sg13g2_o21ai_1 _20281_ (.B1(_04055_),
    .Y(_04056_),
    .A1(net687),
    .A2(_04050_));
 sg13g2_mux2_1 _20282_ (.A0(_04056_),
    .A1(\top_ihp.wb_coproc.dat_o[16] ),
    .S(net204),
    .X(_02577_));
 sg13g2_inv_1 _20283_ (.Y(_04057_),
    .A(_04005_));
 sg13g2_mux2_1 _20284_ (.A0(_04057_),
    .A1(_04000_),
    .S(net995),
    .X(_04058_));
 sg13g2_mux2_1 _20285_ (.A0(_04009_),
    .A1(_04003_),
    .S(net995),
    .X(_04059_));
 sg13g2_nor2_1 _20286_ (.A(net998),
    .B(_04059_),
    .Y(_04060_));
 sg13g2_a21oi_1 _20287_ (.A1(net998),
    .A2(_04058_),
    .Y(_04061_),
    .B1(_04060_));
 sg13g2_nand3_1 _20288_ (.B(_03814_),
    .C(_03821_),
    .A(_03826_),
    .Y(_04062_));
 sg13g2_buf_2 _20289_ (.A(_04062_),
    .X(_04063_));
 sg13g2_buf_1 _20290_ (.A(\top_ihp.wb_coproc.opa[17] ),
    .X(_04064_));
 sg13g2_nand3_1 _20291_ (.B(_04064_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[17] ),
    .Y(_04065_));
 sg13g2_o21ai_1 _20292_ (.B1(_04065_),
    .Y(_04066_),
    .A1(_04064_),
    .A2(net715));
 sg13g2_a21oi_1 _20293_ (.A1(_04064_),
    .A2(net624),
    .Y(_04067_),
    .B1(\top_ihp.wb_coproc.opb[17] ));
 sg13g2_a21o_1 _20294_ (.A2(_04066_),
    .A1(net716),
    .B1(_04067_),
    .X(_04068_));
 sg13g2_o21ai_1 _20295_ (.B1(_04068_),
    .Y(_04069_),
    .A1(_04061_),
    .A2(_04063_));
 sg13g2_mux2_1 _20296_ (.A0(_04069_),
    .A1(\top_ihp.wb_coproc.dat_o[17] ),
    .S(_03920_),
    .X(_02578_));
 sg13g2_nor2_1 _20297_ (.A(net940),
    .B(_03940_),
    .Y(_04070_));
 sg13g2_a21oi_1 _20298_ (.A1(net897),
    .A2(_03928_),
    .Y(_04071_),
    .B1(_04070_));
 sg13g2_buf_1 _20299_ (.A(\top_ihp.wb_coproc.opa[18] ),
    .X(_04072_));
 sg13g2_nand3_1 _20300_ (.B(_04072_),
    .C(net625),
    .A(\top_ihp.wb_coproc.opb[18] ),
    .Y(_04073_));
 sg13g2_o21ai_1 _20301_ (.B1(_04073_),
    .Y(_04074_),
    .A1(_04072_),
    .A2(net715));
 sg13g2_a21oi_1 _20302_ (.A1(_04072_),
    .A2(_03914_),
    .Y(_04075_),
    .B1(\top_ihp.wb_coproc.opb[18] ));
 sg13g2_a21o_1 _20303_ (.A2(_04074_),
    .A1(net716),
    .B1(_04075_),
    .X(_04076_));
 sg13g2_o21ai_1 _20304_ (.B1(_04076_),
    .Y(_04077_),
    .A1(_04063_),
    .A2(_04071_));
 sg13g2_mux2_1 _20305_ (.A0(_04077_),
    .A1(\top_ihp.wb_coproc.dat_o[18] ),
    .S(net204),
    .X(_02579_));
 sg13g2_and2_1 _20306_ (.A(net998),
    .B(_03967_),
    .X(_04078_));
 sg13g2_a21oi_1 _20307_ (.A1(net897),
    .A2(_03973_),
    .Y(_04079_),
    .B1(_04078_));
 sg13g2_buf_1 _20308_ (.A(\top_ihp.wb_coproc.opa[19] ),
    .X(_04080_));
 sg13g2_nand3_1 _20309_ (.B(_04080_),
    .C(_03908_),
    .A(\top_ihp.wb_coproc.opb[19] ),
    .Y(_04081_));
 sg13g2_o21ai_1 _20310_ (.B1(_04081_),
    .Y(_04082_),
    .A1(_04080_),
    .A2(_03902_));
 sg13g2_buf_1 _20311_ (.A(_03913_),
    .X(_04083_));
 sg13g2_a21oi_1 _20312_ (.A1(_04080_),
    .A2(net621),
    .Y(_04084_),
    .B1(\top_ihp.wb_coproc.opb[19] ));
 sg13g2_a21o_1 _20313_ (.A2(_04082_),
    .A1(_03899_),
    .B1(_04084_),
    .X(_04085_));
 sg13g2_o21ai_1 _20314_ (.B1(_04085_),
    .Y(_04086_),
    .A1(_04063_),
    .A2(_04079_));
 sg13g2_buf_1 _20315_ (.A(_03919_),
    .X(_04087_));
 sg13g2_mux2_1 _20316_ (.A0(_04086_),
    .A1(\top_ihp.wb_coproc.dat_o[19] ),
    .S(net203),
    .X(_02580_));
 sg13g2_mux2_1 _20317_ (.A0(_03834_),
    .A1(_03942_),
    .S(net993),
    .X(_04088_));
 sg13g2_mux2_1 _20318_ (.A0(_04088_),
    .A1(_04008_),
    .S(net991),
    .X(_04089_));
 sg13g2_mux2_1 _20319_ (.A0(_00187_),
    .A1(_00189_),
    .S(net945),
    .X(_04090_));
 sg13g2_mux2_1 _20320_ (.A0(_03852_),
    .A1(_04090_),
    .S(net993),
    .X(_04091_));
 sg13g2_nand2_1 _20321_ (.Y(_04092_),
    .A(net944),
    .B(_00185_));
 sg13g2_o21ai_1 _20322_ (.B1(_04092_),
    .Y(_04093_),
    .A1(_03858_),
    .A2(net944));
 sg13g2_nand2_1 _20323_ (.Y(_04094_),
    .A(net993),
    .B(_04093_));
 sg13g2_nor2_1 _20324_ (.A(net944),
    .B(_00211_),
    .Y(_04095_));
 sg13g2_a21oi_1 _20325_ (.A1(_03859_),
    .A2(net898),
    .Y(_04096_),
    .B1(_04095_));
 sg13g2_nand2_1 _20326_ (.Y(_04097_),
    .A(net899),
    .B(_04096_));
 sg13g2_a21oi_1 _20327_ (.A1(_04094_),
    .A2(_04097_),
    .Y(_04098_),
    .B1(net941));
 sg13g2_a21oi_1 _20328_ (.A1(net942),
    .A2(_04091_),
    .Y(_04099_),
    .B1(_04098_));
 sg13g2_nor2_1 _20329_ (.A(net994),
    .B(_04099_),
    .Y(_04100_));
 sg13g2_a21oi_1 _20330_ (.A1(net946),
    .A2(_04089_),
    .Y(_04101_),
    .B1(_04100_));
 sg13g2_nor2_1 _20331_ (.A(net947),
    .B(_04061_),
    .Y(_04102_));
 sg13g2_a21oi_1 _20332_ (.A1(net947),
    .A2(_04101_),
    .Y(_04103_),
    .B1(_04102_));
 sg13g2_buf_1 _20333_ (.A(_03898_),
    .X(_04104_));
 sg13g2_buf_1 _20334_ (.A(_03901_),
    .X(_04105_));
 sg13g2_buf_1 _20335_ (.A(_03907_),
    .X(_04106_));
 sg13g2_nand3_1 _20336_ (.B(net898),
    .C(net620),
    .A(_03857_),
    .Y(_04107_));
 sg13g2_o21ai_1 _20337_ (.B1(_04107_),
    .Y(_04108_),
    .A1(net898),
    .A2(net711));
 sg13g2_a21oi_1 _20338_ (.A1(net898),
    .A2(net621),
    .Y(_04109_),
    .B1(_03857_));
 sg13g2_a21o_1 _20339_ (.A2(_04108_),
    .A1(net712),
    .B1(_04109_),
    .X(_04110_));
 sg13g2_o21ai_1 _20340_ (.B1(_04110_),
    .Y(_04111_),
    .A1(net687),
    .A2(_04103_));
 sg13g2_mux2_1 _20341_ (.A0(_04111_),
    .A1(\top_ihp.wb_coproc.dat_o[1] ),
    .S(net203),
    .X(_02581_));
 sg13g2_nor2_1 _20342_ (.A(_03855_),
    .B(net940),
    .Y(_04112_));
 sg13g2_a22oi_1 _20343_ (.Y(_04113_),
    .B1(_04112_),
    .B2(_03981_),
    .A2(_03987_),
    .A1(net940));
 sg13g2_buf_1 _20344_ (.A(\top_ihp.wb_coproc.opa[20] ),
    .X(_04114_));
 sg13g2_nand3_1 _20345_ (.B(_04114_),
    .C(_04106_),
    .A(\top_ihp.wb_coproc.opb[20] ),
    .Y(_04115_));
 sg13g2_o21ai_1 _20346_ (.B1(_04115_),
    .Y(_04116_),
    .A1(_04114_),
    .A2(net711));
 sg13g2_a21oi_1 _20347_ (.A1(_04114_),
    .A2(net621),
    .Y(_04117_),
    .B1(\top_ihp.wb_coproc.opb[20] ));
 sg13g2_a21o_1 _20348_ (.A2(_04116_),
    .A1(net712),
    .B1(_04117_),
    .X(_04118_));
 sg13g2_o21ai_1 _20349_ (.B1(_04118_),
    .Y(_04119_),
    .A1(_04063_),
    .A2(_04113_));
 sg13g2_mux2_1 _20350_ (.A0(_04119_),
    .A1(\top_ihp.wb_coproc.dat_o[20] ),
    .S(net203),
    .X(_02582_));
 sg13g2_nor2_1 _20351_ (.A(_03829_),
    .B(_04006_),
    .Y(_04120_));
 sg13g2_a21oi_1 _20352_ (.A1(net998),
    .A2(_04001_),
    .Y(_04121_),
    .B1(_04120_));
 sg13g2_buf_1 _20353_ (.A(\top_ihp.wb_coproc.opa[21] ),
    .X(_04122_));
 sg13g2_nand3_1 _20354_ (.B(_04122_),
    .C(net620),
    .A(\top_ihp.wb_coproc.opb[21] ),
    .Y(_04123_));
 sg13g2_o21ai_1 _20355_ (.B1(_04123_),
    .Y(_04124_),
    .A1(_04122_),
    .A2(net711));
 sg13g2_a21oi_1 _20356_ (.A1(_04122_),
    .A2(net621),
    .Y(_04125_),
    .B1(\top_ihp.wb_coproc.opb[21] ));
 sg13g2_a21o_1 _20357_ (.A2(_04124_),
    .A1(net712),
    .B1(_04125_),
    .X(_04126_));
 sg13g2_o21ai_1 _20358_ (.B1(_04126_),
    .Y(_04127_),
    .A1(_04063_),
    .A2(_04121_));
 sg13g2_mux2_1 _20359_ (.A0(_04127_),
    .A1(\top_ihp.wb_coproc.dat_o[21] ),
    .S(net203),
    .X(_02583_));
 sg13g2_nor2_1 _20360_ (.A(net1033),
    .B(_03823_),
    .Y(_04128_));
 sg13g2_nand2_1 _20361_ (.Y(_04129_),
    .A(_04025_),
    .B(_04112_));
 sg13g2_o21ai_1 _20362_ (.B1(_04129_),
    .Y(_04130_),
    .A1(net994),
    .A2(_04027_));
 sg13g2_buf_1 _20363_ (.A(\top_ihp.wb_coproc.opa[22] ),
    .X(_04131_));
 sg13g2_nand3_1 _20364_ (.B(_04131_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[22] ),
    .Y(_04132_));
 sg13g2_o21ai_1 _20365_ (.B1(_04132_),
    .Y(_04133_),
    .A1(_04131_),
    .A2(net713));
 sg13g2_a21oi_1 _20366_ (.A1(_04131_),
    .A2(net622),
    .Y(_04134_),
    .B1(\top_ihp.wb_coproc.opb[22] ));
 sg13g2_a21oi_1 _20367_ (.A1(net714),
    .A2(_04133_),
    .Y(_04135_),
    .B1(_04134_));
 sg13g2_a21o_1 _20368_ (.A2(_04130_),
    .A1(_04128_),
    .B1(_04135_),
    .X(_04136_));
 sg13g2_mux2_1 _20369_ (.A0(_04136_),
    .A1(\top_ihp.wb_coproc.dat_o[22] ),
    .S(net203),
    .X(_02584_));
 sg13g2_a22oi_1 _20370_ (.Y(_04137_),
    .B1(_04112_),
    .B2(_03965_),
    .A2(_04040_),
    .A1(_03929_));
 sg13g2_buf_1 _20371_ (.A(\top_ihp.wb_coproc.opa[23] ),
    .X(_04138_));
 sg13g2_nand3_1 _20372_ (.B(_04138_),
    .C(net620),
    .A(\top_ihp.wb_coproc.opb[23] ),
    .Y(_04139_));
 sg13g2_o21ai_1 _20373_ (.B1(_04139_),
    .Y(_04140_),
    .A1(_04138_),
    .A2(net711));
 sg13g2_a21oi_1 _20374_ (.A1(_04138_),
    .A2(net621),
    .Y(_04141_),
    .B1(\top_ihp.wb_coproc.opb[23] ));
 sg13g2_a21o_1 _20375_ (.A2(_04140_),
    .A1(net712),
    .B1(_04141_),
    .X(_04142_));
 sg13g2_o21ai_1 _20376_ (.B1(_04142_),
    .Y(_04143_),
    .A1(_04063_),
    .A2(_04137_));
 sg13g2_mux2_1 _20377_ (.A0(_04143_),
    .A1(\top_ihp.wb_coproc.dat_o[23] ),
    .S(net203),
    .X(_02585_));
 sg13g2_nand2_1 _20378_ (.Y(_04144_),
    .A(_00181_),
    .B(_04128_));
 sg13g2_buf_1 _20379_ (.A(\top_ihp.wb_coproc.opa[24] ),
    .X(_04145_));
 sg13g2_nand3_1 _20380_ (.B(_04145_),
    .C(net620),
    .A(\top_ihp.wb_coproc.opb[24] ),
    .Y(_04146_));
 sg13g2_o21ai_1 _20381_ (.B1(_04146_),
    .Y(_04147_),
    .A1(_04145_),
    .A2(net711));
 sg13g2_a21oi_1 _20382_ (.A1(_04145_),
    .A2(net621),
    .Y(_04148_),
    .B1(\top_ihp.wb_coproc.opb[24] ));
 sg13g2_a21o_1 _20383_ (.A2(_04147_),
    .A1(net712),
    .B1(_04148_),
    .X(_04149_));
 sg13g2_o21ai_1 _20384_ (.B1(_04149_),
    .Y(_04150_),
    .A1(_03880_),
    .A2(_04144_));
 sg13g2_mux2_1 _20385_ (.A0(_04150_),
    .A1(\top_ihp.wb_coproc.dat_o[24] ),
    .S(net203),
    .X(_02586_));
 sg13g2_nor2_1 _20386_ (.A(_03830_),
    .B(_04063_),
    .Y(_04151_));
 sg13g2_buf_1 _20387_ (.A(\top_ihp.wb_coproc.opa[25] ),
    .X(_04152_));
 sg13g2_nand3_1 _20388_ (.B(_04152_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[25] ),
    .Y(_04153_));
 sg13g2_o21ai_1 _20389_ (.B1(_04153_),
    .Y(_04154_),
    .A1(_04152_),
    .A2(net713));
 sg13g2_a21oi_1 _20390_ (.A1(_04152_),
    .A2(net622),
    .Y(_04155_),
    .B1(\top_ihp.wb_coproc.opb[25] ));
 sg13g2_a21oi_1 _20391_ (.A1(net714),
    .A2(_04154_),
    .Y(_04156_),
    .B1(_04155_));
 sg13g2_a21o_1 _20392_ (.A2(_04151_),
    .A1(_04058_),
    .B1(_04156_),
    .X(_04157_));
 sg13g2_mux2_1 _20393_ (.A0(_04157_),
    .A1(\top_ihp.wb_coproc.dat_o[25] ),
    .S(net203),
    .X(_02587_));
 sg13g2_nor3_1 _20394_ (.A(net946),
    .B(_03940_),
    .C(_04063_),
    .Y(_04158_));
 sg13g2_buf_1 _20395_ (.A(\top_ihp.wb_coproc.opa[26] ),
    .X(_04159_));
 sg13g2_nand3_1 _20396_ (.B(_04159_),
    .C(_03907_),
    .A(\top_ihp.wb_coproc.opb[26] ),
    .Y(_04160_));
 sg13g2_o21ai_1 _20397_ (.B1(_04160_),
    .Y(_04161_),
    .A1(_04159_),
    .A2(_03901_));
 sg13g2_a21oi_1 _20398_ (.A1(_04159_),
    .A2(_03913_),
    .Y(_04162_),
    .B1(\top_ihp.wb_coproc.opb[26] ));
 sg13g2_a21oi_1 _20399_ (.A1(_03898_),
    .A2(_04161_),
    .Y(_04163_),
    .B1(_04162_));
 sg13g2_or2_1 _20400_ (.X(_04164_),
    .B(_04163_),
    .A(_04158_));
 sg13g2_mux2_1 _20401_ (.A0(_04164_),
    .A1(\top_ihp.wb_coproc.dat_o[26] ),
    .S(_04087_),
    .X(_02588_));
 sg13g2_buf_1 _20402_ (.A(\top_ihp.wb_coproc.opa[27] ),
    .X(_04165_));
 sg13g2_nand3_1 _20403_ (.B(_04165_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[27] ),
    .Y(_04166_));
 sg13g2_o21ai_1 _20404_ (.B1(_04166_),
    .Y(_04167_),
    .A1(_04165_),
    .A2(net713));
 sg13g2_a21oi_1 _20405_ (.A1(_04165_),
    .A2(net622),
    .Y(_04168_),
    .B1(\top_ihp.wb_coproc.opb[27] ));
 sg13g2_a21oi_1 _20406_ (.A1(net714),
    .A2(_04167_),
    .Y(_04169_),
    .B1(_04168_));
 sg13g2_a21o_1 _20407_ (.A2(_04151_),
    .A1(_03967_),
    .B1(_04169_),
    .X(_04170_));
 sg13g2_mux2_1 _20408_ (.A0(_04170_),
    .A1(\top_ihp.wb_coproc.dat_o[27] ),
    .S(_04087_),
    .X(_02589_));
 sg13g2_or2_1 _20409_ (.X(_04171_),
    .B(_04144_),
    .A(net939));
 sg13g2_buf_1 _20410_ (.A(\top_ihp.wb_coproc.opa[28] ),
    .X(_04172_));
 sg13g2_nand3_1 _20411_ (.B(_04172_),
    .C(net620),
    .A(\top_ihp.wb_coproc.opb[28] ),
    .Y(_04173_));
 sg13g2_o21ai_1 _20412_ (.B1(_04173_),
    .Y(_04174_),
    .A1(_04172_),
    .A2(_04105_));
 sg13g2_a21oi_1 _20413_ (.A1(_04172_),
    .A2(_04083_),
    .Y(_04175_),
    .B1(\top_ihp.wb_coproc.opb[28] ));
 sg13g2_a21o_1 _20414_ (.A2(_04174_),
    .A1(_04104_),
    .B1(_04175_),
    .X(_04176_));
 sg13g2_o21ai_1 _20415_ (.B1(_04176_),
    .Y(_04177_),
    .A1(_03878_),
    .A2(_04171_));
 sg13g2_buf_1 _20416_ (.A(_03919_),
    .X(_04178_));
 sg13g2_mux2_1 _20417_ (.A0(_04177_),
    .A1(\top_ihp.wb_coproc.dat_o[28] ),
    .S(_04178_),
    .X(_02590_));
 sg13g2_buf_1 _20418_ (.A(\top_ihp.wb_coproc.opb[29] ),
    .X(_04179_));
 sg13g2_nand3_1 _20419_ (.B(_04179_),
    .C(net620),
    .A(_03960_),
    .Y(_04180_));
 sg13g2_o21ai_1 _20420_ (.B1(_04180_),
    .Y(_04181_),
    .A1(_04179_),
    .A2(net711));
 sg13g2_a21oi_1 _20421_ (.A1(_04179_),
    .A2(net621),
    .Y(_04182_),
    .B1(_03960_));
 sg13g2_a21o_1 _20422_ (.A2(_04181_),
    .A1(net712),
    .B1(_04182_),
    .X(_04183_));
 sg13g2_o21ai_1 _20423_ (.B1(_04183_),
    .Y(_04184_),
    .A1(_04002_),
    .A2(_04144_));
 sg13g2_mux2_1 _20424_ (.A0(_04184_),
    .A1(\top_ihp.wb_coproc.dat_o[29] ),
    .S(net202),
    .X(_02591_));
 sg13g2_mux2_1 _20425_ (.A0(_00188_),
    .A1(_00190_),
    .S(net945),
    .X(_04185_));
 sg13g2_mux2_1 _20426_ (.A0(_04090_),
    .A1(_04185_),
    .S(net993),
    .X(_04186_));
 sg13g2_nand2_1 _20427_ (.Y(_04187_),
    .A(net944),
    .B(_00186_));
 sg13g2_o21ai_1 _20428_ (.B1(_04187_),
    .Y(_04188_),
    .A1(_03859_),
    .A2(net898));
 sg13g2_mux2_1 _20429_ (.A0(_04093_),
    .A1(_04188_),
    .S(net993),
    .X(_04189_));
 sg13g2_nor2b_1 _20430_ (.A(net942),
    .B_N(_04189_),
    .Y(_04190_));
 sg13g2_a21oi_1 _20431_ (.A1(net939),
    .A2(_04186_),
    .Y(_04191_),
    .B1(_04190_));
 sg13g2_nor2_1 _20432_ (.A(net897),
    .B(_03947_),
    .Y(_04192_));
 sg13g2_a21oi_1 _20433_ (.A1(net897),
    .A2(_04191_),
    .Y(_04193_),
    .B1(_04192_));
 sg13g2_mux2_1 _20434_ (.A0(_04071_),
    .A1(_04193_),
    .S(net947),
    .X(_04194_));
 sg13g2_buf_1 _20435_ (.A(\top_ihp.wb_coproc.opa[2] ),
    .X(_04195_));
 sg13g2_nand3_1 _20436_ (.B(_04195_),
    .C(net620),
    .A(net939),
    .Y(_04196_));
 sg13g2_o21ai_1 _20437_ (.B1(_04196_),
    .Y(_04197_),
    .A1(_04195_),
    .A2(net711));
 sg13g2_a21oi_1 _20438_ (.A1(_04195_),
    .A2(net621),
    .Y(_04198_),
    .B1(net939));
 sg13g2_a21o_1 _20439_ (.A2(_04197_),
    .A1(net712),
    .B1(_04198_),
    .X(_04199_));
 sg13g2_o21ai_1 _20440_ (.B1(_04199_),
    .Y(_04200_),
    .A1(net687),
    .A2(_04194_));
 sg13g2_mux2_1 _20441_ (.A0(_04200_),
    .A1(\top_ihp.wb_coproc.dat_o[2] ),
    .S(net202),
    .X(_02592_));
 sg13g2_buf_1 _20442_ (.A(\top_ihp.wb_coproc.opb[30] ),
    .X(_04201_));
 sg13g2_nand3_1 _20443_ (.B(_04201_),
    .C(net620),
    .A(_03870_),
    .Y(_04202_));
 sg13g2_o21ai_1 _20444_ (.B1(_04202_),
    .Y(_04203_),
    .A1(_04201_),
    .A2(_04105_));
 sg13g2_a21oi_1 _20445_ (.A1(_04201_),
    .A2(_04083_),
    .Y(_04204_),
    .B1(_03870_));
 sg13g2_a21o_1 _20446_ (.A2(_04203_),
    .A1(_04104_),
    .B1(_04204_),
    .X(_04205_));
 sg13g2_o21ai_1 _20447_ (.B1(_04205_),
    .Y(_04206_),
    .A1(_03939_),
    .A2(_04171_));
 sg13g2_mux2_1 _20448_ (.A0(_04206_),
    .A1(\top_ihp.wb_coproc.dat_o[30] ),
    .S(_04178_),
    .X(_02593_));
 sg13g2_nor2_1 _20449_ (.A(net939),
    .B(_04144_),
    .Y(_04207_));
 sg13g2_buf_1 _20450_ (.A(\top_ihp.wb_coproc.opb[31] ),
    .X(_04208_));
 sg13g2_nand3_1 _20451_ (.B(_04208_),
    .C(net623),
    .A(_03874_),
    .Y(_04209_));
 sg13g2_o21ai_1 _20452_ (.B1(_04209_),
    .Y(_04210_),
    .A1(_04208_),
    .A2(net713));
 sg13g2_nand2_1 _20453_ (.Y(_04211_),
    .A(_04208_),
    .B(_03914_));
 sg13g2_a22oi_1 _20454_ (.Y(_04212_),
    .B1(_04211_),
    .B2(_03964_),
    .A2(_04210_),
    .A1(net714));
 sg13g2_a21o_1 _20455_ (.A2(_04207_),
    .A1(_03965_),
    .B1(_04212_),
    .X(_04213_));
 sg13g2_mux2_1 _20456_ (.A0(_04213_),
    .A1(\top_ihp.wb_coproc.dat_o[31] ),
    .S(net202),
    .X(_02594_));
 sg13g2_mux2_1 _20457_ (.A0(_03836_),
    .A1(_04185_),
    .S(net899),
    .X(_04214_));
 sg13g2_mux2_1 _20458_ (.A0(_03853_),
    .A1(_04188_),
    .S(net899),
    .X(_04215_));
 sg13g2_nor2b_1 _20459_ (.A(net942),
    .B_N(_04215_),
    .Y(_04216_));
 sg13g2_a21oi_1 _20460_ (.A1(net939),
    .A2(_04214_),
    .Y(_04217_),
    .B1(_04216_));
 sg13g2_nor2_1 _20461_ (.A(_03929_),
    .B(_03959_),
    .Y(_04218_));
 sg13g2_a21oi_1 _20462_ (.A1(net897),
    .A2(_04217_),
    .Y(_04219_),
    .B1(_04218_));
 sg13g2_mux2_1 _20463_ (.A0(_04079_),
    .A1(_04219_),
    .S(net947),
    .X(_04220_));
 sg13g2_buf_1 _20464_ (.A(\top_ihp.wb_coproc.opa[3] ),
    .X(_04221_));
 sg13g2_nand3_1 _20465_ (.B(_04221_),
    .C(_04106_),
    .A(net998),
    .Y(_04222_));
 sg13g2_o21ai_1 _20466_ (.B1(_04222_),
    .Y(_04223_),
    .A1(_04221_),
    .A2(net711));
 sg13g2_a21oi_1 _20467_ (.A1(_04221_),
    .A2(net622),
    .Y(_04224_),
    .B1(net946));
 sg13g2_a21o_1 _20468_ (.A2(_04223_),
    .A1(net712),
    .B1(_04224_),
    .X(_04225_));
 sg13g2_o21ai_1 _20469_ (.B1(_04225_),
    .Y(_04226_),
    .A1(_03824_),
    .A2(_04220_));
 sg13g2_mux2_1 _20470_ (.A0(_04226_),
    .A1(\top_ihp.wb_coproc.dat_o[3] ),
    .S(net202),
    .X(_02595_));
 sg13g2_buf_1 _20471_ (.A(\top_ihp.wb_coproc.opa[4] ),
    .X(_04227_));
 sg13g2_and2_1 _20472_ (.A(net1033),
    .B(_04227_),
    .X(_04228_));
 sg13g2_o21ai_1 _20473_ (.B1(_03898_),
    .Y(_04229_),
    .A1(_03911_),
    .A2(_04228_));
 sg13g2_o21ai_1 _20474_ (.B1(_04229_),
    .Y(_04230_),
    .A1(net990),
    .A2(_04227_));
 sg13g2_nand3_1 _20475_ (.B(_03818_),
    .C(_03905_),
    .A(_04227_),
    .Y(_04231_));
 sg13g2_o21ai_1 _20476_ (.B1(_04231_),
    .Y(_04232_),
    .A1(net717),
    .A2(_04113_));
 sg13g2_nand2b_1 _20477_ (.Y(_04233_),
    .B(net941),
    .A_N(_03841_));
 sg13g2_o21ai_1 _20478_ (.B1(_04233_),
    .Y(_04234_),
    .A1(net942),
    .A2(_03854_));
 sg13g2_nor2_1 _20479_ (.A(net940),
    .B(_03985_),
    .Y(_04235_));
 sg13g2_a21oi_1 _20480_ (.A1(net897),
    .A2(_04234_),
    .Y(_04236_),
    .B1(_04235_));
 sg13g2_nor3_1 _20481_ (.A(net990),
    .B(net717),
    .C(_04236_),
    .Y(_04237_));
 sg13g2_a21oi_1 _20482_ (.A1(net990),
    .A2(_04232_),
    .Y(_04238_),
    .B1(_04237_));
 sg13g2_nand2_1 _20483_ (.Y(_04239_),
    .A(_04230_),
    .B(_04238_));
 sg13g2_mux2_1 _20484_ (.A0(_04239_),
    .A1(\top_ihp.wb_coproc.dat_o[4] ),
    .S(net202),
    .X(_02596_));
 sg13g2_nand2_1 _20485_ (.Y(_04240_),
    .A(_03982_),
    .B(_04088_));
 sg13g2_nand2b_1 _20486_ (.Y(_04241_),
    .B(_04091_),
    .A_N(net942));
 sg13g2_a21oi_1 _20487_ (.A1(_04240_),
    .A2(_04241_),
    .Y(_04242_),
    .B1(net994));
 sg13g2_a21oi_1 _20488_ (.A1(net946),
    .A2(_04010_),
    .Y(_04243_),
    .B1(_04242_));
 sg13g2_nor2_1 _20489_ (.A(_03826_),
    .B(_04121_),
    .Y(_04244_));
 sg13g2_a21oi_1 _20490_ (.A1(net947),
    .A2(_04243_),
    .Y(_04245_),
    .B1(_04244_));
 sg13g2_buf_1 _20491_ (.A(\top_ihp.wb_coproc.opa[5] ),
    .X(_04246_));
 sg13g2_nand3_1 _20492_ (.B(_04246_),
    .C(_04018_),
    .A(\top_ihp.wb_coproc.opb[5] ),
    .Y(_04247_));
 sg13g2_o21ai_1 _20493_ (.B1(_04247_),
    .Y(_04248_),
    .A1(_04246_),
    .A2(_04017_));
 sg13g2_a21oi_1 _20494_ (.A1(_04246_),
    .A2(net622),
    .Y(_04249_),
    .B1(\top_ihp.wb_coproc.opb[5] ));
 sg13g2_a21o_1 _20495_ (.A2(_04248_),
    .A1(net714),
    .B1(_04249_),
    .X(_04250_));
 sg13g2_o21ai_1 _20496_ (.B1(_04250_),
    .Y(_04251_),
    .A1(net717),
    .A2(_04245_));
 sg13g2_mux2_1 _20497_ (.A0(_04251_),
    .A1(\top_ihp.wb_coproc.dat_o[5] ),
    .S(net202),
    .X(_02597_));
 sg13g2_nor2b_1 _20498_ (.A(net941),
    .B_N(_04186_),
    .Y(_04252_));
 sg13g2_a21oi_1 _20499_ (.A1(_03848_),
    .A2(_03943_),
    .Y(_04253_),
    .B1(_04252_));
 sg13g2_nand2_1 _20500_ (.Y(_04254_),
    .A(_03829_),
    .B(_04028_));
 sg13g2_o21ai_1 _20501_ (.B1(_04254_),
    .Y(_04255_),
    .A1(net998),
    .A2(_04253_));
 sg13g2_nor2_1 _20502_ (.A(net990),
    .B(_04255_),
    .Y(_04256_));
 sg13g2_a21oi_1 _20503_ (.A1(net990),
    .A2(_04130_),
    .Y(_04257_),
    .B1(_04256_));
 sg13g2_buf_1 _20504_ (.A(\top_ihp.wb_coproc.opa[6] ),
    .X(_04258_));
 sg13g2_nand3_1 _20505_ (.B(_04258_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[6] ),
    .Y(_04259_));
 sg13g2_o21ai_1 _20506_ (.B1(_04259_),
    .Y(_04260_),
    .A1(_04258_),
    .A2(net713));
 sg13g2_a21oi_1 _20507_ (.A1(_04258_),
    .A2(net622),
    .Y(_04261_),
    .B1(\top_ihp.wb_coproc.opb[6] ));
 sg13g2_a21o_1 _20508_ (.A2(_04260_),
    .A1(net714),
    .B1(_04261_),
    .X(_04262_));
 sg13g2_o21ai_1 _20509_ (.B1(_04262_),
    .Y(_04263_),
    .A1(net717),
    .A2(_04257_));
 sg13g2_mux2_1 _20510_ (.A0(_04263_),
    .A1(\top_ihp.wb_coproc.dat_o[6] ),
    .S(net202),
    .X(_02598_));
 sg13g2_nand2_1 _20511_ (.Y(_04264_),
    .A(_03982_),
    .B(_03957_));
 sg13g2_nand2b_1 _20512_ (.Y(_04265_),
    .B(_04214_),
    .A_N(net942));
 sg13g2_a21oi_1 _20513_ (.A1(_04264_),
    .A2(_04265_),
    .Y(_04266_),
    .B1(net998));
 sg13g2_a21oi_1 _20514_ (.A1(_03850_),
    .A2(_04038_),
    .Y(_04267_),
    .B1(_04266_));
 sg13g2_nand2_1 _20515_ (.Y(_04268_),
    .A(net990),
    .B(_04137_));
 sg13g2_o21ai_1 _20516_ (.B1(_04268_),
    .Y(_04269_),
    .A1(_04026_),
    .A2(_04267_));
 sg13g2_buf_1 _20517_ (.A(\top_ihp.wb_coproc.opa[7] ),
    .X(_04270_));
 sg13g2_nand3_1 _20518_ (.B(_04270_),
    .C(_04018_),
    .A(\top_ihp.wb_coproc.opb[7] ),
    .Y(_04271_));
 sg13g2_o21ai_1 _20519_ (.B1(_04271_),
    .Y(_04272_),
    .A1(_04270_),
    .A2(_04017_));
 sg13g2_a21oi_1 _20520_ (.A1(_04270_),
    .A2(net622),
    .Y(_04273_),
    .B1(\top_ihp.wb_coproc.opb[7] ));
 sg13g2_a21o_1 _20521_ (.A2(_04272_),
    .A1(net714),
    .B1(_04273_),
    .X(_04274_));
 sg13g2_o21ai_1 _20522_ (.B1(_04274_),
    .Y(_04275_),
    .A1(net717),
    .A2(_04269_));
 sg13g2_mux2_1 _20523_ (.A0(_04275_),
    .A1(\top_ihp.wb_coproc.dat_o[7] ),
    .S(net202),
    .X(_02599_));
 sg13g2_or2_1 _20524_ (.X(_04276_),
    .B(_03887_),
    .A(net940));
 sg13g2_o21ai_1 _20525_ (.B1(_04276_),
    .Y(_04277_),
    .A1(net994),
    .A2(_03849_));
 sg13g2_nor2_1 _20526_ (.A(_03880_),
    .B(_03983_),
    .Y(_04278_));
 sg13g2_a21oi_1 _20527_ (.A1(net947),
    .A2(_04277_),
    .Y(_04279_),
    .B1(_04278_));
 sg13g2_buf_1 _20528_ (.A(\top_ihp.wb_coproc.opa[8] ),
    .X(_04280_));
 sg13g2_nand3_1 _20529_ (.B(_04280_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[8] ),
    .Y(_04281_));
 sg13g2_o21ai_1 _20530_ (.B1(_04281_),
    .Y(_04282_),
    .A1(_04280_),
    .A2(net713));
 sg13g2_a21oi_1 _20531_ (.A1(_04280_),
    .A2(_04021_),
    .Y(_04283_),
    .B1(\top_ihp.wb_coproc.opb[8] ));
 sg13g2_a21o_1 _20532_ (.A2(_04282_),
    .A1(_04015_),
    .B1(_04283_),
    .X(_04284_));
 sg13g2_o21ai_1 _20533_ (.B1(_04284_),
    .Y(_04285_),
    .A1(net717),
    .A2(_04279_));
 sg13g2_mux2_1 _20534_ (.A0(_04285_),
    .A1(\top_ihp.wb_coproc.dat_o[8] ),
    .S(_03919_),
    .X(_02600_));
 sg13g2_nor2_1 _20535_ (.A(_04026_),
    .B(_04059_),
    .Y(_04286_));
 sg13g2_nor2_1 _20536_ (.A(_03825_),
    .B(_04089_),
    .Y(_04287_));
 sg13g2_a21oi_1 _20537_ (.A1(_03825_),
    .A2(_04058_),
    .Y(_04288_),
    .B1(_04287_));
 sg13g2_nor2_1 _20538_ (.A(net946),
    .B(_04288_),
    .Y(_04289_));
 sg13g2_a21oi_1 _20539_ (.A1(net946),
    .A2(_04286_),
    .Y(_04290_),
    .B1(_04289_));
 sg13g2_buf_1 _20540_ (.A(\top_ihp.wb_coproc.opa[9] ),
    .X(_04291_));
 sg13g2_nand3_1 _20541_ (.B(_04291_),
    .C(net623),
    .A(\top_ihp.wb_coproc.opb[9] ),
    .Y(_04292_));
 sg13g2_o21ai_1 _20542_ (.B1(_04292_),
    .Y(_04293_),
    .A1(_04291_),
    .A2(net713));
 sg13g2_a21oi_1 _20543_ (.A1(_04291_),
    .A2(_04021_),
    .Y(_04294_),
    .B1(\top_ihp.wb_coproc.opb[9] ));
 sg13g2_a21o_1 _20544_ (.A2(_04293_),
    .A1(_04015_),
    .B1(_04294_),
    .X(_04295_));
 sg13g2_o21ai_1 _20545_ (.B1(_04295_),
    .Y(_04296_),
    .A1(net717),
    .A2(_04290_));
 sg13g2_mux2_1 _20546_ (.A0(_04296_),
    .A1(\top_ihp.wb_coproc.dat_o[9] ),
    .S(_03919_),
    .X(_02601_));
 sg13g2_nand2_1 _20547_ (.Y(_04297_),
    .A(net831),
    .B(net832));
 sg13g2_nand3_1 _20548_ (.B(net1046),
    .C(net831),
    .A(_08420_),
    .Y(_04298_));
 sg13g2_o21ai_1 _20549_ (.B1(_04298_),
    .Y(_04299_),
    .A1(_08602_),
    .A2(_04297_));
 sg13g2_nor2_1 _20550_ (.A(_08598_),
    .B(_03818_),
    .Y(_04300_));
 sg13g2_nand4_1 _20551_ (.B(_03820_),
    .C(_04299_),
    .A(_03894_),
    .Y(_04301_),
    .D(_04300_));
 sg13g2_buf_2 _20552_ (.A(_04301_),
    .X(_04302_));
 sg13g2_buf_1 _20553_ (.A(_04302_),
    .X(_04303_));
 sg13g2_mux2_1 _20554_ (.A0(net1034),
    .A1(_03856_),
    .S(net201),
    .X(_02602_));
 sg13g2_mux2_1 _20555_ (.A0(_03757_),
    .A1(_03951_),
    .S(net201),
    .X(_02603_));
 sg13g2_mux2_1 _20556_ (.A0(_03758_),
    .A1(_03975_),
    .S(net201),
    .X(_02604_));
 sg13g2_mux2_1 _20557_ (.A0(_03760_),
    .A1(_03991_),
    .S(net201),
    .X(_02605_));
 sg13g2_mux2_1 _20558_ (.A0(_03763_),
    .A1(_04016_),
    .S(_04303_),
    .X(_02606_));
 sg13g2_mux2_1 _20559_ (.A0(_03765_),
    .A1(_04032_),
    .S(net201),
    .X(_02607_));
 sg13g2_mux2_1 _20560_ (.A0(_03767_),
    .A1(_04044_),
    .S(_04303_),
    .X(_02608_));
 sg13g2_mux2_1 _20561_ (.A0(_03768_),
    .A1(_04051_),
    .S(net201),
    .X(_02609_));
 sg13g2_mux2_1 _20562_ (.A0(_03770_),
    .A1(_04064_),
    .S(net201),
    .X(_02610_));
 sg13g2_mux2_1 _20563_ (.A0(_03772_),
    .A1(_04072_),
    .S(net201),
    .X(_02611_));
 sg13g2_buf_1 _20564_ (.A(_04302_),
    .X(_04304_));
 sg13g2_mux2_1 _20565_ (.A0(_03774_),
    .A1(_04080_),
    .S(_04304_),
    .X(_02612_));
 sg13g2_mux2_1 _20566_ (.A0(_03776_),
    .A1(_03857_),
    .S(net200),
    .X(_02613_));
 sg13g2_mux2_1 _20567_ (.A0(_03778_),
    .A1(_04114_),
    .S(net200),
    .X(_02614_));
 sg13g2_mux2_1 _20568_ (.A0(_03780_),
    .A1(_04122_),
    .S(net200),
    .X(_02615_));
 sg13g2_mux2_1 _20569_ (.A0(_03782_),
    .A1(_04131_),
    .S(net200),
    .X(_02616_));
 sg13g2_mux2_1 _20570_ (.A0(_03784_),
    .A1(_04138_),
    .S(net200),
    .X(_02617_));
 sg13g2_mux2_1 _20571_ (.A0(_03786_),
    .A1(_04145_),
    .S(net200),
    .X(_02618_));
 sg13g2_mux2_1 _20572_ (.A0(_03787_),
    .A1(_04152_),
    .S(_04304_),
    .X(_02619_));
 sg13g2_mux2_1 _20573_ (.A0(_03788_),
    .A1(_04159_),
    .S(net200),
    .X(_02620_));
 sg13g2_mux2_1 _20574_ (.A0(_03789_),
    .A1(_04165_),
    .S(net200),
    .X(_02621_));
 sg13g2_buf_1 _20575_ (.A(_04302_),
    .X(_04305_));
 sg13g2_mux2_1 _20576_ (.A0(_03790_),
    .A1(_04172_),
    .S(net199),
    .X(_02622_));
 sg13g2_mux2_1 _20577_ (.A0(_03792_),
    .A1(_03960_),
    .S(net199),
    .X(_02623_));
 sg13g2_mux2_1 _20578_ (.A0(_03793_),
    .A1(_04195_),
    .S(net199),
    .X(_02624_));
 sg13g2_mux2_1 _20579_ (.A0(_03795_),
    .A1(_03870_),
    .S(net199),
    .X(_02625_));
 sg13g2_mux2_1 _20580_ (.A0(_03797_),
    .A1(_03874_),
    .S(net199),
    .X(_02626_));
 sg13g2_mux2_1 _20581_ (.A0(_03798_),
    .A1(_04221_),
    .S(net199),
    .X(_02627_));
 sg13g2_mux2_1 _20582_ (.A0(_03799_),
    .A1(_04227_),
    .S(net199),
    .X(_02628_));
 sg13g2_mux2_1 _20583_ (.A0(_03800_),
    .A1(_04246_),
    .S(_04305_),
    .X(_02629_));
 sg13g2_mux2_1 _20584_ (.A0(_03801_),
    .A1(_04258_),
    .S(net199),
    .X(_02630_));
 sg13g2_mux2_1 _20585_ (.A0(_03802_),
    .A1(_04270_),
    .S(_04305_),
    .X(_02631_));
 sg13g2_mux2_1 _20586_ (.A0(_03804_),
    .A1(_04280_),
    .S(_04302_),
    .X(_02632_));
 sg13g2_mux2_1 _20587_ (.A0(_03806_),
    .A1(_04291_),
    .S(_04302_),
    .X(_02633_));
 sg13g2_nand3_1 _20588_ (.B(_04299_),
    .C(_04300_),
    .A(_03905_),
    .Y(_04306_));
 sg13g2_buf_2 _20589_ (.A(_04306_),
    .X(_04307_));
 sg13g2_buf_1 _20590_ (.A(_04307_),
    .X(_04308_));
 sg13g2_mux2_1 _20591_ (.A0(net1034),
    .A1(_03860_),
    .S(net198),
    .X(_02634_));
 sg13g2_mux2_1 _20592_ (.A0(_03757_),
    .A1(\top_ihp.wb_coproc.opb[10] ),
    .S(net198),
    .X(_02635_));
 sg13g2_mux2_1 _20593_ (.A0(_03758_),
    .A1(\top_ihp.wb_coproc.opb[11] ),
    .S(net198),
    .X(_02636_));
 sg13g2_mux2_1 _20594_ (.A0(_03760_),
    .A1(\top_ihp.wb_coproc.opb[12] ),
    .S(net198),
    .X(_02637_));
 sg13g2_mux2_1 _20595_ (.A0(_03763_),
    .A1(\top_ihp.wb_coproc.opb[13] ),
    .S(_04308_),
    .X(_02638_));
 sg13g2_mux2_1 _20596_ (.A0(_03765_),
    .A1(\top_ihp.wb_coproc.opb[14] ),
    .S(net198),
    .X(_02639_));
 sg13g2_mux2_1 _20597_ (.A0(_03767_),
    .A1(\top_ihp.wb_coproc.opb[15] ),
    .S(net198),
    .X(_02640_));
 sg13g2_mux2_1 _20598_ (.A0(_03768_),
    .A1(\top_ihp.wb_coproc.opb[16] ),
    .S(net198),
    .X(_02641_));
 sg13g2_mux2_1 _20599_ (.A0(_03770_),
    .A1(\top_ihp.wb_coproc.opb[17] ),
    .S(net198),
    .X(_02642_));
 sg13g2_mux2_1 _20600_ (.A0(_03772_),
    .A1(\top_ihp.wb_coproc.opb[18] ),
    .S(_04308_),
    .X(_02643_));
 sg13g2_buf_1 _20601_ (.A(_04307_),
    .X(_04309_));
 sg13g2_mux2_1 _20602_ (.A0(_03774_),
    .A1(\top_ihp.wb_coproc.opb[19] ),
    .S(net197),
    .X(_02644_));
 sg13g2_mux2_1 _20603_ (.A0(_03776_),
    .A1(net898),
    .S(net197),
    .X(_02645_));
 sg13g2_mux2_1 _20604_ (.A0(_03778_),
    .A1(\top_ihp.wb_coproc.opb[20] ),
    .S(net197),
    .X(_02646_));
 sg13g2_mux2_1 _20605_ (.A0(_03780_),
    .A1(\top_ihp.wb_coproc.opb[21] ),
    .S(net197),
    .X(_02647_));
 sg13g2_mux2_1 _20606_ (.A0(_03782_),
    .A1(\top_ihp.wb_coproc.opb[22] ),
    .S(_04309_),
    .X(_02648_));
 sg13g2_mux2_1 _20607_ (.A0(_03784_),
    .A1(\top_ihp.wb_coproc.opb[23] ),
    .S(net197),
    .X(_02649_));
 sg13g2_mux2_1 _20608_ (.A0(_03786_),
    .A1(\top_ihp.wb_coproc.opb[24] ),
    .S(_04309_),
    .X(_02650_));
 sg13g2_mux2_1 _20609_ (.A0(_03787_),
    .A1(\top_ihp.wb_coproc.opb[25] ),
    .S(net197),
    .X(_02651_));
 sg13g2_mux2_1 _20610_ (.A0(_03788_),
    .A1(\top_ihp.wb_coproc.opb[26] ),
    .S(net197),
    .X(_02652_));
 sg13g2_mux2_1 _20611_ (.A0(_03789_),
    .A1(\top_ihp.wb_coproc.opb[27] ),
    .S(net197),
    .X(_02653_));
 sg13g2_buf_1 _20612_ (.A(_04307_),
    .X(_04310_));
 sg13g2_mux2_1 _20613_ (.A0(_03790_),
    .A1(\top_ihp.wb_coproc.opb[28] ),
    .S(net196),
    .X(_02654_));
 sg13g2_mux2_1 _20614_ (.A0(_03792_),
    .A1(_04179_),
    .S(net196),
    .X(_02655_));
 sg13g2_mux2_1 _20615_ (.A0(_03793_),
    .A1(net939),
    .S(_04310_),
    .X(_02656_));
 sg13g2_mux2_1 _20616_ (.A0(_03795_),
    .A1(_04201_),
    .S(_04310_),
    .X(_02657_));
 sg13g2_mux2_1 _20617_ (.A0(_03797_),
    .A1(_04208_),
    .S(net196),
    .X(_02658_));
 sg13g2_mux2_1 _20618_ (.A0(_03798_),
    .A1(_03830_),
    .S(net196),
    .X(_02659_));
 sg13g2_mux2_1 _20619_ (.A0(_03799_),
    .A1(net990),
    .S(net196),
    .X(_02660_));
 sg13g2_mux2_1 _20620_ (.A0(_03800_),
    .A1(\top_ihp.wb_coproc.opb[5] ),
    .S(net196),
    .X(_02661_));
 sg13g2_mux2_1 _20621_ (.A0(_03801_),
    .A1(\top_ihp.wb_coproc.opb[6] ),
    .S(net196),
    .X(_02662_));
 sg13g2_mux2_1 _20622_ (.A0(_03802_),
    .A1(\top_ihp.wb_coproc.opb[7] ),
    .S(net196),
    .X(_02663_));
 sg13g2_mux2_1 _20623_ (.A0(_03804_),
    .A1(\top_ihp.wb_coproc.opb[8] ),
    .S(_04307_),
    .X(_02664_));
 sg13g2_mux2_1 _20624_ (.A0(_03806_),
    .A1(\top_ihp.wb_coproc.opb[9] ),
    .S(_04307_),
    .X(_02665_));
 sg13g2_inv_1 _20625_ (.Y(_04311_),
    .A(_00264_));
 sg13g2_nand2_1 _20626_ (.Y(_04312_),
    .A(_08948_),
    .B(net1023));
 sg13g2_nand2_1 _20627_ (.Y(_04313_),
    .A(net1022),
    .B(_08953_));
 sg13g2_nand2b_1 _20628_ (.Y(_04314_),
    .B(_04313_),
    .A_N(_04312_));
 sg13g2_buf_1 _20629_ (.A(_04314_),
    .X(_04315_));
 sg13g2_buf_1 _20630_ (.A(\top_ihp.wb_emem.bit_counter[0] ),
    .X(_04316_));
 sg13g2_inv_1 _20631_ (.Y(_04317_),
    .A(_08948_));
 sg13g2_buf_1 _20632_ (.A(_04317_),
    .X(_04318_));
 sg13g2_inv_1 _20633_ (.Y(_04319_),
    .A(net1023));
 sg13g2_nand2_1 _20634_ (.Y(_04320_),
    .A(net896),
    .B(_04319_));
 sg13g2_nand3_1 _20635_ (.B(_04320_),
    .C(_04315_),
    .A(_04316_),
    .Y(_04321_));
 sg13g2_o21ai_1 _20636_ (.B1(_04321_),
    .Y(_02666_),
    .A1(_04311_),
    .A2(_04315_));
 sg13g2_buf_1 _20637_ (.A(\top_ihp.wb_emem.bit_counter[1] ),
    .X(_04322_));
 sg13g2_nor2_1 _20638_ (.A(net891),
    .B(_04312_),
    .Y(_04323_));
 sg13g2_buf_2 _20639_ (.A(_04323_),
    .X(_04324_));
 sg13g2_nand2_1 _20640_ (.Y(_04325_),
    .A(_04316_),
    .B(_04324_));
 sg13g2_nor2_2 _20641_ (.A(net879),
    .B(_04324_),
    .Y(_04326_));
 sg13g2_nor2_1 _20642_ (.A(_04316_),
    .B(_04315_),
    .Y(_04327_));
 sg13g2_o21ai_1 _20643_ (.B1(_04322_),
    .Y(_04328_),
    .A1(_04326_),
    .A2(_04327_));
 sg13g2_o21ai_1 _20644_ (.B1(_04328_),
    .Y(_02667_),
    .A1(_04322_),
    .A2(_04325_));
 sg13g2_nand3_1 _20645_ (.B(_04316_),
    .C(_04324_),
    .A(_04322_),
    .Y(_04329_));
 sg13g2_xor2_1 _20646_ (.B(_04329_),
    .A(\top_ihp.wb_emem.bit_counter[2] ),
    .X(_04330_));
 sg13g2_nor2_1 _20647_ (.A(net879),
    .B(_04330_),
    .Y(_02668_));
 sg13g2_buf_1 _20648_ (.A(\top_ihp.wb_emem.bit_counter[3] ),
    .X(_04331_));
 sg13g2_nand4_1 _20649_ (.B(_04316_),
    .C(\top_ihp.wb_emem.bit_counter[2] ),
    .A(_04322_),
    .Y(_04332_),
    .D(_04324_));
 sg13g2_buf_1 _20650_ (.A(_04332_),
    .X(_04333_));
 sg13g2_nand3_1 _20651_ (.B(_04320_),
    .C(_04333_),
    .A(_04331_),
    .Y(_04334_));
 sg13g2_o21ai_1 _20652_ (.B1(_04334_),
    .Y(_02669_),
    .A1(_04331_),
    .A2(_04333_));
 sg13g2_buf_2 _20653_ (.A(\top_ihp.wb_emem.bit_counter[4] ),
    .X(_04335_));
 sg13g2_and4_1 _20654_ (.A(_04322_),
    .B(_04316_),
    .C(\top_ihp.wb_emem.bit_counter[2] ),
    .D(_04331_),
    .X(_04336_));
 sg13g2_buf_1 _20655_ (.A(_04336_),
    .X(_04337_));
 sg13g2_nand2_1 _20656_ (.Y(_04338_),
    .A(_04324_),
    .B(_04337_));
 sg13g2_nor2_1 _20657_ (.A(_04315_),
    .B(_04337_),
    .Y(_04339_));
 sg13g2_o21ai_1 _20658_ (.B1(_04335_),
    .Y(_04340_),
    .A1(_04326_),
    .A2(_04339_));
 sg13g2_o21ai_1 _20659_ (.B1(_04340_),
    .Y(_02670_),
    .A1(_04335_),
    .A2(_04338_));
 sg13g2_buf_1 _20660_ (.A(\top_ihp.wb_emem.bit_counter[5] ),
    .X(_04341_));
 sg13g2_and2_1 _20661_ (.A(_04335_),
    .B(_04337_),
    .X(_04342_));
 sg13g2_buf_1 _20662_ (.A(_04342_),
    .X(_04343_));
 sg13g2_nand2_1 _20663_ (.Y(_04344_),
    .A(_04324_),
    .B(_04343_));
 sg13g2_nor2_1 _20664_ (.A(_04315_),
    .B(_04343_),
    .Y(_04345_));
 sg13g2_o21ai_1 _20665_ (.B1(_04341_),
    .Y(_04346_),
    .A1(_04326_),
    .A2(_04345_));
 sg13g2_o21ai_1 _20666_ (.B1(_04346_),
    .Y(_02671_),
    .A1(_04341_),
    .A2(_04344_));
 sg13g2_buf_1 _20667_ (.A(\top_ihp.wb_emem.bit_counter[6] ),
    .X(_04347_));
 sg13g2_nand3_1 _20668_ (.B(_04324_),
    .C(_04343_),
    .A(_04341_),
    .Y(_04348_));
 sg13g2_a21oi_1 _20669_ (.A1(_04341_),
    .A2(_04343_),
    .Y(_04349_),
    .B1(_04315_));
 sg13g2_o21ai_1 _20670_ (.B1(_04347_),
    .Y(_04350_),
    .A1(_04326_),
    .A2(_04349_));
 sg13g2_o21ai_1 _20671_ (.B1(_04350_),
    .Y(_02672_),
    .A1(_04347_),
    .A2(_04348_));
 sg13g2_nand2_1 _20672_ (.Y(_04351_),
    .A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(_04320_));
 sg13g2_nand4_1 _20673_ (.B(_04347_),
    .C(_04324_),
    .A(_04341_),
    .Y(_04352_),
    .D(_04343_));
 sg13g2_mux2_1 _20674_ (.A0(\top_ihp.wb_emem.bit_counter[7] ),
    .A1(_04351_),
    .S(_04352_),
    .X(_04353_));
 sg13g2_inv_1 _20675_ (.Y(_02673_),
    .A(_04353_));
 sg13g2_a21oi_1 _20676_ (.A1(_04319_),
    .A2(net891),
    .Y(_04354_),
    .B1(_08948_));
 sg13g2_buf_1 _20677_ (.A(_04354_),
    .X(_04355_));
 sg13g2_buf_1 _20678_ (.A(_04355_),
    .X(_04356_));
 sg13g2_buf_1 _20679_ (.A(_04356_),
    .X(_04357_));
 sg13g2_nand2_1 _20680_ (.Y(_04358_),
    .A(net879),
    .B(_08965_));
 sg13g2_buf_1 _20681_ (.A(_04358_),
    .X(_04359_));
 sg13g2_buf_1 _20682_ (.A(_04359_),
    .X(_04360_));
 sg13g2_nand2_1 _20683_ (.Y(_04361_),
    .A(net4),
    .B(net820));
 sg13g2_nor2_1 _20684_ (.A(_04320_),
    .B(_04313_),
    .Y(_04362_));
 sg13g2_buf_1 _20685_ (.A(_04362_),
    .X(_04363_));
 sg13g2_buf_1 _20686_ (.A(net843),
    .X(_04364_));
 sg13g2_nand3_1 _20687_ (.B(net797),
    .C(net819),
    .A(_03786_),
    .Y(_04365_));
 sg13g2_buf_1 _20688_ (.A(_04355_),
    .X(_04366_));
 sg13g2_a21oi_1 _20689_ (.A1(_04361_),
    .A2(_04365_),
    .Y(_04367_),
    .B1(net818));
 sg13g2_a21o_1 _20690_ (.A2(net789),
    .A1(\top_ihp.wb_dati_ram[24] ),
    .B1(_04367_),
    .X(_02674_));
 sg13g2_nand2_1 _20691_ (.Y(_04368_),
    .A(\top_ihp.wb_dati_ram[17] ),
    .B(net820));
 sg13g2_nand3_1 _20692_ (.B(net797),
    .C(net819),
    .A(_03772_),
    .Y(_04369_));
 sg13g2_a21oi_1 _20693_ (.A1(_04368_),
    .A2(_04369_),
    .Y(_04370_),
    .B1(net818));
 sg13g2_a21o_1 _20694_ (.A2(net789),
    .A1(\top_ihp.wb_dati_ram[18] ),
    .B1(_04370_),
    .X(_02675_));
 sg13g2_nand2_1 _20695_ (.Y(_04371_),
    .A(\top_ihp.wb_dati_ram[18] ),
    .B(net820));
 sg13g2_nand3_1 _20696_ (.B(_08441_),
    .C(net819),
    .A(_03774_),
    .Y(_04372_));
 sg13g2_a21oi_1 _20697_ (.A1(_04371_),
    .A2(_04372_),
    .Y(_04373_),
    .B1(_04366_));
 sg13g2_a21o_1 _20698_ (.A2(_04357_),
    .A1(\top_ihp.wb_dati_ram[19] ),
    .B1(_04373_),
    .X(_02676_));
 sg13g2_nand2_1 _20699_ (.Y(_04374_),
    .A(\top_ihp.wb_dati_ram[19] ),
    .B(net820));
 sg13g2_buf_1 _20700_ (.A(net831),
    .X(_04375_));
 sg13g2_nand3_1 _20701_ (.B(net788),
    .C(net819),
    .A(_03778_),
    .Y(_04376_));
 sg13g2_a21oi_1 _20702_ (.A1(_04374_),
    .A2(_04376_),
    .Y(_04377_),
    .B1(net818));
 sg13g2_a21o_1 _20703_ (.A2(net789),
    .A1(\top_ihp.wb_dati_ram[20] ),
    .B1(_04377_),
    .X(_02677_));
 sg13g2_nand2_1 _20704_ (.Y(_04378_),
    .A(\top_ihp.wb_dati_ram[20] ),
    .B(net820));
 sg13g2_nand3_1 _20705_ (.B(net788),
    .C(net819),
    .A(_03780_),
    .Y(_04379_));
 sg13g2_a21oi_1 _20706_ (.A1(_04378_),
    .A2(_04379_),
    .Y(_04380_),
    .B1(_04366_));
 sg13g2_a21o_1 _20707_ (.A2(net789),
    .A1(\top_ihp.wb_dati_ram[21] ),
    .B1(_04380_),
    .X(_02678_));
 sg13g2_buf_1 _20708_ (.A(_04356_),
    .X(_04381_));
 sg13g2_nand2_1 _20709_ (.Y(_04382_),
    .A(\top_ihp.wb_dati_ram[21] ),
    .B(net820));
 sg13g2_nand3_1 _20710_ (.B(net788),
    .C(net819),
    .A(_03782_),
    .Y(_04383_));
 sg13g2_a21oi_1 _20711_ (.A1(_04382_),
    .A2(_04383_),
    .Y(_04384_),
    .B1(net818));
 sg13g2_a21o_1 _20712_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[22] ),
    .B1(_04384_),
    .X(_02679_));
 sg13g2_nand2_1 _20713_ (.Y(_04385_),
    .A(\top_ihp.wb_dati_ram[22] ),
    .B(_04360_));
 sg13g2_nand3_1 _20714_ (.B(_04375_),
    .C(net819),
    .A(_03784_),
    .Y(_04386_));
 sg13g2_buf_1 _20715_ (.A(_04356_),
    .X(_04387_));
 sg13g2_a21oi_1 _20716_ (.A1(_04385_),
    .A2(_04386_),
    .Y(_04388_),
    .B1(net786));
 sg13g2_a21o_1 _20717_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[23] ),
    .B1(_04388_),
    .X(_02680_));
 sg13g2_nand2_1 _20718_ (.Y(_04389_),
    .A(\top_ihp.wb_dati_ram[23] ),
    .B(_04360_));
 sg13g2_nand3_1 _20719_ (.B(_04375_),
    .C(_04364_),
    .A(_03804_),
    .Y(_04390_));
 sg13g2_a21oi_1 _20720_ (.A1(_04389_),
    .A2(_04390_),
    .Y(_04391_),
    .B1(_04387_));
 sg13g2_a21o_1 _20721_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[8] ),
    .B1(_04391_),
    .X(_02681_));
 sg13g2_buf_1 _20722_ (.A(net844),
    .X(_04392_));
 sg13g2_nand2_1 _20723_ (.Y(_04393_),
    .A(\top_ihp.wb_dati_ram[8] ),
    .B(net817));
 sg13g2_buf_1 _20724_ (.A(net843),
    .X(_04394_));
 sg13g2_nand3_1 _20725_ (.B(net788),
    .C(net816),
    .A(_03806_),
    .Y(_04395_));
 sg13g2_a21oi_1 _20726_ (.A1(_04393_),
    .A2(_04395_),
    .Y(_04396_),
    .B1(net786));
 sg13g2_a21o_1 _20727_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[9] ),
    .B1(_04396_),
    .X(_02682_));
 sg13g2_nand2_1 _20728_ (.Y(_04397_),
    .A(\top_ihp.wb_dati_ram[9] ),
    .B(net817));
 sg13g2_nand3_1 _20729_ (.B(net788),
    .C(net816),
    .A(_03757_),
    .Y(_04398_));
 sg13g2_a21oi_1 _20730_ (.A1(_04397_),
    .A2(_04398_),
    .Y(_04399_),
    .B1(net786));
 sg13g2_a21o_1 _20731_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[10] ),
    .B1(_04399_),
    .X(_02683_));
 sg13g2_nand2_1 _20732_ (.Y(_04400_),
    .A(\top_ihp.wb_dati_ram[10] ),
    .B(net817));
 sg13g2_nand3_1 _20733_ (.B(net788),
    .C(net816),
    .A(_03758_),
    .Y(_04401_));
 sg13g2_a21oi_1 _20734_ (.A1(_04400_),
    .A2(_04401_),
    .Y(_04402_),
    .B1(net786));
 sg13g2_a21o_1 _20735_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[11] ),
    .B1(_04402_),
    .X(_02684_));
 sg13g2_nand2_1 _20736_ (.Y(_04403_),
    .A(\top_ihp.wb_dati_ram[24] ),
    .B(net817));
 sg13g2_nand3_1 _20737_ (.B(net788),
    .C(_04394_),
    .A(_03787_),
    .Y(_04404_));
 sg13g2_a21oi_1 _20738_ (.A1(_04403_),
    .A2(_04404_),
    .Y(_04405_),
    .B1(net786));
 sg13g2_a21o_1 _20739_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[25] ),
    .B1(_04405_),
    .X(_02685_));
 sg13g2_nand2_1 _20740_ (.Y(_04406_),
    .A(\top_ihp.wb_dati_ram[11] ),
    .B(net817));
 sg13g2_nand3_1 _20741_ (.B(net788),
    .C(net816),
    .A(_03760_),
    .Y(_04407_));
 sg13g2_a21oi_1 _20742_ (.A1(_04406_),
    .A2(_04407_),
    .Y(_04408_),
    .B1(net786));
 sg13g2_a21o_1 _20743_ (.A2(net787),
    .A1(\top_ihp.wb_dati_ram[12] ),
    .B1(_04408_),
    .X(_02686_));
 sg13g2_nand2_1 _20744_ (.Y(_04409_),
    .A(\top_ihp.wb_dati_ram[12] ),
    .B(_04392_));
 sg13g2_buf_1 _20745_ (.A(net831),
    .X(_04410_));
 sg13g2_nand3_1 _20746_ (.B(net785),
    .C(_04394_),
    .A(_03763_),
    .Y(_04411_));
 sg13g2_a21oi_1 _20747_ (.A1(_04409_),
    .A2(_04411_),
    .Y(_04412_),
    .B1(net786));
 sg13g2_a21o_1 _20748_ (.A2(_04381_),
    .A1(\top_ihp.wb_dati_ram[13] ),
    .B1(_04412_),
    .X(_02687_));
 sg13g2_nand2_1 _20749_ (.Y(_04413_),
    .A(\top_ihp.wb_dati_ram[13] ),
    .B(_04392_));
 sg13g2_nand3_1 _20750_ (.B(_04410_),
    .C(net816),
    .A(_03765_),
    .Y(_04414_));
 sg13g2_a21oi_1 _20751_ (.A1(_04413_),
    .A2(_04414_),
    .Y(_04415_),
    .B1(_04387_));
 sg13g2_a21o_1 _20752_ (.A2(_04381_),
    .A1(\top_ihp.wb_dati_ram[14] ),
    .B1(_04415_),
    .X(_02688_));
 sg13g2_buf_1 _20753_ (.A(_04356_),
    .X(_04416_));
 sg13g2_nand2_1 _20754_ (.Y(_04417_),
    .A(\top_ihp.wb_dati_ram[14] ),
    .B(net817));
 sg13g2_nand3_1 _20755_ (.B(_04410_),
    .C(net816),
    .A(_03767_),
    .Y(_04418_));
 sg13g2_a21oi_1 _20756_ (.A1(_04417_),
    .A2(_04418_),
    .Y(_04419_),
    .B1(net786));
 sg13g2_a21o_1 _20757_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[15] ),
    .B1(_04419_),
    .X(_02689_));
 sg13g2_buf_1 _20758_ (.A(net844),
    .X(_04420_));
 sg13g2_and2_1 _20759_ (.A(_03753_),
    .B(_04363_),
    .X(_04421_));
 sg13g2_a22oi_1 _20760_ (.Y(_04422_),
    .B1(_04421_),
    .B2(net797),
    .A2(net815),
    .A1(\top_ihp.wb_dati_ram[15] ));
 sg13g2_buf_1 _20761_ (.A(_04356_),
    .X(_04423_));
 sg13g2_nand2_1 _20762_ (.Y(_04424_),
    .A(\top_ihp.wb_dati_ram[0] ),
    .B(net783));
 sg13g2_o21ai_1 _20763_ (.B1(_04424_),
    .Y(_02690_),
    .A1(_04357_),
    .A2(_04422_));
 sg13g2_nand2_1 _20764_ (.Y(_04425_),
    .A(\top_ihp.wb_dati_ram[0] ),
    .B(net817));
 sg13g2_nand3_1 _20765_ (.B(net785),
    .C(net816),
    .A(_03776_),
    .Y(_04426_));
 sg13g2_buf_1 _20766_ (.A(_04355_),
    .X(_04427_));
 sg13g2_a21oi_1 _20767_ (.A1(_04425_),
    .A2(_04426_),
    .Y(_04428_),
    .B1(net814));
 sg13g2_a21o_1 _20768_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[1] ),
    .B1(_04428_),
    .X(_02691_));
 sg13g2_nand2_1 _20769_ (.Y(_04429_),
    .A(\top_ihp.wb_dati_ram[1] ),
    .B(net817));
 sg13g2_nand3_1 _20770_ (.B(net785),
    .C(net816),
    .A(_03793_),
    .Y(_04430_));
 sg13g2_a21oi_1 _20771_ (.A1(_04429_),
    .A2(_04430_),
    .Y(_04431_),
    .B1(net814));
 sg13g2_a21o_1 _20772_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[2] ),
    .B1(_04431_),
    .X(_02692_));
 sg13g2_buf_1 _20773_ (.A(net844),
    .X(_04432_));
 sg13g2_nand2_1 _20774_ (.Y(_04433_),
    .A(\top_ihp.wb_dati_ram[2] ),
    .B(net813));
 sg13g2_buf_1 _20775_ (.A(net843),
    .X(_04434_));
 sg13g2_nand3_1 _20776_ (.B(net785),
    .C(net812),
    .A(_03798_),
    .Y(_04435_));
 sg13g2_a21oi_1 _20777_ (.A1(_04433_),
    .A2(_04435_),
    .Y(_04436_),
    .B1(net814));
 sg13g2_a21o_1 _20778_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[3] ),
    .B1(_04436_),
    .X(_02693_));
 sg13g2_nand2_1 _20779_ (.Y(_04437_),
    .A(\top_ihp.wb_dati_ram[3] ),
    .B(net813));
 sg13g2_nand3_1 _20780_ (.B(net785),
    .C(net812),
    .A(_03799_),
    .Y(_04438_));
 sg13g2_a21oi_1 _20781_ (.A1(_04437_),
    .A2(_04438_),
    .Y(_04439_),
    .B1(_04427_));
 sg13g2_a21o_1 _20782_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[4] ),
    .B1(_04439_),
    .X(_02694_));
 sg13g2_nand2_1 _20783_ (.Y(_04440_),
    .A(\top_ihp.wb_dati_ram[4] ),
    .B(_04432_));
 sg13g2_nand3_1 _20784_ (.B(net785),
    .C(_04434_),
    .A(_03800_),
    .Y(_04441_));
 sg13g2_a21oi_1 _20785_ (.A1(_04440_),
    .A2(_04441_),
    .Y(_04442_),
    .B1(net814));
 sg13g2_a21o_1 _20786_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[5] ),
    .B1(_04442_),
    .X(_02695_));
 sg13g2_nand2_1 _20787_ (.Y(_04443_),
    .A(\top_ihp.wb_dati_ram[25] ),
    .B(net813));
 sg13g2_nand3_1 _20788_ (.B(net785),
    .C(net812),
    .A(_03788_),
    .Y(_04444_));
 sg13g2_a21oi_1 _20789_ (.A1(_04443_),
    .A2(_04444_),
    .Y(_04445_),
    .B1(net814));
 sg13g2_a21o_1 _20790_ (.A2(_04416_),
    .A1(\top_ihp.wb_dati_ram[26] ),
    .B1(_04445_),
    .X(_02696_));
 sg13g2_nand2_1 _20791_ (.Y(_04446_),
    .A(\top_ihp.wb_dati_ram[5] ),
    .B(_04432_));
 sg13g2_nand3_1 _20792_ (.B(net785),
    .C(_04434_),
    .A(_03801_),
    .Y(_04447_));
 sg13g2_a21oi_1 _20793_ (.A1(_04446_),
    .A2(_04447_),
    .Y(_04448_),
    .B1(_04427_));
 sg13g2_a21o_1 _20794_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[6] ),
    .B1(_04448_),
    .X(_02697_));
 sg13g2_nand2_1 _20795_ (.Y(_04449_),
    .A(\top_ihp.wb_dati_ram[6] ),
    .B(net813));
 sg13g2_nand3_1 _20796_ (.B(net795),
    .C(net812),
    .A(_03802_),
    .Y(_04450_));
 sg13g2_a21oi_1 _20797_ (.A1(_04449_),
    .A2(_04450_),
    .Y(_04451_),
    .B1(net814));
 sg13g2_a21o_1 _20798_ (.A2(net784),
    .A1(\top_ihp.wb_dati_ram[7] ),
    .B1(_04451_),
    .X(_02698_));
 sg13g2_and2_1 _20799_ (.A(\top_ihp.oisc.wb_adr_o[0] ),
    .B(net843),
    .X(_04452_));
 sg13g2_a21oi_1 _20800_ (.A1(\top_ihp.wb_dati_ram[7] ),
    .A2(net815),
    .Y(_04453_),
    .B1(_04452_));
 sg13g2_nand2_1 _20801_ (.Y(_04454_),
    .A(\top_ihp.wb_emem.cmd[32] ),
    .B(_04423_));
 sg13g2_o21ai_1 _20802_ (.B1(_04454_),
    .Y(_02699_),
    .A1(net789),
    .A2(_04453_));
 sg13g2_nor2_1 _20803_ (.A(_08611_),
    .B(_04420_),
    .Y(_04455_));
 sg13g2_a21oi_1 _20804_ (.A1(\top_ihp.wb_emem.cmd[32] ),
    .A2(net815),
    .Y(_04456_),
    .B1(_04455_));
 sg13g2_buf_1 _20805_ (.A(_04356_),
    .X(_04457_));
 sg13g2_nand2_1 _20806_ (.Y(_04458_),
    .A(\top_ihp.wb_emem.cmd[33] ),
    .B(net782));
 sg13g2_o21ai_1 _20807_ (.B1(_04458_),
    .Y(_02700_),
    .A1(net789),
    .A2(_04456_));
 sg13g2_nor2_1 _20808_ (.A(net820),
    .B(_03810_),
    .Y(_04459_));
 sg13g2_a21oi_1 _20809_ (.A1(\top_ihp.wb_emem.cmd[33] ),
    .A2(_04420_),
    .Y(_04460_),
    .B1(_04459_));
 sg13g2_nand2_1 _20810_ (.Y(_04461_),
    .A(\top_ihp.wb_emem.cmd[34] ),
    .B(_04457_));
 sg13g2_o21ai_1 _20811_ (.B1(_04461_),
    .Y(_02701_),
    .A1(net789),
    .A2(_04460_));
 sg13g2_inv_1 _20812_ (.Y(_04462_),
    .A(\top_ihp.wb_emem.cmd[35] ));
 sg13g2_o21ai_1 _20813_ (.B1(net896),
    .Y(_04463_),
    .A1(net1023),
    .A2(_04313_));
 sg13g2_nand2_1 _20814_ (.Y(_04464_),
    .A(\top_ihp.wb_emem.cmd[34] ),
    .B(net844));
 sg13g2_o21ai_1 _20815_ (.B1(_04464_),
    .Y(_04465_),
    .A1(net820),
    .A2(_03820_));
 sg13g2_nand2_1 _20816_ (.Y(_04466_),
    .A(_04463_),
    .B(_04465_));
 sg13g2_o21ai_1 _20817_ (.B1(_04466_),
    .Y(_02702_),
    .A1(_04462_),
    .A2(_04463_));
 sg13g2_buf_1 _20818_ (.A(_04355_),
    .X(_04467_));
 sg13g2_a221oi_1 _20819_ (.B2(net896),
    .C1(net811),
    .B1(_03895_),
    .A1(_04462_),
    .Y(_04468_),
    .A2(net815));
 sg13g2_a21o_1 _20820_ (.A2(_04416_),
    .A1(\top_ihp.wb_emem.cmd[36] ),
    .B1(_04468_),
    .X(_02703_));
 sg13g2_buf_1 _20821_ (.A(_04356_),
    .X(_04469_));
 sg13g2_inv_1 _20822_ (.Y(_04470_),
    .A(\top_ihp.wb_emem.cmd[36] ));
 sg13g2_a21o_1 _20823_ (.A2(_10603_),
    .A1(net832),
    .B1(_08420_),
    .X(_04471_));
 sg13g2_buf_1 _20824_ (.A(_08424_),
    .X(_04472_));
 sg13g2_nor3_1 _20825_ (.A(_08341_),
    .B(net762),
    .C(_10603_),
    .Y(_04473_));
 sg13g2_a21oi_2 _20826_ (.B1(_04473_),
    .Y(_04474_),
    .A2(_04471_),
    .A1(_08341_));
 sg13g2_a221oi_1 _20827_ (.B2(net896),
    .C1(_04356_),
    .B1(_04474_),
    .A1(_04470_),
    .Y(_04475_),
    .A2(net815));
 sg13g2_a21o_1 _20828_ (.A2(net781),
    .A1(\top_ihp.wb_emem.cmd[37] ),
    .B1(_04475_),
    .X(_02704_));
 sg13g2_buf_1 _20829_ (.A(net819),
    .X(_04476_));
 sg13g2_nand2_1 _20830_ (.Y(_04477_),
    .A(net796),
    .B(_10628_));
 sg13g2_o21ai_1 _20831_ (.B1(net982),
    .Y(_04478_),
    .A1(net798),
    .A2(_10628_));
 sg13g2_nand2_1 _20832_ (.Y(_04479_),
    .A(_08345_),
    .B(_04478_));
 sg13g2_o21ai_1 _20833_ (.B1(_04479_),
    .Y(_04480_),
    .A1(_08345_),
    .A2(_04477_));
 sg13g2_nand2_1 _20834_ (.Y(_04481_),
    .A(net780),
    .B(_04480_));
 sg13g2_buf_1 _20835_ (.A(_08948_),
    .X(_04482_));
 sg13g2_buf_1 _20836_ (.A(net938),
    .X(_04483_));
 sg13g2_a22oi_1 _20837_ (.Y(_04484_),
    .B1(\top_ihp.wb_emem.cmd[38] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[37] ),
    .A1(net895));
 sg13g2_nand2_1 _20838_ (.Y(_02705_),
    .A(_04481_),
    .B(_04484_));
 sg13g2_buf_1 _20839_ (.A(net815),
    .X(_04485_));
 sg13g2_a22oi_1 _20840_ (.Y(_04486_),
    .B1(_08609_),
    .B2(_10655_),
    .A2(_08314_),
    .A1(net871));
 sg13g2_buf_1 _20841_ (.A(net938),
    .X(_04487_));
 sg13g2_a22oi_1 _20842_ (.Y(_04488_),
    .B1(\top_ihp.wb_emem.cmd[39] ),
    .B2(net782),
    .A2(\top_ihp.wb_emem.cmd[38] ),
    .A1(net894));
 sg13g2_o21ai_1 _20843_ (.B1(_04488_),
    .Y(_02706_),
    .A1(net779),
    .A2(_04486_));
 sg13g2_nand2_1 _20844_ (.Y(_04489_),
    .A(\top_ihp.wb_dati_ram[26] ),
    .B(net813));
 sg13g2_nand3_1 _20845_ (.B(net795),
    .C(net812),
    .A(_03789_),
    .Y(_04490_));
 sg13g2_a21oi_1 _20846_ (.A1(_04489_),
    .A2(_04490_),
    .Y(_04491_),
    .B1(net814));
 sg13g2_a21o_1 _20847_ (.A2(net781),
    .A1(\top_ihp.wb_dati_ram[27] ),
    .B1(_04491_),
    .X(_02707_));
 sg13g2_xnor2_1 _20848_ (.Y(_04492_),
    .A(_08351_),
    .B(_10667_));
 sg13g2_a21o_1 _20849_ (.A2(_04492_),
    .A1(net832),
    .B1(net934),
    .X(_04493_));
 sg13g2_nor3_1 _20850_ (.A(_08350_),
    .B(net762),
    .C(_04492_),
    .Y(_04494_));
 sg13g2_a21oi_1 _20851_ (.A1(_08350_),
    .A2(_04493_),
    .Y(_04495_),
    .B1(_04494_));
 sg13g2_a22oi_1 _20852_ (.Y(_04496_),
    .B1(\top_ihp.wb_emem.cmd[40] ),
    .B2(net782),
    .A2(\top_ihp.wb_emem.cmd[39] ),
    .A1(net894));
 sg13g2_o21ai_1 _20853_ (.B1(_04496_),
    .Y(_02708_),
    .A1(net779),
    .A2(_04495_));
 sg13g2_xnor2_1 _20854_ (.Y(_04497_),
    .A(_08354_),
    .B(_10680_));
 sg13g2_nand2_1 _20855_ (.Y(_04498_),
    .A(net796),
    .B(_04497_));
 sg13g2_o21ai_1 _20856_ (.B1(_09000_),
    .Y(_04499_),
    .A1(net798),
    .A2(_04497_));
 sg13g2_nand2_1 _20857_ (.Y(_04500_),
    .A(_08353_),
    .B(_04499_));
 sg13g2_o21ai_1 _20858_ (.B1(_04500_),
    .Y(_04501_),
    .A1(_08353_),
    .A2(_04498_));
 sg13g2_nand2_1 _20859_ (.Y(_04502_),
    .A(net780),
    .B(_04501_));
 sg13g2_a22oi_1 _20860_ (.Y(_04503_),
    .B1(\top_ihp.wb_emem.cmd[41] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[40] ),
    .A1(net895));
 sg13g2_nand2_1 _20861_ (.Y(_02709_),
    .A(_04502_),
    .B(_04503_));
 sg13g2_xnor2_1 _20862_ (.Y(_04504_),
    .A(_08263_),
    .B(_10001_));
 sg13g2_nand2_1 _20863_ (.Y(_04505_),
    .A(net796),
    .B(_04504_));
 sg13g2_o21ai_1 _20864_ (.B1(net982),
    .Y(_04506_),
    .A1(net798),
    .A2(_04504_));
 sg13g2_nand2_1 _20865_ (.Y(_04507_),
    .A(net1053),
    .B(_04506_));
 sg13g2_o21ai_1 _20866_ (.B1(_04507_),
    .Y(_04508_),
    .A1(net1053),
    .A2(_04505_));
 sg13g2_nand2_1 _20867_ (.Y(_04509_),
    .A(net780),
    .B(_04508_));
 sg13g2_a22oi_1 _20868_ (.Y(_04510_),
    .B1(\top_ihp.wb_emem.cmd[42] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[41] ),
    .A1(net895));
 sg13g2_nand2_1 _20869_ (.Y(_02710_),
    .A(_04509_),
    .B(_04510_));
 sg13g2_nand2_1 _20870_ (.Y(_04511_),
    .A(net796),
    .B(_10033_));
 sg13g2_o21ai_1 _20871_ (.B1(net982),
    .Y(_04512_),
    .A1(net798),
    .A2(_10033_));
 sg13g2_nand2_1 _20872_ (.Y(_04513_),
    .A(net1030),
    .B(_04512_));
 sg13g2_o21ai_1 _20873_ (.B1(_04513_),
    .Y(_04514_),
    .A1(net1030),
    .A2(_04511_));
 sg13g2_nand2_1 _20874_ (.Y(_04515_),
    .A(net780),
    .B(_04514_));
 sg13g2_a22oi_1 _20875_ (.Y(_04516_),
    .B1(\top_ihp.wb_emem.cmd[43] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[42] ),
    .A1(_04483_));
 sg13g2_nand2_1 _20876_ (.Y(_02711_),
    .A(_04515_),
    .B(_04516_));
 sg13g2_nand2_1 _20877_ (.Y(_04517_),
    .A(_03727_),
    .B(_08252_));
 sg13g2_o21ai_1 _20878_ (.B1(_04517_),
    .Y(_04518_),
    .A1(net762),
    .A2(_10084_));
 sg13g2_nand2_1 _20879_ (.Y(_04519_),
    .A(_04476_),
    .B(_04518_));
 sg13g2_a22oi_1 _20880_ (.Y(_04520_),
    .B1(\top_ihp.wb_emem.cmd[44] ),
    .B2(_04423_),
    .A2(\top_ihp.wb_emem.cmd[43] ),
    .A1(_04483_));
 sg13g2_nand2_1 _20881_ (.Y(_02712_),
    .A(_04519_),
    .B(_04520_));
 sg13g2_a22oi_1 _20882_ (.Y(_04521_),
    .B1(net796),
    .B2(_10114_),
    .A2(net1055),
    .A1(net871));
 sg13g2_a22oi_1 _20883_ (.Y(_04522_),
    .B1(\top_ihp.wb_emem.cmd[45] ),
    .B2(net782),
    .A2(\top_ihp.wb_emem.cmd[44] ),
    .A1(net894));
 sg13g2_o21ai_1 _20884_ (.B1(_04522_),
    .Y(_02713_),
    .A1(net779),
    .A2(_04521_));
 sg13g2_xnor2_1 _20885_ (.Y(_04523_),
    .A(_08452_),
    .B(_10147_));
 sg13g2_a21o_1 _20886_ (.A2(_04523_),
    .A1(_08418_),
    .B1(net934),
    .X(_04524_));
 sg13g2_nor3_1 _20887_ (.A(net1051),
    .B(net762),
    .C(_04523_),
    .Y(_04525_));
 sg13g2_a21oi_1 _20888_ (.A1(net1051),
    .A2(_04524_),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_a22oi_1 _20889_ (.Y(_04527_),
    .B1(\top_ihp.wb_emem.cmd[46] ),
    .B2(_04457_),
    .A2(\top_ihp.wb_emem.cmd[45] ),
    .A1(net894));
 sg13g2_o21ai_1 _20890_ (.B1(_04527_),
    .Y(_02714_),
    .A1(net779),
    .A2(_04526_));
 sg13g2_xnor2_1 _20891_ (.Y(_04528_),
    .A(_08279_),
    .B(_08487_));
 sg13g2_nor2_1 _20892_ (.A(_08287_),
    .B(net762),
    .Y(_04529_));
 sg13g2_o21ai_1 _20893_ (.B1(net982),
    .Y(_04530_),
    .A1(net798),
    .A2(_04528_));
 sg13g2_a22oi_1 _20894_ (.Y(_04531_),
    .B1(_04530_),
    .B2(_08287_),
    .A2(_04529_),
    .A1(_04528_));
 sg13g2_a22oi_1 _20895_ (.Y(_04532_),
    .B1(\top_ihp.wb_emem.cmd[47] ),
    .B2(net782),
    .A2(\top_ihp.wb_emem.cmd[46] ),
    .A1(net894));
 sg13g2_o21ai_1 _20896_ (.B1(_04532_),
    .Y(_02715_),
    .A1(net779),
    .A2(_04531_));
 sg13g2_a22oi_1 _20897_ (.Y(_04533_),
    .B1(net796),
    .B2(_10194_),
    .A2(_08282_),
    .A1(net871));
 sg13g2_nor2_1 _20898_ (.A(_04318_),
    .B(\top_ihp.wb_emem.cmd[47] ),
    .Y(_04534_));
 sg13g2_a221oi_1 _20899_ (.B2(net780),
    .C1(_04534_),
    .B1(_04533_),
    .A1(_00340_),
    .Y(_04535_),
    .A2(net811));
 sg13g2_inv_1 _20900_ (.Y(_02716_),
    .A(_04535_));
 sg13g2_a22oi_1 _20901_ (.Y(_04536_),
    .B1(_08609_),
    .B2(_10217_),
    .A2(net1052),
    .A1(net871));
 sg13g2_a22oi_1 _20902_ (.Y(_04537_),
    .B1(\top_ihp.wb_emem.cmd[49] ),
    .B2(net782),
    .A2(\top_ihp.wb_emem.cmd[48] ),
    .A1(net894));
 sg13g2_o21ai_1 _20903_ (.B1(_04537_),
    .Y(_02717_),
    .A1(net779),
    .A2(_04536_));
 sg13g2_nand2_1 _20904_ (.Y(_04538_),
    .A(\top_ihp.wb_dati_ram[27] ),
    .B(net813));
 sg13g2_nand3_1 _20905_ (.B(net795),
    .C(net812),
    .A(_03790_),
    .Y(_04539_));
 sg13g2_a21oi_1 _20906_ (.A1(_04538_),
    .A2(_04539_),
    .Y(_04540_),
    .B1(net814));
 sg13g2_a21o_1 _20907_ (.A2(net781),
    .A1(\top_ihp.wb_dati_ram[28] ),
    .B1(_04540_),
    .X(_02718_));
 sg13g2_xnor2_1 _20908_ (.Y(_04541_),
    .A(_08514_),
    .B(_10227_));
 sg13g2_o21ai_1 _20909_ (.B1(net982),
    .Y(_04542_),
    .A1(net762),
    .A2(_04541_));
 sg13g2_nand2_1 _20910_ (.Y(_04543_),
    .A(net1059),
    .B(_04542_));
 sg13g2_nand3_1 _20911_ (.B(_08548_),
    .C(_04541_),
    .A(_03771_),
    .Y(_04544_));
 sg13g2_nand2_1 _20912_ (.Y(_04545_),
    .A(_04543_),
    .B(_04544_));
 sg13g2_nand2_1 _20913_ (.Y(_04546_),
    .A(_04476_),
    .B(_04545_));
 sg13g2_a22oi_1 _20914_ (.Y(_04547_),
    .B1(\top_ihp.wb_emem.cmd[50] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[49] ),
    .A1(_04487_));
 sg13g2_nand2_1 _20915_ (.Y(_02719_),
    .A(_04546_),
    .B(_04547_));
 sg13g2_o21ai_1 _20916_ (.B1(_04364_),
    .Y(_04548_),
    .A1(_09000_),
    .A2(_08224_));
 sg13g2_o21ai_1 _20917_ (.B1(_08639_),
    .Y(_04549_),
    .A1(_08494_),
    .A2(_08647_));
 sg13g2_xnor2_1 _20918_ (.Y(_04550_),
    .A(_09677_),
    .B(_04549_));
 sg13g2_nor2_1 _20919_ (.A(net762),
    .B(_04550_),
    .Y(_04551_));
 sg13g2_inv_1 _20920_ (.Y(_04552_),
    .A(\top_ihp.wb_emem.cmd[50] ));
 sg13g2_a22oi_1 _20921_ (.Y(_04553_),
    .B1(_00341_),
    .B2(net782),
    .A2(_04552_),
    .A1(net894));
 sg13g2_o21ai_1 _20922_ (.B1(_04553_),
    .Y(_02720_),
    .A1(_04548_),
    .A2(_04551_));
 sg13g2_nand2_1 _20923_ (.Y(_04554_),
    .A(net871),
    .B(net1056));
 sg13g2_o21ai_1 _20924_ (.B1(_04554_),
    .Y(_04555_),
    .A1(_04472_),
    .A2(_10326_));
 sg13g2_inv_1 _20925_ (.Y(_04556_),
    .A(\top_ihp.wb_emem.cmd[51] ));
 sg13g2_a22oi_1 _20926_ (.Y(_04557_),
    .B1(_00342_),
    .B2(net818),
    .A2(_04556_),
    .A1(_04487_));
 sg13g2_o21ai_1 _20927_ (.B1(_04557_),
    .Y(_02721_),
    .A1(net779),
    .A2(_04555_));
 sg13g2_a22oi_1 _20928_ (.Y(_04558_),
    .B1(_08548_),
    .B2(_10346_),
    .A2(_08235_),
    .A1(net871));
 sg13g2_a22oi_1 _20929_ (.Y(_04559_),
    .B1(\top_ihp.wb_emem.cmd[53] ),
    .B2(net818),
    .A2(\top_ihp.wb_emem.cmd[52] ),
    .A1(_04482_));
 sg13g2_o21ai_1 _20930_ (.B1(_04559_),
    .Y(_02722_),
    .A1(net779),
    .A2(_04558_));
 sg13g2_xnor2_1 _20931_ (.Y(_04560_),
    .A(_08523_),
    .B(_08378_));
 sg13g2_nor2_1 _20932_ (.A(_08391_),
    .B(_04472_),
    .Y(_04561_));
 sg13g2_o21ai_1 _20933_ (.B1(net982),
    .Y(_04562_),
    .A1(net798),
    .A2(_04560_));
 sg13g2_a22oi_1 _20934_ (.Y(_04563_),
    .B1(_04562_),
    .B2(_08391_),
    .A2(_04561_),
    .A1(_04560_));
 sg13g2_a22oi_1 _20935_ (.Y(_04564_),
    .B1(\top_ihp.wb_emem.cmd[54] ),
    .B2(net818),
    .A2(\top_ihp.wb_emem.cmd[53] ),
    .A1(net938));
 sg13g2_o21ai_1 _20936_ (.B1(_04564_),
    .Y(_02723_),
    .A1(_04485_),
    .A2(_04563_));
 sg13g2_xnor2_1 _20937_ (.Y(_04565_),
    .A(_08395_),
    .B(_10382_));
 sg13g2_a21o_1 _20938_ (.A2(_04565_),
    .A1(net796),
    .B1(net871),
    .X(_04566_));
 sg13g2_nor3_1 _20939_ (.A(net1047),
    .B(net762),
    .C(_04565_),
    .Y(_04567_));
 sg13g2_a21o_1 _20940_ (.A2(_04566_),
    .A1(net1047),
    .B1(_04567_),
    .X(_04568_));
 sg13g2_inv_1 _20941_ (.Y(_04569_),
    .A(\top_ihp.wb_emem.cmd[54] ));
 sg13g2_a22oi_1 _20942_ (.Y(_04570_),
    .B1(_00343_),
    .B2(net818),
    .A2(_04569_),
    .A1(_04482_));
 sg13g2_o21ai_1 _20943_ (.B1(_04570_),
    .Y(_02724_),
    .A1(_04485_),
    .A2(_04568_));
 sg13g2_nor2_1 _20944_ (.A(net797),
    .B(net815),
    .Y(_04571_));
 sg13g2_a21oi_1 _20945_ (.A1(\top_ihp.wb_emem.cmd[55] ),
    .A2(net815),
    .Y(_04572_),
    .B1(_04571_));
 sg13g2_nand2_1 _20946_ (.Y(_04573_),
    .A(\top_ihp.wb_emem.cmd[56] ),
    .B(net782));
 sg13g2_o21ai_1 _20947_ (.B1(_04573_),
    .Y(_02725_),
    .A1(net789),
    .A2(_04572_));
 sg13g2_inv_1 _20948_ (.Y(_04574_),
    .A(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_a22oi_1 _20949_ (.Y(_04575_),
    .B1(_00344_),
    .B2(net781),
    .A2(_04574_),
    .A1(net895));
 sg13g2_inv_1 _20950_ (.Y(_02726_),
    .A(_04575_));
 sg13g2_inv_1 _20951_ (.Y(_04576_),
    .A(\top_ihp.wb_emem.cmd[57] ));
 sg13g2_a221oi_1 _20952_ (.B2(net811),
    .C1(net780),
    .B1(_00345_),
    .A1(net938),
    .Y(_04577_),
    .A2(_04576_));
 sg13g2_inv_1 _20953_ (.Y(_02727_),
    .A(_04577_));
 sg13g2_a22oi_1 _20954_ (.Y(_04578_),
    .B1(\top_ihp.wb_emem.cmd[59] ),
    .B2(net781),
    .A2(\top_ihp.wb_emem.cmd[58] ),
    .A1(net895));
 sg13g2_inv_1 _20955_ (.Y(_02728_),
    .A(_04578_));
 sg13g2_nand2_1 _20956_ (.Y(_04579_),
    .A(\top_ihp.wb_dati_ram[28] ),
    .B(net813));
 sg13g2_nand3_1 _20957_ (.B(net795),
    .C(net812),
    .A(_03792_),
    .Y(_04580_));
 sg13g2_a21oi_1 _20958_ (.A1(_04579_),
    .A2(_04580_),
    .Y(_04581_),
    .B1(_04467_));
 sg13g2_a21o_1 _20959_ (.A2(net781),
    .A1(\top_ihp.wb_dati_ram[29] ),
    .B1(_04581_),
    .X(_02729_));
 sg13g2_a22oi_1 _20960_ (.Y(_04582_),
    .B1(\top_ihp.wb_emem.cmd[60] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[59] ),
    .A1(net895));
 sg13g2_inv_1 _20961_ (.Y(_02730_),
    .A(_04582_));
 sg13g2_inv_1 _20962_ (.Y(_04583_),
    .A(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_a221oi_1 _20963_ (.B2(net811),
    .C1(net780),
    .B1(_00346_),
    .A1(net938),
    .Y(_04584_),
    .A2(_04583_));
 sg13g2_inv_1 _20964_ (.Y(_02731_),
    .A(_04584_));
 sg13g2_inv_1 _20965_ (.Y(_04585_),
    .A(\top_ihp.wb_emem.cmd[61] ));
 sg13g2_a221oi_1 _20966_ (.B2(net811),
    .C1(net780),
    .B1(_00347_),
    .A1(net938),
    .Y(_04586_),
    .A2(_04585_));
 sg13g2_inv_1 _20967_ (.Y(_02732_),
    .A(_04586_));
 sg13g2_a22oi_1 _20968_ (.Y(_04587_),
    .B1(\top_ihp.wb_emem.cmd[63] ),
    .B2(net783),
    .A2(\top_ihp.wb_emem.cmd[62] ),
    .A1(net895));
 sg13g2_inv_1 _20969_ (.Y(_02733_),
    .A(_04587_));
 sg13g2_nand2_1 _20970_ (.Y(_04588_),
    .A(\top_ihp.wb_dati_ram[29] ),
    .B(net813));
 sg13g2_nand3_1 _20971_ (.B(_08581_),
    .C(net812),
    .A(_03795_),
    .Y(_04589_));
 sg13g2_a21oi_1 _20972_ (.A1(_04588_),
    .A2(_04589_),
    .Y(_04590_),
    .B1(net811));
 sg13g2_a21o_1 _20973_ (.A2(_04469_),
    .A1(\top_ihp.wb_dati_ram[30] ),
    .B1(_04590_),
    .X(_02734_));
 sg13g2_nand2_1 _20974_ (.Y(_04591_),
    .A(\top_ihp.wb_dati_ram[30] ),
    .B(net844));
 sg13g2_nand3_1 _20975_ (.B(_08581_),
    .C(net843),
    .A(_03797_),
    .Y(_04592_));
 sg13g2_a21oi_1 _20976_ (.A1(_04591_),
    .A2(_04592_),
    .Y(_04593_),
    .B1(_04467_));
 sg13g2_a21o_1 _20977_ (.A2(_04469_),
    .A1(\top_ihp.wb_dati_ram[31] ),
    .B1(_04593_),
    .X(_02735_));
 sg13g2_nand2_1 _20978_ (.Y(_04594_),
    .A(\top_ihp.wb_dati_ram[31] ),
    .B(net844));
 sg13g2_nand3_1 _20979_ (.B(net795),
    .C(net843),
    .A(_03768_),
    .Y(_04595_));
 sg13g2_a21oi_1 _20980_ (.A1(_04594_),
    .A2(_04595_),
    .Y(_04596_),
    .B1(net811));
 sg13g2_a21o_1 _20981_ (.A2(net781),
    .A1(\top_ihp.wb_dati_ram[16] ),
    .B1(_04596_),
    .X(_02736_));
 sg13g2_nand2_1 _20982_ (.Y(_04597_),
    .A(\top_ihp.wb_dati_ram[16] ),
    .B(net844));
 sg13g2_nand3_1 _20983_ (.B(net795),
    .C(net843),
    .A(_03770_),
    .Y(_04598_));
 sg13g2_a21oi_1 _20984_ (.A1(_04597_),
    .A2(_04598_),
    .Y(_04599_),
    .B1(net811));
 sg13g2_a21o_1 _20985_ (.A2(net781),
    .A1(\top_ihp.wb_dati_ram[17] ),
    .B1(_04599_),
    .X(_02737_));
 sg13g2_buf_1 _20986_ (.A(\top_ihp.wb_emem.nbits[3] ),
    .X(_04600_));
 sg13g2_xnor2_1 _20987_ (.Y(_04601_),
    .A(_04341_),
    .B(\top_ihp.wb_emem.nbits[5] ));
 sg13g2_buf_1 _20988_ (.A(\top_ihp.wb_emem.nbits[4] ),
    .X(_04602_));
 sg13g2_nor2b_1 _20989_ (.A(_04335_),
    .B_N(_04602_),
    .Y(_04603_));
 sg13g2_nor2_1 _20990_ (.A(_04602_),
    .B(_04601_),
    .Y(_04604_));
 sg13g2_a22oi_1 _20991_ (.Y(_04605_),
    .B1(_04604_),
    .B2(_04335_),
    .A2(_04603_),
    .A1(_04601_));
 sg13g2_nor2_1 _20992_ (.A(_04600_),
    .B(_04605_),
    .Y(_04606_));
 sg13g2_xnor2_1 _20993_ (.Y(_04607_),
    .A(_04335_),
    .B(_04602_));
 sg13g2_nand3_1 _20994_ (.B(_04601_),
    .C(_04607_),
    .A(_04600_),
    .Y(_04608_));
 sg13g2_nor2_1 _20995_ (.A(_04331_),
    .B(_04608_),
    .Y(_04609_));
 sg13g2_a21oi_1 _20996_ (.A1(_04331_),
    .A2(_04606_),
    .Y(_04610_),
    .B1(_04609_));
 sg13g2_nor3_1 _20997_ (.A(_04600_),
    .B(_04602_),
    .C(\top_ihp.wb_emem.nbits[5] ),
    .Y(_04611_));
 sg13g2_nor2b_1 _20998_ (.A(_04611_),
    .B_N(\top_ihp.wb_emem.nbits[6] ),
    .Y(_04612_));
 sg13g2_nor2b_1 _20999_ (.A(\top_ihp.wb_emem.nbits[6] ),
    .B_N(_04611_),
    .Y(_04613_));
 sg13g2_nor3_1 _21000_ (.A(_04347_),
    .B(_04612_),
    .C(_04613_),
    .Y(_04614_));
 sg13g2_a21oi_1 _21001_ (.A1(_04347_),
    .A2(_04612_),
    .Y(_04615_),
    .B1(_04614_));
 sg13g2_nor4_1 _21002_ (.A(\top_ihp.wb_emem.bit_counter[7] ),
    .B(_04333_),
    .C(_04610_),
    .D(_04615_),
    .Y(_04616_));
 sg13g2_a21o_1 _21003_ (.A2(_04326_),
    .A1(net1021),
    .B1(_04616_),
    .X(_02738_));
 sg13g2_buf_2 _21004_ (.A(\top_ihp.wb_emem.last_wait ),
    .X(_04617_));
 sg13g2_inv_1 _21005_ (.Y(_04618_),
    .A(_04617_));
 sg13g2_xor2_1 _21006_ (.B(_08953_),
    .A(_08952_),
    .X(_04619_));
 sg13g2_and2_2 _21007_ (.A(net879),
    .B(_04619_),
    .X(_04620_));
 sg13g2_buf_2 _21008_ (.A(_04620_),
    .X(_04621_));
 sg13g2_inv_1 _21009_ (.Y(_04622_),
    .A(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_buf_1 _21010_ (.A(\top_ihp.wb_emem.wait_counter[1] ),
    .X(_04623_));
 sg13g2_buf_1 _21011_ (.A(\top_ihp.wb_emem.wait_counter[0] ),
    .X(_04624_));
 sg13g2_nand3_1 _21012_ (.B(_04624_),
    .C(\top_ihp.wb_emem.wait_counter[2] ),
    .A(_04623_),
    .Y(_04625_));
 sg13g2_nor2_1 _21013_ (.A(_04622_),
    .B(_04625_),
    .Y(_04626_));
 sg13g2_buf_1 _21014_ (.A(\top_ihp.wb_emem.wait_counter[5] ),
    .X(_04627_));
 sg13g2_buf_1 _21015_ (.A(\top_ihp.wb_emem.wait_counter[4] ),
    .X(_04628_));
 sg13g2_buf_1 _21016_ (.A(\top_ihp.wb_emem.wait_counter[6] ),
    .X(_04629_));
 sg13g2_nor4_1 _21017_ (.A(_04627_),
    .B(_04628_),
    .C(\top_ihp.wb_emem.wait_counter[7] ),
    .D(_04629_),
    .Y(_04630_));
 sg13g2_nand3_1 _21018_ (.B(_04630_),
    .C(_04621_),
    .A(_04626_),
    .Y(_04631_));
 sg13g2_o21ai_1 _21019_ (.B1(_04631_),
    .Y(_02739_),
    .A1(_04618_),
    .A2(_04621_));
 sg13g2_inv_1 _21020_ (.Y(_04632_),
    .A(_04600_));
 sg13g2_nand2b_1 _21021_ (.Y(_04633_),
    .B(_08953_),
    .A_N(net1022));
 sg13g2_nand3_1 _21022_ (.B(_09818_),
    .C(_04633_),
    .A(_09663_),
    .Y(_04634_));
 sg13g2_buf_1 _21023_ (.A(_04634_),
    .X(_04635_));
 sg13g2_and2_1 _21024_ (.A(_09663_),
    .B(net843),
    .X(_04636_));
 sg13g2_buf_1 _21025_ (.A(_04636_),
    .X(_04637_));
 sg13g2_nand3_1 _21026_ (.B(net797),
    .C(_09807_),
    .A(_08659_),
    .Y(_04638_));
 sg13g2_a22oi_1 _21027_ (.Y(_02740_),
    .B1(_04637_),
    .B2(_04638_),
    .A2(_04635_),
    .A1(_04632_));
 sg13g2_o21ai_1 _21028_ (.B1(_08615_),
    .Y(_04639_),
    .A1(_08414_),
    .A2(_08416_));
 sg13g2_nor2_1 _21029_ (.A(net951),
    .B(_08660_),
    .Y(_04640_));
 sg13g2_and3_1 _21030_ (.X(_04641_),
    .A(net999),
    .B(_04639_),
    .C(_04640_));
 sg13g2_buf_1 _21031_ (.A(_04641_),
    .X(_04642_));
 sg13g2_buf_1 _21032_ (.A(net778),
    .X(_04643_));
 sg13g2_nand3_1 _21033_ (.B(_04637_),
    .C(_04643_),
    .A(net797),
    .Y(_04644_));
 sg13g2_nand2_1 _21034_ (.Y(_04645_),
    .A(_04602_),
    .B(_04635_));
 sg13g2_nand2_1 _21035_ (.Y(_02741_),
    .A(_04644_),
    .B(_04645_));
 sg13g2_nand3_1 _21036_ (.B(_04637_),
    .C(_04640_),
    .A(net797),
    .Y(_04646_));
 sg13g2_nand2_1 _21037_ (.Y(_04647_),
    .A(\top_ihp.wb_emem.nbits[5] ),
    .B(_04635_));
 sg13g2_nand2_1 _21038_ (.Y(_02742_),
    .A(_04646_),
    .B(_04647_));
 sg13g2_nand2_1 _21039_ (.Y(_04648_),
    .A(net797),
    .B(_04640_));
 sg13g2_and2_1 _21040_ (.A(\top_ihp.wb_emem.nbits[6] ),
    .B(_04635_),
    .X(_04649_));
 sg13g2_a21o_1 _21041_ (.A2(_04648_),
    .A1(_04637_),
    .B1(_04649_),
    .X(_02743_));
 sg13g2_inv_1 _21042_ (.Y(_04650_),
    .A(_04633_));
 sg13g2_nor2_1 _21043_ (.A(_08949_),
    .B(_04617_),
    .Y(_04651_));
 sg13g2_nand3_1 _21044_ (.B(_10523_),
    .C(_10525_),
    .A(net832),
    .Y(_04652_));
 sg13g2_a21oi_1 _21045_ (.A1(net934),
    .A2(_09673_),
    .Y(_04653_),
    .B1(net844));
 sg13g2_a21oi_1 _21046_ (.A1(net1023),
    .A2(net1021),
    .Y(_04654_),
    .B1(net896));
 sg13g2_a221oi_1 _21047_ (.B2(_04653_),
    .C1(_04654_),
    .B1(_04652_),
    .A1(_04650_),
    .Y(_04655_),
    .A2(_04651_));
 sg13g2_buf_1 _21048_ (.A(_04655_),
    .X(_04656_));
 sg13g2_inv_1 _21049_ (.Y(_04657_),
    .A(_08953_));
 sg13g2_nor2_1 _21050_ (.A(_08948_),
    .B(_04319_),
    .Y(_04658_));
 sg13g2_nand2_1 _21051_ (.Y(_04659_),
    .A(_04657_),
    .B(_04658_));
 sg13g2_o21ai_1 _21052_ (.B1(_04659_),
    .Y(_04660_),
    .A1(_04657_),
    .A2(net1023));
 sg13g2_and3_1 _21053_ (.X(_04661_),
    .A(net938),
    .B(_04319_),
    .C(_04617_));
 sg13g2_a21o_1 _21054_ (.A2(_04660_),
    .A1(net1022),
    .B1(_04661_),
    .X(_04662_));
 sg13g2_a21o_1 _21055_ (.A2(_04617_),
    .A1(_08953_),
    .B1(net1023),
    .X(_04663_));
 sg13g2_a21oi_1 _21056_ (.A1(net896),
    .A2(_04663_),
    .Y(_04664_),
    .B1(net1022));
 sg13g2_a21oi_1 _21057_ (.A1(_04656_),
    .A2(_04662_),
    .Y(_02744_),
    .B1(_04664_));
 sg13g2_a21o_1 _21058_ (.A2(_04658_),
    .A1(net1022),
    .B1(_08953_),
    .X(_02745_));
 sg13g2_nand2b_1 _21059_ (.Y(_04665_),
    .B(net1022),
    .A_N(_04617_));
 sg13g2_o21ai_1 _21060_ (.B1(net1023),
    .Y(_04666_),
    .A1(net896),
    .A2(net1021));
 sg13g2_o21ai_1 _21061_ (.B1(_04666_),
    .Y(_04667_),
    .A1(net938),
    .A2(_04665_));
 sg13g2_a21oi_1 _21062_ (.A1(_04319_),
    .A2(_04656_),
    .Y(_04668_),
    .B1(net894));
 sg13g2_a221oi_1 _21063_ (.B2(_04657_),
    .C1(_04668_),
    .B1(_04667_),
    .A1(_04650_),
    .Y(_02746_),
    .A2(_04656_));
 sg13g2_a21oi_1 _21064_ (.A1(net1022),
    .A2(_04651_),
    .Y(_04669_),
    .B1(_04658_));
 sg13g2_nand2_1 _21065_ (.Y(_04670_),
    .A(net896),
    .B(_04650_));
 sg13g2_mux2_1 _21066_ (.A0(_08949_),
    .A1(_04670_),
    .S(_04656_),
    .X(_04671_));
 sg13g2_o21ai_1 _21067_ (.B1(_04671_),
    .Y(_04672_),
    .A1(_08953_),
    .A2(_04669_));
 sg13g2_inv_1 _21068_ (.Y(_02747_),
    .A(_04672_));
 sg13g2_inv_1 _21069_ (.Y(_04673_),
    .A(_00265_));
 sg13g2_nand2_2 _21070_ (.Y(_04674_),
    .A(_09818_),
    .B(_04619_));
 sg13g2_buf_1 _21071_ (.A(_04674_),
    .X(_04675_));
 sg13g2_nand2b_2 _21072_ (.Y(_04676_),
    .B(_04657_),
    .A_N(_04312_));
 sg13g2_buf_1 _21073_ (.A(_04676_),
    .X(_04677_));
 sg13g2_nand3_1 _21074_ (.B(_04675_),
    .C(_04677_),
    .A(_04624_),
    .Y(_04678_));
 sg13g2_o21ai_1 _21075_ (.B1(_04678_),
    .Y(_02748_),
    .A1(_04673_),
    .A2(net842));
 sg13g2_nand2_1 _21076_ (.Y(_04679_),
    .A(_04624_),
    .B(_04621_));
 sg13g2_and2_1 _21077_ (.A(net842),
    .B(_04677_),
    .X(_04680_));
 sg13g2_buf_1 _21078_ (.A(_04680_),
    .X(_04681_));
 sg13g2_nor2_1 _21079_ (.A(_04624_),
    .B(net842),
    .Y(_04682_));
 sg13g2_o21ai_1 _21080_ (.B1(_04623_),
    .Y(_04683_),
    .A1(_04681_),
    .A2(_04682_));
 sg13g2_o21ai_1 _21081_ (.B1(_04683_),
    .Y(_02749_),
    .A1(_04623_),
    .A2(_04679_));
 sg13g2_nand3_1 _21082_ (.B(_04624_),
    .C(_04621_),
    .A(_04623_),
    .Y(_04684_));
 sg13g2_a21oi_1 _21083_ (.A1(_04623_),
    .A2(_04624_),
    .Y(_04685_),
    .B1(net842));
 sg13g2_o21ai_1 _21084_ (.B1(\top_ihp.wb_emem.wait_counter[2] ),
    .Y(_04686_),
    .A1(_04681_),
    .A2(_04685_));
 sg13g2_o21ai_1 _21085_ (.B1(_04686_),
    .Y(_02750_),
    .A1(\top_ihp.wb_emem.wait_counter[2] ),
    .A2(_04684_));
 sg13g2_xnor2_1 _21086_ (.Y(_04687_),
    .A(_04622_),
    .B(_04625_));
 sg13g2_nand3_1 _21087_ (.B(_04675_),
    .C(_04677_),
    .A(\top_ihp.wb_emem.wait_counter[3] ),
    .Y(_04688_));
 sg13g2_o21ai_1 _21088_ (.B1(_04688_),
    .Y(_02751_),
    .A1(net842),
    .A2(_04687_));
 sg13g2_nand2_1 _21089_ (.Y(_04689_),
    .A(_04626_),
    .B(_04621_));
 sg13g2_nor2_1 _21090_ (.A(_04626_),
    .B(net842),
    .Y(_04690_));
 sg13g2_o21ai_1 _21091_ (.B1(_04628_),
    .Y(_04691_),
    .A1(_04681_),
    .A2(_04690_));
 sg13g2_o21ai_1 _21092_ (.B1(_04691_),
    .Y(_02752_),
    .A1(_04628_),
    .A2(_04689_));
 sg13g2_and2_1 _21093_ (.A(_04628_),
    .B(_04626_),
    .X(_04692_));
 sg13g2_buf_1 _21094_ (.A(_04692_),
    .X(_04693_));
 sg13g2_nand2_1 _21095_ (.Y(_04694_),
    .A(_04621_),
    .B(_04693_));
 sg13g2_nor2_1 _21096_ (.A(net842),
    .B(_04693_),
    .Y(_04695_));
 sg13g2_o21ai_1 _21097_ (.B1(_04627_),
    .Y(_04696_),
    .A1(_04681_),
    .A2(_04695_));
 sg13g2_o21ai_1 _21098_ (.B1(_04696_),
    .Y(_02753_),
    .A1(_04627_),
    .A2(_04694_));
 sg13g2_nand3_1 _21099_ (.B(_04621_),
    .C(_04693_),
    .A(_04627_),
    .Y(_04697_));
 sg13g2_a21oi_1 _21100_ (.A1(_04627_),
    .A2(_04693_),
    .Y(_04698_),
    .B1(net842));
 sg13g2_o21ai_1 _21101_ (.B1(_04629_),
    .Y(_04699_),
    .A1(_04681_),
    .A2(_04698_));
 sg13g2_o21ai_1 _21102_ (.B1(_04699_),
    .Y(_02754_),
    .A1(_04629_),
    .A2(_04697_));
 sg13g2_nand2_1 _21103_ (.Y(_04700_),
    .A(\top_ihp.wb_emem.wait_counter[7] ),
    .B(_04677_));
 sg13g2_nand4_1 _21104_ (.B(_04629_),
    .C(_04621_),
    .A(_04627_),
    .Y(_04701_),
    .D(_04693_));
 sg13g2_mux2_1 _21105_ (.A0(\top_ihp.wb_emem.wait_counter[7] ),
    .A1(_04700_),
    .S(_04701_),
    .X(_04702_));
 sg13g2_inv_1 _21106_ (.Y(_02755_),
    .A(_04702_));
 sg13g2_mux4_1 _21107_ (.S0(\top_ihp.oisc.wb_adr_o[0] ),
    .A0(net6),
    .A1(net7),
    .A2(net8),
    .A3(net9),
    .S1(\top_ihp.oisc.wb_adr_o[1] ),
    .X(_04703_));
 sg13g2_nand3b_1 _21108_ (.B(_08543_),
    .C(_08213_),
    .Y(_04704_),
    .A_N(_08542_));
 sg13g2_mux2_1 _21109_ (.A0(_04703_),
    .A1(\top_ihp.wb_dati_gpio[0] ),
    .S(_04704_),
    .X(_02756_));
 sg13g2_nand2_1 _21110_ (.Y(_04705_),
    .A(_08543_),
    .B(_08440_));
 sg13g2_nor3_1 _21111_ (.A(_08542_),
    .B(_03813_),
    .C(_04705_),
    .Y(_04706_));
 sg13g2_mux2_1 _21112_ (.A0(\top_ihp.gpio_o_1 ),
    .A1(net1034),
    .S(_04706_),
    .X(_02757_));
 sg13g2_nand2_1 _21113_ (.Y(_04707_),
    .A(_08611_),
    .B(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_mux2_1 _21114_ (.A0(net1034),
    .A1(\top_ihp.gpio_o_2 ),
    .S(_04707_),
    .X(_04708_));
 sg13g2_inv_1 _21115_ (.Y(_04709_),
    .A(_04708_));
 sg13g2_nor2_1 _21116_ (.A(_08542_),
    .B(_04705_),
    .Y(_04710_));
 sg13g2_mux2_1 _21117_ (.A0(_00348_),
    .A1(_04709_),
    .S(_04710_),
    .X(_02758_));
 sg13g2_inv_1 _21118_ (.Y(_04711_),
    .A(_00222_));
 sg13g2_nor4_1 _21119_ (.A(_08542_),
    .B(_08611_),
    .C(\top_ihp.oisc.wb_adr_o[0] ),
    .D(_04705_),
    .Y(_04712_));
 sg13g2_mux2_1 _21120_ (.A0(\top_ihp.gpio_o_3 ),
    .A1(_04711_),
    .S(_04712_),
    .X(_02759_));
 sg13g2_nand2_1 _21121_ (.Y(_04713_),
    .A(\top_ihp.oisc.wb_adr_o[1] ),
    .B(\top_ihp.oisc.wb_adr_o[0] ));
 sg13g2_mux2_1 _21122_ (.A0(net1034),
    .A1(\top_ihp.gpio_o_4 ),
    .S(_04713_),
    .X(_04714_));
 sg13g2_inv_1 _21123_ (.Y(_04715_),
    .A(_04714_));
 sg13g2_mux2_1 _21124_ (.A0(_00349_),
    .A1(_04715_),
    .S(_04710_),
    .X(_02760_));
 sg13g2_nor3_1 _21125_ (.A(net1026),
    .B(_08439_),
    .C(_08613_),
    .Y(_04716_));
 sg13g2_nor3_1 _21126_ (.A(_09693_),
    .B(_08439_),
    .C(_08613_),
    .Y(_04717_));
 sg13g2_mux2_1 _21127_ (.A0(_04716_),
    .A1(_04717_),
    .S(_08578_),
    .X(_04718_));
 sg13g2_buf_1 _21128_ (.A(_04718_),
    .X(_04719_));
 sg13g2_o21ai_1 _21129_ (.B1(_08544_),
    .Y(_04720_),
    .A1(_08439_),
    .A2(_08547_));
 sg13g2_buf_1 _21130_ (.A(_04720_),
    .X(_04721_));
 sg13g2_or2_1 _21131_ (.X(_04722_),
    .B(_08589_),
    .A(net953));
 sg13g2_buf_1 _21132_ (.A(_04722_),
    .X(_04723_));
 sg13g2_o21ai_1 _21133_ (.B1(net866),
    .Y(_04724_),
    .A1(_04719_),
    .A2(_04721_));
 sg13g2_buf_1 _21134_ (.A(_04724_),
    .X(_04725_));
 sg13g2_nor2_1 _21135_ (.A(net953),
    .B(_08589_),
    .Y(_04726_));
 sg13g2_buf_1 _21136_ (.A(_04726_),
    .X(_04727_));
 sg13g2_nand2b_1 _21137_ (.Y(_04728_),
    .B(_04727_),
    .A_N(_08544_));
 sg13g2_o21ai_1 _21138_ (.B1(_04728_),
    .Y(_04729_),
    .A1(_04719_),
    .A2(_04721_));
 sg13g2_buf_1 _21139_ (.A(_04729_),
    .X(_04730_));
 sg13g2_buf_1 _21140_ (.A(_04730_),
    .X(_04731_));
 sg13g2_nand2_1 _21141_ (.Y(_04732_),
    .A(_08586_),
    .B(net619));
 sg13g2_o21ai_1 _21142_ (.B1(_04732_),
    .Y(_02761_),
    .A1(_08586_),
    .A2(net686));
 sg13g2_buf_1 _21143_ (.A(_04730_),
    .X(_04733_));
 sg13g2_buf_1 _21144_ (.A(net618),
    .X(_04734_));
 sg13g2_inv_1 _21145_ (.Y(_04735_),
    .A(_08591_));
 sg13g2_a21oi_1 _21146_ (.A1(net953),
    .A2(_04735_),
    .Y(_04736_),
    .B1(_08589_));
 sg13g2_nand2b_1 _21147_ (.Y(_04737_),
    .B(_08592_),
    .A_N(_04736_));
 sg13g2_nor2b_1 _21148_ (.A(_04736_),
    .B_N(_08586_),
    .Y(_04738_));
 sg13g2_o21ai_1 _21149_ (.B1(_08585_),
    .Y(_04739_),
    .A1(net618),
    .A2(_04738_));
 sg13g2_o21ai_1 _21150_ (.B1(_04739_),
    .Y(_02762_),
    .A1(net461),
    .A2(_04737_));
 sg13g2_o21ai_1 _21151_ (.B1(_08583_),
    .Y(_04740_),
    .A1(_08586_),
    .A2(_08585_));
 sg13g2_nor3_1 _21152_ (.A(_08586_),
    .B(_08585_),
    .C(_08583_),
    .Y(_04741_));
 sg13g2_nand2b_1 _21153_ (.Y(_04742_),
    .B(_04741_),
    .A_N(_04730_));
 sg13g2_a21o_1 _21154_ (.A2(_08596_),
    .A1(_08591_),
    .B1(_04736_),
    .X(_04743_));
 sg13g2_buf_1 _21155_ (.A(_04743_),
    .X(_04744_));
 sg13g2_a21oi_1 _21156_ (.A1(_04740_),
    .A2(_04742_),
    .Y(_04745_),
    .B1(_04744_));
 sg13g2_a21o_1 _21157_ (.A2(net619),
    .A1(_08583_),
    .B1(_04745_),
    .X(_02763_));
 sg13g2_nor2_1 _21158_ (.A(_04719_),
    .B(_04721_),
    .Y(_04746_));
 sg13g2_nor2b_1 _21159_ (.A(_04746_),
    .B_N(_04728_),
    .Y(_04747_));
 sg13g2_buf_2 _21160_ (.A(_04747_),
    .X(_04748_));
 sg13g2_o21ai_1 _21161_ (.B1(_04748_),
    .Y(_04749_),
    .A1(_04744_),
    .A2(_04741_));
 sg13g2_nor2b_1 _21162_ (.A(\top_ihp.wb_imem.bits_left[3] ),
    .B_N(_04741_),
    .Y(_04750_));
 sg13g2_nand2b_1 _21163_ (.Y(_04751_),
    .B(_04750_),
    .A_N(_04730_));
 sg13g2_nor2_1 _21164_ (.A(_04744_),
    .B(_04751_),
    .Y(_04752_));
 sg13g2_a21o_1 _21165_ (.A2(_04749_),
    .A1(\top_ihp.wb_imem.bits_left[3] ),
    .B1(_04752_),
    .X(_02764_));
 sg13g2_o21ai_1 _21166_ (.B1(_04748_),
    .Y(_04753_),
    .A1(_04744_),
    .A2(_04750_));
 sg13g2_mux2_1 _21167_ (.A0(_04752_),
    .A1(_04753_),
    .S(\top_ihp.wb_imem.bits_left[4] ),
    .X(_02765_));
 sg13g2_buf_1 _21168_ (.A(_04727_),
    .X(_04754_));
 sg13g2_nor2_1 _21169_ (.A(net862),
    .B(net857),
    .Y(_04755_));
 sg13g2_a21oi_1 _21170_ (.A1(_08597_),
    .A2(_04755_),
    .Y(_04756_),
    .B1(net618));
 sg13g2_o21ai_1 _21171_ (.B1(\top_ihp.wb_imem.bits_left[5] ),
    .Y(_04757_),
    .A1(\top_ihp.wb_imem.bits_left[4] ),
    .A2(_04751_));
 sg13g2_nand2b_1 _21172_ (.Y(_02766_),
    .B(_04757_),
    .A_N(_04756_));
 sg13g2_buf_1 _21173_ (.A(_04727_),
    .X(_04758_));
 sg13g2_a22oi_1 _21174_ (.Y(_04759_),
    .B1(\top_ihp.oisc.wb_adr_o[0] ),
    .B2(net856),
    .A2(net3),
    .A1(net953));
 sg13g2_nand2_1 _21175_ (.Y(_04760_),
    .A(\top_ihp.wb_dati_rom[24] ),
    .B(net619));
 sg13g2_o21ai_1 _21176_ (.B1(_04760_),
    .Y(_02767_),
    .A1(_04734_),
    .A2(_04759_));
 sg13g2_and2_1 _21177_ (.A(\top_ihp.wb_dati_rom[17] ),
    .B(net866),
    .X(_04761_));
 sg13g2_a21oi_1 _21178_ (.A1(_04508_),
    .A2(net856),
    .Y(_04762_),
    .B1(_04761_));
 sg13g2_nand2_1 _21179_ (.Y(_04763_),
    .A(\top_ihp.wb_dati_rom[18] ),
    .B(net619));
 sg13g2_o21ai_1 _21180_ (.B1(_04763_),
    .Y(_02768_),
    .A1(net461),
    .A2(_04762_));
 sg13g2_and2_1 _21181_ (.A(\top_ihp.wb_dati_rom[18] ),
    .B(net866),
    .X(_04764_));
 sg13g2_a21oi_1 _21182_ (.A1(_04514_),
    .A2(net856),
    .Y(_04765_),
    .B1(_04764_));
 sg13g2_nand2_1 _21183_ (.Y(_04766_),
    .A(\top_ihp.wb_dati_rom[19] ),
    .B(net619));
 sg13g2_o21ai_1 _21184_ (.B1(_04766_),
    .Y(_02769_),
    .A1(net461),
    .A2(_04765_));
 sg13g2_and2_1 _21185_ (.A(\top_ihp.wb_dati_rom[19] ),
    .B(net866),
    .X(_04767_));
 sg13g2_a21oi_1 _21186_ (.A1(_04518_),
    .A2(net856),
    .Y(_04768_),
    .B1(_04767_));
 sg13g2_buf_1 _21187_ (.A(_04730_),
    .X(_04769_));
 sg13g2_nand2_1 _21188_ (.Y(_04770_),
    .A(\top_ihp.wb_dati_rom[20] ),
    .B(net617));
 sg13g2_o21ai_1 _21189_ (.B1(_04770_),
    .Y(_02770_),
    .A1(net461),
    .A2(_04768_));
 sg13g2_buf_1 _21190_ (.A(_04723_),
    .X(_04771_));
 sg13g2_buf_1 _21191_ (.A(net866),
    .X(_04772_));
 sg13g2_nor2_1 _21192_ (.A(_04521_),
    .B(net854),
    .Y(_04773_));
 sg13g2_a21oi_1 _21193_ (.A1(\top_ihp.wb_dati_rom[20] ),
    .A2(net855),
    .Y(_04774_),
    .B1(_04773_));
 sg13g2_nand2_1 _21194_ (.Y(_04775_),
    .A(\top_ihp.wb_dati_rom[21] ),
    .B(net617));
 sg13g2_o21ai_1 _21195_ (.B1(_04775_),
    .Y(_02771_),
    .A1(net461),
    .A2(_04774_));
 sg13g2_nor2_1 _21196_ (.A(_04526_),
    .B(net854),
    .Y(_04776_));
 sg13g2_a21oi_1 _21197_ (.A1(\top_ihp.wb_dati_rom[21] ),
    .A2(net855),
    .Y(_04777_),
    .B1(_04776_));
 sg13g2_nand2_1 _21198_ (.Y(_04778_),
    .A(\top_ihp.wb_dati_rom[22] ),
    .B(net617));
 sg13g2_o21ai_1 _21199_ (.B1(_04778_),
    .Y(_02772_),
    .A1(net461),
    .A2(_04777_));
 sg13g2_nand2_1 _21200_ (.Y(_04779_),
    .A(_04531_),
    .B(_04754_));
 sg13g2_o21ai_1 _21201_ (.B1(_04779_),
    .Y(_04780_),
    .A1(\top_ihp.wb_dati_rom[22] ),
    .A2(_04754_));
 sg13g2_nand2_1 _21202_ (.Y(_04781_),
    .A(\top_ihp.wb_dati_rom[23] ),
    .B(net617));
 sg13g2_o21ai_1 _21203_ (.B1(_04781_),
    .Y(_02773_),
    .A1(net461),
    .A2(_04780_));
 sg13g2_buf_1 _21204_ (.A(net618),
    .X(_04782_));
 sg13g2_nor2_1 _21205_ (.A(_04533_),
    .B(net854),
    .Y(_04783_));
 sg13g2_a21oi_1 _21206_ (.A1(\top_ihp.wb_dati_rom[23] ),
    .A2(net855),
    .Y(_04784_),
    .B1(_04783_));
 sg13g2_nand2_1 _21207_ (.Y(_04785_),
    .A(\top_ihp.wb_dati_rom[8] ),
    .B(net617));
 sg13g2_o21ai_1 _21208_ (.B1(_04785_),
    .Y(_02774_),
    .A1(net460),
    .A2(_04784_));
 sg13g2_nand2_1 _21209_ (.Y(_04786_),
    .A(_04536_),
    .B(net857));
 sg13g2_o21ai_1 _21210_ (.B1(_04786_),
    .Y(_04787_),
    .A1(\top_ihp.wb_dati_rom[8] ),
    .A2(net857));
 sg13g2_nand2_1 _21211_ (.Y(_04788_),
    .A(\top_ihp.wb_dati_rom[9] ),
    .B(net617));
 sg13g2_o21ai_1 _21212_ (.B1(_04788_),
    .Y(_02775_),
    .A1(net460),
    .A2(_04787_));
 sg13g2_and2_1 _21213_ (.A(\top_ihp.wb_dati_rom[9] ),
    .B(net866),
    .X(_04789_));
 sg13g2_a21oi_1 _21214_ (.A1(_04545_),
    .A2(net856),
    .Y(_04790_),
    .B1(_04789_));
 sg13g2_nand2_1 _21215_ (.Y(_04791_),
    .A(\top_ihp.wb_dati_rom[10] ),
    .B(net617));
 sg13g2_o21ai_1 _21216_ (.B1(_04791_),
    .Y(_02776_),
    .A1(net460),
    .A2(_04790_));
 sg13g2_a21oi_1 _21217_ (.A1(net871),
    .A2(net1058),
    .Y(_04792_),
    .B1(_04551_));
 sg13g2_nor2_1 _21218_ (.A(\top_ihp.wb_dati_rom[10] ),
    .B(_04727_),
    .Y(_04793_));
 sg13g2_a21oi_1 _21219_ (.A1(net856),
    .A2(_04792_),
    .Y(_04794_),
    .B1(_04793_));
 sg13g2_mux2_1 _21220_ (.A0(\top_ihp.wb_dati_rom[11] ),
    .A1(_04794_),
    .S(_04748_),
    .X(_02777_));
 sg13g2_nor2_1 _21221_ (.A(_08611_),
    .B(net854),
    .Y(_04795_));
 sg13g2_a21oi_1 _21222_ (.A1(\top_ihp.wb_dati_rom[24] ),
    .A2(net855),
    .Y(_04796_),
    .B1(_04795_));
 sg13g2_nand2_1 _21223_ (.Y(_04797_),
    .A(\top_ihp.wb_dati_rom[25] ),
    .B(_04769_));
 sg13g2_o21ai_1 _21224_ (.B1(_04797_),
    .Y(_02778_),
    .A1(net460),
    .A2(_04796_));
 sg13g2_nand2b_1 _21225_ (.Y(_04798_),
    .B(net854),
    .A_N(\top_ihp.wb_dati_rom[11] ));
 sg13g2_o21ai_1 _21226_ (.B1(_04798_),
    .Y(_04799_),
    .A1(_04555_),
    .A2(net855));
 sg13g2_nand2_1 _21227_ (.Y(_04800_),
    .A(\top_ihp.wb_dati_rom[12] ),
    .B(net617));
 sg13g2_o21ai_1 _21228_ (.B1(_04800_),
    .Y(_02779_),
    .A1(_04782_),
    .A2(_04799_));
 sg13g2_nor2_1 _21229_ (.A(_04558_),
    .B(_04772_),
    .Y(_04801_));
 sg13g2_a21oi_1 _21230_ (.A1(\top_ihp.wb_dati_rom[12] ),
    .A2(_04771_),
    .Y(_04802_),
    .B1(_04801_));
 sg13g2_nand2_1 _21231_ (.Y(_04803_),
    .A(\top_ihp.wb_dati_rom[13] ),
    .B(_04769_));
 sg13g2_o21ai_1 _21232_ (.B1(_04803_),
    .Y(_02780_),
    .A1(_04782_),
    .A2(_04802_));
 sg13g2_inv_1 _21233_ (.Y(_04804_),
    .A(\top_ihp.wb_dati_rom[14] ));
 sg13g2_a21oi_1 _21234_ (.A1(_04563_),
    .A2(net857),
    .Y(_04805_),
    .B1(net618));
 sg13g2_o21ai_1 _21235_ (.B1(_04805_),
    .Y(_04806_),
    .A1(\top_ihp.wb_dati_rom[13] ),
    .A2(_04758_));
 sg13g2_o21ai_1 _21236_ (.B1(_04806_),
    .Y(_02781_),
    .A1(_04804_),
    .A2(_04748_));
 sg13g2_and2_1 _21237_ (.A(\top_ihp.wb_dati_rom[14] ),
    .B(_04723_),
    .X(_04807_));
 sg13g2_a21oi_1 _21238_ (.A1(_04568_),
    .A2(_04758_),
    .Y(_04808_),
    .B1(_04807_));
 sg13g2_buf_1 _21239_ (.A(_04730_),
    .X(_04809_));
 sg13g2_nand2_1 _21240_ (.Y(_04810_),
    .A(\top_ihp.wb_dati_rom[15] ),
    .B(_04809_));
 sg13g2_o21ai_1 _21241_ (.B1(_04810_),
    .Y(_02782_),
    .A1(net460),
    .A2(_04808_));
 sg13g2_inv_1 _21242_ (.Y(_04811_),
    .A(\top_ihp.wb_dati_rom[0] ));
 sg13g2_nor2_1 _21243_ (.A(\top_ihp.wb_dati_rom[15] ),
    .B(net686),
    .Y(_04812_));
 sg13g2_a21oi_1 _21244_ (.A1(_04811_),
    .A2(_04734_),
    .Y(_02783_),
    .B1(_04812_));
 sg13g2_inv_1 _21245_ (.Y(_04813_),
    .A(\top_ihp.wb_dati_rom[1] ));
 sg13g2_nor2_1 _21246_ (.A(\top_ihp.wb_dati_rom[0] ),
    .B(_04725_),
    .Y(_04814_));
 sg13g2_a21oi_1 _21247_ (.A1(_04813_),
    .A2(net461),
    .Y(_02784_),
    .B1(_04814_));
 sg13g2_nand2_1 _21248_ (.Y(_04815_),
    .A(\top_ihp.wb_dati_rom[2] ),
    .B(net616));
 sg13g2_o21ai_1 _21249_ (.B1(_04815_),
    .Y(_02785_),
    .A1(_04813_),
    .A2(net686));
 sg13g2_inv_1 _21250_ (.Y(_04816_),
    .A(\top_ihp.wb_dati_rom[2] ));
 sg13g2_nand2_1 _21251_ (.Y(_04817_),
    .A(\top_ihp.wb_dati_rom[3] ),
    .B(net616));
 sg13g2_o21ai_1 _21252_ (.B1(_04817_),
    .Y(_02786_),
    .A1(_04816_),
    .A2(net686));
 sg13g2_inv_1 _21253_ (.Y(_04818_),
    .A(\top_ihp.wb_dati_rom[3] ));
 sg13g2_nand2_1 _21254_ (.Y(_04819_),
    .A(\top_ihp.wb_dati_rom[4] ),
    .B(net616));
 sg13g2_o21ai_1 _21255_ (.B1(_04819_),
    .Y(_02787_),
    .A1(_04818_),
    .A2(net686));
 sg13g2_inv_1 _21256_ (.Y(_04820_),
    .A(\top_ihp.wb_dati_rom[4] ));
 sg13g2_nand2_1 _21257_ (.Y(_04821_),
    .A(\top_ihp.wb_dati_rom[5] ),
    .B(net616));
 sg13g2_o21ai_1 _21258_ (.B1(_04821_),
    .Y(_02788_),
    .A1(_04820_),
    .A2(net686));
 sg13g2_nor2_1 _21259_ (.A(_03810_),
    .B(_04772_),
    .Y(_04822_));
 sg13g2_a21oi_1 _21260_ (.A1(\top_ihp.wb_dati_rom[25] ),
    .A2(_04771_),
    .Y(_04823_),
    .B1(_04822_));
 sg13g2_nand2_1 _21261_ (.Y(_04824_),
    .A(\top_ihp.wb_dati_rom[26] ),
    .B(net616));
 sg13g2_o21ai_1 _21262_ (.B1(_04824_),
    .Y(_02789_),
    .A1(net460),
    .A2(_04823_));
 sg13g2_inv_1 _21263_ (.Y(_04825_),
    .A(\top_ihp.wb_dati_rom[5] ));
 sg13g2_nand2_1 _21264_ (.Y(_04826_),
    .A(\top_ihp.wb_dati_rom[6] ),
    .B(net616));
 sg13g2_o21ai_1 _21265_ (.B1(_04826_),
    .Y(_02790_),
    .A1(_04825_),
    .A2(net686));
 sg13g2_inv_1 _21266_ (.Y(_04827_),
    .A(\top_ihp.wb_dati_rom[6] ));
 sg13g2_nand2_1 _21267_ (.Y(_04828_),
    .A(\top_ihp.wb_dati_rom[7] ),
    .B(net616));
 sg13g2_o21ai_1 _21268_ (.B1(_04828_),
    .Y(_02791_),
    .A1(_04827_),
    .A2(net686));
 sg13g2_nand2_1 _21269_ (.Y(_04829_),
    .A(_03820_),
    .B(net857));
 sg13g2_o21ai_1 _21270_ (.B1(_04829_),
    .Y(_04830_),
    .A1(\top_ihp.wb_dati_rom[26] ),
    .A2(net857));
 sg13g2_nand2_1 _21271_ (.Y(_04831_),
    .A(\top_ihp.wb_dati_rom[27] ),
    .B(_04809_));
 sg13g2_o21ai_1 _21272_ (.B1(_04831_),
    .Y(_02792_),
    .A1(net460),
    .A2(_04830_));
 sg13g2_nor2_1 _21273_ (.A(_03895_),
    .B(net854),
    .Y(_04832_));
 sg13g2_a21oi_1 _21274_ (.A1(\top_ihp.wb_dati_rom[27] ),
    .A2(net855),
    .Y(_04833_),
    .B1(_04832_));
 sg13g2_nand2_1 _21275_ (.Y(_04834_),
    .A(\top_ihp.wb_dati_rom[28] ),
    .B(net616));
 sg13g2_o21ai_1 _21276_ (.B1(_04834_),
    .Y(_02793_),
    .A1(net460),
    .A2(_04833_));
 sg13g2_nor2_1 _21277_ (.A(_04474_),
    .B(net854),
    .Y(_04835_));
 sg13g2_a21oi_1 _21278_ (.A1(\top_ihp.wb_dati_rom[28] ),
    .A2(net855),
    .Y(_04836_),
    .B1(_04835_));
 sg13g2_nand2_1 _21279_ (.Y(_04837_),
    .A(\top_ihp.wb_dati_rom[29] ),
    .B(_04733_));
 sg13g2_o21ai_1 _21280_ (.B1(_04837_),
    .Y(_02794_),
    .A1(net619),
    .A2(_04836_));
 sg13g2_and2_1 _21281_ (.A(\top_ihp.wb_dati_rom[29] ),
    .B(net866),
    .X(_04838_));
 sg13g2_a21oi_1 _21282_ (.A1(_04480_),
    .A2(net856),
    .Y(_04839_),
    .B1(_04838_));
 sg13g2_nand2_1 _21283_ (.Y(_04840_),
    .A(\top_ihp.wb_dati_rom[30] ),
    .B(net618));
 sg13g2_o21ai_1 _21284_ (.B1(_04840_),
    .Y(_02795_),
    .A1(net619),
    .A2(_04839_));
 sg13g2_nor2_1 _21285_ (.A(_04486_),
    .B(net854),
    .Y(_04841_));
 sg13g2_a21oi_1 _21286_ (.A1(\top_ihp.wb_dati_rom[30] ),
    .A2(net855),
    .Y(_04842_),
    .B1(_04841_));
 sg13g2_nand2_1 _21287_ (.Y(_04843_),
    .A(\top_ihp.wb_dati_rom[31] ),
    .B(_04733_));
 sg13g2_o21ai_1 _21288_ (.B1(_04843_),
    .Y(_02796_),
    .A1(net619),
    .A2(_04842_));
 sg13g2_nand2_1 _21289_ (.Y(_04844_),
    .A(_04495_),
    .B(net857));
 sg13g2_o21ai_1 _21290_ (.B1(_04844_),
    .Y(_04845_),
    .A1(\top_ihp.wb_dati_rom[31] ),
    .A2(net857));
 sg13g2_nand2_1 _21291_ (.Y(_04846_),
    .A(\top_ihp.wb_dati_rom[16] ),
    .B(net618));
 sg13g2_o21ai_1 _21292_ (.B1(_04846_),
    .Y(_02797_),
    .A1(_04731_),
    .A2(_04845_));
 sg13g2_and2_1 _21293_ (.A(\top_ihp.wb_dati_rom[16] ),
    .B(net866),
    .X(_04847_));
 sg13g2_a21oi_1 _21294_ (.A1(_04501_),
    .A2(net856),
    .Y(_04848_),
    .B1(_04847_));
 sg13g2_nand2_1 _21295_ (.Y(_04849_),
    .A(\top_ihp.wb_dati_rom[17] ),
    .B(net618));
 sg13g2_o21ai_1 _21296_ (.B1(_04849_),
    .Y(_02798_),
    .A1(_04731_),
    .A2(_04848_));
 sg13g2_nor2b_1 _21297_ (.A(net862),
    .B_N(_00350_),
    .Y(_04850_));
 sg13g2_nand2_1 _21298_ (.Y(_04851_),
    .A(_08591_),
    .B(net862));
 sg13g2_nor2_1 _21299_ (.A(_04746_),
    .B(_04851_),
    .Y(_04852_));
 sg13g2_o21ai_1 _21300_ (.B1(net953),
    .Y(_04853_),
    .A1(_04850_),
    .A2(_04852_));
 sg13g2_inv_1 _21301_ (.Y(_04854_),
    .A(net953));
 sg13g2_nand4_1 _21302_ (.B(_08544_),
    .C(_08591_),
    .A(_04854_),
    .Y(_04855_),
    .D(_08582_));
 sg13g2_nor2_1 _21303_ (.A(net953),
    .B(_08544_),
    .Y(_04856_));
 sg13g2_o21ai_1 _21304_ (.B1(_00350_),
    .Y(_04857_),
    .A1(_04746_),
    .A2(_04856_));
 sg13g2_nand3_1 _21305_ (.B(_04855_),
    .C(_04857_),
    .A(_04853_),
    .Y(_02799_));
 sg13g2_nor3_1 _21306_ (.A(net1031),
    .B(_08213_),
    .C(_08613_),
    .Y(_04858_));
 sg13g2_and3_1 _21307_ (.X(_04859_),
    .A(net1031),
    .B(_08439_),
    .C(_08609_));
 sg13g2_mux2_1 _21308_ (.A0(_04858_),
    .A1(_04859_),
    .S(_08411_),
    .X(_04860_));
 sg13g2_nand2_1 _21309_ (.Y(_04861_),
    .A(net984),
    .B(net1031));
 sg13g2_o21ai_1 _21310_ (.B1(_00096_),
    .Y(_04862_),
    .A1(_08213_),
    .A2(_04861_));
 sg13g2_buf_1 _21311_ (.A(_08215_),
    .X(_04863_));
 sg13g2_nor3_1 _21312_ (.A(_08428_),
    .B(net937),
    .C(_08434_),
    .Y(_04864_));
 sg13g2_o21ai_1 _21313_ (.B1(_04864_),
    .Y(_04865_),
    .A1(_04860_),
    .A2(_04862_));
 sg13g2_nor2_2 _21314_ (.A(_04860_),
    .B(_04862_),
    .Y(_04866_));
 sg13g2_a21o_1 _21315_ (.A2(_08434_),
    .A1(_08214_),
    .B1(_04866_),
    .X(_04867_));
 sg13g2_buf_8 _21316_ (.A(_04867_),
    .X(_04868_));
 sg13g2_buf_8 _21317_ (.A(_04868_),
    .X(_04869_));
 sg13g2_nand2_1 _21318_ (.Y(_04870_),
    .A(_08428_),
    .B(net459));
 sg13g2_nand2_1 _21319_ (.Y(_02800_),
    .A(_04865_),
    .B(_04870_));
 sg13g2_nor2_1 _21320_ (.A(_08428_),
    .B(_08434_),
    .Y(_04871_));
 sg13g2_nor2_1 _21321_ (.A(net937),
    .B(_04871_),
    .Y(_04872_));
 sg13g2_o21ai_1 _21322_ (.B1(_08429_),
    .Y(_04873_),
    .A1(_04866_),
    .A2(_04872_));
 sg13g2_o21ai_1 _21323_ (.B1(_04873_),
    .Y(_02801_),
    .A1(_08429_),
    .A2(_04865_));
 sg13g2_buf_1 _21324_ (.A(_04868_),
    .X(_04874_));
 sg13g2_nor3_1 _21325_ (.A(_08428_),
    .B(_08429_),
    .C(\top_ihp.wb_spi.bits_left[2] ),
    .Y(_04875_));
 sg13g2_nand2_1 _21326_ (.Y(_04876_),
    .A(_08436_),
    .B(_04875_));
 sg13g2_buf_8 _21327_ (.A(_04868_),
    .X(_04877_));
 sg13g2_o21ai_1 _21328_ (.B1(_08214_),
    .Y(_04878_),
    .A1(_08428_),
    .A2(_08429_));
 sg13g2_inv_1 _21329_ (.Y(_04879_),
    .A(_04878_));
 sg13g2_o21ai_1 _21330_ (.B1(\top_ihp.wb_spi.bits_left[2] ),
    .Y(_04880_),
    .A1(_04877_),
    .A2(_04879_));
 sg13g2_o21ai_1 _21331_ (.B1(_04880_),
    .Y(_02802_),
    .A1(net458),
    .A2(_04876_));
 sg13g2_and3_1 _21332_ (.X(_04881_),
    .A(_08659_),
    .B(_09807_),
    .C(_04639_));
 sg13g2_buf_1 _21333_ (.A(_04881_),
    .X(_04882_));
 sg13g2_a21oi_1 _21334_ (.A1(_08428_),
    .A2(_08431_),
    .Y(_04883_),
    .B1(_08215_));
 sg13g2_nor2b_1 _21335_ (.A(\top_ihp.wb_spi.bits_left[3] ),
    .B_N(_04875_),
    .Y(_04884_));
 sg13g2_a22oi_1 _21336_ (.Y(_04885_),
    .B1(_04883_),
    .B2(_04884_),
    .A2(_04882_),
    .A1(net937));
 sg13g2_nor2b_1 _21337_ (.A(_04875_),
    .B_N(_04883_),
    .Y(_04886_));
 sg13g2_o21ai_1 _21338_ (.B1(\top_ihp.wb_spi.bits_left[3] ),
    .Y(_04887_),
    .A1(_04877_),
    .A2(_04886_));
 sg13g2_o21ai_1 _21339_ (.B1(_04887_),
    .Y(_02803_),
    .A1(net458),
    .A2(_04885_));
 sg13g2_nor2_1 _21340_ (.A(_08428_),
    .B(net937),
    .Y(_04888_));
 sg13g2_a22oi_1 _21341_ (.Y(_04889_),
    .B1(_04888_),
    .B2(_08430_),
    .A2(net761),
    .A1(_04863_));
 sg13g2_nor2b_1 _21342_ (.A(_08434_),
    .B_N(_04884_),
    .Y(_04890_));
 sg13g2_nor2_1 _21343_ (.A(net937),
    .B(_04890_),
    .Y(_04891_));
 sg13g2_o21ai_1 _21344_ (.B1(\top_ihp.wb_spi.bits_left[4] ),
    .Y(_04892_),
    .A1(_04866_),
    .A2(_04891_));
 sg13g2_o21ai_1 _21345_ (.B1(_04892_),
    .Y(_02804_),
    .A1(net458),
    .A2(_04889_));
 sg13g2_nand2_1 _21346_ (.Y(_04893_),
    .A(net950),
    .B(_08659_));
 sg13g2_o21ai_1 _21347_ (.B1(_04639_),
    .Y(_04894_),
    .A1(net999),
    .A2(_04893_));
 sg13g2_buf_1 _21348_ (.A(_04894_),
    .X(_04895_));
 sg13g2_buf_1 _21349_ (.A(_04895_),
    .X(_04896_));
 sg13g2_buf_1 _21350_ (.A(net760),
    .X(_04897_));
 sg13g2_a22oi_1 _21351_ (.Y(_04898_),
    .B1(net746),
    .B2(net937),
    .A2(_04864_),
    .A1(_08431_));
 sg13g2_a21oi_1 _21352_ (.A1(_08430_),
    .A2(_04871_),
    .Y(_04899_),
    .B1(net937));
 sg13g2_o21ai_1 _21353_ (.B1(\top_ihp.wb_spi.bits_left[5] ),
    .Y(_04900_),
    .A1(_04866_),
    .A2(_04899_));
 sg13g2_o21ai_1 _21354_ (.B1(_04900_),
    .Y(_02805_),
    .A1(_04866_),
    .A2(_04898_));
 sg13g2_buf_1 _21355_ (.A(_08214_),
    .X(_04901_));
 sg13g2_buf_1 _21356_ (.A(_08214_),
    .X(_04902_));
 sg13g2_nor2_1 _21357_ (.A(_04902_),
    .B(_00222_),
    .Y(_04903_));
 sg13g2_a22oi_1 _21358_ (.Y(_04904_),
    .B1(net746),
    .B2(_04903_),
    .A2(net5),
    .A1(net989));
 sg13g2_nand2_1 _21359_ (.Y(_04905_),
    .A(\top_ihp.wb_dati_spi[0] ),
    .B(net459));
 sg13g2_o21ai_1 _21360_ (.B1(_04905_),
    .Y(_02806_),
    .A1(net458),
    .A2(_04904_));
 sg13g2_buf_1 _21361_ (.A(_08214_),
    .X(_04906_));
 sg13g2_nor2b_1 _21362_ (.A(net987),
    .B_N(_03757_),
    .Y(_04907_));
 sg13g2_a22oi_1 _21363_ (.Y(_04908_),
    .B1(_04897_),
    .B2(_04907_),
    .A2(\top_ihp.wb_dati_spi[9] ),
    .A1(net989));
 sg13g2_nand2_1 _21364_ (.Y(_04909_),
    .A(\top_ihp.wb_dati_spi[10] ),
    .B(net459));
 sg13g2_o21ai_1 _21365_ (.B1(_04909_),
    .Y(_02807_),
    .A1(net458),
    .A2(_04908_));
 sg13g2_nor2b_1 _21366_ (.A(net987),
    .B_N(_03758_),
    .Y(_04910_));
 sg13g2_a22oi_1 _21367_ (.Y(_04911_),
    .B1(net746),
    .B2(_04910_),
    .A2(\top_ihp.wb_dati_spi[10] ),
    .A1(net989));
 sg13g2_nand2_1 _21368_ (.Y(_04912_),
    .A(\top_ihp.wb_dati_spi[11] ),
    .B(_04869_));
 sg13g2_o21ai_1 _21369_ (.B1(_04912_),
    .Y(_02808_),
    .A1(net458),
    .A2(_04911_));
 sg13g2_nor2b_1 _21370_ (.A(_04906_),
    .B_N(_03760_),
    .Y(_04913_));
 sg13g2_a22oi_1 _21371_ (.Y(_04914_),
    .B1(net746),
    .B2(_04913_),
    .A2(\top_ihp.wb_dati_spi[11] ),
    .A1(net989));
 sg13g2_nand2_1 _21372_ (.Y(_04915_),
    .A(\top_ihp.wb_dati_spi[12] ),
    .B(_04869_));
 sg13g2_o21ai_1 _21373_ (.B1(_04915_),
    .Y(_02809_),
    .A1(_04874_),
    .A2(_04914_));
 sg13g2_nor2b_1 _21374_ (.A(_04906_),
    .B_N(_03763_),
    .Y(_04916_));
 sg13g2_a22oi_1 _21375_ (.Y(_04917_),
    .B1(_04897_),
    .B2(_04916_),
    .A2(\top_ihp.wb_dati_spi[12] ),
    .A1(net989));
 sg13g2_buf_8 _21376_ (.A(_04868_),
    .X(_04918_));
 sg13g2_nand2_1 _21377_ (.Y(_04919_),
    .A(\top_ihp.wb_dati_spi[13] ),
    .B(net456));
 sg13g2_o21ai_1 _21378_ (.B1(_04919_),
    .Y(_02810_),
    .A1(_04874_),
    .A2(_04917_));
 sg13g2_buf_1 _21379_ (.A(_08214_),
    .X(_04920_));
 sg13g2_nor2b_1 _21380_ (.A(net986),
    .B_N(_03765_),
    .Y(_04921_));
 sg13g2_a22oi_1 _21381_ (.Y(_04922_),
    .B1(net746),
    .B2(_04921_),
    .A2(\top_ihp.wb_dati_spi[13] ),
    .A1(_04901_));
 sg13g2_nand2_1 _21382_ (.Y(_04923_),
    .A(\top_ihp.wb_dati_spi[14] ),
    .B(_04918_));
 sg13g2_o21ai_1 _21383_ (.B1(_04923_),
    .Y(_02811_),
    .A1(net458),
    .A2(_04922_));
 sg13g2_nor2b_1 _21384_ (.A(_04920_),
    .B_N(_03767_),
    .Y(_04924_));
 sg13g2_a22oi_1 _21385_ (.Y(_04925_),
    .B1(net746),
    .B2(_04924_),
    .A2(\top_ihp.wb_dati_spi[14] ),
    .A1(_04901_));
 sg13g2_nand2_1 _21386_ (.Y(_04926_),
    .A(\top_ihp.wb_dati_spi[15] ),
    .B(_04918_));
 sg13g2_o21ai_1 _21387_ (.B1(_04926_),
    .Y(_02812_),
    .A1(net458),
    .A2(_04925_));
 sg13g2_nor2_1 _21388_ (.A(net937),
    .B(\top_ihp.wb_dati_spi[15] ),
    .Y(_04927_));
 sg13g2_a221oi_1 _21389_ (.B2(_03768_),
    .C1(_08435_),
    .B1(_04896_),
    .A1(_04711_),
    .Y(_04928_),
    .A2(net761));
 sg13g2_nor3_1 _21390_ (.A(net457),
    .B(_04927_),
    .C(_04928_),
    .Y(_04929_));
 sg13g2_a21o_1 _21391_ (.A2(net459),
    .A1(\top_ihp.wb_dati_spi[16] ),
    .B1(_04929_),
    .X(_02813_));
 sg13g2_buf_1 _21392_ (.A(_04868_),
    .X(_04930_));
 sg13g2_inv_1 _21393_ (.Y(_04931_),
    .A(_00223_));
 sg13g2_a22oi_1 _21394_ (.Y(_04932_),
    .B1(net760),
    .B2(_03770_),
    .A2(net761),
    .A1(_04931_));
 sg13g2_nor2_1 _21395_ (.A(net986),
    .B(_04932_),
    .Y(_04933_));
 sg13g2_a21oi_1 _21396_ (.A1(net983),
    .A2(\top_ihp.wb_dati_spi[16] ),
    .Y(_04934_),
    .B1(_04933_));
 sg13g2_nand2_1 _21397_ (.Y(_04935_),
    .A(\top_ihp.wb_dati_spi[17] ),
    .B(net456));
 sg13g2_o21ai_1 _21398_ (.B1(_04935_),
    .Y(_02814_),
    .A1(net455),
    .A2(_04934_));
 sg13g2_inv_1 _21399_ (.Y(_04936_),
    .A(_00224_));
 sg13g2_buf_1 _21400_ (.A(_04895_),
    .X(_04937_));
 sg13g2_a22oi_1 _21401_ (.Y(_04938_),
    .B1(net759),
    .B2(_03772_),
    .A2(net761),
    .A1(_04936_));
 sg13g2_nor2_1 _21402_ (.A(net986),
    .B(_04938_),
    .Y(_04939_));
 sg13g2_a21oi_1 _21403_ (.A1(net983),
    .A2(\top_ihp.wb_dati_spi[17] ),
    .Y(_04940_),
    .B1(_04939_));
 sg13g2_nand2_1 _21404_ (.Y(_04941_),
    .A(\top_ihp.wb_dati_spi[18] ),
    .B(net456));
 sg13g2_o21ai_1 _21405_ (.B1(_04941_),
    .Y(_02815_),
    .A1(net455),
    .A2(_04940_));
 sg13g2_inv_1 _21406_ (.Y(_04942_),
    .A(_00225_));
 sg13g2_a22oi_1 _21407_ (.Y(_04943_),
    .B1(net759),
    .B2(_03774_),
    .A2(net761),
    .A1(_04942_));
 sg13g2_nor2_1 _21408_ (.A(net986),
    .B(_04943_),
    .Y(_04944_));
 sg13g2_a21oi_1 _21409_ (.A1(net983),
    .A2(\top_ihp.wb_dati_spi[18] ),
    .Y(_04945_),
    .B1(_04944_));
 sg13g2_nand2_1 _21410_ (.Y(_04946_),
    .A(\top_ihp.wb_dati_spi[19] ),
    .B(net456));
 sg13g2_o21ai_1 _21411_ (.B1(_04946_),
    .Y(_02816_),
    .A1(net455),
    .A2(_04945_));
 sg13g2_nor2_1 _21412_ (.A(net1027),
    .B(_00223_),
    .Y(_04947_));
 sg13g2_a22oi_1 _21413_ (.Y(_04948_),
    .B1(net746),
    .B2(_04947_),
    .A2(\top_ihp.wb_dati_spi[0] ),
    .A1(net989));
 sg13g2_nand2_1 _21414_ (.Y(_04949_),
    .A(\top_ihp.wb_dati_spi[1] ),
    .B(net456));
 sg13g2_o21ai_1 _21415_ (.B1(_04949_),
    .Y(_02817_),
    .A1(net455),
    .A2(_04948_));
 sg13g2_inv_1 _21416_ (.Y(_04950_),
    .A(_00226_));
 sg13g2_a22oi_1 _21417_ (.Y(_04951_),
    .B1(net759),
    .B2(_03778_),
    .A2(net761),
    .A1(_04950_));
 sg13g2_nor2_1 _21418_ (.A(net986),
    .B(_04951_),
    .Y(_04952_));
 sg13g2_a21oi_1 _21419_ (.A1(net983),
    .A2(\top_ihp.wb_dati_spi[19] ),
    .Y(_04953_),
    .B1(_04952_));
 sg13g2_nand2_1 _21420_ (.Y(_04954_),
    .A(\top_ihp.wb_dati_spi[20] ),
    .B(net456));
 sg13g2_o21ai_1 _21421_ (.B1(_04954_),
    .Y(_02818_),
    .A1(net455),
    .A2(_04953_));
 sg13g2_inv_1 _21422_ (.Y(_04955_),
    .A(_00227_));
 sg13g2_a22oi_1 _21423_ (.Y(_04956_),
    .B1(net759),
    .B2(_03780_),
    .A2(net761),
    .A1(_04955_));
 sg13g2_nor2_1 _21424_ (.A(net986),
    .B(_04956_),
    .Y(_04957_));
 sg13g2_a21oi_1 _21425_ (.A1(_08436_),
    .A2(\top_ihp.wb_dati_spi[20] ),
    .Y(_04958_),
    .B1(_04957_));
 sg13g2_nand2_1 _21426_ (.Y(_04959_),
    .A(\top_ihp.wb_dati_spi[21] ),
    .B(net456));
 sg13g2_o21ai_1 _21427_ (.B1(_04959_),
    .Y(_02819_),
    .A1(net455),
    .A2(_04958_));
 sg13g2_buf_1 _21428_ (.A(_08435_),
    .X(_04960_));
 sg13g2_inv_1 _21429_ (.Y(_04961_),
    .A(_00228_));
 sg13g2_a22oi_1 _21430_ (.Y(_04962_),
    .B1(net759),
    .B2(_03782_),
    .A2(_04643_),
    .A1(_04961_));
 sg13g2_nor2_1 _21431_ (.A(net986),
    .B(_04962_),
    .Y(_04963_));
 sg13g2_a21oi_1 _21432_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[21] ),
    .Y(_04964_),
    .B1(_04963_));
 sg13g2_nand2_1 _21433_ (.Y(_04965_),
    .A(\top_ihp.wb_dati_spi[22] ),
    .B(net456));
 sg13g2_o21ai_1 _21434_ (.B1(_04965_),
    .Y(_02820_),
    .A1(net455),
    .A2(_04964_));
 sg13g2_inv_1 _21435_ (.Y(_04966_),
    .A(_00229_));
 sg13g2_a22oi_1 _21436_ (.Y(_04967_),
    .B1(net759),
    .B2(_03784_),
    .A2(net761),
    .A1(_04966_));
 sg13g2_nor2_1 _21437_ (.A(_04902_),
    .B(_04967_),
    .Y(_04968_));
 sg13g2_a21oi_1 _21438_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[22] ),
    .Y(_04969_),
    .B1(_04968_));
 sg13g2_buf_8 _21439_ (.A(_04868_),
    .X(_04970_));
 sg13g2_nand2_1 _21440_ (.Y(_04971_),
    .A(\top_ihp.wb_dati_spi[23] ),
    .B(_04970_));
 sg13g2_o21ai_1 _21441_ (.B1(_04971_),
    .Y(_02821_),
    .A1(_04930_),
    .A2(_04969_));
 sg13g2_nand2_1 _21442_ (.Y(_04972_),
    .A(_03786_),
    .B(_04937_));
 sg13g2_a22oi_1 _21443_ (.Y(_04973_),
    .B1(net777),
    .B2(net1034),
    .A2(net778),
    .A1(_03804_));
 sg13g2_a21oi_1 _21444_ (.A1(_04972_),
    .A2(_04973_),
    .Y(_04974_),
    .B1(net988));
 sg13g2_a21oi_1 _21445_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[23] ),
    .Y(_04975_),
    .B1(_04974_));
 sg13g2_nand2_1 _21446_ (.Y(_04976_),
    .A(\top_ihp.wb_dati_spi[24] ),
    .B(net454));
 sg13g2_o21ai_1 _21447_ (.B1(_04976_),
    .Y(_02822_),
    .A1(net455),
    .A2(_04975_));
 sg13g2_nand2_1 _21448_ (.Y(_04977_),
    .A(_03787_),
    .B(net759));
 sg13g2_a22oi_1 _21449_ (.Y(_04978_),
    .B1(net777),
    .B2(_03776_),
    .A2(net778),
    .A1(_03806_));
 sg13g2_a21oi_1 _21450_ (.A1(_04977_),
    .A2(_04978_),
    .Y(_04979_),
    .B1(net988));
 sg13g2_a21oi_1 _21451_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[24] ),
    .Y(_04980_),
    .B1(_04979_));
 sg13g2_nand2_1 _21452_ (.Y(_04981_),
    .A(\top_ihp.wb_dati_spi[25] ),
    .B(net454));
 sg13g2_o21ai_1 _21453_ (.B1(_04981_),
    .Y(_02823_),
    .A1(_04930_),
    .A2(_04980_));
 sg13g2_buf_1 _21454_ (.A(_04868_),
    .X(_04982_));
 sg13g2_nand2_1 _21455_ (.Y(_04983_),
    .A(_03788_),
    .B(_04937_));
 sg13g2_a22oi_1 _21456_ (.Y(_04984_),
    .B1(net777),
    .B2(_03793_),
    .A2(net778),
    .A1(_03757_));
 sg13g2_a21oi_1 _21457_ (.A1(_04983_),
    .A2(_04984_),
    .Y(_04985_),
    .B1(net988));
 sg13g2_a21oi_1 _21458_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[25] ),
    .Y(_04986_),
    .B1(_04985_));
 sg13g2_nand2_1 _21459_ (.Y(_04987_),
    .A(\top_ihp.wb_dati_spi[26] ),
    .B(net454));
 sg13g2_o21ai_1 _21460_ (.B1(_04987_),
    .Y(_02824_),
    .A1(net453),
    .A2(_04986_));
 sg13g2_nand2_1 _21461_ (.Y(_04988_),
    .A(_03789_),
    .B(net759));
 sg13g2_a22oi_1 _21462_ (.Y(_04989_),
    .B1(net777),
    .B2(_03798_),
    .A2(net778),
    .A1(_03758_));
 sg13g2_a21oi_1 _21463_ (.A1(_04988_),
    .A2(_04989_),
    .Y(_04990_),
    .B1(net988));
 sg13g2_a21oi_1 _21464_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[26] ),
    .Y(_04991_),
    .B1(_04990_));
 sg13g2_nand2_1 _21465_ (.Y(_04992_),
    .A(\top_ihp.wb_dati_spi[27] ),
    .B(net454));
 sg13g2_o21ai_1 _21466_ (.B1(_04992_),
    .Y(_02825_),
    .A1(net453),
    .A2(_04991_));
 sg13g2_nand2_1 _21467_ (.Y(_04993_),
    .A(_03790_),
    .B(_04895_));
 sg13g2_a22oi_1 _21468_ (.Y(_04994_),
    .B1(net777),
    .B2(_03799_),
    .A2(net778),
    .A1(_03760_));
 sg13g2_a21oi_1 _21469_ (.A1(_04993_),
    .A2(_04994_),
    .Y(_04995_),
    .B1(net988));
 sg13g2_a21oi_1 _21470_ (.A1(_04960_),
    .A2(\top_ihp.wb_dati_spi[27] ),
    .Y(_04996_),
    .B1(_04995_));
 sg13g2_nand2_1 _21471_ (.Y(_04997_),
    .A(\top_ihp.wb_dati_spi[28] ),
    .B(net454));
 sg13g2_o21ai_1 _21472_ (.B1(_04997_),
    .Y(_02826_),
    .A1(_04982_),
    .A2(_04996_));
 sg13g2_nand2_1 _21473_ (.Y(_04998_),
    .A(_03792_),
    .B(_04895_));
 sg13g2_a22oi_1 _21474_ (.Y(_04999_),
    .B1(net777),
    .B2(_03800_),
    .A2(net778),
    .A1(_03763_));
 sg13g2_a21oi_1 _21475_ (.A1(_04998_),
    .A2(_04999_),
    .Y(_05000_),
    .B1(net988));
 sg13g2_a21oi_1 _21476_ (.A1(_04960_),
    .A2(\top_ihp.wb_dati_spi[28] ),
    .Y(_05001_),
    .B1(_05000_));
 sg13g2_nand2_1 _21477_ (.Y(_05002_),
    .A(\top_ihp.wb_dati_spi[29] ),
    .B(_04970_));
 sg13g2_o21ai_1 _21478_ (.B1(_05002_),
    .Y(_02827_),
    .A1(_04982_),
    .A2(_05001_));
 sg13g2_nor2_1 _21479_ (.A(net1027),
    .B(_00224_),
    .Y(_05003_));
 sg13g2_a22oi_1 _21480_ (.Y(_05004_),
    .B1(net746),
    .B2(_05003_),
    .A2(\top_ihp.wb_dati_spi[1] ),
    .A1(net989));
 sg13g2_nand2_1 _21481_ (.Y(_05005_),
    .A(\top_ihp.wb_dati_spi[2] ),
    .B(net454));
 sg13g2_o21ai_1 _21482_ (.B1(_05005_),
    .Y(_02828_),
    .A1(net453),
    .A2(_05004_));
 sg13g2_nand2_1 _21483_ (.Y(_05006_),
    .A(_03795_),
    .B(_04895_));
 sg13g2_a22oi_1 _21484_ (.Y(_05007_),
    .B1(net777),
    .B2(_03801_),
    .A2(_04642_),
    .A1(_03765_));
 sg13g2_a21oi_1 _21485_ (.A1(_05006_),
    .A2(_05007_),
    .Y(_05008_),
    .B1(net988));
 sg13g2_a21oi_1 _21486_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[29] ),
    .Y(_05009_),
    .B1(_05008_));
 sg13g2_nand2_1 _21487_ (.Y(_05010_),
    .A(\top_ihp.wb_dati_spi[30] ),
    .B(net454));
 sg13g2_o21ai_1 _21488_ (.B1(_05010_),
    .Y(_02829_),
    .A1(net453),
    .A2(_05009_));
 sg13g2_nand2_1 _21489_ (.Y(_05011_),
    .A(_03797_),
    .B(_04895_));
 sg13g2_a22oi_1 _21490_ (.Y(_05012_),
    .B1(net777),
    .B2(_03802_),
    .A2(net778),
    .A1(_03767_));
 sg13g2_a21oi_1 _21491_ (.A1(_05011_),
    .A2(_05012_),
    .Y(_05013_),
    .B1(net988));
 sg13g2_a21oi_1 _21492_ (.A1(net936),
    .A2(\top_ihp.wb_dati_spi[30] ),
    .Y(_05014_),
    .B1(_05013_));
 sg13g2_nand2_1 _21493_ (.Y(_05015_),
    .A(\top_ihp.wb_dati_spi[31] ),
    .B(net454));
 sg13g2_o21ai_1 _21494_ (.B1(_05015_),
    .Y(_02830_),
    .A1(net453),
    .A2(_05014_));
 sg13g2_nor2_1 _21495_ (.A(net1027),
    .B(_00225_),
    .Y(_05016_));
 sg13g2_a22oi_1 _21496_ (.Y(_05017_),
    .B1(net760),
    .B2(_05016_),
    .A2(\top_ihp.wb_dati_spi[2] ),
    .A1(net989));
 sg13g2_nand2_1 _21497_ (.Y(_05018_),
    .A(\top_ihp.wb_dati_spi[3] ),
    .B(net457));
 sg13g2_o21ai_1 _21498_ (.B1(_05018_),
    .Y(_02831_),
    .A1(net453),
    .A2(_05017_));
 sg13g2_nor2_1 _21499_ (.A(net1027),
    .B(_00226_),
    .Y(_05019_));
 sg13g2_a22oi_1 _21500_ (.Y(_05020_),
    .B1(net760),
    .B2(_05019_),
    .A2(\top_ihp.wb_dati_spi[3] ),
    .A1(net987));
 sg13g2_nand2_1 _21501_ (.Y(_05021_),
    .A(\top_ihp.wb_dati_spi[4] ),
    .B(net457));
 sg13g2_o21ai_1 _21502_ (.B1(_05021_),
    .Y(_02832_),
    .A1(net453),
    .A2(_05020_));
 sg13g2_nor2_1 _21503_ (.A(net1027),
    .B(_00227_),
    .Y(_05022_));
 sg13g2_a22oi_1 _21504_ (.Y(_05023_),
    .B1(net760),
    .B2(_05022_),
    .A2(\top_ihp.wb_dati_spi[4] ),
    .A1(net987));
 sg13g2_nand2_1 _21505_ (.Y(_05024_),
    .A(\top_ihp.wb_dati_spi[5] ),
    .B(net457));
 sg13g2_o21ai_1 _21506_ (.B1(_05024_),
    .Y(_02833_),
    .A1(net453),
    .A2(_05023_));
 sg13g2_nor2_1 _21507_ (.A(net1027),
    .B(_00228_),
    .Y(_05025_));
 sg13g2_a22oi_1 _21508_ (.Y(_05026_),
    .B1(net760),
    .B2(_05025_),
    .A2(\top_ihp.wb_dati_spi[5] ),
    .A1(net987));
 sg13g2_nand2_1 _21509_ (.Y(_05027_),
    .A(\top_ihp.wb_dati_spi[6] ),
    .B(net457));
 sg13g2_o21ai_1 _21510_ (.B1(_05027_),
    .Y(_02834_),
    .A1(net459),
    .A2(_05026_));
 sg13g2_nor2_1 _21511_ (.A(net1027),
    .B(_00229_),
    .Y(_05028_));
 sg13g2_a22oi_1 _21512_ (.Y(_05029_),
    .B1(net760),
    .B2(_05028_),
    .A2(\top_ihp.wb_dati_spi[6] ),
    .A1(net987));
 sg13g2_nand2_1 _21513_ (.Y(_05030_),
    .A(\top_ihp.wb_dati_spi[7] ),
    .B(net457));
 sg13g2_o21ai_1 _21514_ (.B1(_05030_),
    .Y(_02835_),
    .A1(net459),
    .A2(_05029_));
 sg13g2_nor2b_1 _21515_ (.A(net986),
    .B_N(_03804_),
    .Y(_05031_));
 sg13g2_a22oi_1 _21516_ (.Y(_05032_),
    .B1(net760),
    .B2(_05031_),
    .A2(\top_ihp.wb_dati_spi[7] ),
    .A1(net987));
 sg13g2_nand2_1 _21517_ (.Y(_05033_),
    .A(\top_ihp.wb_dati_spi[8] ),
    .B(net457));
 sg13g2_o21ai_1 _21518_ (.B1(_05033_),
    .Y(_02836_),
    .A1(net459),
    .A2(_05032_));
 sg13g2_nor2b_1 _21519_ (.A(_04920_),
    .B_N(_03806_),
    .Y(_05034_));
 sg13g2_a22oi_1 _21520_ (.Y(_05035_),
    .B1(_04896_),
    .B2(_05034_),
    .A2(\top_ihp.wb_dati_spi[8] ),
    .A1(net987));
 sg13g2_nand2_1 _21521_ (.Y(_05036_),
    .A(\top_ihp.wb_dati_spi[9] ),
    .B(net457));
 sg13g2_o21ai_1 _21522_ (.B1(_05036_),
    .Y(_02837_),
    .A1(net459),
    .A2(_05035_));
 sg13g2_nor2_1 _21523_ (.A(net983),
    .B(_03818_),
    .Y(_05037_));
 sg13g2_and2_1 _21524_ (.A(_00096_),
    .B(_08213_),
    .X(_05038_));
 sg13g2_a22oi_1 _21525_ (.Y(_05039_),
    .B1(_05038_),
    .B2(_08426_),
    .A2(_08442_),
    .A1(_08427_));
 sg13g2_buf_1 _21526_ (.A(_05039_),
    .X(_05040_));
 sg13g2_mux2_1 _21527_ (.A0(_00351_),
    .A1(_05037_),
    .S(_05040_),
    .X(_02838_));
 sg13g2_and2_1 _21528_ (.A(_04863_),
    .B(_04474_),
    .X(_05041_));
 sg13g2_mux2_1 _21529_ (.A0(_00352_),
    .A1(_05041_),
    .S(_05040_),
    .X(_02839_));
 sg13g2_nor2_1 _21530_ (.A(net983),
    .B(_04480_),
    .Y(_05042_));
 sg13g2_mux2_1 _21531_ (.A0(_00353_),
    .A1(_05042_),
    .S(_05040_),
    .X(_02840_));
 sg13g2_buf_1 _21532_ (.A(\top_ihp.wb_uart.state[1] ),
    .X(_05043_));
 sg13g2_nor2b_1 _21533_ (.A(_05043_),
    .B_N(\top_ihp.wb_uart.state[0] ),
    .Y(_05044_));
 sg13g2_a22oi_1 _21534_ (.Y(_05045_),
    .B1(\top_ihp.wb_uart.tx_ready ),
    .B2(_05044_),
    .A2(\top_ihp.wb_uart.rx_ready ),
    .A1(_05043_));
 sg13g2_nor2_1 _21535_ (.A(_09663_),
    .B(_09860_),
    .Y(_05046_));
 sg13g2_a21oi_1 _21536_ (.A1(_09663_),
    .A2(_05045_),
    .Y(_02841_),
    .B1(_05046_));
 sg13g2_inv_1 _21537_ (.Y(_05047_),
    .A(\top_ihp.wb_uart.rx_ready ));
 sg13g2_nand3_1 _21538_ (.B(\top_ihp.wb_uart.state[0] ),
    .C(_05047_),
    .A(_05043_),
    .Y(_05048_));
 sg13g2_nor2_1 _21539_ (.A(_05043_),
    .B(\top_ihp.wb_uart.state[0] ),
    .Y(_05049_));
 sg13g2_nand2_1 _21540_ (.Y(_05050_),
    .A(_08813_),
    .B(_05049_));
 sg13g2_nand2b_1 _21541_ (.Y(_05051_),
    .B(_05044_),
    .A_N(\top_ihp.wb_uart.tx_ready ));
 sg13g2_nand3_1 _21542_ (.B(_05050_),
    .C(_05051_),
    .A(_05048_),
    .Y(_02842_));
 sg13g2_nor2b_1 _21543_ (.A(\top_ihp.wb_uart.rx_ready ),
    .B_N(_05043_),
    .Y(_05052_));
 sg13g2_a21o_1 _21544_ (.A2(_05049_),
    .A1(_08667_),
    .B1(_05052_),
    .X(_02843_));
 sg13g2_xnor2_1 _21545_ (.Y(_05053_),
    .A(net1044),
    .B(_08707_));
 sg13g2_nor2_1 _21546_ (.A(_08722_),
    .B(_05053_),
    .Y(_02844_));
 sg13g2_nand2_1 _21547_ (.Y(_05054_),
    .A(net1044),
    .B(_08707_));
 sg13g2_xor2_1 _21548_ (.B(_05054_),
    .A(net1043),
    .X(_05055_));
 sg13g2_nor2_1 _21549_ (.A(_08722_),
    .B(_05055_),
    .Y(_02845_));
 sg13g2_nand3_1 _21550_ (.B(net1043),
    .C(_08707_),
    .A(net1044),
    .Y(_05056_));
 sg13g2_xor2_1 _21551_ (.B(_05056_),
    .A(net1042),
    .X(_05057_));
 sg13g2_nor2_1 _21552_ (.A(_08722_),
    .B(_05057_),
    .Y(_02846_));
 sg13g2_inv_1 _21553_ (.Y(_05058_),
    .A(_00220_));
 sg13g2_nand4_1 _21554_ (.B(net1042),
    .C(_05058_),
    .A(net1043),
    .Y(_05059_),
    .D(_08707_));
 sg13g2_xor2_1 _21555_ (.B(_05059_),
    .A(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ),
    .X(_05060_));
 sg13g2_nor2_1 _21556_ (.A(_08722_),
    .B(_05060_),
    .Y(_02847_));
 sg13g2_inv_2 _21557_ (.Y(_05061_),
    .A(_08722_));
 sg13g2_and2_1 _21558_ (.A(_08703_),
    .B(_08702_),
    .X(_05062_));
 sg13g2_nor3_1 _21559_ (.A(_08694_),
    .B(_08686_),
    .C(_08692_),
    .Y(_05063_));
 sg13g2_inv_1 _21560_ (.Y(_05064_),
    .A(_08695_));
 sg13g2_nand4_1 _21561_ (.B(_08698_),
    .C(_08699_),
    .A(_08697_),
    .Y(_05065_),
    .D(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ));
 sg13g2_nor3_1 _21562_ (.A(_05064_),
    .B(_08704_),
    .C(_05065_),
    .Y(_05066_));
 sg13g2_nand4_1 _21563_ (.B(_05062_),
    .C(_05063_),
    .A(_05061_),
    .Y(_05067_),
    .D(_05066_));
 sg13g2_buf_1 _21564_ (.A(_05067_),
    .X(_05068_));
 sg13g2_or4_1 _21565_ (.A(net1044),
    .B(net1043),
    .C(net1042),
    .D(_05068_),
    .X(_05069_));
 sg13g2_nand2_1 _21566_ (.Y(_05070_),
    .A(_00220_),
    .B(net1060));
 sg13g2_nand2_1 _21567_ (.Y(_05071_),
    .A(\top_ihp.wb_dati_uart[0] ),
    .B(_05069_));
 sg13g2_o21ai_1 _21568_ (.B1(_05071_),
    .Y(_02848_),
    .A1(_05069_),
    .A2(_05070_));
 sg13g2_inv_1 _21569_ (.Y(_05072_),
    .A(net1044));
 sg13g2_nor4_1 _21570_ (.A(_05072_),
    .B(net1043),
    .C(net1042),
    .D(_05068_),
    .Y(_05073_));
 sg13g2_mux2_1 _21571_ (.A0(\top_ihp.wb_dati_uart[1] ),
    .A1(net1060),
    .S(_05073_),
    .X(_02849_));
 sg13g2_nor2_1 _21572_ (.A(net1044),
    .B(_05068_),
    .Y(_05074_));
 sg13g2_nand3b_1 _21573_ (.B(_05074_),
    .C(net1043),
    .Y(_05075_),
    .A_N(net1042));
 sg13g2_mux2_1 _21574_ (.A0(net1060),
    .A1(\top_ihp.wb_dati_uart[2] ),
    .S(_05075_),
    .X(_02850_));
 sg13g2_nand2_1 _21575_ (.Y(_05076_),
    .A(net1044),
    .B(net1043));
 sg13g2_nor3_1 _21576_ (.A(net1042),
    .B(_05076_),
    .C(_05068_),
    .Y(_05077_));
 sg13g2_mux2_1 _21577_ (.A0(\top_ihp.wb_dati_uart[3] ),
    .A1(net1060),
    .S(_05077_),
    .X(_02851_));
 sg13g2_nor2_1 _21578_ (.A(net1042),
    .B(_05076_),
    .Y(_05078_));
 sg13g2_nor2b_1 _21579_ (.A(_08709_),
    .B_N(_08710_),
    .Y(_05079_));
 sg13g2_and2_1 _21580_ (.A(_05072_),
    .B(_05079_),
    .X(_05080_));
 sg13g2_o21ai_1 _21581_ (.B1(_00220_),
    .Y(_05081_),
    .A1(_05078_),
    .A2(_05080_));
 sg13g2_o21ai_1 _21582_ (.B1(\top_ihp.wb_dati_uart[4] ),
    .Y(_05082_),
    .A1(_05068_),
    .A2(_05081_));
 sg13g2_nand3_1 _21583_ (.B(_05074_),
    .C(_05079_),
    .A(net1060),
    .Y(_05083_));
 sg13g2_nand2_1 _21584_ (.Y(_02852_),
    .A(_05082_),
    .B(_05083_));
 sg13g2_inv_1 _21585_ (.Y(_05084_),
    .A(_05068_));
 sg13g2_nand3_1 _21586_ (.B(_05084_),
    .C(_05079_),
    .A(_08708_),
    .Y(_05085_));
 sg13g2_mux2_1 _21587_ (.A0(_08669_),
    .A1(_10607_),
    .S(_05085_),
    .X(_02853_));
 sg13g2_nand3_1 _21588_ (.B(_08710_),
    .C(_05074_),
    .A(_08709_),
    .Y(_05086_));
 sg13g2_mux2_1 _21589_ (.A0(net1060),
    .A1(\top_ihp.wb_dati_uart[6] ),
    .S(_05086_),
    .X(_02854_));
 sg13g2_nor2_1 _21590_ (.A(_08712_),
    .B(_05068_),
    .Y(_05087_));
 sg13g2_mux2_1 _21591_ (.A0(\top_ihp.wb_dati_uart[7] ),
    .A1(_08669_),
    .S(_05087_),
    .X(_02855_));
 sg13g2_a21oi_1 _21592_ (.A1(_08697_),
    .A2(_00097_),
    .Y(_05088_),
    .B1(_08745_));
 sg13g2_a21o_1 _21593_ (.A2(_05088_),
    .A1(_08704_),
    .B1(_05066_),
    .X(_05089_));
 sg13g2_a22oi_1 _21594_ (.Y(_05090_),
    .B1(_05089_),
    .B2(_05062_),
    .A2(_05088_),
    .A1(_05065_));
 sg13g2_nand2_2 _21595_ (.Y(_05091_),
    .A(_05063_),
    .B(_05090_));
 sg13g2_a21oi_1 _21596_ (.A1(_08620_),
    .A2(_08719_),
    .Y(_05092_),
    .B1(_05047_));
 sg13g2_a21o_1 _21597_ (.A2(_05091_),
    .A1(_08720_),
    .B1(_05092_),
    .X(_02856_));
 sg13g2_xnor2_1 _21598_ (.Y(_05093_),
    .A(_08818_),
    .B(_08849_));
 sg13g2_nor2_1 _21599_ (.A(_08853_),
    .B(_05093_),
    .Y(_02857_));
 sg13g2_nand2_1 _21600_ (.Y(_05094_),
    .A(_08818_),
    .B(_08849_));
 sg13g2_xor2_1 _21601_ (.B(_05094_),
    .A(_08819_),
    .X(_05095_));
 sg13g2_nor2_1 _21602_ (.A(_08853_),
    .B(_05095_),
    .Y(_02858_));
 sg13g2_o21ai_1 _21603_ (.B1(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .Y(_05096_),
    .A1(_08834_),
    .A2(_08847_));
 sg13g2_nand2_1 _21604_ (.Y(_05097_),
    .A(_08818_),
    .B(_08819_));
 sg13g2_xor2_1 _21605_ (.B(_05097_),
    .A(_00221_),
    .X(_05098_));
 sg13g2_nand2_1 _21606_ (.Y(_05099_),
    .A(_08849_),
    .B(_05098_));
 sg13g2_a21oi_1 _21607_ (.A1(_05096_),
    .A2(_05099_),
    .Y(_02859_),
    .B1(_08853_));
 sg13g2_xor2_1 _21608_ (.B(_08850_),
    .A(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ),
    .X(_05100_));
 sg13g2_nor2_1 _21609_ (.A(_08853_),
    .B(_05100_),
    .Y(_02860_));
 sg13g2_mux2_1 _21610_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .A1(net1034),
    .S(_08859_),
    .X(_02861_));
 sg13g2_mux2_1 _21611_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .A1(_03776_),
    .S(net593),
    .X(_02862_));
 sg13g2_mux2_1 _21612_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .A1(_03793_),
    .S(net593),
    .X(_02863_));
 sg13g2_mux2_1 _21613_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .A1(_03798_),
    .S(net593),
    .X(_02864_));
 sg13g2_mux2_1 _21614_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .A1(_03799_),
    .S(net593),
    .X(_02865_));
 sg13g2_mux2_1 _21615_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .A1(_03800_),
    .S(net593),
    .X(_02866_));
 sg13g2_mux2_1 _21616_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .A1(_03801_),
    .S(net593),
    .X(_02867_));
 sg13g2_mux2_1 _21617_ (.A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .A1(_03802_),
    .S(_08859_),
    .X(_02868_));
 sg13g2_inv_1 _21618_ (.Y(_05101_),
    .A(_08814_));
 sg13g2_nor2_1 _21619_ (.A(_05101_),
    .B(_08854_),
    .Y(_05102_));
 sg13g2_nor3_1 _21620_ (.A(\top_ihp.wb_uart.tx_ready ),
    .B(_08816_),
    .C(_05102_),
    .Y(_05103_));
 sg13g2_nor2_1 _21621_ (.A(net593),
    .B(_05103_),
    .Y(_02869_));
 sg13g2_nand2_1 _21622_ (.Y(_05104_),
    .A(_10098_),
    .B(_10131_));
 sg13g2_nor2_2 _21623_ (.A(_10071_),
    .B(_10131_),
    .Y(_05105_));
 sg13g2_nand2_1 _21624_ (.Y(_05106_),
    .A(net731),
    .B(_05105_));
 sg13g2_nor2_1 _21625_ (.A(_10470_),
    .B(_10474_),
    .Y(_05107_));
 sg13g2_a21oi_1 _21626_ (.A1(net1001),
    .A2(\top_ihp.wb_dati_uart[2] ),
    .Y(_05108_),
    .B1(_05107_));
 sg13g2_buf_1 _21627_ (.A(_05108_),
    .X(_05109_));
 sg13g2_nor2b_1 _21628_ (.A(\top_ihp.wb_dati_uart[4] ),
    .B_N(net1001),
    .Y(_05110_));
 sg13g2_nor3_1 _21629_ (.A(_10470_),
    .B(_10581_),
    .C(_10611_),
    .Y(_05111_));
 sg13g2_a21o_1 _21630_ (.A2(_05110_),
    .A1(_10607_),
    .B1(_05111_),
    .X(_05112_));
 sg13g2_buf_2 _21631_ (.A(_05112_),
    .X(_05113_));
 sg13g2_nand2_1 _21632_ (.Y(_05114_),
    .A(net738),
    .B(_05113_));
 sg13g2_a21oi_1 _21633_ (.A1(_05104_),
    .A2(_05106_),
    .Y(_05115_),
    .B1(_05114_));
 sg13g2_or2_1 _21634_ (.X(_05116_),
    .B(_10583_),
    .A(net749));
 sg13g2_buf_2 _21635_ (.A(_05116_),
    .X(_05117_));
 sg13g2_buf_1 _21636_ (.A(_10071_),
    .X(_05118_));
 sg13g2_buf_1 _21637_ (.A(_10133_),
    .X(_05119_));
 sg13g2_nor2_1 _21638_ (.A(net727),
    .B(net726),
    .Y(_05120_));
 sg13g2_a21oi_1 _21639_ (.A1(net727),
    .A2(_05104_),
    .Y(_05121_),
    .B1(_05120_));
 sg13g2_nor2_1 _21640_ (.A(_05117_),
    .B(_05121_),
    .Y(_05122_));
 sg13g2_nand2_1 _21641_ (.Y(_05123_),
    .A(_10637_),
    .B(_05113_));
 sg13g2_inv_1 _21642_ (.Y(_05124_),
    .A(_10637_));
 sg13g2_nand2_2 _21643_ (.Y(_05125_),
    .A(_10071_),
    .B(_10097_));
 sg13g2_a21oi_1 _21644_ (.A1(_10614_),
    .A2(_05125_),
    .Y(_05126_),
    .B1(_05117_));
 sg13g2_nand3_1 _21645_ (.B(_05124_),
    .C(_05126_),
    .A(_10139_),
    .Y(_05127_));
 sg13g2_a21o_1 _21646_ (.A2(_05127_),
    .A1(_05123_),
    .B1(_10544_),
    .X(_05128_));
 sg13g2_buf_2 _21647_ (.A(_05128_),
    .X(_05129_));
 sg13g2_buf_1 _21648_ (.A(_05129_),
    .X(_05130_));
 sg13g2_mux2_1 _21649_ (.A0(_05115_),
    .A1(_05122_),
    .S(net340),
    .X(_05131_));
 sg13g2_buf_1 _21650_ (.A(net747),
    .X(_05132_));
 sg13g2_mux2_1 _21651_ (.A0(\top_ihp.oisc.decoder.decoded[0] ),
    .A1(_05131_),
    .S(net737),
    .X(_00357_));
 sg13g2_and2_1 _21652_ (.A(_10544_),
    .B(_10637_),
    .X(_05133_));
 sg13g2_nor2_1 _21653_ (.A(_10544_),
    .B(_10637_),
    .Y(_05134_));
 sg13g2_a22oi_1 _21654_ (.Y(_05135_),
    .B1(_05134_),
    .B2(net730),
    .A2(_05133_),
    .A1(_05113_));
 sg13g2_buf_1 _21655_ (.A(_05135_),
    .X(_05136_));
 sg13g2_or2_1 _21656_ (.X(_05137_),
    .B(_05136_),
    .A(net738));
 sg13g2_buf_2 _21657_ (.A(_05137_),
    .X(_05138_));
 sg13g2_inv_1 _21658_ (.Y(_05139_),
    .A(_10071_));
 sg13g2_nor2_1 _21659_ (.A(net738),
    .B(_05136_),
    .Y(_05140_));
 sg13g2_nor2_1 _21660_ (.A(_05139_),
    .B(_05140_),
    .Y(_05141_));
 sg13g2_buf_1 _21661_ (.A(_10098_),
    .X(_05142_));
 sg13g2_a221oi_1 _21662_ (.B2(net725),
    .C1(_05114_),
    .B1(_05141_),
    .A1(_10131_),
    .Y(_05143_),
    .A2(_05138_));
 sg13g2_nand2_1 _21663_ (.Y(_05144_),
    .A(net340),
    .B(_05143_));
 sg13g2_nand2_1 _21664_ (.Y(_05145_),
    .A(_08201_),
    .B(net750));
 sg13g2_o21ai_1 _21665_ (.B1(_05145_),
    .Y(_00358_),
    .A1(net751),
    .A2(_05144_));
 sg13g2_buf_1 _21666_ (.A(net763),
    .X(_05146_));
 sg13g2_buf_1 _21667_ (.A(net749),
    .X(_05147_));
 sg13g2_buf_1 _21668_ (.A(_10614_),
    .X(_05148_));
 sg13g2_o21ai_1 _21669_ (.B1(net710),
    .Y(_05149_),
    .A1(net731),
    .A2(_05105_));
 sg13g2_nor4_1 _21670_ (.A(net763),
    .B(net736),
    .C(net730),
    .D(_05149_),
    .Y(_05150_));
 sg13g2_a21o_1 _21671_ (.A2(net745),
    .A1(_08415_),
    .B1(_05150_),
    .X(_00359_));
 sg13g2_nor2_1 _21672_ (.A(net726),
    .B(_05140_),
    .Y(_05151_));
 sg13g2_nor2_1 _21673_ (.A(_05117_),
    .B(_05125_),
    .Y(_05152_));
 sg13g2_a21oi_2 _21674_ (.B1(_05129_),
    .Y(_05153_),
    .A2(_05152_),
    .A1(_05151_));
 sg13g2_buf_1 _21675_ (.A(_10583_),
    .X(_05154_));
 sg13g2_nor2_1 _21676_ (.A(net736),
    .B(net735),
    .Y(_05155_));
 sg13g2_nor2_1 _21677_ (.A(net738),
    .B(net730),
    .Y(_05156_));
 sg13g2_a21oi_1 _21678_ (.A1(_05106_),
    .A2(_05138_),
    .Y(_05157_),
    .B1(net710));
 sg13g2_o21ai_1 _21679_ (.B1(_05157_),
    .Y(_05158_),
    .A1(_05155_),
    .A2(_05156_));
 sg13g2_nand2_1 _21680_ (.Y(_05159_),
    .A(_10583_),
    .B(net710));
 sg13g2_a21oi_2 _21681_ (.B1(net738),
    .Y(_05160_),
    .A2(_05136_),
    .A1(_05106_));
 sg13g2_and2_1 _21682_ (.A(net735),
    .B(_05149_),
    .X(_05161_));
 sg13g2_o21ai_1 _21683_ (.B1(net340),
    .Y(_05162_),
    .A1(_05147_),
    .A2(_05161_));
 sg13g2_a21oi_1 _21684_ (.A1(_05159_),
    .A2(_05160_),
    .Y(_05163_),
    .B1(_05162_));
 sg13g2_a21oi_1 _21685_ (.A1(_05153_),
    .A2(_05158_),
    .Y(_05164_),
    .B1(_05163_));
 sg13g2_mux2_1 _21686_ (.A0(_09893_),
    .A1(_05164_),
    .S(net737),
    .X(_00360_));
 sg13g2_nand2_1 _21687_ (.Y(_05165_),
    .A(net727),
    .B(net710));
 sg13g2_o21ai_1 _21688_ (.B1(net731),
    .Y(_05166_),
    .A1(_05109_),
    .A2(_05105_));
 sg13g2_a221oi_1 _21689_ (.B2(_05138_),
    .C1(net735),
    .B1(_05166_),
    .A1(net738),
    .Y(_05167_),
    .A2(_05165_));
 sg13g2_o21ai_1 _21690_ (.B1(_05167_),
    .Y(_05168_),
    .A1(net340),
    .A2(_05151_));
 sg13g2_and2_1 _21691_ (.A(net747),
    .B(_05168_),
    .X(_05169_));
 sg13g2_a22oi_1 _21692_ (.Y(_00361_),
    .B1(_05144_),
    .B2(_05169_),
    .A2(net751),
    .A1(_09799_));
 sg13g2_nor2_1 _21693_ (.A(_05147_),
    .B(net710),
    .Y(_05170_));
 sg13g2_a21oi_1 _21694_ (.A1(net730),
    .A2(_05125_),
    .Y(_05171_),
    .B1(net726));
 sg13g2_nand2_1 _21695_ (.Y(_05172_),
    .A(net731),
    .B(_10133_));
 sg13g2_nor2_1 _21696_ (.A(_05139_),
    .B(_10583_),
    .Y(_05173_));
 sg13g2_nor2_1 _21697_ (.A(_05172_),
    .B(_05173_),
    .Y(_05174_));
 sg13g2_nor3_1 _21698_ (.A(_05129_),
    .B(_05171_),
    .C(_05174_),
    .Y(_05175_));
 sg13g2_a21oi_1 _21699_ (.A1(_05154_),
    .A2(net340),
    .Y(_05176_),
    .B1(_05175_));
 sg13g2_a22oi_1 _21700_ (.Y(_05177_),
    .B1(_05170_),
    .B2(_05176_),
    .A2(_05160_),
    .A1(net730));
 sg13g2_nand2_1 _21701_ (.Y(_05178_),
    .A(net1004),
    .B(net750));
 sg13g2_o21ai_1 _21702_ (.B1(_05178_),
    .Y(_00362_),
    .A1(net751),
    .A2(_05177_));
 sg13g2_nand2_1 _21703_ (.Y(_05179_),
    .A(_05113_),
    .B(_05160_));
 sg13g2_nand3_1 _21704_ (.B(net340),
    .C(_05179_),
    .A(_03736_),
    .Y(_05180_));
 sg13g2_nor2_1 _21705_ (.A(_05126_),
    .B(_05180_),
    .Y(_05181_));
 sg13g2_nor2_1 _21706_ (.A(_09797_),
    .B(net747),
    .Y(_05182_));
 sg13g2_buf_1 _21707_ (.A(net763),
    .X(_05183_));
 sg13g2_or3_1 _21708_ (.A(net749),
    .B(net710),
    .C(_05106_),
    .X(_05184_));
 sg13g2_buf_1 _21709_ (.A(_05184_),
    .X(_05185_));
 sg13g2_o21ai_1 _21710_ (.B1(_05153_),
    .Y(_05186_),
    .A1(net735),
    .A2(_05185_));
 sg13g2_nor2_1 _21711_ (.A(net744),
    .B(_05186_),
    .Y(_05187_));
 sg13g2_nor3_1 _21712_ (.A(_05181_),
    .B(_05182_),
    .C(_05187_),
    .Y(_00363_));
 sg13g2_nor2_1 _21713_ (.A(net726),
    .B(net736),
    .Y(_05188_));
 sg13g2_o21ai_1 _21714_ (.B1(_05113_),
    .Y(_05189_),
    .A1(_05160_),
    .A2(_05188_));
 sg13g2_or2_1 _21715_ (.X(_05190_),
    .B(_10637_),
    .A(_10544_));
 sg13g2_nand2_1 _21716_ (.Y(_05191_),
    .A(net730),
    .B(_05148_));
 sg13g2_o21ai_1 _21717_ (.B1(net749),
    .Y(_05192_),
    .A1(_05190_),
    .A2(_05191_));
 sg13g2_nand2_1 _21718_ (.Y(_05193_),
    .A(_10544_),
    .B(_10637_));
 sg13g2_o21ai_1 _21719_ (.B1(net749),
    .Y(_05194_),
    .A1(net710),
    .A2(_05193_));
 sg13g2_a21oi_1 _21720_ (.A1(_10607_),
    .A2(_05110_),
    .Y(_05195_),
    .B1(_05111_));
 sg13g2_nand3_1 _21721_ (.B(_10586_),
    .C(_10614_),
    .A(net749),
    .Y(_05196_));
 sg13g2_a21oi_1 _21722_ (.A1(_05195_),
    .A2(_05196_),
    .Y(_05197_),
    .B1(_05118_));
 sg13g2_a221oi_1 _21723_ (.B2(net735),
    .C1(_05197_),
    .B1(_05194_),
    .A1(_05118_),
    .Y(_05198_),
    .A2(_05192_));
 sg13g2_a21o_1 _21724_ (.A2(_05138_),
    .A1(_05172_),
    .B1(_05198_),
    .X(_05199_));
 sg13g2_a21oi_1 _21725_ (.A1(net731),
    .A2(_05148_),
    .Y(_05200_),
    .B1(net730));
 sg13g2_nor2_1 _21726_ (.A(_10133_),
    .B(_05200_),
    .Y(_05201_));
 sg13g2_a21oi_1 _21727_ (.A1(net725),
    .A2(_05105_),
    .Y(_05202_),
    .B1(_05201_));
 sg13g2_o21ai_1 _21728_ (.B1(_05129_),
    .Y(_05203_),
    .A1(net736),
    .A2(_05202_));
 sg13g2_inv_1 _21729_ (.Y(_05204_),
    .A(_05203_));
 sg13g2_a221oi_1 _21730_ (.B2(_05204_),
    .C1(net763),
    .B1(_05199_),
    .A1(_05153_),
    .Y(_05205_),
    .A2(_05189_));
 sg13g2_a21o_1 _21731_ (.A2(net745),
    .A1(\top_ihp.oisc.decoder.decoded[1] ),
    .B1(_05205_),
    .X(_00364_));
 sg13g2_inv_1 _21732_ (.Y(_05206_),
    .A(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_nor4_1 _21733_ (.A(_05139_),
    .B(_05119_),
    .C(net749),
    .D(_05195_),
    .Y(_05207_));
 sg13g2_nor3_1 _21734_ (.A(net763),
    .B(_05129_),
    .C(_05207_),
    .Y(_05208_));
 sg13g2_nand2_1 _21735_ (.Y(_05209_),
    .A(_03736_),
    .B(_05130_));
 sg13g2_o21ai_1 _21736_ (.B1(_05159_),
    .Y(_05210_),
    .A1(_05139_),
    .A2(_10583_));
 sg13g2_nand4_1 _21737_ (.B(_10131_),
    .C(_05138_),
    .A(net731),
    .Y(_05211_),
    .D(_05210_));
 sg13g2_nand3_1 _21738_ (.B(net735),
    .C(_05105_),
    .A(_05142_),
    .Y(_05212_));
 sg13g2_a21oi_1 _21739_ (.A1(_05211_),
    .A2(_05212_),
    .Y(_05213_),
    .B1(net736));
 sg13g2_o21ai_1 _21740_ (.B1(net738),
    .Y(_05214_),
    .A1(net727),
    .A2(_05154_));
 sg13g2_a21o_1 _21741_ (.A2(net736),
    .A1(net727),
    .B1(_05172_),
    .X(_05215_));
 sg13g2_a22oi_1 _21742_ (.Y(_05216_),
    .B1(_05215_),
    .B2(_05138_),
    .A2(_05214_),
    .A1(_05196_));
 sg13g2_nor3_1 _21743_ (.A(_05209_),
    .B(_05213_),
    .C(_05216_),
    .Y(_05217_));
 sg13g2_a221oi_1 _21744_ (.B2(_05208_),
    .C1(_05217_),
    .B1(_05185_),
    .A1(_05206_),
    .Y(_00365_),
    .A2(net750));
 sg13g2_a22oi_1 _21745_ (.Y(_05218_),
    .B1(_05141_),
    .B2(_10097_),
    .A2(net725),
    .A1(_05139_));
 sg13g2_nand3_1 _21746_ (.B(net738),
    .C(_05113_),
    .A(_10131_),
    .Y(_05219_));
 sg13g2_o21ai_1 _21747_ (.B1(_05179_),
    .Y(_05220_),
    .A1(_05218_),
    .A2(_05219_));
 sg13g2_a21oi_1 _21748_ (.A1(_10131_),
    .A2(net735),
    .Y(_05221_),
    .B1(net727));
 sg13g2_o21ai_1 _21749_ (.B1(_10583_),
    .Y(_05222_),
    .A1(_10133_),
    .A2(net710));
 sg13g2_nor2_1 _21750_ (.A(net725),
    .B(_05222_),
    .Y(_05223_));
 sg13g2_a21oi_1 _21751_ (.A1(_05142_),
    .A2(_05221_),
    .Y(_05224_),
    .B1(_05223_));
 sg13g2_o21ai_1 _21752_ (.B1(_05130_),
    .Y(_05225_),
    .A1(net736),
    .A2(_05224_));
 sg13g2_o21ai_1 _21753_ (.B1(_05225_),
    .Y(_05226_),
    .A1(net340),
    .A2(_05220_));
 sg13g2_nand2_1 _21754_ (.Y(_05227_),
    .A(\top_ihp.oisc.decoder.decoded[3] ),
    .B(net750));
 sg13g2_o21ai_1 _21755_ (.B1(_05227_),
    .Y(_00366_),
    .A1(net751),
    .A2(_05226_));
 sg13g2_inv_1 _21756_ (.Y(_05228_),
    .A(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_a21oi_1 _21757_ (.A1(net727),
    .A2(_10131_),
    .Y(_05229_),
    .B1(net725));
 sg13g2_nor2_1 _21758_ (.A(_05117_),
    .B(_05229_),
    .Y(_05230_));
 sg13g2_nand2_1 _21759_ (.Y(_05231_),
    .A(net735),
    .B(_05157_));
 sg13g2_nor3_1 _21760_ (.A(net725),
    .B(net726),
    .C(net736),
    .Y(_05232_));
 sg13g2_o21ai_1 _21761_ (.B1(_05232_),
    .Y(_05233_),
    .A1(_05113_),
    .A2(_05173_));
 sg13g2_nand3_1 _21762_ (.B(_05231_),
    .C(_05233_),
    .A(_05208_),
    .Y(_05234_));
 sg13g2_o21ai_1 _21763_ (.B1(_05234_),
    .Y(_05235_),
    .A1(_05180_),
    .A2(_05230_));
 sg13g2_a21oi_1 _21764_ (.A1(_05228_),
    .A2(net751),
    .Y(_00367_),
    .B1(_05235_));
 sg13g2_inv_1 _21765_ (.Y(_05236_),
    .A(_05151_));
 sg13g2_o21ai_1 _21766_ (.B1(_05125_),
    .Y(_05237_),
    .A1(net727),
    .A2(_05236_));
 sg13g2_a21oi_1 _21767_ (.A1(_05155_),
    .A2(_05237_),
    .Y(_05238_),
    .B1(_05209_));
 sg13g2_nor2_1 _21768_ (.A(\top_ihp.oisc.decoder.decoded[5] ),
    .B(net747),
    .Y(_05239_));
 sg13g2_o21ai_1 _21769_ (.B1(_05153_),
    .Y(_05240_),
    .A1(net730),
    .A2(_05185_));
 sg13g2_nor2_1 _21770_ (.A(net744),
    .B(_05240_),
    .Y(_05241_));
 sg13g2_nor3_1 _21771_ (.A(_05238_),
    .B(_05239_),
    .C(_05241_),
    .Y(_00368_));
 sg13g2_a21oi_1 _21772_ (.A1(net726),
    .A2(_05125_),
    .Y(_05242_),
    .B1(_05114_));
 sg13g2_a21oi_1 _21773_ (.A1(net725),
    .A2(net726),
    .Y(_05243_),
    .B1(_05120_));
 sg13g2_nor2_1 _21774_ (.A(_05117_),
    .B(_05243_),
    .Y(_05244_));
 sg13g2_mux2_1 _21775_ (.A0(_05242_),
    .A1(_05244_),
    .S(net340),
    .X(_05245_));
 sg13g2_mux2_1 _21776_ (.A0(\top_ihp.oisc.decoder.decoded[6] ),
    .A1(_05245_),
    .S(net737),
    .X(_00369_));
 sg13g2_a21oi_1 _21777_ (.A1(net725),
    .A2(net726),
    .Y(_05246_),
    .B1(_05141_));
 sg13g2_nor4_1 _21778_ (.A(net763),
    .B(_05117_),
    .C(_05153_),
    .D(_05246_),
    .Y(_05247_));
 sg13g2_a21o_1 _21779_ (.A2(net750),
    .A1(\top_ihp.oisc.decoder.decoded[7] ),
    .B1(_05247_),
    .X(_00370_));
 sg13g2_nand2_1 _21780_ (.Y(_05248_),
    .A(_09902_),
    .B(_08982_));
 sg13g2_o21ai_1 _21781_ (.B1(_05248_),
    .Y(_00371_),
    .A1(_08981_),
    .A2(_09987_));
 sg13g2_mux2_1 _21782_ (.A0(_09919_),
    .A1(_10018_),
    .S(net737),
    .X(_00372_));
 sg13g2_nand2_1 _21783_ (.Y(_05249_),
    .A(_09999_),
    .B(net750));
 sg13g2_o21ai_1 _21784_ (.B1(_05249_),
    .Y(_00373_),
    .A1(net751),
    .A2(_05139_));
 sg13g2_nand2_1 _21785_ (.Y(_05250_),
    .A(_10092_),
    .B(net750));
 sg13g2_o21ai_1 _21786_ (.B1(_05250_),
    .Y(_00374_),
    .A1(_08981_),
    .A2(net731));
 sg13g2_nand2_1 _21787_ (.Y(_05251_),
    .A(_09968_),
    .B(net750));
 sg13g2_o21ai_1 _21788_ (.B1(_05251_),
    .Y(_00375_),
    .A1(net751),
    .A2(_05119_));
 sg13g2_nand2_1 _21789_ (.Y(_05252_),
    .A(\top_ihp.oisc.decoder.instruction[16] ),
    .B(net744));
 sg13g2_o21ai_1 _21790_ (.B1(_05252_),
    .Y(_00376_),
    .A1(net745),
    .A2(_09868_));
 sg13g2_nand2_1 _21791_ (.Y(_05253_),
    .A(\top_ihp.oisc.decoder.instruction[17] ),
    .B(net744));
 sg13g2_o21ai_1 _21792_ (.B1(_05253_),
    .Y(_00377_),
    .A1(net745),
    .A2(_10215_));
 sg13g2_nand2_1 _21793_ (.Y(_05254_),
    .A(\top_ihp.oisc.decoder.instruction[18] ),
    .B(net744));
 sg13g2_o21ai_1 _21794_ (.B1(_05254_),
    .Y(_00378_),
    .A1(net745),
    .A2(_10235_));
 sg13g2_nand2_1 _21795_ (.Y(_05255_),
    .A(\top_ihp.oisc.decoder.instruction[19] ),
    .B(_05183_));
 sg13g2_o21ai_1 _21796_ (.B1(_05255_),
    .Y(_00379_),
    .A1(_05146_),
    .A2(_10257_));
 sg13g2_mux2_1 _21797_ (.A0(_09796_),
    .A1(_10338_),
    .S(net737),
    .X(_00380_));
 sg13g2_mux2_1 _21798_ (.A0(_10279_),
    .A1(_10352_),
    .S(net737),
    .X(_00381_));
 sg13g2_mux2_1 _21799_ (.A0(_10374_),
    .A1(_10370_),
    .S(net737),
    .X(_00382_));
 sg13g2_nand2_1 _21800_ (.Y(_05256_),
    .A(_10387_),
    .B(_05183_));
 sg13g2_o21ai_1 _21801_ (.B1(_05256_),
    .Y(_00383_),
    .A1(_05146_),
    .A2(_09967_));
 sg13g2_mux2_1 _21802_ (.A0(_10395_),
    .A1(_09836_),
    .S(net737),
    .X(_00384_));
 sg13g2_mux2_1 _21803_ (.A0(_10418_),
    .A1(_10295_),
    .S(_05132_),
    .X(_00385_));
 sg13g2_nand2_1 _21804_ (.Y(_05257_),
    .A(_10435_),
    .B(net744));
 sg13g2_o21ai_1 _21805_ (.B1(_05257_),
    .Y(_00386_),
    .A1(net745),
    .A2(_09996_));
 sg13g2_mux2_1 _21806_ (.A0(\top_ihp.oisc.decoder.instruction[27] ),
    .A1(_10025_),
    .S(_05132_),
    .X(_00387_));
 sg13g2_mux2_1 _21807_ (.A0(\top_ihp.oisc.decoder.instruction[28] ),
    .A1(_10077_),
    .S(_03737_),
    .X(_00388_));
 sg13g2_mux2_1 _21808_ (.A0(\top_ihp.oisc.decoder.instruction[29] ),
    .A1(_10106_),
    .S(_03737_),
    .X(_00389_));
 sg13g2_mux2_1 _21809_ (.A0(\top_ihp.oisc.decoder.instruction[30] ),
    .A1(_10139_),
    .S(net747),
    .X(_00390_));
 sg13g2_nor2_1 _21810_ (.A(net906),
    .B(_10512_),
    .Y(_05258_));
 sg13g2_mux2_1 _21811_ (.A0(_10043_),
    .A1(_05258_),
    .S(net747),
    .X(_00391_));
 sg13g2_mux2_1 _21812_ (.A0(_09794_),
    .A1(_10650_),
    .S(net747),
    .X(_00392_));
 sg13g2_nand2_1 _21813_ (.Y(_05259_),
    .A(_09930_),
    .B(net744));
 sg13g2_o21ai_1 _21814_ (.B1(_05259_),
    .Y(_00393_),
    .A1(net745),
    .A2(_09842_));
 sg13g2_nand2_1 _21815_ (.Y(_05260_),
    .A(_09906_),
    .B(net744));
 sg13g2_o21ai_1 _21816_ (.B1(_05260_),
    .Y(_00394_),
    .A1(net745),
    .A2(_10303_));
 sg13g2_inv_2 _21817_ (.Y(_05261_),
    .A(_09923_));
 sg13g2_nand2_1 _21818_ (.Y(_05262_),
    .A(_09933_),
    .B(_08987_));
 sg13g2_nand3b_1 _21819_ (.B(net1036),
    .C(_09797_),
    .Y(_05263_),
    .A_N(_09803_));
 sg13g2_buf_2 _21820_ (.A(_05263_),
    .X(_05264_));
 sg13g2_nand3b_1 _21821_ (.B(_05264_),
    .C(net1037),
    .Y(_05265_),
    .A_N(_00234_));
 sg13g2_o21ai_1 _21822_ (.B1(_05265_),
    .Y(_05266_),
    .A1(_09366_),
    .A2(_05262_));
 sg13g2_buf_2 _21823_ (.A(_05266_),
    .X(_05267_));
 sg13g2_a21oi_1 _21824_ (.A1(_08412_),
    .A2(_08978_),
    .Y(_05268_),
    .B1(_05267_));
 sg13g2_a21oi_2 _21825_ (.B1(_05268_),
    .Y(_05269_),
    .A2(_10215_),
    .A1(_03736_));
 sg13g2_nand2_1 _21826_ (.Y(_05270_),
    .A(_05261_),
    .B(_05269_));
 sg13g2_buf_2 _21827_ (.A(_05270_),
    .X(_05271_));
 sg13g2_buf_8 _21828_ (.A(_05271_),
    .X(_05272_));
 sg13g2_inv_2 _21829_ (.Y(_05273_),
    .A(\top_ihp.oisc.micro_op[12] ));
 sg13g2_nand3_1 _21830_ (.B(_09796_),
    .C(_05264_),
    .A(net1037),
    .Y(_05274_));
 sg13g2_buf_2 _21831_ (.A(_05274_),
    .X(_05275_));
 sg13g2_o21ai_1 _21832_ (.B1(_05275_),
    .Y(_05276_),
    .A1(_05273_),
    .A2(_05262_));
 sg13g2_a21oi_1 _21833_ (.A1(_08412_),
    .A2(net793),
    .Y(_05277_),
    .B1(_05276_));
 sg13g2_a21o_1 _21834_ (.A2(_03736_),
    .A1(_08972_),
    .B1(_05277_),
    .X(_05278_));
 sg13g2_buf_2 _21835_ (.A(_05278_),
    .X(_05279_));
 sg13g2_nand2_1 _21836_ (.Y(_05280_),
    .A(_05261_),
    .B(_05279_));
 sg13g2_buf_8 _21837_ (.A(_05280_),
    .X(_05281_));
 sg13g2_buf_8 _21838_ (.A(_05281_),
    .X(_05282_));
 sg13g2_nor2_1 _21839_ (.A(_09782_),
    .B(_08991_),
    .Y(_05283_));
 sg13g2_buf_2 _21840_ (.A(_05283_),
    .X(_05284_));
 sg13g2_nor2_1 _21841_ (.A(_09913_),
    .B(_00236_),
    .Y(_05285_));
 sg13g2_nand2_2 _21842_ (.Y(_05286_),
    .A(_05264_),
    .B(_05285_));
 sg13g2_nor3_1 _21843_ (.A(_09923_),
    .B(_05284_),
    .C(_05286_),
    .Y(_05287_));
 sg13g2_nand3_1 _21844_ (.B(_05261_),
    .C(net793),
    .A(net1028),
    .Y(_05288_));
 sg13g2_nor2_1 _21845_ (.A(_10257_),
    .B(_05288_),
    .Y(_05289_));
 sg13g2_a21oi_1 _21846_ (.A1(_08980_),
    .A2(_05287_),
    .Y(_05290_),
    .B1(_05289_));
 sg13g2_buf_2 _21847_ (.A(_05290_),
    .X(_05291_));
 sg13g2_buf_2 _21848_ (.A(_05291_),
    .X(_05292_));
 sg13g2_inv_1 _21849_ (.Y(_05293_),
    .A(_00235_));
 sg13g2_and2_1 _21850_ (.A(net1037),
    .B(_05264_),
    .X(_05294_));
 sg13g2_buf_1 _21851_ (.A(_05294_),
    .X(_05295_));
 sg13g2_a22oi_1 _21852_ (.Y(_05296_),
    .B1(_05284_),
    .B2(\top_ihp.oisc.micro_op[15] ),
    .A2(_05295_),
    .A1(_05293_));
 sg13g2_mux2_1 _21853_ (.A0(_10235_),
    .A1(_05296_),
    .S(_08979_),
    .X(_05297_));
 sg13g2_buf_2 _21854_ (.A(_05297_),
    .X(_05298_));
 sg13g2_nor2_1 _21855_ (.A(net1000),
    .B(_05298_),
    .Y(_05299_));
 sg13g2_buf_2 _21856_ (.A(_05299_),
    .X(_05300_));
 sg13g2_inv_1 _21857_ (.Y(_05301_),
    .A(_00233_));
 sg13g2_a22oi_1 _21858_ (.Y(_05302_),
    .B1(_05284_),
    .B2(\top_ihp.oisc.micro_op[13] ),
    .A2(_05295_),
    .A1(_05301_));
 sg13g2_buf_2 _21859_ (.A(_05302_),
    .X(_05303_));
 sg13g2_mux2_1 _21860_ (.A0(_09868_),
    .A1(net841),
    .S(_08980_),
    .X(_05304_));
 sg13g2_or2_1 _21861_ (.X(_05305_),
    .B(_05304_),
    .A(_09923_));
 sg13g2_buf_8 _21862_ (.A(_05305_),
    .X(_05306_));
 sg13g2_nand2_1 _21863_ (.Y(_05307_),
    .A(_05300_),
    .B(_05306_));
 sg13g2_buf_2 _21864_ (.A(_05307_),
    .X(_05308_));
 sg13g2_nor4_2 _21865_ (.A(net709),
    .B(net685),
    .C(net708),
    .Y(_05309_),
    .D(_05308_));
 sg13g2_buf_8 _21866_ (.A(_05309_),
    .X(_05310_));
 sg13g2_buf_8 _21867_ (.A(net452),
    .X(_05311_));
 sg13g2_a21o_1 _21868_ (.A2(_10215_),
    .A1(_03736_),
    .B1(_05268_),
    .X(_05312_));
 sg13g2_buf_2 _21869_ (.A(_05312_),
    .X(_05313_));
 sg13g2_nor2_1 _21870_ (.A(_09923_),
    .B(_05313_),
    .Y(_05314_));
 sg13g2_buf_2 _21871_ (.A(_05314_),
    .X(_05315_));
 sg13g2_nand2_1 _21872_ (.Y(_05316_),
    .A(_05315_),
    .B(_05300_));
 sg13g2_buf_2 _21873_ (.A(_05316_),
    .X(_05317_));
 sg13g2_a21oi_1 _21874_ (.A1(_08972_),
    .A2(_03736_),
    .Y(_05318_),
    .B1(_05277_));
 sg13g2_buf_2 _21875_ (.A(_05318_),
    .X(_05319_));
 sg13g2_nor2_2 _21876_ (.A(net1000),
    .B(_05319_),
    .Y(_05320_));
 sg13g2_a21oi_1 _21877_ (.A1(net1028),
    .A2(net793),
    .Y(_05321_),
    .B1(_05284_));
 sg13g2_a22oi_1 _21878_ (.Y(_05322_),
    .B1(_05286_),
    .B2(_05321_),
    .A2(_10257_),
    .A1(_03736_));
 sg13g2_nor2_2 _21879_ (.A(net1000),
    .B(_05322_),
    .Y(_05323_));
 sg13g2_nand3_1 _21880_ (.B(_05306_),
    .C(_05323_),
    .A(_05320_),
    .Y(_05324_));
 sg13g2_buf_2 _21881_ (.A(_05324_),
    .X(_05325_));
 sg13g2_nor2_2 _21882_ (.A(_05317_),
    .B(_05325_),
    .Y(_05326_));
 sg13g2_buf_8 _21883_ (.A(_05326_),
    .X(_05327_));
 sg13g2_buf_8 _21884_ (.A(net338),
    .X(_05328_));
 sg13g2_or2_1 _21885_ (.X(_05329_),
    .B(_05322_),
    .A(net1000));
 sg13g2_buf_1 _21886_ (.A(_05329_),
    .X(_05330_));
 sg13g2_buf_1 _21887_ (.A(_05330_),
    .X(_05331_));
 sg13g2_or2_1 _21888_ (.X(_05332_),
    .B(_05298_),
    .A(_09923_));
 sg13g2_buf_8 _21889_ (.A(_05332_),
    .X(_05333_));
 sg13g2_nand2_1 _21890_ (.Y(_05334_),
    .A(_05315_),
    .B(_05333_));
 sg13g2_buf_2 _21891_ (.A(_05334_),
    .X(_05335_));
 sg13g2_nor4_1 _21892_ (.A(_05281_),
    .B(_05306_),
    .C(net707),
    .D(_05335_),
    .Y(_05336_));
 sg13g2_buf_1 _21893_ (.A(_05336_),
    .X(_05337_));
 sg13g2_buf_1 _21894_ (.A(_05337_),
    .X(_05338_));
 sg13g2_and2_1 _21895_ (.A(\top_ihp.oisc.regs[38][0] ),
    .B(net194),
    .X(_05339_));
 sg13g2_a221oi_1 _21896_ (.B2(\top_ihp.oisc.regs[44][0] ),
    .C1(_05339_),
    .B1(net195),
    .A1(\top_ihp.oisc.regs[60][0] ),
    .Y(_05340_),
    .A2(net339));
 sg13g2_buf_8 _21897_ (.A(_05315_),
    .X(_05341_));
 sg13g2_buf_8 _21898_ (.A(net684),
    .X(_05342_));
 sg13g2_buf_8 _21899_ (.A(_05300_),
    .X(_05343_));
 sg13g2_buf_8 _21900_ (.A(net706),
    .X(_05344_));
 sg13g2_nand2_1 _21901_ (.Y(_05345_),
    .A(_05273_),
    .B(_05275_));
 sg13g2_and2_1 _21902_ (.A(_05264_),
    .B(_05285_),
    .X(_05346_));
 sg13g2_buf_1 _21903_ (.A(_05346_),
    .X(_05347_));
 sg13g2_nand3_1 _21904_ (.B(_05284_),
    .C(_05347_),
    .A(_05261_),
    .Y(_05348_));
 sg13g2_buf_1 _21905_ (.A(_05348_),
    .X(_05349_));
 sg13g2_a21o_1 _21906_ (.A2(net793),
    .A1(net1028),
    .B1(_05349_),
    .X(_05350_));
 sg13g2_buf_1 _21907_ (.A(_05350_),
    .X(_05351_));
 sg13g2_nor2_1 _21908_ (.A(_05345_),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_buf_1 _21909_ (.A(_05352_),
    .X(_05353_));
 sg13g2_nand2_1 _21910_ (.Y(_05354_),
    .A(net841),
    .B(net724));
 sg13g2_buf_2 _21911_ (.A(_05354_),
    .X(_05355_));
 sg13g2_nor3_1 _21912_ (.A(net615),
    .B(net683),
    .C(_05355_),
    .Y(_05356_));
 sg13g2_buf_2 _21913_ (.A(_05356_),
    .X(_05357_));
 sg13g2_buf_8 _21914_ (.A(_05320_),
    .X(_05358_));
 sg13g2_buf_8 _21915_ (.A(net705),
    .X(_05359_));
 sg13g2_buf_8 _21916_ (.A(net682),
    .X(_05360_));
 sg13g2_mux2_1 _21917_ (.A0(\top_ihp.oisc.regs[15][0] ),
    .A1(\top_ihp.oisc.regs[14][0] ),
    .S(net614),
    .X(_05361_));
 sg13g2_buf_8 _21918_ (.A(_05333_),
    .X(_05362_));
 sg13g2_buf_2 _21919_ (.A(net704),
    .X(_05363_));
 sg13g2_a21oi_1 _21920_ (.A1(_08413_),
    .A2(net793),
    .Y(_05364_),
    .B1(_05262_));
 sg13g2_buf_1 _21921_ (.A(_05364_),
    .X(_05365_));
 sg13g2_nor2_1 _21922_ (.A(_09923_),
    .B(_05347_),
    .Y(_05366_));
 sg13g2_nand3_1 _21923_ (.B(net743),
    .C(_05366_),
    .A(_05267_),
    .Y(_05367_));
 sg13g2_buf_2 _21924_ (.A(_05367_),
    .X(_05368_));
 sg13g2_inv_1 _21925_ (.Y(_05369_),
    .A(\top_ihp.oisc.micro_op[13] ));
 sg13g2_nand3_1 _21926_ (.B(_05301_),
    .C(_05264_),
    .A(net1037),
    .Y(_05370_));
 sg13g2_o21ai_1 _21927_ (.B1(_05370_),
    .Y(_05371_),
    .A1(_05369_),
    .A2(_05262_));
 sg13g2_buf_1 _21928_ (.A(_05371_),
    .X(_05372_));
 sg13g2_buf_2 _21929_ (.A(_05372_),
    .X(_05373_));
 sg13g2_nand2b_1 _21930_ (.Y(_05374_),
    .B(net840),
    .A_N(_05368_));
 sg13g2_buf_2 _21931_ (.A(_05374_),
    .X(_05375_));
 sg13g2_nor2_2 _21932_ (.A(_05363_),
    .B(_05375_),
    .Y(_05376_));
 sg13g2_a22oi_1 _21933_ (.Y(_05377_),
    .B1(_05361_),
    .B2(_05376_),
    .A2(_05357_),
    .A1(\top_ihp.oisc.regs[16][0] ));
 sg13g2_or2_1 _21934_ (.X(_05378_),
    .B(_05368_),
    .A(net840));
 sg13g2_buf_2 _21935_ (.A(_05378_),
    .X(_05379_));
 sg13g2_nor3_1 _21936_ (.A(net705),
    .B(net706),
    .C(_05379_),
    .Y(_05380_));
 sg13g2_buf_2 _21937_ (.A(_05380_),
    .X(_05381_));
 sg13g2_buf_1 _21938_ (.A(_05381_),
    .X(_05382_));
 sg13g2_nor3_1 _21939_ (.A(net705),
    .B(net683),
    .C(_05375_),
    .Y(_05383_));
 sg13g2_buf_1 _21940_ (.A(_05383_),
    .X(_05384_));
 sg13g2_a22oi_1 _21941_ (.Y(_05385_),
    .B1(net451),
    .B2(\top_ihp.oisc.regs[7][0] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][0] ));
 sg13g2_buf_8 _21942_ (.A(_05281_),
    .X(_05386_));
 sg13g2_nor3_1 _21943_ (.A(net680),
    .B(net683),
    .C(_05375_),
    .Y(_05387_));
 sg13g2_buf_1 _21944_ (.A(_05387_),
    .X(_05388_));
 sg13g2_nor3_1 _21945_ (.A(net709),
    .B(net683),
    .C(_05355_),
    .Y(_05389_));
 sg13g2_buf_1 _21946_ (.A(_05389_),
    .X(_05390_));
 sg13g2_a22oi_1 _21947_ (.Y(_05391_),
    .B1(net449),
    .B2(\top_ihp.oisc.regs[20][0] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[6][0] ));
 sg13g2_nor3_1 _21948_ (.A(_05267_),
    .B(_05347_),
    .C(_05372_),
    .Y(_05392_));
 sg13g2_a21oi_2 _21949_ (.B1(net948),
    .Y(_05393_),
    .A2(_05392_),
    .A1(net743));
 sg13g2_nor3_1 _21950_ (.A(_05281_),
    .B(_05333_),
    .C(_05393_),
    .Y(_05394_));
 sg13g2_buf_2 _21951_ (.A(_05394_),
    .X(_05395_));
 sg13g2_nor3_2 _21952_ (.A(net680),
    .B(net704),
    .C(_05379_),
    .Y(_05396_));
 sg13g2_buf_1 _21953_ (.A(_05396_),
    .X(_05397_));
 sg13g2_a22oi_1 _21954_ (.Y(_05398_),
    .B1(net448),
    .B2(\top_ihp.oisc.regs[12][0] ),
    .A2(_05395_),
    .A1(\top_ihp.oisc.regs[8][0] ));
 sg13g2_nand4_1 _21955_ (.B(_05385_),
    .C(_05391_),
    .A(_05377_),
    .Y(_05399_),
    .D(_05398_));
 sg13g2_buf_8 _21956_ (.A(_05333_),
    .X(_05400_));
 sg13g2_nor3_1 _21957_ (.A(net705),
    .B(net703),
    .C(_05379_),
    .Y(_05401_));
 sg13g2_buf_2 _21958_ (.A(_05401_),
    .X(_05402_));
 sg13g2_buf_1 _21959_ (.A(_05402_),
    .X(_05403_));
 sg13g2_buf_8 _21960_ (.A(_05282_),
    .X(_05404_));
 sg13g2_and2_1 _21961_ (.A(_05372_),
    .B(_05366_),
    .X(_05405_));
 sg13g2_and2_1 _21962_ (.A(net743),
    .B(_05405_),
    .X(_05406_));
 sg13g2_buf_2 _21963_ (.A(_05406_),
    .X(_05407_));
 sg13g2_nand2b_1 _21964_ (.Y(_05408_),
    .B(_05407_),
    .A_N(_05267_));
 sg13g2_buf_2 _21965_ (.A(_05408_),
    .X(_05409_));
 sg13g2_nor2_1 _21966_ (.A(net613),
    .B(_05409_),
    .Y(_05410_));
 sg13g2_mux2_1 _21967_ (.A0(\top_ihp.oisc.regs[10][0] ),
    .A1(\top_ihp.oisc.regs[2][0] ),
    .S(net681),
    .X(_05411_));
 sg13g2_a22oi_1 _21968_ (.Y(_05412_),
    .B1(_05410_),
    .B2(_05411_),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[13][0] ));
 sg13g2_nor3_1 _21969_ (.A(net705),
    .B(_05333_),
    .C(_05393_),
    .Y(_05413_));
 sg13g2_buf_2 _21970_ (.A(_05413_),
    .X(_05414_));
 sg13g2_buf_1 _21971_ (.A(_05414_),
    .X(_05415_));
 sg13g2_a21oi_1 _21972_ (.A1(_05313_),
    .A2(_05298_),
    .Y(_05416_),
    .B1(net1000));
 sg13g2_buf_1 _21973_ (.A(_05416_),
    .X(_05417_));
 sg13g2_nand2_1 _21974_ (.Y(_05418_),
    .A(net840),
    .B(net724));
 sg13g2_buf_2 _21975_ (.A(_05418_),
    .X(_05419_));
 sg13g2_nor2_1 _21976_ (.A(net702),
    .B(_05419_),
    .Y(_05420_));
 sg13g2_buf_1 _21977_ (.A(_05420_),
    .X(_05421_));
 sg13g2_buf_1 _21978_ (.A(_05421_),
    .X(_05422_));
 sg13g2_a22oi_1 _21979_ (.Y(_05423_),
    .B1(net335),
    .B2(\top_ihp.oisc.regs[18][0] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[9][0] ));
 sg13g2_nand2_1 _21980_ (.Y(_05424_),
    .A(_05412_),
    .B(_05423_));
 sg13g2_a21oi_1 _21981_ (.A1(_05298_),
    .A2(_05304_),
    .Y(_05425_),
    .B1(_09924_));
 sg13g2_buf_1 _21982_ (.A(_05425_),
    .X(_05426_));
 sg13g2_nand3_1 _21983_ (.B(_05279_),
    .C(_05323_),
    .A(_05271_),
    .Y(_05427_));
 sg13g2_buf_1 _21984_ (.A(_05427_),
    .X(_05428_));
 sg13g2_nor2_2 _21985_ (.A(net723),
    .B(_05428_),
    .Y(_05429_));
 sg13g2_buf_8 _21986_ (.A(_05429_),
    .X(_05430_));
 sg13g2_nand2_1 _21987_ (.Y(_05431_),
    .A(\top_ihp.oisc.regs[32][0] ),
    .B(_05430_));
 sg13g2_a221oi_1 _21988_ (.B2(_05273_),
    .C1(_05349_),
    .B1(_05275_),
    .A1(net984),
    .Y(_05432_),
    .A2(_09003_));
 sg13g2_buf_1 _21989_ (.A(_05432_),
    .X(_05433_));
 sg13g2_nand2_2 _21990_ (.Y(_05434_),
    .A(net840),
    .B(net742));
 sg13g2_nor2_1 _21991_ (.A(net702),
    .B(_05434_),
    .Y(_05435_));
 sg13g2_buf_2 _21992_ (.A(_05435_),
    .X(_05436_));
 sg13g2_buf_1 _21993_ (.A(_05436_),
    .X(_05437_));
 sg13g2_a22oi_1 _21994_ (.Y(_05438_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[19][0] ),
    .A2(net739),
    .A1(_08321_));
 sg13g2_and2_1 _21995_ (.A(net840),
    .B(net742),
    .X(_05439_));
 sg13g2_buf_2 _21996_ (.A(_05439_),
    .X(_05440_));
 sg13g2_nor3_1 _21997_ (.A(net1000),
    .B(_05269_),
    .C(_05298_),
    .Y(_05441_));
 sg13g2_buf_2 _21998_ (.A(_05441_),
    .X(_05442_));
 sg13g2_and2_1 _21999_ (.A(_05440_),
    .B(_05442_),
    .X(_05443_));
 sg13g2_buf_2 _22000_ (.A(_05443_),
    .X(_05444_));
 sg13g2_a21oi_2 _22001_ (.B1(_05349_),
    .Y(_05445_),
    .A2(net793),
    .A1(net984));
 sg13g2_and2_1 _22002_ (.A(_05273_),
    .B(_05275_),
    .X(_05446_));
 sg13g2_nor2_1 _22003_ (.A(_05373_),
    .B(_05446_),
    .Y(_05447_));
 sg13g2_nand2_1 _22004_ (.Y(_05448_),
    .A(_05445_),
    .B(_05447_));
 sg13g2_nor3_1 _22005_ (.A(net709),
    .B(net706),
    .C(_05448_),
    .Y(_05449_));
 sg13g2_buf_2 _22006_ (.A(_05449_),
    .X(_05450_));
 sg13g2_buf_1 _22007_ (.A(_05450_),
    .X(_05451_));
 sg13g2_a22oi_1 _22008_ (.Y(_05452_),
    .B1(net444),
    .B2(\top_ihp.oisc.regs[21][0] ),
    .A2(_05444_),
    .A1(\top_ihp.oisc.regs[27][0] ));
 sg13g2_nor3_1 _22009_ (.A(net682),
    .B(net704),
    .C(_05409_),
    .Y(_05453_));
 sg13g2_buf_1 _22010_ (.A(_05453_),
    .X(_05454_));
 sg13g2_nor3_2 _22011_ (.A(_05313_),
    .B(_05362_),
    .C(_05355_),
    .Y(_05455_));
 sg13g2_buf_1 _22012_ (.A(_05455_),
    .X(_05456_));
 sg13g2_a22oi_1 _22013_ (.Y(_05457_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[28][0] ),
    .A2(_05454_),
    .A1(\top_ihp.oisc.regs[11][0] ));
 sg13g2_nand4_1 _22014_ (.B(_05438_),
    .C(_05452_),
    .A(_05431_),
    .Y(_05458_),
    .D(_05457_));
 sg13g2_nor4_1 _22015_ (.A(net684),
    .B(net705),
    .C(net708),
    .D(net723),
    .Y(_05459_));
 sg13g2_buf_1 _22016_ (.A(_05459_),
    .X(_05460_));
 sg13g2_nor2_1 _22017_ (.A(_05271_),
    .B(_05281_),
    .Y(_05461_));
 sg13g2_buf_2 _22018_ (.A(_05461_),
    .X(_05462_));
 sg13g2_nor3_2 _22019_ (.A(_05291_),
    .B(_05333_),
    .C(_05306_),
    .Y(_05463_));
 sg13g2_and2_1 _22020_ (.A(_05462_),
    .B(_05463_),
    .X(_05464_));
 sg13g2_buf_2 _22021_ (.A(_05464_),
    .X(_05465_));
 sg13g2_buf_1 _22022_ (.A(_05465_),
    .X(_05466_));
 sg13g2_a22oi_1 _22023_ (.Y(_05467_),
    .B1(net193),
    .B2(\top_ihp.oisc.regs[62][0] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][0] ));
 sg13g2_nand2_1 _22024_ (.Y(_05468_),
    .A(_05315_),
    .B(_05319_));
 sg13g2_buf_8 _22025_ (.A(_05468_),
    .X(_05469_));
 sg13g2_nor3_1 _22026_ (.A(net707),
    .B(net612),
    .C(net723),
    .Y(_05470_));
 sg13g2_buf_2 _22027_ (.A(_05470_),
    .X(_05471_));
 sg13g2_buf_1 _22028_ (.A(_05471_),
    .X(_05472_));
 sg13g2_nor2_1 _22029_ (.A(_09924_),
    .B(_05304_),
    .Y(_05473_));
 sg13g2_buf_2 _22030_ (.A(_05473_),
    .X(_05474_));
 sg13g2_nand2_1 _22031_ (.Y(_05475_),
    .A(_05300_),
    .B(_05474_));
 sg13g2_nand2_2 _22032_ (.Y(_05476_),
    .A(_05271_),
    .B(_05319_));
 sg13g2_nor3_1 _22033_ (.A(net707),
    .B(_05475_),
    .C(_05476_),
    .Y(_05477_));
 sg13g2_buf_2 _22034_ (.A(_05477_),
    .X(_05478_));
 sg13g2_buf_8 _22035_ (.A(_05478_),
    .X(_05479_));
 sg13g2_a22oi_1 _22036_ (.Y(_05480_),
    .B1(net440),
    .B2(\top_ihp.oisc.regs[43][0] ),
    .A2(_05472_),
    .A1(\top_ihp.oisc.regs[37][0] ));
 sg13g2_nand2_1 _22037_ (.Y(_05481_),
    .A(_05467_),
    .B(_05480_));
 sg13g2_nor4_1 _22038_ (.A(_05399_),
    .B(_05424_),
    .C(_05458_),
    .D(_05481_),
    .Y(_05482_));
 sg13g2_nor2_1 _22039_ (.A(_05428_),
    .B(_05475_),
    .Y(_05483_));
 sg13g2_buf_2 _22040_ (.A(_05483_),
    .X(_05484_));
 sg13g2_buf_8 _22041_ (.A(_05484_),
    .X(_05485_));
 sg13g2_buf_1 _22042_ (.A(net334),
    .X(_05486_));
 sg13g2_nor3_1 _22043_ (.A(_05358_),
    .B(net706),
    .C(_05393_),
    .Y(_05487_));
 sg13g2_buf_2 _22044_ (.A(_05487_),
    .X(_05488_));
 sg13g2_buf_8 _22045_ (.A(_05488_),
    .X(_05489_));
 sg13g2_nand2_1 _22046_ (.Y(_05490_),
    .A(\top_ihp.oisc.regs[1][0] ),
    .B(net439));
 sg13g2_nand2_1 _22047_ (.Y(_05491_),
    .A(_05271_),
    .B(_05300_));
 sg13g2_nor2_1 _22048_ (.A(_05419_),
    .B(_05491_),
    .Y(_05492_));
 sg13g2_buf_2 _22049_ (.A(_05492_),
    .X(_05493_));
 sg13g2_buf_1 _22050_ (.A(_05493_),
    .X(_05494_));
 sg13g2_nor3_2 _22051_ (.A(net709),
    .B(_05344_),
    .C(_05434_),
    .Y(_05495_));
 sg13g2_buf_8 _22052_ (.A(_05495_),
    .X(_05496_));
 sg13g2_a22oi_1 _22053_ (.Y(_05497_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][0] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[26][0] ));
 sg13g2_nand2_1 _22054_ (.Y(_05498_),
    .A(_05281_),
    .B(_05333_));
 sg13g2_nor2_1 _22055_ (.A(_05498_),
    .B(_05409_),
    .Y(_05499_));
 sg13g2_buf_2 _22056_ (.A(_05499_),
    .X(_05500_));
 sg13g2_buf_8 _22057_ (.A(_05500_),
    .X(_05501_));
 sg13g2_nor3_1 _22058_ (.A(net709),
    .B(net703),
    .C(_05434_),
    .Y(_05502_));
 sg13g2_buf_1 _22059_ (.A(_05502_),
    .X(_05503_));
 sg13g2_buf_2 _22060_ (.A(net611),
    .X(_05504_));
 sg13g2_a22oi_1 _22061_ (.Y(_05505_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[31][0] ),
    .A2(net332),
    .A1(\top_ihp.oisc.regs[3][0] ));
 sg13g2_nor3_1 _22062_ (.A(net680),
    .B(net683),
    .C(_05379_),
    .Y(_05506_));
 sg13g2_buf_1 _22063_ (.A(_05506_),
    .X(_05507_));
 sg13g2_buf_2 _22064_ (.A(_05491_),
    .X(_05508_));
 sg13g2_buf_1 _22065_ (.A(_05448_),
    .X(_05509_));
 sg13g2_nor2_2 _22066_ (.A(net679),
    .B(net734),
    .Y(_05510_));
 sg13g2_a22oi_1 _22067_ (.Y(_05511_),
    .B1(_05510_),
    .B2(\top_ihp.oisc.regs[25][0] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[4][0] ));
 sg13g2_nand4_1 _22068_ (.B(_05497_),
    .C(_05505_),
    .A(_05490_),
    .Y(_05512_),
    .D(_05511_));
 sg13g2_a21oi_1 _22069_ (.A1(\top_ihp.oisc.regs[42][0] ),
    .A2(_05486_),
    .Y(_05513_),
    .B1(_05512_));
 sg13g2_nand2_1 _22070_ (.Y(_05514_),
    .A(_05333_),
    .B(_05474_));
 sg13g2_nor4_1 _22071_ (.A(net709),
    .B(net685),
    .C(net708),
    .D(_05514_),
    .Y(_05515_));
 sg13g2_buf_2 _22072_ (.A(_05515_),
    .X(_05516_));
 sg13g2_nand2_1 _22073_ (.Y(_05517_),
    .A(_05300_),
    .B(_05323_));
 sg13g2_buf_2 _22074_ (.A(_05517_),
    .X(_05518_));
 sg13g2_nor4_2 _22075_ (.A(net684),
    .B(_05319_),
    .C(_05474_),
    .Y(_05519_),
    .D(_05518_));
 sg13g2_buf_1 _22076_ (.A(_05519_),
    .X(_05520_));
 sg13g2_a22oi_1 _22077_ (.Y(_05521_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[40][0] ),
    .A2(_05516_),
    .A1(\top_ihp.oisc.regs[54][0] ));
 sg13g2_nor4_1 _22078_ (.A(net685),
    .B(_05291_),
    .C(_05306_),
    .D(net702),
    .Y(_05522_));
 sg13g2_buf_2 _22079_ (.A(_05522_),
    .X(_05523_));
 sg13g2_nor3_1 _22080_ (.A(_05474_),
    .B(_05518_),
    .C(net612),
    .Y(_05524_));
 sg13g2_buf_2 _22081_ (.A(_05524_),
    .X(_05525_));
 sg13g2_a22oi_1 _22082_ (.Y(_05526_),
    .B1(_05525_),
    .B2(\top_ihp.oisc.regs[45][0] ),
    .A2(_05523_),
    .A1(\top_ihp.oisc.regs[50][0] ));
 sg13g2_nor4_1 _22083_ (.A(net684),
    .B(net705),
    .C(_05330_),
    .D(net723),
    .Y(_05527_));
 sg13g2_buf_2 _22084_ (.A(_05527_),
    .X(_05528_));
 sg13g2_buf_1 _22085_ (.A(_05292_),
    .X(_05529_));
 sg13g2_buf_8 _22086_ (.A(_05306_),
    .X(_05530_));
 sg13g2_nand2_2 _22087_ (.Y(_05531_),
    .A(net682),
    .B(net701));
 sg13g2_nor3_2 _22088_ (.A(net678),
    .B(_05531_),
    .C(_05335_),
    .Y(_05532_));
 sg13g2_a22oi_1 _22089_ (.Y(_05533_),
    .B1(_05532_),
    .B2(\top_ihp.oisc.regs[52][0] ),
    .A2(_05528_),
    .A1(\top_ihp.oisc.regs[33][0] ));
 sg13g2_nor2_1 _22090_ (.A(_05271_),
    .B(_05279_),
    .Y(_05534_));
 sg13g2_buf_2 _22091_ (.A(_05534_),
    .X(_05535_));
 sg13g2_and2_1 _22092_ (.A(_05535_),
    .B(_05463_),
    .X(_05536_));
 sg13g2_buf_2 _22093_ (.A(_05536_),
    .X(_05537_));
 sg13g2_nor4_1 _22094_ (.A(_05291_),
    .B(net706),
    .C(_05306_),
    .D(net612),
    .Y(_05538_));
 sg13g2_buf_2 _22095_ (.A(_05538_),
    .X(_05539_));
 sg13g2_a22oi_1 _22096_ (.Y(_05540_),
    .B1(_05539_),
    .B2(\top_ihp.oisc.regs[55][0] ),
    .A2(_05537_),
    .A1(\top_ihp.oisc.regs[63][0] ));
 sg13g2_nand4_1 _22097_ (.B(_05526_),
    .C(_05533_),
    .A(_05521_),
    .Y(_05541_),
    .D(_05540_));
 sg13g2_nor3_1 _22098_ (.A(net708),
    .B(_05308_),
    .C(net612),
    .Y(_05542_));
 sg13g2_buf_2 _22099_ (.A(_05542_),
    .X(_05543_));
 sg13g2_nor4_2 _22100_ (.A(net684),
    .B(net685),
    .C(net708),
    .Y(_05544_),
    .D(_05475_));
 sg13g2_a22oi_1 _22101_ (.Y(_05545_),
    .B1(_05544_),
    .B2(\top_ihp.oisc.regs[58][0] ),
    .A2(_05543_),
    .A1(\top_ihp.oisc.regs[61][0] ));
 sg13g2_o21ai_1 _22102_ (.B1(_05287_),
    .Y(_05546_),
    .A1(_08615_),
    .A2(_03720_));
 sg13g2_o21ai_1 _22103_ (.B1(_05546_),
    .Y(_05547_),
    .A1(_10257_),
    .A2(_05288_));
 sg13g2_buf_2 _22104_ (.A(_05547_),
    .X(_05548_));
 sg13g2_o21ai_1 _22105_ (.B1(_05548_),
    .Y(_05549_),
    .A1(net948),
    .A2(_05313_));
 sg13g2_nor3_1 _22106_ (.A(net680),
    .B(net723),
    .C(_05549_),
    .Y(_05550_));
 sg13g2_buf_2 _22107_ (.A(_05550_),
    .X(_05551_));
 sg13g2_nor4_1 _22108_ (.A(net706),
    .B(_05306_),
    .C(net707),
    .D(net612),
    .Y(_05552_));
 sg13g2_buf_2 _22109_ (.A(_05552_),
    .X(_05553_));
 sg13g2_a22oi_1 _22110_ (.Y(_05554_),
    .B1(_05553_),
    .B2(\top_ihp.oisc.regs[39][0] ),
    .A2(_05551_),
    .A1(\top_ihp.oisc.regs[48][0] ));
 sg13g2_nor2_1 _22111_ (.A(_05315_),
    .B(_05320_),
    .Y(_05555_));
 sg13g2_buf_2 _22112_ (.A(_05555_),
    .X(_05556_));
 sg13g2_and2_1 _22113_ (.A(_05556_),
    .B(_05463_),
    .X(_05557_));
 sg13g2_buf_1 _22114_ (.A(_05557_),
    .X(_05558_));
 sg13g2_nor3_1 _22115_ (.A(net707),
    .B(_05476_),
    .C(_05514_),
    .Y(_05559_));
 sg13g2_buf_2 _22116_ (.A(_05559_),
    .X(_05560_));
 sg13g2_a22oi_1 _22117_ (.Y(_05561_),
    .B1(_05560_),
    .B2(\top_ihp.oisc.regs[35][0] ),
    .A2(_05558_),
    .A1(\top_ihp.oisc.regs[59][0] ));
 sg13g2_nor2_1 _22118_ (.A(_05428_),
    .B(_05514_),
    .Y(_05562_));
 sg13g2_buf_2 _22119_ (.A(_05562_),
    .X(_05563_));
 sg13g2_buf_8 _22120_ (.A(net709),
    .X(_05564_));
 sg13g2_buf_8 _22121_ (.A(net677),
    .X(_05565_));
 sg13g2_buf_8 _22122_ (.A(net706),
    .X(_05566_));
 sg13g2_nand2_1 _22123_ (.Y(_05567_),
    .A(_05446_),
    .B(_05445_));
 sg13g2_buf_2 _22124_ (.A(_05567_),
    .X(_05568_));
 sg13g2_nor2_1 _22125_ (.A(net840),
    .B(_05568_),
    .Y(_05569_));
 sg13g2_buf_2 _22126_ (.A(_05569_),
    .X(_05570_));
 sg13g2_nand3_1 _22127_ (.B(net676),
    .C(_05570_),
    .A(\top_ihp.oisc.regs[24][0] ),
    .Y(_05571_));
 sg13g2_buf_8 _22128_ (.A(net703),
    .X(_05572_));
 sg13g2_and2_1 _22129_ (.A(_05445_),
    .B(_05447_),
    .X(_05573_));
 sg13g2_buf_1 _22130_ (.A(_05573_),
    .X(_05574_));
 sg13g2_buf_1 _22131_ (.A(_05574_),
    .X(_05575_));
 sg13g2_nand3_1 _22132_ (.B(net675),
    .C(net722),
    .A(\top_ihp.oisc.regs[17][0] ),
    .Y(_05576_));
 sg13g2_nand3_1 _22133_ (.B(_05571_),
    .C(_05576_),
    .A(_05565_),
    .Y(_05577_));
 sg13g2_buf_8 _22134_ (.A(net615),
    .X(_05578_));
 sg13g2_nor2_1 _22135_ (.A(net841),
    .B(_05345_),
    .Y(_05579_));
 sg13g2_a22oi_1 _22136_ (.Y(_05580_),
    .B1(_05579_),
    .B2(\top_ihp.oisc.regs[30][0] ),
    .A2(_05447_),
    .A1(\top_ihp.oisc.regs[29][0] ));
 sg13g2_nand3b_1 _22137_ (.B(_05445_),
    .C(net676),
    .Y(_05581_),
    .A_N(_05580_));
 sg13g2_nor3_1 _22138_ (.A(net841),
    .B(_05345_),
    .C(_05351_),
    .Y(_05582_));
 sg13g2_nand3_1 _22139_ (.B(_05572_),
    .C(_05582_),
    .A(\top_ihp.oisc.regs[22][0] ),
    .Y(_05583_));
 sg13g2_nand3_1 _22140_ (.B(_05581_),
    .C(_05583_),
    .A(_05578_),
    .Y(_05584_));
 sg13g2_a22oi_1 _22141_ (.Y(_05585_),
    .B1(_05577_),
    .B2(_05584_),
    .A2(_05563_),
    .A1(\top_ihp.oisc.regs[34][0] ));
 sg13g2_nand4_1 _22142_ (.B(_05554_),
    .C(_05561_),
    .A(_05545_),
    .Y(_05586_),
    .D(_05585_));
 sg13g2_nor3_1 _22143_ (.A(net701),
    .B(_05518_),
    .C(net612),
    .Y(_05587_));
 sg13g2_buf_2 _22144_ (.A(_05587_),
    .X(_05588_));
 sg13g2_nor4_1 _22145_ (.A(net705),
    .B(_05400_),
    .C(_05474_),
    .D(_05549_),
    .Y(_05589_));
 sg13g2_buf_1 _22146_ (.A(_05589_),
    .X(_05590_));
 sg13g2_a22oi_1 _22147_ (.Y(_05591_),
    .B1(_05590_),
    .B2(\top_ihp.oisc.regs[57][0] ),
    .A2(_05588_),
    .A1(\top_ihp.oisc.regs[47][0] ));
 sg13g2_nor3_1 _22148_ (.A(net708),
    .B(net612),
    .C(net723),
    .Y(_05592_));
 sg13g2_buf_2 _22149_ (.A(_05592_),
    .X(_05593_));
 sg13g2_nor2_1 _22150_ (.A(_05325_),
    .B(_05335_),
    .Y(_05594_));
 sg13g2_buf_1 _22151_ (.A(_05594_),
    .X(_05595_));
 sg13g2_a22oi_1 _22152_ (.Y(_05596_),
    .B1(_05595_),
    .B2(\top_ihp.oisc.regs[36][0] ),
    .A2(_05593_),
    .A1(\top_ihp.oisc.regs[53][0] ));
 sg13g2_nor3_1 _22153_ (.A(net682),
    .B(_05514_),
    .C(_05549_),
    .Y(_05597_));
 sg13g2_buf_2 _22154_ (.A(_05597_),
    .X(_05598_));
 sg13g2_buf_8 _22155_ (.A(_05474_),
    .X(_05599_));
 sg13g2_nor4_2 _22156_ (.A(net615),
    .B(net614),
    .C(net700),
    .Y(_05600_),
    .D(_05518_));
 sg13g2_a22oi_1 _22157_ (.Y(_05601_),
    .B1(_05600_),
    .B2(\top_ihp.oisc.regs[41][0] ),
    .A2(_05598_),
    .A1(\top_ihp.oisc.regs[51][0] ));
 sg13g2_nor4_1 _22158_ (.A(net685),
    .B(net701),
    .C(_05317_),
    .D(net707),
    .Y(_05602_));
 sg13g2_buf_2 _22159_ (.A(_05602_),
    .X(_05603_));
 sg13g2_nor4_1 _22160_ (.A(net684),
    .B(net685),
    .C(net708),
    .D(_05308_),
    .Y(_05604_));
 sg13g2_buf_4 _22161_ (.X(_05605_),
    .A(_05604_));
 sg13g2_a22oi_1 _22162_ (.Y(_05606_),
    .B1(_05605_),
    .B2(\top_ihp.oisc.regs[56][0] ),
    .A2(_05603_),
    .A1(\top_ihp.oisc.regs[46][0] ));
 sg13g2_nand4_1 _22163_ (.B(_05596_),
    .C(_05601_),
    .A(_05591_),
    .Y(_05607_),
    .D(_05606_));
 sg13g2_a21o_1 _22164_ (.A2(net743),
    .A1(_05286_),
    .B1(net948),
    .X(_05608_));
 sg13g2_buf_1 _22165_ (.A(_05608_),
    .X(_05609_));
 sg13g2_nand2_2 _22166_ (.Y(_05610_),
    .A(net701),
    .B(_05609_));
 sg13g2_nor4_2 _22167_ (.A(net613),
    .B(_05535_),
    .C(_05610_),
    .Y(_05611_),
    .D(net702));
 sg13g2_buf_8 _22168_ (.A(_05611_),
    .X(_05612_));
 sg13g2_nor4_1 _22169_ (.A(_05541_),
    .B(_05586_),
    .C(_05607_),
    .D(net331),
    .Y(_05613_));
 sg13g2_and4_1 _22170_ (.A(_05340_),
    .B(_05482_),
    .C(_05513_),
    .D(_05613_),
    .X(_05614_));
 sg13g2_inv_1 _22171_ (.Y(_05615_),
    .A(\top_ihp.oisc.regs[0][0] ));
 sg13g2_buf_1 _22172_ (.A(_05611_),
    .X(_05616_));
 sg13g2_nand2_1 _22173_ (.Y(_05617_),
    .A(net677),
    .B(_05323_));
 sg13g2_nor2_1 _22174_ (.A(net948),
    .B(net743),
    .Y(_05618_));
 sg13g2_o21ai_1 _22175_ (.B1(_05618_),
    .Y(_05619_),
    .A1(_05426_),
    .A2(_05617_));
 sg13g2_nor2_1 _22176_ (.A(_05609_),
    .B(_05528_),
    .Y(_05620_));
 sg13g2_a21o_1 _22177_ (.A2(_05620_),
    .A1(_05619_),
    .B1(net739),
    .X(_05621_));
 sg13g2_buf_1 _22178_ (.A(_05621_),
    .X(_05622_));
 sg13g2_buf_1 _22179_ (.A(_05622_),
    .X(_05623_));
 sg13g2_a21oi_1 _22180_ (.A1(_05615_),
    .A2(net330),
    .Y(_05624_),
    .B1(net34));
 sg13g2_a21oi_1 _22181_ (.A1(_08321_),
    .A2(net718),
    .Y(_05625_),
    .B1(_05624_));
 sg13g2_nor2_1 _22182_ (.A(_05614_),
    .B(_05625_),
    .Y(_00420_));
 sg13g2_buf_2 _22183_ (.A(_05612_),
    .X(_05626_));
 sg13g2_buf_8 _22184_ (.A(_05523_),
    .X(_05627_));
 sg13g2_buf_1 _22185_ (.A(net329),
    .X(_05628_));
 sg13g2_nand2_1 _22186_ (.Y(_05629_),
    .A(\top_ihp.oisc.regs[50][10] ),
    .B(net189));
 sg13g2_buf_2 _22187_ (.A(_05543_),
    .X(_05630_));
 sg13g2_a22oi_1 _22188_ (.Y(_05631_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][10] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][10] ));
 sg13g2_buf_1 _22189_ (.A(_05337_),
    .X(_05632_));
 sg13g2_buf_8 _22190_ (.A(_05528_),
    .X(_05633_));
 sg13g2_buf_1 _22191_ (.A(net328),
    .X(_05634_));
 sg13g2_a22oi_1 _22192_ (.Y(_05635_),
    .B1(net186),
    .B2(\top_ihp.oisc.regs[33][10] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][10] ));
 sg13g2_buf_1 _22193_ (.A(_05558_),
    .X(_05636_));
 sg13g2_buf_8 _22194_ (.A(net185),
    .X(_05637_));
 sg13g2_a22oi_1 _22195_ (.Y(_05638_),
    .B1(net78),
    .B2(\top_ihp.oisc.regs[59][10] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[42][10] ));
 sg13g2_nand4_1 _22196_ (.B(_05631_),
    .C(_05635_),
    .A(_05629_),
    .Y(_05639_),
    .D(_05638_));
 sg13g2_buf_2 _22197_ (.A(net441),
    .X(_05640_));
 sg13g2_buf_8 _22198_ (.A(_05598_),
    .X(_05641_));
 sg13g2_buf_8 _22199_ (.A(net326),
    .X(_05642_));
 sg13g2_a22oi_1 _22200_ (.Y(_05643_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][10] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][10] ));
 sg13g2_buf_8 _22201_ (.A(_05560_),
    .X(_05644_));
 sg13g2_buf_8 _22202_ (.A(net433),
    .X(_05645_));
 sg13g2_buf_2 _22203_ (.A(net609),
    .X(_05646_));
 sg13g2_a22oi_1 _22204_ (.Y(_05647_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][10] ),
    .A2(net325),
    .A1(\top_ihp.oisc.regs[35][10] ));
 sg13g2_buf_8 _22205_ (.A(_05537_),
    .X(_05648_));
 sg13g2_buf_2 _22206_ (.A(_05648_),
    .X(_05649_));
 sg13g2_a22oi_1 _22207_ (.Y(_05650_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[63][10] ),
    .A2(_05430_),
    .A1(\top_ihp.oisc.regs[32][10] ));
 sg13g2_buf_8 _22208_ (.A(_05539_),
    .X(_05651_));
 sg13g2_buf_1 _22209_ (.A(net182),
    .X(_05652_));
 sg13g2_nor3_2 _22210_ (.A(_05474_),
    .B(_05518_),
    .C(_05476_),
    .Y(_05653_));
 sg13g2_buf_8 _22211_ (.A(_05653_),
    .X(_05654_));
 sg13g2_buf_2 _22212_ (.A(_05654_),
    .X(_05655_));
 sg13g2_a22oi_1 _22213_ (.Y(_05656_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][10] ),
    .A2(net77),
    .A1(\top_ihp.oisc.regs[55][10] ));
 sg13g2_nand4_1 _22214_ (.B(_05647_),
    .C(_05650_),
    .A(_05643_),
    .Y(_05657_),
    .D(_05656_));
 sg13g2_buf_8 _22215_ (.A(_05588_),
    .X(_05658_));
 sg13g2_buf_2 _22216_ (.A(net181),
    .X(_05659_));
 sg13g2_a22oi_1 _22217_ (.Y(_05660_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][10] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][10] ));
 sg13g2_buf_2 _22218_ (.A(_05525_),
    .X(_05661_));
 sg13g2_buf_8 _22219_ (.A(_05544_),
    .X(_05662_));
 sg13g2_buf_8 _22220_ (.A(net430),
    .X(_05663_));
 sg13g2_a22oi_1 _22221_ (.Y(_05664_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][10] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[45][10] ));
 sg13g2_buf_8 _22222_ (.A(_05516_),
    .X(_05665_));
 sg13g2_buf_8 _22223_ (.A(net321),
    .X(_05666_));
 sg13g2_a22oi_1 _22224_ (.Y(_05667_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[54][10] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][10] ));
 sg13g2_buf_8 _22225_ (.A(net193),
    .X(_05668_));
 sg13g2_buf_2 _22226_ (.A(_05603_),
    .X(_05669_));
 sg13g2_a22oi_1 _22227_ (.Y(_05670_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][10] ),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][10] ));
 sg13g2_nand4_1 _22228_ (.B(_05664_),
    .C(_05667_),
    .A(_05660_),
    .Y(_05671_),
    .D(_05670_));
 sg13g2_nor4_2 _22229_ (.A(net190),
    .B(_05639_),
    .C(_05657_),
    .Y(_05672_),
    .D(_05671_));
 sg13g2_inv_1 _22230_ (.Y(_05673_),
    .A(\top_ihp.oisc.regs[36][10] ));
 sg13g2_buf_1 _22231_ (.A(net676),
    .X(_05674_));
 sg13g2_nor3_1 _22232_ (.A(_05673_),
    .B(net608),
    .C(_05325_),
    .Y(_05675_));
 sg13g2_buf_8 _22233_ (.A(net676),
    .X(_05676_));
 sg13g2_nand2_1 _22234_ (.Y(_05677_),
    .A(\top_ihp.oisc.regs[31][10] ),
    .B(net607));
 sg13g2_buf_1 _22235_ (.A(net704),
    .X(_05678_));
 sg13g2_nand2_1 _22236_ (.Y(_05679_),
    .A(\top_ihp.oisc.regs[23][10] ),
    .B(net674));
 sg13g2_a21oi_1 _22237_ (.A1(_05677_),
    .A2(_05679_),
    .Y(_05680_),
    .B1(_05434_));
 sg13g2_buf_1 _22238_ (.A(net434),
    .X(_05681_));
 sg13g2_o21ai_1 _22239_ (.B1(net320),
    .Y(_05682_),
    .A1(_05675_),
    .A2(_05680_));
 sg13g2_buf_1 _22240_ (.A(_05395_),
    .X(_05683_));
 sg13g2_nor3_1 _22241_ (.A(net684),
    .B(net683),
    .C(_05509_),
    .Y(_05684_));
 sg13g2_buf_1 _22242_ (.A(_05684_),
    .X(_05685_));
 sg13g2_buf_1 _22243_ (.A(net428),
    .X(_05686_));
 sg13g2_a22oi_1 _22244_ (.Y(_05687_),
    .B1(_05686_),
    .B2(\top_ihp.oisc.regs[17][10] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[8][10] ));
 sg13g2_buf_1 _22245_ (.A(net443),
    .X(_05688_));
 sg13g2_a22oi_1 _22246_ (.Y(_05689_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][10] ),
    .A2(net444),
    .A1(\top_ihp.oisc.regs[21][10] ));
 sg13g2_nor3_1 _22247_ (.A(_05282_),
    .B(_05343_),
    .C(_05409_),
    .Y(_05690_));
 sg13g2_buf_2 _22248_ (.A(_05690_),
    .X(_05691_));
 sg13g2_mux2_1 _22249_ (.A0(\top_ihp.oisc.regs[30][10] ),
    .A1(\top_ihp.oisc.regs[22][10] ),
    .S(net703),
    .X(_05692_));
 sg13g2_and4_1 _22250_ (.A(net615),
    .B(net700),
    .C(net724),
    .D(_05692_),
    .X(_05693_));
 sg13g2_a221oi_1 _22251_ (.B2(\top_ihp.oisc.regs[2][10] ),
    .C1(_05693_),
    .B1(_05691_),
    .A1(\top_ihp.oisc.regs[4][10] ),
    .Y(_05694_),
    .A2(_05506_));
 sg13g2_a22oi_1 _22252_ (.Y(_05695_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[6][10] ),
    .A2(_05381_),
    .A1(\top_ihp.oisc.regs[5][10] ));
 sg13g2_buf_2 _22253_ (.A(net681),
    .X(_05696_));
 sg13g2_mux2_1 _22254_ (.A0(\top_ihp.oisc.regs[7][10] ),
    .A1(\top_ihp.oisc.regs[3][10] ),
    .S(_05564_),
    .X(_05697_));
 sg13g2_nand2_1 _22255_ (.Y(_05698_),
    .A(_05365_),
    .B(_05405_));
 sg13g2_buf_2 _22256_ (.A(_05698_),
    .X(_05699_));
 sg13g2_nor2_2 _22257_ (.A(net614),
    .B(_05699_),
    .Y(_05700_));
 sg13g2_nand3_1 _22258_ (.B(_05697_),
    .C(_05700_),
    .A(net606),
    .Y(_05701_));
 sg13g2_nand2_1 _22259_ (.Y(_05702_),
    .A(\top_ihp.oisc.regs[26][10] ),
    .B(_05493_));
 sg13g2_and4_1 _22260_ (.A(_05694_),
    .B(_05695_),
    .C(_05701_),
    .D(_05702_),
    .X(_05703_));
 sg13g2_nand4_1 _22261_ (.B(_05687_),
    .C(_05689_),
    .A(_05682_),
    .Y(_05704_),
    .D(_05703_));
 sg13g2_buf_1 _22262_ (.A(net439),
    .X(_05705_));
 sg13g2_mux2_1 _22263_ (.A0(\top_ihp.oisc.regs[28][10] ),
    .A1(\top_ihp.oisc.regs[20][10] ),
    .S(net606),
    .X(_05706_));
 sg13g2_nor2_2 _22264_ (.A(net610),
    .B(_05355_),
    .Y(_05707_));
 sg13g2_a22oi_1 _22265_ (.Y(_05708_),
    .B1(_05706_),
    .B2(_05707_),
    .A2(net317),
    .A1(\top_ihp.oisc.regs[1][10] ));
 sg13g2_buf_2 _22266_ (.A(_05436_),
    .X(_05709_));
 sg13g2_buf_2 _22267_ (.A(_05444_),
    .X(_05710_));
 sg13g2_a22oi_1 _22268_ (.Y(_05711_),
    .B1(net605),
    .B2(\top_ihp.oisc.regs[27][10] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[19][10] ));
 sg13g2_buf_2 _22269_ (.A(_05357_),
    .X(_05712_));
 sg13g2_nor3_1 _22270_ (.A(_05341_),
    .B(net703),
    .C(_05448_),
    .Y(_05713_));
 sg13g2_buf_1 _22271_ (.A(_05713_),
    .X(_05714_));
 sg13g2_buf_2 _22272_ (.A(net426),
    .X(_05715_));
 sg13g2_a22oi_1 _22273_ (.Y(_05716_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][10] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][10] ));
 sg13g2_buf_1 _22274_ (.A(net335),
    .X(_05717_));
 sg13g2_nor3_1 _22275_ (.A(_05358_),
    .B(_05400_),
    .C(_05375_),
    .Y(_05718_));
 sg13g2_buf_2 _22276_ (.A(_05718_),
    .X(_05719_));
 sg13g2_buf_1 _22277_ (.A(_05719_),
    .X(_05720_));
 sg13g2_a22oi_1 _22278_ (.Y(_05721_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][10] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][10] ));
 sg13g2_nand4_1 _22279_ (.B(_05711_),
    .C(_05716_),
    .A(_05708_),
    .Y(_05722_),
    .D(_05721_));
 sg13g2_buf_1 _22280_ (.A(net447),
    .X(_05723_));
 sg13g2_nor3_1 _22281_ (.A(net677),
    .B(_05362_),
    .C(net734),
    .Y(_05724_));
 sg13g2_buf_1 _22282_ (.A(_05724_),
    .X(_05725_));
 sg13g2_a22oi_1 _22283_ (.Y(_05726_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][10] ),
    .A2(net314),
    .A1(\top_ihp.oisc.regs[9][10] ));
 sg13g2_buf_1 _22284_ (.A(net448),
    .X(_05727_));
 sg13g2_nor3_2 _22285_ (.A(net680),
    .B(net704),
    .C(_05409_),
    .Y(_05728_));
 sg13g2_buf_8 _22286_ (.A(_05728_),
    .X(_05729_));
 sg13g2_buf_1 _22287_ (.A(net424),
    .X(_05730_));
 sg13g2_a22oi_1 _22288_ (.Y(_05731_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][10] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][10] ));
 sg13g2_buf_1 _22289_ (.A(net336),
    .X(_05732_));
 sg13g2_nor3_2 _22290_ (.A(net685),
    .B(net703),
    .C(_05375_),
    .Y(_05733_));
 sg13g2_buf_1 _22291_ (.A(_05733_),
    .X(_05734_));
 sg13g2_a22oi_1 _22292_ (.Y(_05735_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[14][10] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[13][10] ));
 sg13g2_nor3_2 _22293_ (.A(net434),
    .B(_05308_),
    .C(_05568_),
    .Y(_05736_));
 sg13g2_a22oi_1 _22294_ (.Y(_05737_),
    .B1(_05736_),
    .B2(\top_ihp.oisc.regs[24][10] ),
    .A2(_03716_),
    .A1(net1053));
 sg13g2_nand4_1 _22295_ (.B(_05731_),
    .C(_05735_),
    .A(_05726_),
    .Y(_05738_),
    .D(_05737_));
 sg13g2_buf_8 _22296_ (.A(net192),
    .X(_05739_));
 sg13g2_nor4_1 _22297_ (.A(net709),
    .B(net685),
    .C(_05292_),
    .D(net723),
    .Y(_05740_));
 sg13g2_buf_2 _22298_ (.A(_05740_),
    .X(_05741_));
 sg13g2_buf_1 _22299_ (.A(_05741_),
    .X(_05742_));
 sg13g2_a22oi_1 _22300_ (.Y(_05743_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][10] ),
    .A2(net74),
    .A1(\top_ihp.oisc.regs[37][10] ));
 sg13g2_buf_2 _22301_ (.A(_05551_),
    .X(_05744_));
 sg13g2_buf_8 _22302_ (.A(_05605_),
    .X(_05745_));
 sg13g2_a22oi_1 _22303_ (.Y(_05746_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][10] ),
    .A2(net310),
    .A1(\top_ihp.oisc.regs[48][10] ));
 sg13g2_buf_1 _22304_ (.A(_05553_),
    .X(_05747_));
 sg13g2_buf_8 _22305_ (.A(_05593_),
    .X(_05748_));
 sg13g2_buf_2 _22306_ (.A(net173),
    .X(_05749_));
 sg13g2_a22oi_1 _22307_ (.Y(_05750_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][10] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[39][10] ));
 sg13g2_buf_8 _22308_ (.A(net435),
    .X(_05751_));
 sg13g2_buf_2 _22309_ (.A(_05563_),
    .X(_05752_));
 sg13g2_a22oi_1 _22310_ (.Y(_05753_),
    .B1(net307),
    .B2(\top_ihp.oisc.regs[34][10] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][10] ));
 sg13g2_nand4_1 _22311_ (.B(_05746_),
    .C(_05750_),
    .A(_05743_),
    .Y(_05754_),
    .D(_05753_));
 sg13g2_nor4_1 _22312_ (.A(_05704_),
    .B(_05722_),
    .C(_05738_),
    .D(_05754_),
    .Y(_05755_));
 sg13g2_a21oi_1 _22313_ (.A1(_00251_),
    .A2(net330),
    .Y(_05756_),
    .B1(net34));
 sg13g2_a21oi_1 _22314_ (.A1(_08262_),
    .A2(net718),
    .Y(_05757_),
    .B1(_05756_));
 sg13g2_a21oi_1 _22315_ (.A1(_05672_),
    .A2(_05755_),
    .Y(_00421_),
    .B1(_05757_));
 sg13g2_buf_8 _22316_ (.A(_05563_),
    .X(_05758_));
 sg13g2_buf_1 _22317_ (.A(_05598_),
    .X(_05759_));
 sg13g2_a22oi_1 _22318_ (.Y(_05760_),
    .B1(_05759_),
    .B2(\top_ihp.oisc.regs[51][11] ),
    .A2(net306),
    .A1(\top_ihp.oisc.regs[34][11] ));
 sg13g2_buf_1 _22319_ (.A(_05471_),
    .X(_05761_));
 sg13g2_buf_8 _22320_ (.A(net430),
    .X(_05762_));
 sg13g2_a22oi_1 _22321_ (.Y(_05763_),
    .B1(net304),
    .B2(\top_ihp.oisc.regs[58][11] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][11] ));
 sg13g2_nor3_1 _22322_ (.A(net678),
    .B(net723),
    .C(_05476_),
    .Y(_05764_));
 sg13g2_buf_2 _22323_ (.A(_05764_),
    .X(_05765_));
 sg13g2_a22oi_1 _22324_ (.Y(_05766_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[49][11] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][11] ));
 sg13g2_buf_1 _22325_ (.A(net338),
    .X(_05767_));
 sg13g2_buf_2 _22326_ (.A(_05595_),
    .X(_05768_));
 sg13g2_a22oi_1 _22327_ (.Y(_05769_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[36][11] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][11] ));
 sg13g2_nand4_1 _22328_ (.B(_05763_),
    .C(_05766_),
    .A(_05760_),
    .Y(_05770_),
    .D(_05769_));
 sg13g2_buf_8 _22329_ (.A(_05603_),
    .X(_05771_));
 sg13g2_buf_2 _22330_ (.A(net431),
    .X(_05772_));
 sg13g2_a22oi_1 _22331_ (.Y(_05773_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][11] ),
    .A2(net169),
    .A1(\top_ihp.oisc.regs[46][11] ));
 sg13g2_buf_8 _22332_ (.A(net446),
    .X(_05774_));
 sg13g2_a22oi_1 _22333_ (.Y(_05775_),
    .B1(net302),
    .B2(\top_ihp.oisc.regs[32][11] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][11] ));
 sg13g2_buf_2 _22334_ (.A(net609),
    .X(_05776_));
 sg13g2_a22oi_1 _22335_ (.Y(_05777_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][11] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[42][11] ));
 sg13g2_buf_8 _22336_ (.A(_05665_),
    .X(_05778_));
 sg13g2_buf_8 _22337_ (.A(_05605_),
    .X(_05779_));
 sg13g2_a22oi_1 _22338_ (.Y(_05780_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][11] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][11] ));
 sg13g2_nand4_1 _22339_ (.B(_05775_),
    .C(_05777_),
    .A(_05773_),
    .Y(_05781_),
    .D(_05780_));
 sg13g2_buf_1 _22340_ (.A(net433),
    .X(_05782_));
 sg13g2_a22oi_1 _22341_ (.Y(_05783_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][11] ),
    .A2(_05782_),
    .A1(\top_ihp.oisc.regs[35][11] ));
 sg13g2_buf_8 _22342_ (.A(net329),
    .X(_05784_));
 sg13g2_a22oi_1 _22343_ (.Y(_05785_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[63][11] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][11] ));
 sg13g2_buf_1 _22344_ (.A(net173),
    .X(_05786_));
 sg13g2_a22oi_1 _22345_ (.Y(_05787_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][11] ),
    .A2(net72),
    .A1(\top_ihp.oisc.regs[53][11] ));
 sg13g2_buf_8 _22346_ (.A(net440),
    .X(_05788_));
 sg13g2_buf_1 _22347_ (.A(net328),
    .X(_05789_));
 sg13g2_a22oi_1 _22348_ (.Y(_05790_),
    .B1(_05789_),
    .B2(\top_ihp.oisc.regs[33][11] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][11] ));
 sg13g2_nand4_1 _22349_ (.B(_05785_),
    .C(_05787_),
    .A(_05783_),
    .Y(_05791_),
    .D(_05790_));
 sg13g2_nor4_1 _22350_ (.A(net190),
    .B(_05770_),
    .C(_05781_),
    .D(_05791_),
    .Y(_05792_));
 sg13g2_a22oi_1 _22351_ (.Y(_05793_),
    .B1(net78),
    .B2(\top_ihp.oisc.regs[59][11] ),
    .A2(net193),
    .A1(\top_ihp.oisc.regs[62][11] ));
 sg13g2_a22oi_1 _22352_ (.Y(_05794_),
    .B1(net174),
    .B2(\top_ihp.oisc.regs[39][11] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][11] ));
 sg13g2_buf_8 _22353_ (.A(_05525_),
    .X(_05795_));
 sg13g2_buf_2 _22354_ (.A(_05551_),
    .X(_05796_));
 sg13g2_a22oi_1 _22355_ (.Y(_05797_),
    .B1(net298),
    .B2(\top_ihp.oisc.regs[48][11] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][11] ));
 sg13g2_nor2_1 _22356_ (.A(_05272_),
    .B(_05344_),
    .Y(_05798_));
 sg13g2_buf_1 _22357_ (.A(_05798_),
    .X(_05799_));
 sg13g2_a22oi_1 _22358_ (.Y(_05800_),
    .B1(_05442_),
    .B2(\top_ihp.oisc.regs[24][11] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[20][11] ));
 sg13g2_inv_1 _22359_ (.Y(_05801_),
    .A(_05800_));
 sg13g2_buf_1 _22360_ (.A(_05570_),
    .X(_05802_));
 sg13g2_a22oi_1 _22361_ (.Y(_05803_),
    .B1(_05801_),
    .B2(net673),
    .A2(_05520_),
    .A1(\top_ihp.oisc.regs[40][11] ));
 sg13g2_nand4_1 _22362_ (.B(_05794_),
    .C(_05797_),
    .A(_05793_),
    .Y(_05804_),
    .D(_05803_));
 sg13g2_mux2_1 _22363_ (.A0(\top_ihp.oisc.regs[29][11] ),
    .A1(\top_ihp.oisc.regs[21][11] ),
    .S(net606),
    .X(_05805_));
 sg13g2_buf_1 _22364_ (.A(net677),
    .X(_05806_));
 sg13g2_nor2_2 _22365_ (.A(_05806_),
    .B(net734),
    .Y(_05807_));
 sg13g2_a22oi_1 _22366_ (.Y(_05808_),
    .B1(_05805_),
    .B2(_05807_),
    .A2(net317),
    .A1(\top_ihp.oisc.regs[1][11] ));
 sg13g2_buf_1 _22367_ (.A(_05381_),
    .X(_05809_));
 sg13g2_buf_1 _22368_ (.A(_05442_),
    .X(_05810_));
 sg13g2_a22oi_1 _22369_ (.Y(_05811_),
    .B1(_05284_),
    .B2(\top_ihp.oisc.micro_op[12] ),
    .A2(_05295_),
    .A1(_09796_));
 sg13g2_and4_1 _22370_ (.A(_05811_),
    .B(net841),
    .C(net743),
    .D(_05366_),
    .X(_05812_));
 sg13g2_buf_2 _22371_ (.A(_05812_),
    .X(_05813_));
 sg13g2_and2_1 _22372_ (.A(net699),
    .B(_05813_),
    .X(_05814_));
 sg13g2_a22oi_1 _22373_ (.Y(_05815_),
    .B1(_05814_),
    .B2(\top_ihp.oisc.regs[8][11] ),
    .A2(net297),
    .A1(\top_ihp.oisc.regs[5][11] ));
 sg13g2_nor2_1 _22374_ (.A(_05317_),
    .B(_05419_),
    .Y(_05816_));
 sg13g2_buf_2 _22375_ (.A(_05816_),
    .X(_05817_));
 sg13g2_buf_1 _22376_ (.A(_05817_),
    .X(_05818_));
 sg13g2_a22oi_1 _22377_ (.Y(_05819_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][11] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[10][11] ));
 sg13g2_buf_2 _22378_ (.A(_05444_),
    .X(_05820_));
 sg13g2_buf_1 _22379_ (.A(net442),
    .X(_05821_));
 sg13g2_a22oi_1 _22380_ (.Y(_05822_),
    .B1(net296),
    .B2(\top_ihp.oisc.regs[28][11] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][11] ));
 sg13g2_nand4_1 _22381_ (.B(_05815_),
    .C(_05819_),
    .A(_05808_),
    .Y(_05823_),
    .D(_05822_));
 sg13g2_nor2_1 _22382_ (.A(_05276_),
    .B(_05699_),
    .Y(_05824_));
 sg13g2_buf_2 _22383_ (.A(_05824_),
    .X(_05825_));
 sg13g2_nand3_1 _22384_ (.B(_05799_),
    .C(_05825_),
    .A(\top_ihp.oisc.regs[6][11] ),
    .Y(_05826_));
 sg13g2_nand2_1 _22385_ (.Y(_05827_),
    .A(\top_ihp.oisc.regs[26][11] ),
    .B(net333));
 sg13g2_buf_8 _22386_ (.A(_05691_),
    .X(_05828_));
 sg13g2_buf_1 _22387_ (.A(net295),
    .X(_05829_));
 sg13g2_a22oi_1 _22388_ (.Y(_05830_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][11] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[9][11] ));
 sg13g2_buf_8 _22389_ (.A(_05543_),
    .X(_05831_));
 sg13g2_buf_1 _22390_ (.A(net674),
    .X(_05832_));
 sg13g2_a22oi_1 _22391_ (.Y(_05833_),
    .B1(_05556_),
    .B2(\top_ihp.oisc.regs[11][11] ),
    .A2(_05462_),
    .A1(\top_ihp.oisc.regs[14][11] ));
 sg13g2_nor3_1 _22392_ (.A(net602),
    .B(_05699_),
    .C(_05833_),
    .Y(_05834_));
 sg13g2_a21oi_1 _22393_ (.A1(\top_ihp.oisc.regs[61][11] ),
    .A2(net162),
    .Y(_05835_),
    .B1(_05834_));
 sg13g2_nand4_1 _22394_ (.B(_05827_),
    .C(_05830_),
    .A(_05826_),
    .Y(_05836_),
    .D(_05835_));
 sg13g2_a22oi_1 _22395_ (.Y(_05837_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][11] ),
    .A2(_05357_),
    .A1(\top_ihp.oisc.regs[16][11] ));
 sg13g2_nor3_1 _22396_ (.A(_05272_),
    .B(_05343_),
    .C(_05419_),
    .Y(_05838_));
 sg13g2_buf_2 _22397_ (.A(_05838_),
    .X(_05839_));
 sg13g2_a22oi_1 _22398_ (.Y(_05840_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][11] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[31][11] ));
 sg13g2_a22oi_1 _22399_ (.Y(_05841_),
    .B1(net332),
    .B2(\top_ihp.oisc.regs[3][11] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[18][11] ));
 sg13g2_a22oi_1 _22400_ (.Y(_05842_),
    .B1(net445),
    .B2(\top_ihp.oisc.regs[19][11] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[7][11] ));
 sg13g2_and4_1 _22401_ (.A(_05837_),
    .B(_05840_),
    .C(_05841_),
    .D(_05842_),
    .X(_05843_));
 sg13g2_nor2_1 _22402_ (.A(_05279_),
    .B(net703),
    .Y(_05844_));
 sg13g2_buf_1 _22403_ (.A(_05844_),
    .X(_05845_));
 sg13g2_mux2_1 _22404_ (.A0(\top_ihp.oisc.regs[12][11] ),
    .A1(\top_ihp.oisc.regs[4][11] ),
    .S(net674),
    .X(_05846_));
 sg13g2_buf_8 _22405_ (.A(net614),
    .X(_05847_));
 sg13g2_a22oi_1 _22406_ (.Y(_05848_),
    .B1(_05846_),
    .B2(net420),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[13][11] ));
 sg13g2_nor2_1 _22407_ (.A(_05373_),
    .B(_05368_),
    .Y(_05849_));
 sg13g2_buf_2 _22408_ (.A(_05849_),
    .X(_05850_));
 sg13g2_buf_2 _22409_ (.A(_05850_),
    .X(_05851_));
 sg13g2_nand2b_1 _22410_ (.Y(_05852_),
    .B(net600),
    .A_N(_05848_));
 sg13g2_a22oi_1 _22411_ (.Y(_05853_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][11] ),
    .A2(net316),
    .A1(\top_ihp.oisc.regs[25][11] ));
 sg13g2_a22oi_1 _22412_ (.Y(_05854_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][11] ),
    .A2(_03716_),
    .A1(_08260_));
 sg13g2_nand4_1 _22413_ (.B(_05852_),
    .C(_05853_),
    .A(_05843_),
    .Y(_05855_),
    .D(_05854_));
 sg13g2_nor4_1 _22414_ (.A(_05804_),
    .B(_05823_),
    .C(_05836_),
    .D(_05855_),
    .Y(_05856_));
 sg13g2_a21oi_1 _22415_ (.A1(_00252_),
    .A2(net330),
    .Y(_05857_),
    .B1(net34));
 sg13g2_a21oi_1 _22416_ (.A1(_08260_),
    .A2(_03733_),
    .Y(_05858_),
    .B1(_05857_));
 sg13g2_a21oi_1 _22417_ (.A1(_05792_),
    .A2(_05856_),
    .Y(_00422_),
    .B1(_05858_));
 sg13g2_buf_8 _22418_ (.A(net436),
    .X(_05859_));
 sg13g2_a22oi_1 _22419_ (.Y(_05860_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[14][12] ),
    .A2(net294),
    .A1(\top_ihp.oisc.regs[4][12] ));
 sg13g2_buf_2 _22420_ (.A(net449),
    .X(_05861_));
 sg13g2_a22oi_1 _22421_ (.Y(_05862_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][12] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][12] ));
 sg13g2_nor2_2 _22422_ (.A(_05335_),
    .B(net734),
    .Y(_05863_));
 sg13g2_a22oi_1 _22423_ (.Y(_05864_),
    .B1(_05863_),
    .B2(\top_ihp.oisc.regs[21][12] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[17][12] ));
 sg13g2_a22oi_1 _22424_ (.Y(_05865_),
    .B1(net317),
    .B2(\top_ihp.oisc.regs[1][12] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[9][12] ));
 sg13g2_nand4_1 _22425_ (.B(_05862_),
    .C(_05864_),
    .A(_05860_),
    .Y(_05866_),
    .D(_05865_));
 sg13g2_a22oi_1 _22426_ (.Y(_05867_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[13][12] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][12] ));
 sg13g2_a22oi_1 _22427_ (.Y(_05868_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][12] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[19][12] ));
 sg13g2_a22oi_1 _22428_ (.Y(_05869_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[45][12] ),
    .A2(_05751_),
    .A1(\top_ihp.oisc.regs[40][12] ));
 sg13g2_nand3_1 _22429_ (.B(_05868_),
    .C(_05869_),
    .A(_05867_),
    .Y(_05870_));
 sg13g2_buf_1 _22430_ (.A(_05440_),
    .X(_05871_));
 sg13g2_a22oi_1 _22431_ (.Y(_05872_),
    .B1(_05825_),
    .B2(\top_ihp.oisc.regs[10][12] ),
    .A2(net698),
    .A1(\top_ihp.oisc.regs[27][12] ));
 sg13g2_nand2_1 _22432_ (.Y(_05873_),
    .A(_08252_),
    .B(net748));
 sg13g2_o21ai_1 _22433_ (.B1(_05873_),
    .Y(_05874_),
    .A1(net679),
    .A2(_05872_));
 sg13g2_a221oi_1 _22434_ (.B2(\top_ihp.oisc.regs[50][12] ),
    .C1(_05874_),
    .B1(_05627_),
    .A1(\top_ihp.oisc.regs[8][12] ),
    .Y(_05875_),
    .A2(net429));
 sg13g2_buf_8 _22435_ (.A(net450),
    .X(_05876_));
 sg13g2_nand2_1 _22436_ (.Y(_05877_),
    .A(\top_ihp.oisc.regs[28][12] ),
    .B(_05455_));
 sg13g2_buf_1 _22437_ (.A(net615),
    .X(_05878_));
 sg13g2_nor2_1 _22438_ (.A(net675),
    .B(net701),
    .Y(_05879_));
 sg13g2_nand4_1 _22439_ (.B(net419),
    .C(net742),
    .A(\top_ihp.oisc.regs[31][12] ),
    .Y(_05880_),
    .D(_05879_));
 sg13g2_nand2_1 _22440_ (.Y(_05881_),
    .A(_05877_),
    .B(_05880_));
 sg13g2_a221oi_1 _22441_ (.B2(\top_ihp.oisc.regs[25][12] ),
    .C1(_05881_),
    .B1(_05510_),
    .A1(\top_ihp.oisc.regs[6][12] ),
    .Y(_05882_),
    .A2(net292));
 sg13g2_a22oi_1 _22442_ (.Y(_05883_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][12] ),
    .A2(_05658_),
    .A1(\top_ihp.oisc.regs[47][12] ));
 sg13g2_nor3_2 _22443_ (.A(net608),
    .B(net612),
    .C(_05699_),
    .Y(_05884_));
 sg13g2_a22oi_1 _22444_ (.Y(_05885_),
    .B1(_05884_),
    .B2(\top_ihp.oisc.regs[7][12] ),
    .A2(_05651_),
    .A1(\top_ihp.oisc.regs[55][12] ));
 sg13g2_nand4_1 _22445_ (.B(_05882_),
    .C(_05883_),
    .A(_05875_),
    .Y(_05886_),
    .D(_05885_));
 sg13g2_buf_1 _22446_ (.A(net610),
    .X(_05887_));
 sg13g2_mux2_1 _22447_ (.A0(\top_ihp.oisc.regs[22][12] ),
    .A1(\top_ihp.oisc.regs[18][12] ),
    .S(net418),
    .X(_05888_));
 sg13g2_buf_1 _22448_ (.A(_05572_),
    .X(_05889_));
 sg13g2_buf_8 _22449_ (.A(net599),
    .X(_05890_));
 sg13g2_a22oi_1 _22450_ (.Y(_05891_),
    .B1(_05888_),
    .B2(net417),
    .A2(net699),
    .A1(\top_ihp.oisc.regs[26][12] ));
 sg13g2_buf_1 _22451_ (.A(net434),
    .X(_05892_));
 sg13g2_nor3_1 _22452_ (.A(_05811_),
    .B(_05347_),
    .C(net840),
    .Y(_05893_));
 sg13g2_a21o_1 _22453_ (.A2(_05893_),
    .A1(net743),
    .B1(net948),
    .X(_05894_));
 sg13g2_buf_2 _22454_ (.A(_05894_),
    .X(_05895_));
 sg13g2_nand3_1 _22455_ (.B(_05892_),
    .C(_05895_),
    .A(\top_ihp.oisc.regs[5][12] ),
    .Y(_05896_));
 sg13g2_nand3_1 _22456_ (.B(net418),
    .C(_05700_),
    .A(\top_ihp.oisc.regs[3][12] ),
    .Y(_05897_));
 sg13g2_nand2_1 _22457_ (.Y(_05898_),
    .A(_05896_),
    .B(_05897_));
 sg13g2_nor2_1 _22458_ (.A(net684),
    .B(net706),
    .Y(_05899_));
 sg13g2_buf_1 _22459_ (.A(_05899_),
    .X(_05900_));
 sg13g2_buf_2 _22460_ (.A(_05900_),
    .X(_05901_));
 sg13g2_nand3_1 _22461_ (.B(net420),
    .C(net290),
    .A(\top_ihp.oisc.regs[2][12] ),
    .Y(_05902_));
 sg13g2_nand3_1 _22462_ (.B(net608),
    .C(_05535_),
    .A(\top_ihp.oisc.regs[15][12] ),
    .Y(_05903_));
 sg13g2_nand2_1 _22463_ (.Y(_05904_),
    .A(_05902_),
    .B(_05903_));
 sg13g2_a22oi_1 _22464_ (.Y(_05905_),
    .B1(_05904_),
    .B2(_05407_),
    .A2(_05898_),
    .A1(net417));
 sg13g2_o21ai_1 _22465_ (.B1(_05905_),
    .Y(_05906_),
    .A1(_05419_),
    .A2(_05891_));
 sg13g2_nor4_1 _22466_ (.A(_05866_),
    .B(_05870_),
    .C(_05886_),
    .D(_05906_),
    .Y(_05907_));
 sg13g2_a22oi_1 _22467_ (.Y(_05908_),
    .B1(net186),
    .B2(\top_ihp.oisc.regs[33][12] ),
    .A2(_05472_),
    .A1(\top_ihp.oisc.regs[37][12] ));
 sg13g2_buf_1 _22468_ (.A(_05595_),
    .X(_05909_));
 sg13g2_a22oi_1 _22469_ (.Y(_05910_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][12] ),
    .A2(net306),
    .A1(\top_ihp.oisc.regs[34][12] ));
 sg13g2_a22oi_1 _22470_ (.Y(_05911_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[35][12] ),
    .A2(_05310_),
    .A1(\top_ihp.oisc.regs[60][12] ));
 sg13g2_a22oi_1 _22471_ (.Y(_05912_),
    .B1(net334),
    .B2(\top_ihp.oisc.regs[42][12] ),
    .A2(_05460_),
    .A1(\top_ihp.oisc.regs[49][12] ));
 sg13g2_nand4_1 _22472_ (.B(_05910_),
    .C(_05911_),
    .A(_05908_),
    .Y(_05913_),
    .D(_05912_));
 sg13g2_buf_1 _22473_ (.A(net614),
    .X(_05914_));
 sg13g2_a21oi_2 _22474_ (.B1(_03728_),
    .Y(_05915_),
    .A2(net743),
    .A1(_05286_));
 sg13g2_nor2_1 _22475_ (.A(net700),
    .B(_05915_),
    .Y(_05916_));
 sg13g2_nand4_1 _22476_ (.B(_05469_),
    .C(_05916_),
    .A(net416),
    .Y(_05917_),
    .D(_05900_));
 sg13g2_buf_2 _22477_ (.A(_05917_),
    .X(_05918_));
 sg13g2_a22oi_1 _22478_ (.Y(_05919_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][12] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][12] ));
 sg13g2_a22oi_1 _22479_ (.Y(_05920_),
    .B1(net72),
    .B2(\top_ihp.oisc.regs[53][12] ),
    .A2(net78),
    .A1(\top_ihp.oisc.regs[59][12] ));
 sg13g2_nand3_1 _22480_ (.B(_05919_),
    .C(_05920_),
    .A(_05918_),
    .Y(_05921_));
 sg13g2_buf_1 _22481_ (.A(net324),
    .X(_05922_));
 sg13g2_a22oi_1 _22482_ (.Y(_05923_),
    .B1(net174),
    .B2(\top_ihp.oisc.regs[39][12] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[63][12] ));
 sg13g2_nand2_1 _22483_ (.Y(_05924_),
    .A(\top_ihp.oisc.regs[58][12] ),
    .B(net304));
 sg13g2_a22oi_1 _22484_ (.Y(_05925_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][12] ),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][12] ));
 sg13g2_buf_2 _22485_ (.A(_05741_),
    .X(_05926_));
 sg13g2_a22oi_1 _22486_ (.Y(_05927_),
    .B1(_05926_),
    .B2(\top_ihp.oisc.regs[52][12] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][12] ));
 sg13g2_nand4_1 _22487_ (.B(_05924_),
    .C(_05925_),
    .A(_05923_),
    .Y(_05928_),
    .D(_05927_));
 sg13g2_a22oi_1 _22488_ (.Y(_05929_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][12] ),
    .A2(_05669_),
    .A1(\top_ihp.oisc.regs[46][12] ));
 sg13g2_a22oi_1 _22489_ (.Y(_05930_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[54][12] ),
    .A2(_05788_),
    .A1(\top_ihp.oisc.regs[43][12] ));
 sg13g2_buf_1 _22490_ (.A(_05676_),
    .X(_05931_));
 sg13g2_buf_2 _22491_ (.A(net722),
    .X(_05932_));
 sg13g2_nand3_1 _22492_ (.B(net419),
    .C(net697),
    .A(\top_ihp.oisc.regs[29][12] ),
    .Y(_05933_));
 sg13g2_buf_1 _22493_ (.A(_05570_),
    .X(_05934_));
 sg13g2_nand3_1 _22494_ (.B(net604),
    .C(net672),
    .A(\top_ihp.oisc.regs[24][12] ),
    .Y(_05935_));
 sg13g2_nand3_1 _22495_ (.B(_05933_),
    .C(_05935_),
    .A(net415),
    .Y(_05936_));
 sg13g2_nand3_1 _22496_ (.B(net419),
    .C(_05871_),
    .A(\top_ihp.oisc.regs[23][12] ),
    .Y(_05937_));
 sg13g2_buf_1 _22497_ (.A(net677),
    .X(_05938_));
 sg13g2_nand3_1 _22498_ (.B(net598),
    .C(net673),
    .A(\top_ihp.oisc.regs[16][12] ),
    .Y(_05939_));
 sg13g2_nand3_1 _22499_ (.B(_05937_),
    .C(_05939_),
    .A(net602),
    .Y(_05940_));
 sg13g2_a22oi_1 _22500_ (.Y(_05941_),
    .B1(_05936_),
    .B2(_05940_),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][12] ));
 sg13g2_a22oi_1 _22501_ (.Y(_05942_),
    .B1(net302),
    .B2(\top_ihp.oisc.regs[32][12] ),
    .A2(_05338_),
    .A1(\top_ihp.oisc.regs[38][12] ));
 sg13g2_nand4_1 _22502_ (.B(_05930_),
    .C(_05941_),
    .A(_05929_),
    .Y(_05943_),
    .D(_05942_));
 sg13g2_nor4_1 _22503_ (.A(_05913_),
    .B(_05921_),
    .C(_05928_),
    .D(_05943_),
    .Y(_05944_));
 sg13g2_buf_1 _22504_ (.A(net331),
    .X(_05945_));
 sg13g2_buf_1 _22505_ (.A(_05622_),
    .X(_05946_));
 sg13g2_a21o_1 _22506_ (.A2(net159),
    .A1(_00253_),
    .B1(net33),
    .X(_05947_));
 sg13g2_a22oi_1 _22507_ (.Y(_00423_),
    .B1(_05947_),
    .B2(_05873_),
    .A2(_05944_),
    .A1(_05907_));
 sg13g2_buf_1 _22508_ (.A(net331),
    .X(_05948_));
 sg13g2_a22oi_1 _22509_ (.Y(_05949_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][13] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[33][13] ));
 sg13g2_nor2_1 _22510_ (.A(net676),
    .B(_05355_),
    .Y(_05950_));
 sg13g2_nand2_1 _22511_ (.Y(_05951_),
    .A(\top_ihp.oisc.regs[16][13] ),
    .B(_05950_));
 sg13g2_nand4_1 _22512_ (.B(_05878_),
    .C(net724),
    .A(\top_ihp.oisc.regs[30][13] ),
    .Y(_05952_),
    .D(_05879_));
 sg13g2_o21ai_1 _22513_ (.B1(_05952_),
    .Y(_05953_),
    .A1(net320),
    .A2(_05951_));
 sg13g2_a21oi_1 _22514_ (.A1(\top_ihp.oisc.regs[37][13] ),
    .A2(_05761_),
    .Y(_05954_),
    .B1(_05953_));
 sg13g2_nor3_2 _22515_ (.A(net678),
    .B(_05531_),
    .C(net679),
    .Y(_05955_));
 sg13g2_buf_1 _22516_ (.A(net613),
    .X(_05956_));
 sg13g2_nor3_2 _22517_ (.A(net414),
    .B(_05610_),
    .C(_05508_),
    .Y(_05957_));
 sg13g2_a22oi_1 _22518_ (.Y(_05958_),
    .B1(_05957_),
    .B2(\top_ihp.oisc.regs[8][13] ),
    .A2(_05955_),
    .A1(\top_ihp.oisc.regs[56][13] ));
 sg13g2_nor3_1 _22519_ (.A(net599),
    .B(_05469_),
    .C(_05699_),
    .Y(_05959_));
 sg13g2_nand2_1 _22520_ (.Y(_05960_),
    .A(\top_ihp.oisc.regs[15][13] ),
    .B(_05959_));
 sg13g2_nand4_1 _22521_ (.B(_05954_),
    .C(_05958_),
    .A(_05949_),
    .Y(_05961_),
    .D(_05960_));
 sg13g2_a22oi_1 _22522_ (.Y(_05962_),
    .B1(_05742_),
    .B2(\top_ihp.oisc.regs[52][13] ),
    .A2(net181),
    .A1(\top_ihp.oisc.regs[47][13] ));
 sg13g2_a22oi_1 _22523_ (.Y(_05963_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][13] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][13] ));
 sg13g2_a22oi_1 _22524_ (.Y(_05964_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][13] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][13] ));
 sg13g2_a22oi_1 _22525_ (.Y(_05965_),
    .B1(net310),
    .B2(\top_ihp.oisc.regs[48][13] ),
    .A2(net193),
    .A1(\top_ihp.oisc.regs[62][13] ));
 sg13g2_nand4_1 _22526_ (.B(_05963_),
    .C(_05964_),
    .A(_05962_),
    .Y(_05966_),
    .D(_05965_));
 sg13g2_a22oi_1 _22527_ (.Y(_05967_),
    .B1(_05663_),
    .B2(\top_ihp.oisc.regs[58][13] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][13] ));
 sg13g2_buf_1 _22528_ (.A(net435),
    .X(_05968_));
 sg13g2_a22oi_1 _22529_ (.Y(_05969_),
    .B1(net288),
    .B2(\top_ihp.oisc.regs[40][13] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][13] ));
 sg13g2_buf_1 _22530_ (.A(_05337_),
    .X(_05970_));
 sg13g2_a22oi_1 _22531_ (.Y(_05971_),
    .B1(_05666_),
    .B2(\top_ihp.oisc.regs[54][13] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][13] ));
 sg13g2_a22oi_1 _22532_ (.Y(_05972_),
    .B1(_05747_),
    .B2(\top_ihp.oisc.regs[39][13] ),
    .A2(_05922_),
    .A1(\top_ihp.oisc.regs[63][13] ));
 sg13g2_nand4_1 _22533_ (.B(_05969_),
    .C(_05971_),
    .A(_05967_),
    .Y(_05973_),
    .D(_05972_));
 sg13g2_nor4_1 _22534_ (.A(net158),
    .B(_05961_),
    .C(_05966_),
    .D(_05973_),
    .Y(_05974_));
 sg13g2_buf_8 _22535_ (.A(_05479_),
    .X(_05975_));
 sg13g2_a22oi_1 _22536_ (.Y(_05976_),
    .B1(_05772_),
    .B2(\top_ihp.oisc.regs[41][13] ),
    .A2(_05975_),
    .A1(\top_ihp.oisc.regs[43][13] ));
 sg13g2_a22oi_1 _22537_ (.Y(_05977_),
    .B1(_05774_),
    .B2(\top_ihp.oisc.regs[32][13] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][13] ));
 sg13g2_buf_2 _22538_ (.A(_05595_),
    .X(_05978_));
 sg13g2_a22oi_1 _22539_ (.Y(_05979_),
    .B1(_05978_),
    .B2(\top_ihp.oisc.regs[36][13] ),
    .A2(net73),
    .A1(\top_ihp.oisc.regs[53][13] ));
 sg13g2_buf_8 _22540_ (.A(net185),
    .X(_05980_));
 sg13g2_a22oi_1 _22541_ (.Y(_05981_),
    .B1(_05980_),
    .B2(\top_ihp.oisc.regs[59][13] ),
    .A2(_05486_),
    .A1(\top_ihp.oisc.regs[42][13] ));
 sg13g2_nand4_1 _22542_ (.B(_05977_),
    .C(_05979_),
    .A(_05976_),
    .Y(_05982_),
    .D(_05981_));
 sg13g2_a22oi_1 _22543_ (.Y(_05983_),
    .B1(_05736_),
    .B2(\top_ihp.oisc.regs[24][13] ),
    .A2(net424),
    .A1(\top_ihp.oisc.regs[10][13] ));
 sg13g2_a22oi_1 _22544_ (.Y(_05984_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[25][13] ),
    .A2(_05450_),
    .A1(\top_ihp.oisc.regs[21][13] ));
 sg13g2_a22oi_1 _22545_ (.Y(_05985_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][13] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[7][13] ));
 sg13g2_a22oi_1 _22546_ (.Y(_05986_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[28][13] ),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][13] ));
 sg13g2_nand4_1 _22547_ (.B(_05984_),
    .C(_05985_),
    .A(_05983_),
    .Y(_05987_),
    .D(_05986_));
 sg13g2_nor2_1 _22548_ (.A(_05529_),
    .B(net700),
    .Y(_05988_));
 sg13g2_and4_1 _22549_ (.A(\top_ihp.oisc.regs[57][13] ),
    .B(net613),
    .C(_05442_),
    .D(_05988_),
    .X(_05989_));
 sg13g2_a21oi_1 _22550_ (.A1(\top_ihp.oisc.regs[18][13] ),
    .A2(net335),
    .Y(_05990_),
    .B1(_05989_));
 sg13g2_a22oi_1 _22551_ (.Y(_05991_),
    .B1(net611),
    .B2(\top_ihp.oisc.regs[31][13] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[6][13] ));
 sg13g2_a22oi_1 _22552_ (.Y(_05992_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][13] ),
    .A2(_05436_),
    .A1(\top_ihp.oisc.regs[19][13] ));
 sg13g2_nand3_1 _22553_ (.B(net614),
    .C(_05850_),
    .A(\top_ihp.oisc.regs[12][13] ),
    .Y(_05993_));
 sg13g2_nor2_1 _22554_ (.A(_05267_),
    .B(_05699_),
    .Y(_05994_));
 sg13g2_buf_1 _22555_ (.A(_05994_),
    .X(_05995_));
 sg13g2_nand3_1 _22556_ (.B(net613),
    .C(_05995_),
    .A(\top_ihp.oisc.regs[11][13] ),
    .Y(_05996_));
 sg13g2_nand2_1 _22557_ (.Y(_05997_),
    .A(_05993_),
    .B(_05996_));
 sg13g2_buf_1 _22558_ (.A(net607),
    .X(_05998_));
 sg13g2_a22oi_1 _22559_ (.Y(_05999_),
    .B1(_05997_),
    .B2(net413),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[4][13] ));
 sg13g2_nand4_1 _22560_ (.B(_05991_),
    .C(_05992_),
    .A(_05990_),
    .Y(_06000_),
    .D(_05999_));
 sg13g2_a22oi_1 _22561_ (.Y(_06001_),
    .B1(net295),
    .B2(\top_ihp.oisc.regs[2][13] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[26][13] ));
 sg13g2_nor2_2 _22562_ (.A(net680),
    .B(net683),
    .Y(_06002_));
 sg13g2_buf_1 _22563_ (.A(net700),
    .X(_06003_));
 sg13g2_nor2_1 _22564_ (.A(net615),
    .B(net707),
    .Y(_06004_));
 sg13g2_and3_1 _22565_ (.X(_06005_),
    .A(\top_ihp.oisc.regs[34][13] ),
    .B(net671),
    .C(_06004_));
 sg13g2_a22oi_1 _22566_ (.Y(_06006_),
    .B1(_06002_),
    .B2(_06005_),
    .A2(_05444_),
    .A1(\top_ihp.oisc.regs[27][13] ));
 sg13g2_a22oi_1 _22567_ (.Y(_06007_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][13] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[17][13] ));
 sg13g2_nor3_1 _22568_ (.A(net948),
    .B(_05313_),
    .C(_05298_),
    .Y(_06008_));
 sg13g2_buf_2 _22569_ (.A(_06008_),
    .X(_06009_));
 sg13g2_and2_1 _22570_ (.A(net696),
    .B(_05895_),
    .X(_06010_));
 sg13g2_a22oi_1 _22571_ (.Y(_06011_),
    .B1(_06010_),
    .B2(\top_ihp.oisc.regs[13][13] ),
    .A2(_05488_),
    .A1(\top_ihp.oisc.regs[1][13] ));
 sg13g2_nand4_1 _22572_ (.B(_06006_),
    .C(_06007_),
    .A(_06001_),
    .Y(_06012_),
    .D(_06011_));
 sg13g2_nand2_1 _22573_ (.Y(_06013_),
    .A(\top_ihp.oisc.regs[3][13] ),
    .B(net332));
 sg13g2_nor2_1 _22574_ (.A(net614),
    .B(net671),
    .Y(_06014_));
 sg13g2_nand4_1 _22575_ (.B(_05548_),
    .C(net290),
    .A(\top_ihp.oisc.regs[49][13] ),
    .Y(_06015_),
    .D(_06014_));
 sg13g2_nor2_1 _22576_ (.A(net682),
    .B(net683),
    .Y(_06016_));
 sg13g2_buf_2 _22577_ (.A(_06016_),
    .X(_06017_));
 sg13g2_nand3_1 _22578_ (.B(_06017_),
    .C(_05850_),
    .A(\top_ihp.oisc.regs[5][13] ),
    .Y(_06018_));
 sg13g2_nand2_1 _22579_ (.Y(_06019_),
    .A(_08256_),
    .B(net748));
 sg13g2_nor2_1 _22580_ (.A(net841),
    .B(_05368_),
    .Y(_06020_));
 sg13g2_buf_1 _22581_ (.A(_06020_),
    .X(_06021_));
 sg13g2_nor2_1 _22582_ (.A(net680),
    .B(net704),
    .Y(_06022_));
 sg13g2_nand3_1 _22583_ (.B(net670),
    .C(_06022_),
    .A(\top_ihp.oisc.regs[14][13] ),
    .Y(_06023_));
 sg13g2_and3_1 _22584_ (.X(_06024_),
    .A(_06018_),
    .B(_06019_),
    .C(_06023_));
 sg13g2_a22oi_1 _22585_ (.Y(_06025_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][13] ),
    .A2(net329),
    .A1(\top_ihp.oisc.regs[50][13] ));
 sg13g2_nand4_1 _22586_ (.B(_06015_),
    .C(_06024_),
    .A(_06013_),
    .Y(_06026_),
    .D(_06025_));
 sg13g2_nor4_1 _22587_ (.A(_05987_),
    .B(_06000_),
    .C(_06012_),
    .D(_06026_),
    .Y(_06027_));
 sg13g2_nor2b_1 _22588_ (.A(_05982_),
    .B_N(_06027_),
    .Y(_06028_));
 sg13g2_a21o_1 _22589_ (.A2(net159),
    .A1(_00254_),
    .B1(net33),
    .X(_06029_));
 sg13g2_a22oi_1 _22590_ (.Y(_00424_),
    .B1(_06029_),
    .B2(_06019_),
    .A2(_06028_),
    .A1(_05974_));
 sg13g2_a21oi_1 _22591_ (.A1(_00255_),
    .A2(net330),
    .Y(_06030_),
    .B1(_05623_));
 sg13g2_a21oi_1 _22592_ (.A1(_08285_),
    .A2(net718),
    .Y(_06031_),
    .B1(_06030_));
 sg13g2_and2_1 _22593_ (.A(\top_ihp.oisc.regs[48][14] ),
    .B(net310),
    .X(_06032_));
 sg13g2_a221oi_1 _22594_ (.B2(\top_ihp.oisc.regs[58][14] ),
    .C1(_06032_),
    .B1(_05663_),
    .A1(\top_ihp.oisc.regs[33][14] ),
    .Y(_06033_),
    .A2(net166));
 sg13g2_a22oi_1 _22595_ (.Y(_06034_),
    .B1(net165),
    .B2(\top_ihp.oisc.regs[45][14] ),
    .A2(_05484_),
    .A1(\top_ihp.oisc.regs[42][14] ));
 sg13g2_buf_8 _22596_ (.A(_05553_),
    .X(_06035_));
 sg13g2_a22oi_1 _22597_ (.Y(_06036_),
    .B1(net155),
    .B2(\top_ihp.oisc.regs[39][14] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[44][14] ));
 sg13g2_a22oi_1 _22598_ (.Y(_06037_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][14] ),
    .A2(_05478_),
    .A1(\top_ihp.oisc.regs[43][14] ));
 sg13g2_a22oi_1 _22599_ (.Y(_06038_),
    .B1(net329),
    .B2(\top_ihp.oisc.regs[50][14] ),
    .A2(_05465_),
    .A1(\top_ihp.oisc.regs[62][14] ));
 sg13g2_nand4_1 _22600_ (.B(_06036_),
    .C(_06037_),
    .A(_06034_),
    .Y(_06039_),
    .D(_06038_));
 sg13g2_a22oi_1 _22601_ (.Y(_06040_),
    .B1(_05741_),
    .B2(\top_ihp.oisc.regs[52][14] ),
    .A2(_05593_),
    .A1(\top_ihp.oisc.regs[53][14] ));
 sg13g2_a22oi_1 _22602_ (.Y(_06041_),
    .B1(_05337_),
    .B2(\top_ihp.oisc.regs[38][14] ),
    .A2(_05309_),
    .A1(\top_ihp.oisc.regs[60][14] ));
 sg13g2_a22oi_1 _22603_ (.Y(_06042_),
    .B1(net321),
    .B2(\top_ihp.oisc.regs[54][14] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][14] ));
 sg13g2_a22oi_1 _22604_ (.Y(_06043_),
    .B1(_05605_),
    .B2(\top_ihp.oisc.regs[56][14] ),
    .A2(_05560_),
    .A1(\top_ihp.oisc.regs[35][14] ));
 sg13g2_nand4_1 _22605_ (.B(_06041_),
    .C(_06042_),
    .A(_06040_),
    .Y(_06044_),
    .D(_06043_));
 sg13g2_a22oi_1 _22606_ (.Y(_06045_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[46][14] ),
    .A2(_05758_),
    .A1(\top_ihp.oisc.regs[34][14] ));
 sg13g2_nor4_1 _22607_ (.A(net682),
    .B(net678),
    .C(net700),
    .D(net702),
    .Y(_06046_));
 sg13g2_buf_2 _22608_ (.A(_06046_),
    .X(_06047_));
 sg13g2_a22oi_1 _22609_ (.Y(_06048_),
    .B1(_06047_),
    .B2(\top_ihp.oisc.regs[49][14] ),
    .A2(_05598_),
    .A1(\top_ihp.oisc.regs[51][14] ));
 sg13g2_a22oi_1 _22610_ (.Y(_06049_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[47][14] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][14] ));
 sg13g2_a22oi_1 _22611_ (.Y(_06050_),
    .B1(_05520_),
    .B2(\top_ihp.oisc.regs[40][14] ),
    .A2(_05471_),
    .A1(\top_ihp.oisc.regs[37][14] ));
 sg13g2_nand4_1 _22612_ (.B(_06048_),
    .C(_06049_),
    .A(_06045_),
    .Y(_06051_),
    .D(_06050_));
 sg13g2_nor4_1 _22613_ (.A(_05612_),
    .B(_06039_),
    .C(_06044_),
    .D(_06051_),
    .Y(_06052_));
 sg13g2_buf_1 _22614_ (.A(net610),
    .X(_06053_));
 sg13g2_nand4_1 _22615_ (.B(net412),
    .C(net601),
    .A(\top_ihp.oisc.regs[57][14] ),
    .Y(_06054_),
    .D(_05988_));
 sg13g2_nand3_1 _22616_ (.B(net434),
    .C(net722),
    .A(\top_ihp.oisc.regs[29][14] ),
    .Y(_06055_));
 sg13g2_buf_1 _22617_ (.A(_05582_),
    .X(_06056_));
 sg13g2_nand3_1 _22618_ (.B(net610),
    .C(net721),
    .A(\top_ihp.oisc.regs[26][14] ),
    .Y(_06057_));
 sg13g2_nand2_1 _22619_ (.Y(_06058_),
    .A(_06055_),
    .B(_06057_));
 sg13g2_and2_1 _22620_ (.A(_06009_),
    .B(_05353_),
    .X(_06059_));
 sg13g2_mux2_1 _22621_ (.A0(\top_ihp.oisc.regs[30][14] ),
    .A1(\top_ihp.oisc.regs[28][14] ),
    .S(net841),
    .X(_06060_));
 sg13g2_a22oi_1 _22622_ (.Y(_06061_),
    .B1(_06059_),
    .B2(_06060_),
    .A2(_06058_),
    .A1(net413));
 sg13g2_a22oi_1 _22623_ (.Y(_06062_),
    .B1(net295),
    .B2(\top_ihp.oisc.regs[2][14] ),
    .A2(net438),
    .A1(\top_ihp.oisc.regs[23][14] ));
 sg13g2_a22oi_1 _22624_ (.Y(_06063_),
    .B1(net611),
    .B2(\top_ihp.oisc.regs[31][14] ),
    .A2(net332),
    .A1(\top_ihp.oisc.regs[3][14] ));
 sg13g2_nand4_1 _22625_ (.B(_06061_),
    .C(_06062_),
    .A(_06054_),
    .Y(_06064_),
    .D(_06063_));
 sg13g2_a221oi_1 _22626_ (.B2(\top_ihp.oisc.regs[6][14] ),
    .C1(_06064_),
    .B1(net292),
    .A1(_08285_),
    .Y(_06065_),
    .A2(net728));
 sg13g2_buf_1 _22627_ (.A(_05839_),
    .X(_06066_));
 sg13g2_a22oi_1 _22628_ (.Y(_06067_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][14] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[11][14] ));
 sg13g2_a22oi_1 _22629_ (.Y(_06068_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[4][14] ),
    .A2(_05357_),
    .A1(\top_ihp.oisc.regs[16][14] ));
 sg13g2_a22oi_1 _22630_ (.Y(_06069_),
    .B1(_05729_),
    .B2(\top_ihp.oisc.regs[10][14] ),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][14] ));
 sg13g2_buf_1 _22631_ (.A(_05395_),
    .X(_06070_));
 sg13g2_a22oi_1 _22632_ (.Y(_06071_),
    .B1(_05451_),
    .B2(\top_ihp.oisc.regs[21][14] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[8][14] ));
 sg13g2_nand4_1 _22633_ (.B(_06068_),
    .C(_06069_),
    .A(_06067_),
    .Y(_06072_),
    .D(_06071_));
 sg13g2_nand3_1 _22634_ (.B(net607),
    .C(_05440_),
    .A(\top_ihp.oisc.regs[27][14] ),
    .Y(_06073_));
 sg13g2_nand3_1 _22635_ (.B(net674),
    .C(_06056_),
    .A(\top_ihp.oisc.regs[18][14] ),
    .Y(_06074_));
 sg13g2_a21o_1 _22636_ (.A2(_06074_),
    .A1(_06073_),
    .B1(net291),
    .X(_06075_));
 sg13g2_nand3_1 _22637_ (.B(_05535_),
    .C(_05463_),
    .A(\top_ihp.oisc.regs[63][14] ),
    .Y(_06076_));
 sg13g2_a22oi_1 _22638_ (.Y(_06077_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[17][14] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[7][14] ));
 sg13g2_nand3_1 _22639_ (.B(_06076_),
    .C(_06077_),
    .A(_06075_),
    .Y(_06078_));
 sg13g2_a22oi_1 _22640_ (.Y(_06079_),
    .B1(_05734_),
    .B2(\top_ihp.oisc.regs[14][14] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[13][14] ));
 sg13g2_a22oi_1 _22641_ (.Y(_06080_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[15][14] ),
    .A2(_05436_),
    .A1(\top_ihp.oisc.regs[19][14] ));
 sg13g2_a22oi_1 _22642_ (.Y(_06081_),
    .B1(net448),
    .B2(\top_ihp.oisc.regs[12][14] ),
    .A2(net449),
    .A1(\top_ihp.oisc.regs[20][14] ));
 sg13g2_nor3_1 _22643_ (.A(_05341_),
    .B(net703),
    .C(_05355_),
    .Y(_06082_));
 sg13g2_buf_2 _22644_ (.A(_06082_),
    .X(_06083_));
 sg13g2_a22oi_1 _22645_ (.Y(_06084_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][14] ),
    .A2(_05714_),
    .A1(\top_ihp.oisc.regs[25][14] ));
 sg13g2_nand4_1 _22646_ (.B(_06080_),
    .C(_06081_),
    .A(_06079_),
    .Y(_06085_),
    .D(_06084_));
 sg13g2_a22oi_1 _22647_ (.Y(_06086_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[1][14] ),
    .A2(_05382_),
    .A1(\top_ihp.oisc.regs[5][14] ));
 sg13g2_nand2_1 _22648_ (.Y(_06087_),
    .A(\top_ihp.oisc.regs[36][14] ),
    .B(net161));
 sg13g2_a22oi_1 _22649_ (.Y(_06088_),
    .B1(_05636_),
    .B2(\top_ihp.oisc.regs[59][14] ),
    .A2(_05651_),
    .A1(\top_ihp.oisc.regs[55][14] ));
 sg13g2_nand3_1 _22650_ (.B(_06087_),
    .C(_06088_),
    .A(_06086_),
    .Y(_06089_));
 sg13g2_nor4_1 _22651_ (.A(_06072_),
    .B(_06078_),
    .C(_06085_),
    .D(_06089_),
    .Y(_06090_));
 sg13g2_nand4_1 _22652_ (.B(_06052_),
    .C(_06065_),
    .A(_06033_),
    .Y(_06091_),
    .D(_06090_));
 sg13g2_nor2b_1 _22653_ (.A(_06031_),
    .B_N(_06091_),
    .Y(_00425_));
 sg13g2_a22oi_1 _22654_ (.Y(_06092_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][15] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][15] ));
 sg13g2_a22oi_1 _22655_ (.Y(_06093_),
    .B1(_05652_),
    .B2(\top_ihp.oisc.regs[55][15] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][15] ));
 sg13g2_a22oi_1 _22656_ (.Y(_06094_),
    .B1(net155),
    .B2(\top_ihp.oisc.regs[39][15] ),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][15] ));
 sg13g2_a22oi_1 _22657_ (.Y(_06095_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][15] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][15] ));
 sg13g2_nand4_1 _22658_ (.B(_06093_),
    .C(_06094_),
    .A(_06092_),
    .Y(_06096_),
    .D(_06095_));
 sg13g2_a22oi_1 _22659_ (.Y(_06097_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][15] ),
    .A2(net304),
    .A1(\top_ihp.oisc.regs[58][15] ));
 sg13g2_a22oi_1 _22660_ (.Y(_06098_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][15] ),
    .A2(_05644_),
    .A1(\top_ihp.oisc.regs[35][15] ));
 sg13g2_a22oi_1 _22661_ (.Y(_06099_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][15] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[11][15] ));
 sg13g2_a22oi_1 _22662_ (.Y(_06100_),
    .B1(net428),
    .B2(\top_ihp.oisc.regs[17][15] ),
    .A2(_05415_),
    .A1(\top_ihp.oisc.regs[9][15] ));
 sg13g2_and2_1 _22663_ (.A(_06099_),
    .B(_06100_),
    .X(_06101_));
 sg13g2_nand2_1 _22664_ (.Y(_06102_),
    .A(_08287_),
    .B(net748));
 sg13g2_nand3_1 _22665_ (.B(net696),
    .C(_05825_),
    .A(\top_ihp.oisc.regs[14][15] ),
    .Y(_06103_));
 sg13g2_nand2_1 _22666_ (.Y(_06104_),
    .A(_06102_),
    .B(_06103_));
 sg13g2_a221oi_1 _22667_ (.B2(\top_ihp.oisc.regs[22][15] ),
    .C1(_06104_),
    .B1(net286),
    .A1(\top_ihp.oisc.regs[62][15] ),
    .Y(_06105_),
    .A2(net193));
 sg13g2_nand4_1 _22668_ (.B(_06098_),
    .C(_06101_),
    .A(_06097_),
    .Y(_06106_),
    .D(_06105_));
 sg13g2_a22oi_1 _22669_ (.Y(_06107_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][15] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][15] ));
 sg13g2_buf_8 _22670_ (.A(net452),
    .X(_06108_));
 sg13g2_a22oi_1 _22671_ (.Y(_06109_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][15] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][15] ));
 sg13g2_a22oi_1 _22672_ (.Y(_06110_),
    .B1(_05789_),
    .B2(\top_ihp.oisc.regs[33][15] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][15] ));
 sg13g2_a22oi_1 _22673_ (.Y(_06111_),
    .B1(net308),
    .B2(\top_ihp.oisc.regs[40][15] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[42][15] ));
 sg13g2_nand4_1 _22674_ (.B(_06109_),
    .C(_06110_),
    .A(_06107_),
    .Y(_06112_),
    .D(_06111_));
 sg13g2_buf_2 _22675_ (.A(_05551_),
    .X(_06113_));
 sg13g2_nor3_2 _22676_ (.A(_05531_),
    .B(_05915_),
    .C(net679),
    .Y(_06114_));
 sg13g2_a22oi_1 _22677_ (.Y(_06115_),
    .B1(_06114_),
    .B2(\top_ihp.oisc.regs[8][15] ),
    .A2(net284),
    .A1(\top_ihp.oisc.regs[48][15] ));
 sg13g2_a22oi_1 _22678_ (.Y(_06116_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][15] ),
    .A2(_05768_),
    .A1(\top_ihp.oisc.regs[36][15] ));
 sg13g2_buf_2 _22679_ (.A(_05588_),
    .X(_06117_));
 sg13g2_a22oi_1 _22680_ (.Y(_06118_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][15] ),
    .A2(_05338_),
    .A1(\top_ihp.oisc.regs[38][15] ));
 sg13g2_buf_2 _22681_ (.A(net696),
    .X(_06119_));
 sg13g2_a22oi_1 _22682_ (.Y(_06120_),
    .B1(net290),
    .B2(\top_ihp.oisc.regs[32][15] ),
    .A2(net669),
    .A1(\top_ihp.oisc.regs[44][15] ));
 sg13g2_nor2_1 _22683_ (.A(_05325_),
    .B(_06120_),
    .Y(_06121_));
 sg13g2_a21oi_1 _22684_ (.A1(\top_ihp.oisc.regs[51][15] ),
    .A2(_05759_),
    .Y(_06122_),
    .B1(_06121_));
 sg13g2_nand4_1 _22685_ (.B(_06116_),
    .C(_06118_),
    .A(_06115_),
    .Y(_06123_),
    .D(_06122_));
 sg13g2_nor4_1 _22686_ (.A(_06096_),
    .B(_06106_),
    .C(_06112_),
    .D(_06123_),
    .Y(_06124_));
 sg13g2_a22oi_1 _22687_ (.Y(_06125_),
    .B1(_05440_),
    .B2(\top_ihp.oisc.regs[31][15] ),
    .A2(_05570_),
    .A1(\top_ihp.oisc.regs[28][15] ));
 sg13g2_a221oi_1 _22688_ (.B2(\top_ihp.oisc.regs[25][15] ),
    .C1(net615),
    .B1(net722),
    .A1(\top_ihp.oisc.regs[24][15] ),
    .Y(_06126_),
    .A2(_05570_));
 sg13g2_a21oi_1 _22689_ (.A1(net434),
    .A2(_06125_),
    .Y(_06127_),
    .B1(_06126_));
 sg13g2_a22oi_1 _22690_ (.Y(_06128_),
    .B1(_06127_),
    .B2(_05998_),
    .A2(_05728_),
    .A1(\top_ihp.oisc.regs[10][15] ));
 sg13g2_a22oi_1 _22691_ (.Y(_06129_),
    .B1(_05817_),
    .B2(\top_ihp.oisc.regs[30][15] ),
    .A2(_05450_),
    .A1(\top_ihp.oisc.regs[21][15] ));
 sg13g2_a22oi_1 _22692_ (.Y(_06130_),
    .B1(_05444_),
    .B2(\top_ihp.oisc.regs[27][15] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[6][15] ));
 sg13g2_a22oi_1 _22693_ (.Y(_06131_),
    .B1(_05493_),
    .B2(\top_ihp.oisc.regs[26][15] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][15] ));
 sg13g2_and4_1 _22694_ (.A(_06128_),
    .B(_06129_),
    .C(_06130_),
    .D(_06131_),
    .X(_06132_));
 sg13g2_a22oi_1 _22695_ (.Y(_06133_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[13][15] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][15] ));
 sg13g2_buf_1 _22696_ (.A(net670),
    .X(_06134_));
 sg13g2_mux2_1 _22697_ (.A0(\top_ihp.oisc.regs[15][15] ),
    .A1(\top_ihp.oisc.regs[7][15] ),
    .S(net606),
    .X(_06135_));
 sg13g2_nand3_1 _22698_ (.B(_06134_),
    .C(_06135_),
    .A(net414),
    .Y(_06136_));
 sg13g2_nand3_1 _22699_ (.B(_06133_),
    .C(_06136_),
    .A(_06132_),
    .Y(_06137_));
 sg13g2_buf_1 _22700_ (.A(net438),
    .X(_06138_));
 sg13g2_mux2_1 _22701_ (.A0(\top_ihp.oisc.regs[20][15] ),
    .A1(\top_ihp.oisc.regs[16][15] ),
    .S(net418),
    .X(_06139_));
 sg13g2_a22oi_1 _22702_ (.Y(_06140_),
    .B1(_05950_),
    .B2(_06139_),
    .A2(net283),
    .A1(\top_ihp.oisc.regs[23][15] ));
 sg13g2_a22oi_1 _22703_ (.Y(_06141_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][15] ),
    .A2(_05489_),
    .A1(\top_ihp.oisc.regs[1][15] ));
 sg13g2_and2_1 _22704_ (.A(\top_ihp.oisc.regs[3][15] ),
    .B(_06017_),
    .X(_06142_));
 sg13g2_buf_1 _22705_ (.A(_05995_),
    .X(_06143_));
 sg13g2_a22oi_1 _22706_ (.Y(_06144_),
    .B1(_06142_),
    .B2(net596),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][15] ));
 sg13g2_a22oi_1 _22707_ (.Y(_06145_),
    .B1(net294),
    .B2(\top_ihp.oisc.regs[4][15] ),
    .A2(net445),
    .A1(\top_ihp.oisc.regs[19][15] ));
 sg13g2_nand4_1 _22708_ (.B(_06141_),
    .C(_06144_),
    .A(_06140_),
    .Y(_06146_),
    .D(_06145_));
 sg13g2_nand2_1 _22709_ (.Y(_06147_),
    .A(\top_ihp.oisc.regs[63][15] ),
    .B(net183));
 sg13g2_buf_1 _22710_ (.A(net306),
    .X(_06148_));
 sg13g2_a22oi_1 _22711_ (.Y(_06149_),
    .B1(_05742_),
    .B2(\top_ihp.oisc.regs[52][15] ),
    .A2(_06148_),
    .A1(\top_ihp.oisc.regs[34][15] ));
 sg13g2_nand2_1 _22712_ (.Y(_06150_),
    .A(_06147_),
    .B(_06149_));
 sg13g2_nor4_1 _22713_ (.A(net330),
    .B(_06137_),
    .C(_06146_),
    .D(_06150_),
    .Y(_06151_));
 sg13g2_a21o_1 _22714_ (.A2(net159),
    .A1(_00256_),
    .B1(net33),
    .X(_06152_));
 sg13g2_a22oi_1 _22715_ (.Y(_00426_),
    .B1(_06152_),
    .B2(_06102_),
    .A2(_06151_),
    .A1(_06124_));
 sg13g2_nor2_1 _22716_ (.A(net708),
    .B(net701),
    .Y(_06153_));
 sg13g2_buf_2 _22717_ (.A(_06153_),
    .X(_06154_));
 sg13g2_and4_1 _22718_ (.A(\top_ihp.oisc.regs[50][16] ),
    .B(net420),
    .C(_05901_),
    .D(_06154_),
    .X(_06155_));
 sg13g2_a21oi_1 _22719_ (.A1(\top_ihp.oisc.regs[27][16] ),
    .A2(net605),
    .Y(_06156_),
    .B1(_06155_));
 sg13g2_a22oi_1 _22720_ (.Y(_06157_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][16] ),
    .A2(net319),
    .A1(\top_ihp.oisc.regs[17][16] ));
 sg13g2_buf_2 _22721_ (.A(_06083_),
    .X(_06158_));
 sg13g2_a22oi_1 _22722_ (.Y(_06159_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][16] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[13][16] ));
 sg13g2_buf_2 _22723_ (.A(net721),
    .X(_06160_));
 sg13g2_nand3_1 _22724_ (.B(net608),
    .C(net695),
    .A(\top_ihp.oisc.regs[26][16] ),
    .Y(_06161_));
 sg13g2_buf_1 _22725_ (.A(net681),
    .X(_06162_));
 sg13g2_buf_1 _22726_ (.A(_05440_),
    .X(_06163_));
 sg13g2_nand3_1 _22727_ (.B(net595),
    .C(net694),
    .A(\top_ihp.oisc.regs[19][16] ),
    .Y(_06164_));
 sg13g2_nand2_1 _22728_ (.Y(_06165_),
    .A(_06161_),
    .B(_06164_));
 sg13g2_a22oi_1 _22729_ (.Y(_06166_),
    .B1(_06165_),
    .B2(net412),
    .A2(net294),
    .A1(\top_ihp.oisc.regs[4][16] ));
 sg13g2_nand4_1 _22730_ (.B(_06157_),
    .C(_06159_),
    .A(_06156_),
    .Y(_06167_),
    .D(_06166_));
 sg13g2_nand2_1 _22731_ (.Y(_06168_),
    .A(\top_ihp.oisc.regs[12][16] ),
    .B(net841));
 sg13g2_nand2_1 _22732_ (.Y(_06169_),
    .A(\top_ihp.oisc.regs[14][16] ),
    .B(net840));
 sg13g2_a21oi_1 _22733_ (.A1(_06168_),
    .A2(_06169_),
    .Y(_06170_),
    .B1(_05368_));
 sg13g2_nor2_1 _22734_ (.A(_05308_),
    .B(_05617_),
    .Y(_06171_));
 sg13g2_and3_1 _22735_ (.X(_06172_),
    .A(\top_ihp.oisc.regs[2][16] ),
    .B(net602),
    .C(net596));
 sg13g2_a221oi_1 _22736_ (.B2(\top_ihp.oisc.regs[40][16] ),
    .C1(_06172_),
    .B1(_06171_),
    .A1(net415),
    .Y(_06173_),
    .A2(_06170_));
 sg13g2_nor2_1 _22737_ (.A(net678),
    .B(net679),
    .Y(_06174_));
 sg13g2_nand4_1 _22738_ (.B(net420),
    .C(net671),
    .A(\top_ihp.oisc.regs[58][16] ),
    .Y(_06175_),
    .D(_06174_));
 sg13g2_o21ai_1 _22739_ (.B1(_06175_),
    .Y(_06176_),
    .A1(net414),
    .A2(_06173_));
 sg13g2_nor2_1 _22740_ (.A(_06167_),
    .B(_06176_),
    .Y(_06177_));
 sg13g2_a22oi_1 _22741_ (.Y(_06178_),
    .B1(net290),
    .B2(\top_ihp.oisc.regs[18][16] ),
    .A2(net669),
    .A1(\top_ihp.oisc.regs[30][16] ));
 sg13g2_a22oi_1 _22742_ (.Y(_06179_),
    .B1(_05758_),
    .B2(\top_ihp.oisc.regs[34][16] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][16] ));
 sg13g2_o21ai_1 _22743_ (.B1(_06179_),
    .Y(_06180_),
    .A1(_05419_),
    .A2(_06178_));
 sg13g2_a22oi_1 _22744_ (.Y(_06181_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[10][16] ),
    .A2(net444),
    .A1(\top_ihp.oisc.regs[21][16] ));
 sg13g2_nor2_2 _22745_ (.A(net613),
    .B(net700),
    .Y(_06182_));
 sg13g2_nand3_1 _22746_ (.B(_06182_),
    .C(_06174_),
    .A(\top_ihp.oisc.regs[56][16] ),
    .Y(_06183_));
 sg13g2_a22oi_1 _22747_ (.Y(_06184_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][16] ),
    .A2(_05714_),
    .A1(\top_ihp.oisc.regs[25][16] ));
 sg13g2_nand3_1 _22748_ (.B(_06183_),
    .C(_06184_),
    .A(_06181_),
    .Y(_06185_));
 sg13g2_nor3_1 _22749_ (.A(net331),
    .B(_06180_),
    .C(_06185_),
    .Y(_06186_));
 sg13g2_nand2_1 _22750_ (.Y(_06187_),
    .A(_08282_),
    .B(net739));
 sg13g2_a22oi_1 _22751_ (.Y(_06188_),
    .B1(_05500_),
    .B2(\top_ihp.oisc.regs[3][16] ),
    .A2(_05488_),
    .A1(\top_ihp.oisc.regs[1][16] ));
 sg13g2_a22oi_1 _22752_ (.Y(_06189_),
    .B1(net596),
    .B2(\top_ihp.oisc.regs[11][16] ),
    .A2(net670),
    .A1(\top_ihp.oisc.regs[15][16] ));
 sg13g2_nand2b_1 _22753_ (.Y(_06190_),
    .B(net601),
    .A_N(_06189_));
 sg13g2_a22oi_1 _22754_ (.Y(_06191_),
    .B1(_05456_),
    .B2(\top_ihp.oisc.regs[28][16] ),
    .A2(net449),
    .A1(\top_ihp.oisc.regs[20][16] ));
 sg13g2_nand4_1 _22755_ (.B(_06188_),
    .C(_06190_),
    .A(_06187_),
    .Y(_06192_),
    .D(_06191_));
 sg13g2_a22oi_1 _22756_ (.Y(_06193_),
    .B1(net450),
    .B2(\top_ihp.oisc.regs[6][16] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[7][16] ));
 sg13g2_a22oi_1 _22757_ (.Y(_06194_),
    .B1(net411),
    .B2(\top_ihp.oisc.regs[8][16] ),
    .A2(_05382_),
    .A1(\top_ihp.oisc.regs[5][16] ));
 sg13g2_nand2_1 _22758_ (.Y(_06195_),
    .A(_06193_),
    .B(_06194_));
 sg13g2_a22oi_1 _22759_ (.Y(_06196_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[53][16] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][16] ));
 sg13g2_nor4_2 _22760_ (.A(net613),
    .B(net678),
    .C(net700),
    .Y(_06197_),
    .D(_05317_));
 sg13g2_a22oi_1 _22761_ (.Y(_06198_),
    .B1(_06197_),
    .B2(\top_ihp.oisc.regs[60][16] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][16] ));
 sg13g2_nand2_1 _22762_ (.Y(_06199_),
    .A(_06196_),
    .B(_06198_));
 sg13g2_a22oi_1 _22763_ (.Y(_06200_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][16] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][16] ));
 sg13g2_a22oi_1 _22764_ (.Y(_06201_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[57][16] ),
    .A2(net433),
    .A1(\top_ihp.oisc.regs[35][16] ));
 sg13g2_and2_1 _22765_ (.A(\top_ihp.oisc.regs[9][16] ),
    .B(_05414_),
    .X(_06202_));
 sg13g2_a221oi_1 _22766_ (.B2(\top_ihp.oisc.regs[52][16] ),
    .C1(_06202_),
    .B1(_05741_),
    .A1(\top_ihp.oisc.regs[16][16] ),
    .Y(_06203_),
    .A2(_05357_));
 sg13g2_a22oi_1 _22767_ (.Y(_06204_),
    .B1(_05654_),
    .B2(\top_ihp.oisc.regs[41][16] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[59][16] ));
 sg13g2_nand4_1 _22768_ (.B(_06201_),
    .C(_06203_),
    .A(_06200_),
    .Y(_06205_),
    .D(_06204_));
 sg13g2_nor4_1 _22769_ (.A(_06192_),
    .B(_06195_),
    .C(_06199_),
    .D(_06205_),
    .Y(_06206_));
 sg13g2_a22oi_1 _22770_ (.Y(_06207_),
    .B1(_05771_),
    .B2(\top_ihp.oisc.regs[46][16] ),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][16] ));
 sg13g2_a22oi_1 _22771_ (.Y(_06208_),
    .B1(_06047_),
    .B2(\top_ihp.oisc.regs[49][16] ),
    .A2(_05551_),
    .A1(\top_ihp.oisc.regs[48][16] ));
 sg13g2_a22oi_1 _22772_ (.Y(_06209_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[47][16] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[44][16] ));
 sg13g2_a22oi_1 _22773_ (.Y(_06210_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][16] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][16] ));
 sg13g2_nand4_1 _22774_ (.B(_06208_),
    .C(_06209_),
    .A(_06207_),
    .Y(_06211_),
    .D(_06210_));
 sg13g2_a22oi_1 _22775_ (.Y(_06212_),
    .B1(net328),
    .B2(\top_ihp.oisc.regs[33][16] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][16] ));
 sg13g2_a22oi_1 _22776_ (.Y(_06213_),
    .B1(net155),
    .B2(\top_ihp.oisc.regs[39][16] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][16] ));
 sg13g2_mux2_1 _22777_ (.A0(\top_ihp.oisc.regs[31][16] ),
    .A1(\top_ihp.oisc.regs[23][16] ),
    .S(_05678_),
    .X(_06214_));
 sg13g2_nor2_2 _22778_ (.A(_05806_),
    .B(_05434_),
    .Y(_06215_));
 sg13g2_a22oi_1 _22779_ (.Y(_06216_),
    .B1(_06214_),
    .B2(_06215_),
    .A2(net324),
    .A1(\top_ihp.oisc.regs[63][16] ));
 sg13g2_a22oi_1 _22780_ (.Y(_06217_),
    .B1(_05485_),
    .B2(\top_ihp.oisc.regs[42][16] ),
    .A2(_05466_),
    .A1(\top_ihp.oisc.regs[62][16] ));
 sg13g2_nand4_1 _22781_ (.B(_06213_),
    .C(_06216_),
    .A(_06212_),
    .Y(_06218_),
    .D(_06217_));
 sg13g2_nor2_1 _22782_ (.A(_06211_),
    .B(_06218_),
    .Y(_06219_));
 sg13g2_and3_1 _22783_ (.X(_06220_),
    .A(_06186_),
    .B(_06206_),
    .C(_06219_));
 sg13g2_a21o_1 _22784_ (.A2(net159),
    .A1(_00257_),
    .B1(net33),
    .X(_06221_));
 sg13g2_a22oi_1 _22785_ (.Y(_00427_),
    .B1(_06221_),
    .B2(_06187_),
    .A2(_06220_),
    .A1(_06177_));
 sg13g2_a22oi_1 _22786_ (.Y(_06222_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][17] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[57][17] ));
 sg13g2_a22oi_1 _22787_ (.Y(_06223_),
    .B1(net78),
    .B2(\top_ihp.oisc.regs[59][17] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][17] ));
 sg13g2_a22oi_1 _22788_ (.Y(_06224_),
    .B1(net325),
    .B2(\top_ihp.oisc.regs[35][17] ),
    .A2(net324),
    .A1(\top_ihp.oisc.regs[63][17] ));
 sg13g2_a22oi_1 _22789_ (.Y(_06225_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][17] ),
    .A2(_05632_),
    .A1(\top_ihp.oisc.regs[38][17] ));
 sg13g2_nand4_1 _22790_ (.B(_06223_),
    .C(_06224_),
    .A(_06222_),
    .Y(_06226_),
    .D(_06225_));
 sg13g2_a22oi_1 _22791_ (.Y(_06227_),
    .B1(_05642_),
    .B2(\top_ihp.oisc.regs[51][17] ),
    .A2(net74),
    .A1(\top_ihp.oisc.regs[37][17] ));
 sg13g2_a22oi_1 _22792_ (.Y(_06228_),
    .B1(_05628_),
    .B2(\top_ihp.oisc.regs[50][17] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][17] ));
 sg13g2_a22oi_1 _22793_ (.Y(_06229_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][17] ),
    .A2(_05909_),
    .A1(\top_ihp.oisc.regs[36][17] ));
 sg13g2_a22oi_1 _22794_ (.Y(_06230_),
    .B1(_05968_),
    .B2(\top_ihp.oisc.regs[40][17] ),
    .A2(_05668_),
    .A1(\top_ihp.oisc.regs[62][17] ));
 sg13g2_nand4_1 _22795_ (.B(_06228_),
    .C(_06229_),
    .A(_06227_),
    .Y(_06231_),
    .D(_06230_));
 sg13g2_a22oi_1 _22796_ (.Y(_06232_),
    .B1(_05659_),
    .B2(\top_ihp.oisc.regs[47][17] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[42][17] ));
 sg13g2_buf_1 _22797_ (.A(net165),
    .X(_06233_));
 sg13g2_a22oi_1 _22798_ (.Y(_06234_),
    .B1(net70),
    .B2(\top_ihp.oisc.regs[45][17] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][17] ));
 sg13g2_buf_8 _22799_ (.A(net155),
    .X(_06235_));
 sg13g2_a22oi_1 _22800_ (.Y(_06236_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][17] ),
    .A2(net310),
    .A1(\top_ihp.oisc.regs[48][17] ));
 sg13g2_a22oi_1 _22801_ (.Y(_06237_),
    .B1(_05749_),
    .B2(\top_ihp.oisc.regs[53][17] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[33][17] ));
 sg13g2_nand4_1 _22802_ (.B(_06234_),
    .C(_06236_),
    .A(_06232_),
    .Y(_06238_),
    .D(_06237_));
 sg13g2_nor4_1 _22803_ (.A(net190),
    .B(_06226_),
    .C(_06231_),
    .D(_06238_),
    .Y(_06239_));
 sg13g2_buf_1 _22804_ (.A(_06022_),
    .X(_06240_));
 sg13g2_mux2_1 _22805_ (.A0(\top_ihp.oisc.regs[3][17] ),
    .A1(\top_ihp.oisc.regs[2][17] ),
    .S(net416),
    .X(_06241_));
 sg13g2_a22oi_1 _22806_ (.Y(_06242_),
    .B1(_06241_),
    .B2(net417),
    .A2(net410),
    .A1(\top_ihp.oisc.regs[10][17] ));
 sg13g2_nand2_1 _22807_ (.Y(_06243_),
    .A(\top_ihp.oisc.regs[8][17] ),
    .B(net411));
 sg13g2_mux2_1 _22808_ (.A0(\top_ihp.oisc.regs[28][17] ),
    .A1(\top_ihp.oisc.regs[20][17] ),
    .S(net675),
    .X(_06244_));
 sg13g2_a22oi_1 _22809_ (.Y(_06245_),
    .B1(_06244_),
    .B2(_05707_),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[13][17] ));
 sg13g2_a22oi_1 _22810_ (.Y(_06246_),
    .B1(net443),
    .B2(\top_ihp.oisc.regs[11][17] ),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][17] ));
 sg13g2_a22oi_1 _22811_ (.Y(_06247_),
    .B1(_05450_),
    .B2(\top_ihp.oisc.regs[21][17] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[12][17] ));
 sg13g2_and4_1 _22812_ (.A(_06243_),
    .B(_06245_),
    .C(_06246_),
    .D(_06247_),
    .X(_06248_));
 sg13g2_o21ai_1 _22813_ (.B1(_06248_),
    .Y(_06249_),
    .A1(_05409_),
    .A2(_06242_));
 sg13g2_a22oi_1 _22814_ (.Y(_06250_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][17] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][17] ));
 sg13g2_a22oi_1 _22815_ (.Y(_06251_),
    .B1(_05709_),
    .B2(\top_ihp.oisc.regs[19][17] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][17] ));
 sg13g2_a22oi_1 _22816_ (.Y(_06252_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][17] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][17] ));
 sg13g2_a22oi_1 _22817_ (.Y(_06253_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][17] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[17][17] ));
 sg13g2_nand4_1 _22818_ (.B(_06251_),
    .C(_06252_),
    .A(_06250_),
    .Y(_06254_),
    .D(_06253_));
 sg13g2_a22oi_1 _22819_ (.Y(_06255_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][17] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[31][17] ));
 sg13g2_buf_1 _22820_ (.A(_05384_),
    .X(_06256_));
 sg13g2_a22oi_1 _22821_ (.Y(_06257_),
    .B1(net283),
    .B2(\top_ihp.oisc.regs[23][17] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][17] ));
 sg13g2_a22oi_1 _22822_ (.Y(_06258_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][17] ),
    .A2(net297),
    .A1(\top_ihp.oisc.regs[5][17] ));
 sg13g2_nor4_1 _22823_ (.A(net418),
    .B(net414),
    .C(_05529_),
    .D(net413),
    .Y(_06259_));
 sg13g2_buf_1 _22824_ (.A(net701),
    .X(_06260_));
 sg13g2_mux2_1 _22825_ (.A0(\top_ihp.oisc.regs[54][17] ),
    .A1(\top_ihp.oisc.regs[52][17] ),
    .S(net668),
    .X(_06261_));
 sg13g2_a22oi_1 _22826_ (.Y(_06262_),
    .B1(_06259_),
    .B2(_06261_),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[1][17] ));
 sg13g2_nand4_1 _22827_ (.B(_06257_),
    .C(_06258_),
    .A(_06255_),
    .Y(_06263_),
    .D(_06262_));
 sg13g2_a22oi_1 _22828_ (.Y(_06264_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][17] ),
    .A2(net302),
    .A1(\top_ihp.oisc.regs[32][17] ));
 sg13g2_a22oi_1 _22829_ (.Y(_06265_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][17] ),
    .A2(_05494_),
    .A1(\top_ihp.oisc.regs[26][17] ));
 sg13g2_a22oi_1 _22830_ (.Y(_06266_),
    .B1(_05850_),
    .B2(\top_ihp.oisc.regs[4][17] ),
    .A2(net670),
    .A1(\top_ihp.oisc.regs[6][17] ));
 sg13g2_nor2b_1 _22831_ (.A(_06266_),
    .B_N(_06002_),
    .Y(_06267_));
 sg13g2_a221oi_1 _22832_ (.B2(\top_ihp.oisc.regs[14][17] ),
    .C1(_06267_),
    .B1(_05733_),
    .A1(net1052),
    .Y(_06268_),
    .A2(net739));
 sg13g2_and2_1 _22833_ (.A(_06265_),
    .B(_06268_),
    .X(_06269_));
 sg13g2_a22oi_1 _22834_ (.Y(_06270_),
    .B1(_05655_),
    .B2(\top_ihp.oisc.regs[41][17] ),
    .A2(_06108_),
    .A1(\top_ihp.oisc.regs[60][17] ));
 sg13g2_a22oi_1 _22835_ (.Y(_06271_),
    .B1(net304),
    .B2(\top_ihp.oisc.regs[58][17] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][17] ));
 sg13g2_nand4_1 _22836_ (.B(_06269_),
    .C(_06270_),
    .A(_06264_),
    .Y(_06272_),
    .D(_06271_));
 sg13g2_nor4_1 _22837_ (.A(_06249_),
    .B(_06254_),
    .C(_06263_),
    .D(_06272_),
    .Y(_06273_));
 sg13g2_a21oi_1 _22838_ (.A1(_00258_),
    .A2(net330),
    .Y(_06274_),
    .B1(_05623_));
 sg13g2_a21oi_1 _22839_ (.A1(_08274_),
    .A2(net718),
    .Y(_06275_),
    .B1(_06274_));
 sg13g2_a21oi_1 _22840_ (.A1(_06239_),
    .A2(_06273_),
    .Y(_00428_),
    .B1(_06275_));
 sg13g2_buf_1 _22841_ (.A(net446),
    .X(_06276_));
 sg13g2_a22oi_1 _22842_ (.Y(_06277_),
    .B1(_05669_),
    .B2(\top_ihp.oisc.regs[46][18] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][18] ));
 sg13g2_a22oi_1 _22843_ (.Y(_06278_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[47][18] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][18] ));
 sg13g2_a22oi_1 _22844_ (.Y(_06279_),
    .B1(_05922_),
    .B2(\top_ihp.oisc.regs[63][18] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][18] ));
 sg13g2_a22oi_1 _22845_ (.Y(_06280_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][18] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][18] ));
 sg13g2_nand4_1 _22846_ (.B(_06278_),
    .C(_06279_),
    .A(_06277_),
    .Y(_06281_),
    .D(_06280_));
 sg13g2_a22oi_1 _22847_ (.Y(_06282_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][18] ),
    .A2(_05661_),
    .A1(\top_ihp.oisc.regs[45][18] ));
 sg13g2_a22oi_1 _22848_ (.Y(_06283_),
    .B1(_05978_),
    .B2(\top_ihp.oisc.regs[36][18] ),
    .A2(_05668_),
    .A1(\top_ihp.oisc.regs[62][18] ));
 sg13g2_a22oi_1 _22849_ (.Y(_06284_),
    .B1(_05926_),
    .B2(\top_ihp.oisc.regs[52][18] ),
    .A2(_05662_),
    .A1(\top_ihp.oisc.regs[58][18] ));
 sg13g2_a22oi_1 _22850_ (.Y(_06285_),
    .B1(_05752_),
    .B2(\top_ihp.oisc.regs[34][18] ),
    .A2(net328),
    .A1(\top_ihp.oisc.regs[33][18] ));
 sg13g2_nand4_1 _22851_ (.B(_06283_),
    .C(_06284_),
    .A(_06282_),
    .Y(_06286_),
    .D(_06285_));
 sg13g2_buf_2 _22852_ (.A(_05484_),
    .X(_06287_));
 sg13g2_a22oi_1 _22853_ (.Y(_06288_),
    .B1(_05749_),
    .B2(\top_ihp.oisc.regs[53][18] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][18] ));
 sg13g2_a22oi_1 _22854_ (.Y(_06289_),
    .B1(_06197_),
    .B2(\top_ihp.oisc.regs[60][18] ),
    .A2(_05784_),
    .A1(\top_ihp.oisc.regs[50][18] ));
 sg13g2_nand3_1 _22855_ (.B(net599),
    .C(net600),
    .A(\top_ihp.oisc.regs[5][18] ),
    .Y(_06290_));
 sg13g2_nand3_1 _22856_ (.B(net607),
    .C(net597),
    .A(\top_ihp.oisc.regs[15][18] ),
    .Y(_06291_));
 sg13g2_a21oi_1 _22857_ (.A1(_06290_),
    .A2(_06291_),
    .Y(_06292_),
    .B1(net420));
 sg13g2_a221oi_1 _22858_ (.B2(\top_ihp.oisc.regs[23][18] ),
    .C1(_06292_),
    .B1(net283),
    .A1(\top_ihp.oisc.regs[37][18] ),
    .Y(_06293_),
    .A2(net192));
 sg13g2_buf_2 _22859_ (.A(net182),
    .X(_06294_));
 sg13g2_a22oi_1 _22860_ (.Y(_06295_),
    .B1(net68),
    .B2(\top_ihp.oisc.regs[55][18] ),
    .A2(_05970_),
    .A1(\top_ihp.oisc.regs[38][18] ));
 sg13g2_nand4_1 _22861_ (.B(_06289_),
    .C(_06293_),
    .A(_06288_),
    .Y(_06296_),
    .D(_06295_));
 sg13g2_nor4_1 _22862_ (.A(_05626_),
    .B(_06281_),
    .C(_06286_),
    .D(_06296_),
    .Y(_06297_));
 sg13g2_a22oi_1 _22863_ (.Y(_06298_),
    .B1(_05600_),
    .B2(\top_ihp.oisc.regs[41][18] ),
    .A2(_05641_),
    .A1(\top_ihp.oisc.regs[51][18] ));
 sg13g2_a22oi_1 _22864_ (.Y(_06299_),
    .B1(net298),
    .B2(\top_ihp.oisc.regs[48][18] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][18] ));
 sg13g2_a22oi_1 _22865_ (.Y(_06300_),
    .B1(net325),
    .B2(\top_ihp.oisc.regs[35][18] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[59][18] ));
 sg13g2_a22oi_1 _22866_ (.Y(_06301_),
    .B1(_05640_),
    .B2(\top_ihp.oisc.regs[49][18] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[44][18] ));
 sg13g2_nand4_1 _22867_ (.B(_06299_),
    .C(_06300_),
    .A(_06298_),
    .Y(_06302_),
    .D(_06301_));
 sg13g2_a22oi_1 _22868_ (.Y(_06303_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[10][18] ),
    .A2(_05388_),
    .A1(\top_ihp.oisc.regs[6][18] ));
 sg13g2_a22oi_1 _22869_ (.Y(_06304_),
    .B1(_05500_),
    .B2(\top_ihp.oisc.regs[3][18] ),
    .A2(_05436_),
    .A1(\top_ihp.oisc.regs[19][18] ));
 sg13g2_a22oi_1 _22870_ (.Y(_06305_),
    .B1(net336),
    .B2(\top_ihp.oisc.regs[13][18] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[8][18] ));
 sg13g2_a22oi_1 _22871_ (.Y(_06306_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][18] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[17][18] ));
 sg13g2_and4_1 _22872_ (.A(_06303_),
    .B(_06304_),
    .C(_06305_),
    .D(_06306_),
    .X(_06307_));
 sg13g2_buf_2 _22873_ (.A(net286),
    .X(_06308_));
 sg13g2_a22oi_1 _22874_ (.Y(_06309_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][18] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[27][18] ));
 sg13g2_a22oi_1 _22875_ (.Y(_06310_),
    .B1(_05510_),
    .B2(\top_ihp.oisc.regs[25][18] ),
    .A2(net294),
    .A1(\top_ihp.oisc.regs[4][18] ));
 sg13g2_nand3_1 _22876_ (.B(_06309_),
    .C(_06310_),
    .A(_06307_),
    .Y(_06311_));
 sg13g2_buf_1 _22877_ (.A(net739),
    .X(_06312_));
 sg13g2_nor2_2 _22878_ (.A(net615),
    .B(_05355_),
    .Y(_06313_));
 sg13g2_a22oi_1 _22879_ (.Y(_06314_),
    .B1(_05410_),
    .B2(\top_ihp.oisc.regs[2][18] ),
    .A2(_06313_),
    .A1(\top_ihp.oisc.regs[16][18] ));
 sg13g2_inv_1 _22880_ (.Y(_06315_),
    .A(_06314_));
 sg13g2_a21o_1 _22881_ (.A2(_05392_),
    .A1(_05365_),
    .B1(_03728_),
    .X(_06316_));
 sg13g2_buf_2 _22882_ (.A(_06316_),
    .X(_06317_));
 sg13g2_a22oi_1 _22883_ (.Y(_06318_),
    .B1(_06317_),
    .B2(\top_ihp.oisc.regs[1][18] ),
    .A2(net670),
    .A1(\top_ihp.oisc.regs[7][18] ));
 sg13g2_nand3_1 _22884_ (.B(net597),
    .C(net410),
    .A(\top_ihp.oisc.regs[14][18] ),
    .Y(_06319_));
 sg13g2_o21ai_1 _22885_ (.B1(_06319_),
    .Y(_06320_),
    .A1(_05498_),
    .A2(_06318_));
 sg13g2_a221oi_1 _22886_ (.B2(_06315_),
    .C1(_06320_),
    .B1(net417),
    .A1(_08221_),
    .Y(_06321_),
    .A2(net720));
 sg13g2_nand3_1 _22887_ (.B(_06014_),
    .C(_06174_),
    .A(\top_ihp.oisc.regs[57][18] ),
    .Y(_06322_));
 sg13g2_nand2_1 _22888_ (.Y(_06323_),
    .A(\top_ihp.oisc.regs[21][18] ),
    .B(net444));
 sg13g2_a22oi_1 _22889_ (.Y(_06324_),
    .B1(_05723_),
    .B2(\top_ihp.oisc.regs[9][18] ),
    .A2(_05397_),
    .A1(\top_ihp.oisc.regs[12][18] ));
 sg13g2_nand4_1 _22890_ (.B(_06322_),
    .C(_06323_),
    .A(_06321_),
    .Y(_06325_),
    .D(_06324_));
 sg13g2_a22oi_1 _22891_ (.Y(_06326_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][18] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][18] ));
 sg13g2_a22oi_1 _22892_ (.Y(_06327_),
    .B1(_05725_),
    .B2(\top_ihp.oisc.regs[29][18] ),
    .A2(_05688_),
    .A1(\top_ihp.oisc.regs[11][18] ));
 sg13g2_a22oi_1 _22893_ (.Y(_06328_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[31][18] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[26][18] ));
 sg13g2_a22oi_1 _22894_ (.Y(_06329_),
    .B1(net296),
    .B2(\top_ihp.oisc.regs[28][18] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][18] ));
 sg13g2_nand4_1 _22895_ (.B(_06327_),
    .C(_06328_),
    .A(_06326_),
    .Y(_06330_),
    .D(_06329_));
 sg13g2_nor4_1 _22896_ (.A(_06302_),
    .B(_06311_),
    .C(_06325_),
    .D(_06330_),
    .Y(_06331_));
 sg13g2_a21oi_1 _22897_ (.A1(_00259_),
    .A2(_05616_),
    .Y(_06332_),
    .B1(net34));
 sg13g2_a21oi_1 _22898_ (.A1(_08221_),
    .A2(net718),
    .Y(_06333_),
    .B1(_06332_));
 sg13g2_a21oi_1 _22899_ (.A1(_06297_),
    .A2(_06331_),
    .Y(_00429_),
    .B1(_06333_));
 sg13g2_buf_8 _22900_ (.A(net162),
    .X(_06334_));
 sg13g2_a22oi_1 _22901_ (.Y(_06335_),
    .B1(_06334_),
    .B2(\top_ihp.oisc.regs[61][19] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][19] ));
 sg13g2_a22oi_1 _22902_ (.Y(_06336_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[45][19] ),
    .A2(net193),
    .A1(\top_ihp.oisc.regs[62][19] ));
 sg13g2_a22oi_1 _22903_ (.Y(_06337_),
    .B1(_05658_),
    .B2(\top_ihp.oisc.regs[47][19] ),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][19] ));
 sg13g2_a22oi_1 _22904_ (.Y(_06338_),
    .B1(_05779_),
    .B2(\top_ihp.oisc.regs[56][19] ),
    .A2(_05909_),
    .A1(\top_ihp.oisc.regs[36][19] ));
 sg13g2_nand4_1 _22905_ (.B(_06336_),
    .C(_06337_),
    .A(_06335_),
    .Y(_06339_),
    .D(_06338_));
 sg13g2_a22oi_1 _22906_ (.Y(_06340_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][19] ),
    .A2(net296),
    .A1(\top_ihp.oisc.regs[28][19] ));
 sg13g2_a22oi_1 _22907_ (.Y(_06341_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][19] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][19] ));
 sg13g2_mux2_1 _22908_ (.A0(\top_ihp.oisc.regs[29][19] ),
    .A1(\top_ihp.oisc.regs[21][19] ),
    .S(net606),
    .X(_06342_));
 sg13g2_a22oi_1 _22909_ (.Y(_06343_),
    .B1(_05807_),
    .B2(_06342_),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][19] ));
 sg13g2_a22oi_1 _22910_ (.Y(_06344_),
    .B1(net317),
    .B2(\top_ihp.oisc.regs[1][19] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][19] ));
 sg13g2_nand4_1 _22911_ (.B(_06341_),
    .C(_06343_),
    .A(_06340_),
    .Y(_06345_),
    .D(_06344_));
 sg13g2_a22oi_1 _22912_ (.Y(_06346_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][19] ),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][19] ));
 sg13g2_nand2_1 _22913_ (.Y(_06347_),
    .A(\top_ihp.oisc.regs[38][19] ),
    .B(_05970_));
 sg13g2_nor2_1 _22914_ (.A(_05565_),
    .B(_05599_),
    .Y(_06348_));
 sg13g2_nor2_1 _22915_ (.A(_05578_),
    .B(net668),
    .Y(_06349_));
 sg13g2_a22oi_1 _22916_ (.Y(_06350_),
    .B1(_06349_),
    .B2(\top_ihp.oisc.regs[18][19] ),
    .A2(_06348_),
    .A1(\top_ihp.oisc.regs[20][19] ));
 sg13g2_nor3_2 _22917_ (.A(net413),
    .B(_05568_),
    .C(_06350_),
    .Y(_06351_));
 sg13g2_a21oi_1 _22918_ (.A1(\top_ihp.oisc.regs[42][19] ),
    .A2(net279),
    .Y(_06352_),
    .B1(_06351_));
 sg13g2_nand3_1 _22919_ (.B(_06347_),
    .C(_06352_),
    .A(_06346_),
    .Y(_06353_));
 sg13g2_buf_8 _22920_ (.A(net332),
    .X(_06354_));
 sg13g2_a22oi_1 _22921_ (.Y(_06355_),
    .B1(net294),
    .B2(\top_ihp.oisc.regs[4][19] ),
    .A2(net151),
    .A1(\top_ihp.oisc.regs[3][19] ));
 sg13g2_a22oi_1 _22922_ (.Y(_06356_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][19] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[13][19] ));
 sg13g2_nand3_1 _22923_ (.B(net607),
    .C(net695),
    .A(\top_ihp.oisc.regs[26][19] ),
    .Y(_06357_));
 sg13g2_nand3_1 _22924_ (.B(net674),
    .C(net698),
    .A(\top_ihp.oisc.regs[19][19] ),
    .Y(_06358_));
 sg13g2_a21oi_1 _22925_ (.A1(_06357_),
    .A2(_06358_),
    .Y(_06359_),
    .B1(net320));
 sg13g2_a221oi_1 _22926_ (.B2(\top_ihp.oisc.regs[15][19] ),
    .C1(_06359_),
    .B1(_05719_),
    .A1(\top_ihp.oisc.regs[12][19] ),
    .Y(_06360_),
    .A2(net448));
 sg13g2_mux2_1 _22927_ (.A0(\top_ihp.oisc.regs[31][19] ),
    .A1(\top_ihp.oisc.regs[23][19] ),
    .S(net681),
    .X(_06361_));
 sg13g2_nand3_1 _22928_ (.B(net694),
    .C(_06361_),
    .A(net320),
    .Y(_06362_));
 sg13g2_nand4_1 _22929_ (.B(net412),
    .C(net413),
    .A(\top_ihp.oisc.regs[24][19] ),
    .Y(_06363_),
    .D(net673));
 sg13g2_and2_1 _22930_ (.A(_06362_),
    .B(_06363_),
    .X(_06364_));
 sg13g2_nand4_1 _22931_ (.B(_06356_),
    .C(_06360_),
    .A(_06355_),
    .Y(_06365_),
    .D(_06364_));
 sg13g2_nor4_1 _22932_ (.A(_06339_),
    .B(_06345_),
    .C(_06353_),
    .D(_06365_),
    .Y(_06366_));
 sg13g2_a22oi_1 _22933_ (.Y(_06367_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[57][19] ),
    .A2(_05537_),
    .A1(\top_ihp.oisc.regs[63][19] ));
 sg13g2_a22oi_1 _22934_ (.Y(_06368_),
    .B1(_05627_),
    .B2(\top_ihp.oisc.regs[50][19] ),
    .A2(_05429_),
    .A1(\top_ihp.oisc.regs[32][19] ));
 sg13g2_a22oi_1 _22935_ (.Y(_06369_),
    .B1(_05563_),
    .B2(\top_ihp.oisc.regs[34][19] ),
    .A2(_05539_),
    .A1(\top_ihp.oisc.regs[55][19] ));
 sg13g2_a22oi_1 _22936_ (.Y(_06370_),
    .B1(_05741_),
    .B2(\top_ihp.oisc.regs[52][19] ),
    .A2(_05326_),
    .A1(\top_ihp.oisc.regs[44][19] ));
 sg13g2_nand4_1 _22937_ (.B(_06368_),
    .C(_06369_),
    .A(_06367_),
    .Y(_06371_),
    .D(_06370_));
 sg13g2_a22oi_1 _22938_ (.Y(_06372_),
    .B1(_05553_),
    .B2(\top_ihp.oisc.regs[39][19] ),
    .A2(_05309_),
    .A1(\top_ihp.oisc.regs[60][19] ));
 sg13g2_a22oi_1 _22939_ (.Y(_06373_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[58][19] ),
    .A2(_05460_),
    .A1(\top_ihp.oisc.regs[49][19] ));
 sg13g2_and2_1 _22940_ (.A(\top_ihp.oisc.regs[14][19] ),
    .B(_05733_),
    .X(_06374_));
 sg13g2_a221oi_1 _22941_ (.B2(\top_ihp.oisc.regs[35][19] ),
    .C1(_06374_),
    .B1(_05560_),
    .A1(\top_ihp.oisc.regs[8][19] ),
    .Y(_06375_),
    .A2(_05395_));
 sg13g2_a22oi_1 _22942_ (.Y(_06376_),
    .B1(_05653_),
    .B2(\top_ihp.oisc.regs[41][19] ),
    .A2(_05516_),
    .A1(\top_ihp.oisc.regs[54][19] ));
 sg13g2_nand4_1 _22943_ (.B(_06373_),
    .C(_06375_),
    .A(_06372_),
    .Y(_06377_),
    .D(_06376_));
 sg13g2_or2_1 _22944_ (.X(_06378_),
    .B(_06377_),
    .A(_06371_));
 sg13g2_a22oi_1 _22945_ (.Y(_06379_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][19] ),
    .A2(net319),
    .A1(\top_ihp.oisc.regs[17][19] ));
 sg13g2_a22oi_1 _22946_ (.Y(_06380_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][19] ),
    .A2(net314),
    .A1(\top_ihp.oisc.regs[9][19] ));
 sg13g2_a22oi_1 _22947_ (.Y(_06381_),
    .B1(net297),
    .B2(\top_ihp.oisc.regs[5][19] ),
    .A2(net728),
    .A1(_08223_));
 sg13g2_nand3_1 _22948_ (.B(_06380_),
    .C(_06381_),
    .A(_06379_),
    .Y(_06382_));
 sg13g2_buf_8 _22949_ (.A(net169),
    .X(_06383_));
 sg13g2_nand2_1 _22950_ (.Y(_06384_),
    .A(\top_ihp.oisc.regs[46][19] ),
    .B(net66));
 sg13g2_a22oi_1 _22951_ (.Y(_06385_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][19] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][19] ));
 sg13g2_a22oi_1 _22952_ (.Y(_06386_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][19] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][19] ));
 sg13g2_a22oi_1 _22953_ (.Y(_06387_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][19] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[33][19] ));
 sg13g2_nand4_1 _22954_ (.B(_06385_),
    .C(_06386_),
    .A(_06384_),
    .Y(_06388_),
    .D(_06387_));
 sg13g2_nor4_1 _22955_ (.A(net158),
    .B(_06378_),
    .C(_06382_),
    .D(_06388_),
    .Y(_06389_));
 sg13g2_buf_1 _22956_ (.A(net728),
    .X(_06390_));
 sg13g2_a21oi_1 _22957_ (.A1(_00260_),
    .A2(net330),
    .Y(_06391_),
    .B1(net34));
 sg13g2_a21oi_1 _22958_ (.A1(_08223_),
    .A2(net693),
    .Y(_06392_),
    .B1(_06391_));
 sg13g2_a21oi_1 _22959_ (.A1(_06366_),
    .A2(_06389_),
    .Y(_00430_),
    .B1(_06392_));
 sg13g2_nand2_1 _22960_ (.Y(_06393_),
    .A(\top_ihp.oisc.regs[46][1] ),
    .B(net66));
 sg13g2_a22oi_1 _22961_ (.Y(_06394_),
    .B1(net327),
    .B2(\top_ihp.oisc.regs[49][1] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][1] ));
 sg13g2_a22oi_1 _22962_ (.Y(_06395_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][1] ),
    .A2(net306),
    .A1(\top_ihp.oisc.regs[34][1] ));
 sg13g2_a22oi_1 _22963_ (.Y(_06396_),
    .B1(net77),
    .B2(\top_ihp.oisc.regs[55][1] ),
    .A2(net328),
    .A1(\top_ihp.oisc.regs[33][1] ));
 sg13g2_nand4_1 _22964_ (.B(_06394_),
    .C(_06395_),
    .A(_06393_),
    .Y(_06397_),
    .D(_06396_));
 sg13g2_a22oi_1 _22965_ (.Y(_06398_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[50][1] ),
    .A2(_05751_),
    .A1(\top_ihp.oisc.regs[40][1] ));
 sg13g2_a22oi_1 _22966_ (.Y(_06399_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][1] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[63][1] ));
 sg13g2_a22oi_1 _22967_ (.Y(_06400_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][1] ),
    .A2(net78),
    .A1(\top_ihp.oisc.regs[59][1] ));
 sg13g2_a22oi_1 _22968_ (.Y(_06401_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][1] ),
    .A2(net155),
    .A1(\top_ihp.oisc.regs[39][1] ));
 sg13g2_nand4_1 _22969_ (.B(_06399_),
    .C(_06400_),
    .A(_06398_),
    .Y(_06402_),
    .D(_06401_));
 sg13g2_buf_8 _22970_ (.A(net193),
    .X(_06403_));
 sg13g2_a22oi_1 _22971_ (.Y(_06404_),
    .B1(net67),
    .B2(\top_ihp.oisc.regs[61][1] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][1] ));
 sg13g2_a22oi_1 _22972_ (.Y(_06405_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][1] ),
    .A2(_05328_),
    .A1(\top_ihp.oisc.regs[44][1] ));
 sg13g2_a22oi_1 _22973_ (.Y(_06406_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][1] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][1] ));
 sg13g2_a22oi_1 _22974_ (.Y(_06407_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][1] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][1] ));
 sg13g2_nand4_1 _22975_ (.B(_06405_),
    .C(_06406_),
    .A(_06404_),
    .Y(_06408_),
    .D(_06407_));
 sg13g2_nor4_1 _22976_ (.A(net190),
    .B(_06397_),
    .C(_06402_),
    .D(_06408_),
    .Y(_06409_));
 sg13g2_a22oi_1 _22977_ (.Y(_06410_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[45][1] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][1] ));
 sg13g2_a22oi_1 _22978_ (.Y(_06411_),
    .B1(net333),
    .B2(\top_ihp.oisc.regs[26][1] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][1] ));
 sg13g2_a22oi_1 _22979_ (.Y(_06412_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][1] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][1] ));
 sg13g2_nand4_1 _22980_ (.B(net420),
    .C(net595),
    .A(\top_ihp.oisc.regs[6][1] ),
    .Y(_06413_),
    .D(net597));
 sg13g2_mux2_1 _22981_ (.A0(\top_ihp.oisc.regs[13][1] ),
    .A1(\top_ihp.oisc.regs[5][1] ),
    .S(net675),
    .X(_06414_));
 sg13g2_nand3_1 _22982_ (.B(net600),
    .C(_06414_),
    .A(net414),
    .Y(_06415_));
 sg13g2_and2_1 _22983_ (.A(_06413_),
    .B(_06415_),
    .X(_06416_));
 sg13g2_nand4_1 _22984_ (.B(_06411_),
    .C(_06412_),
    .A(_06410_),
    .Y(_06417_),
    .D(_06416_));
 sg13g2_nor2_1 _22985_ (.A(_05360_),
    .B(_05393_),
    .Y(_06418_));
 sg13g2_mux2_1 _22986_ (.A0(\top_ihp.oisc.regs[9][1] ),
    .A1(\top_ihp.oisc.regs[1][1] ),
    .S(net606),
    .X(_06419_));
 sg13g2_a22oi_1 _22987_ (.Y(_06420_),
    .B1(_06418_),
    .B2(_06419_),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][1] ));
 sg13g2_a22oi_1 _22988_ (.Y(_06421_),
    .B1(net283),
    .B2(\top_ihp.oisc.regs[23][1] ),
    .A2(net445),
    .A1(\top_ihp.oisc.regs[19][1] ));
 sg13g2_a22oi_1 _22989_ (.Y(_06422_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][1] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][1] ));
 sg13g2_a22oi_1 _22990_ (.Y(_06423_),
    .B1(net151),
    .B2(\top_ihp.oisc.regs[3][1] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][1] ));
 sg13g2_nand4_1 _22991_ (.B(_06421_),
    .C(_06422_),
    .A(_06420_),
    .Y(_06424_),
    .D(_06423_));
 sg13g2_mux2_1 _22992_ (.A0(\top_ihp.oisc.regs[29][1] ),
    .A1(\top_ihp.oisc.regs[21][1] ),
    .S(net595),
    .X(_06425_));
 sg13g2_a22oi_1 _22993_ (.Y(_06426_),
    .B1(_06425_),
    .B2(_05807_),
    .A2(_05686_),
    .A1(\top_ihp.oisc.regs[17][1] ));
 sg13g2_a22oi_1 _22994_ (.Y(_06427_),
    .B1(_05715_),
    .B2(\top_ihp.oisc.regs[25][1] ),
    .A2(net296),
    .A1(\top_ihp.oisc.regs[28][1] ));
 sg13g2_mux2_1 _22995_ (.A0(\top_ihp.oisc.regs[15][1] ),
    .A1(\top_ihp.oisc.regs[14][1] ),
    .S(net416),
    .X(_06428_));
 sg13g2_nor2_2 _22996_ (.A(_05566_),
    .B(_05599_),
    .Y(_06429_));
 sg13g2_and4_1 _22997_ (.A(\top_ihp.oisc.regs[53][1] ),
    .B(_05548_),
    .C(_05535_),
    .D(_06429_),
    .X(_06430_));
 sg13g2_a21oi_1 _22998_ (.A1(_05376_),
    .A2(_06428_),
    .Y(_06431_),
    .B1(_06430_));
 sg13g2_nand3_1 _22999_ (.B(net416),
    .C(net596),
    .A(\top_ihp.oisc.regs[2][1] ),
    .Y(_06432_));
 sg13g2_buf_1 _23000_ (.A(net680),
    .X(_06433_));
 sg13g2_nand3_1 _23001_ (.B(net594),
    .C(net597),
    .A(\top_ihp.oisc.regs[7][1] ),
    .Y(_06434_));
 sg13g2_nand2_1 _23002_ (.Y(_06435_),
    .A(_06432_),
    .B(_06434_));
 sg13g2_a22oi_1 _23003_ (.Y(_06436_),
    .B1(_06435_),
    .B2(net417),
    .A2(_06083_),
    .A1(\top_ihp.oisc.regs[24][1] ));
 sg13g2_nand4_1 _23004_ (.B(_06427_),
    .C(_06431_),
    .A(_06426_),
    .Y(_06437_),
    .D(_06436_));
 sg13g2_a22oi_1 _23005_ (.Y(_06438_),
    .B1(net436),
    .B2(\top_ihp.oisc.regs[4][1] ),
    .A2(_05395_),
    .A1(\top_ihp.oisc.regs[8][1] ));
 sg13g2_a22oi_1 _23006_ (.Y(_06439_),
    .B1(_05440_),
    .B2(\top_ihp.oisc.regs[31][1] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[30][1] ));
 sg13g2_inv_1 _23007_ (.Y(_06440_),
    .A(_06439_));
 sg13g2_a22oi_1 _23008_ (.Y(_06441_),
    .B1(net669),
    .B2(_06440_),
    .A2(_03715_),
    .A1(_08317_));
 sg13g2_nand3_1 _23009_ (.B(net601),
    .C(_06143_),
    .A(\top_ihp.oisc.regs[11][1] ),
    .Y(_06442_));
 sg13g2_nand3_1 _23010_ (.B(_06441_),
    .C(_06442_),
    .A(_06438_),
    .Y(_06443_));
 sg13g2_a221oi_1 _23011_ (.B2(\top_ihp.oisc.regs[36][1] ),
    .C1(_06443_),
    .B1(net170),
    .A1(\top_ihp.oisc.regs[37][1] ),
    .Y(_06444_),
    .A2(_05761_));
 sg13g2_a22oi_1 _23012_ (.Y(_06445_),
    .B1(net287),
    .B2(\top_ihp.oisc.regs[43][1] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][1] ));
 sg13g2_a22oi_1 _23013_ (.Y(_06446_),
    .B1(_05772_),
    .B2(\top_ihp.oisc.regs[41][1] ),
    .A2(net304),
    .A1(\top_ihp.oisc.regs[58][1] ));
 sg13g2_nand3_1 _23014_ (.B(_06445_),
    .C(_06446_),
    .A(_06444_),
    .Y(_06447_));
 sg13g2_nor4_1 _23015_ (.A(_06417_),
    .B(_06424_),
    .C(_06437_),
    .D(_06447_),
    .Y(_06448_));
 sg13g2_a21oi_1 _23016_ (.A1(_00242_),
    .A2(net330),
    .Y(_06449_),
    .B1(net34));
 sg13g2_a21oi_1 _23017_ (.A1(_08317_),
    .A2(net693),
    .Y(_06450_),
    .B1(_06449_));
 sg13g2_a21oi_1 _23018_ (.A1(_06409_),
    .A2(_06448_),
    .Y(_00431_),
    .B1(_06450_));
 sg13g2_a22oi_1 _23019_ (.Y(_06451_),
    .B1(_06294_),
    .B2(\top_ihp.oisc.regs[55][20] ),
    .A2(_05788_),
    .A1(\top_ihp.oisc.regs[43][20] ));
 sg13g2_a22oi_1 _23020_ (.Y(_06452_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][20] ),
    .A2(net173),
    .A1(\top_ihp.oisc.regs[53][20] ));
 sg13g2_a22oi_1 _23021_ (.Y(_06453_),
    .B1(_06287_),
    .B2(\top_ihp.oisc.regs[42][20] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][20] ));
 sg13g2_a22oi_1 _23022_ (.Y(_06454_),
    .B1(net186),
    .B2(\top_ihp.oisc.regs[33][20] ),
    .A2(net329),
    .A1(\top_ihp.oisc.regs[50][20] ));
 sg13g2_nand4_1 _23023_ (.B(_06452_),
    .C(_06453_),
    .A(_06451_),
    .Y(_06455_),
    .D(_06454_));
 sg13g2_a22oi_1 _23024_ (.Y(_06456_),
    .B1(_05968_),
    .B2(\top_ihp.oisc.regs[40][20] ),
    .A2(_05767_),
    .A1(\top_ihp.oisc.regs[44][20] ));
 sg13g2_a22oi_1 _23025_ (.Y(_06457_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][20] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[45][20] ));
 sg13g2_a22oi_1 _23026_ (.Y(_06458_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[63][20] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][20] ));
 sg13g2_a22oi_1 _23027_ (.Y(_06459_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][20] ),
    .A2(net306),
    .A1(\top_ihp.oisc.regs[34][20] ));
 sg13g2_nand4_1 _23028_ (.B(_06457_),
    .C(_06458_),
    .A(_06456_),
    .Y(_06460_),
    .D(_06459_));
 sg13g2_a22oi_1 _23029_ (.Y(_06461_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][20] ),
    .A2(net69),
    .A1(\top_ihp.oisc.regs[39][20] ));
 sg13g2_a22oi_1 _23030_ (.Y(_06462_),
    .B1(_05782_),
    .B2(\top_ihp.oisc.regs[35][20] ),
    .A2(net310),
    .A1(\top_ihp.oisc.regs[48][20] ));
 sg13g2_nand2_1 _23031_ (.Y(_06463_),
    .A(\top_ihp.oisc.regs[46][20] ),
    .B(_06383_));
 sg13g2_a22oi_1 _23032_ (.Y(_06464_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][20] ),
    .A2(net304),
    .A1(\top_ihp.oisc.regs[58][20] ));
 sg13g2_nand4_1 _23033_ (.B(_06462_),
    .C(_06463_),
    .A(_06461_),
    .Y(_06465_),
    .D(_06464_));
 sg13g2_nor4_1 _23034_ (.A(net190),
    .B(_06455_),
    .C(_06460_),
    .D(_06465_),
    .Y(_06466_));
 sg13g2_nand2_1 _23035_ (.Y(_06467_),
    .A(\top_ihp.oisc.regs[56][20] ),
    .B(net309));
 sg13g2_a22oi_1 _23036_ (.Y(_06468_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][20] ),
    .A2(net720),
    .A1(_08228_));
 sg13g2_a22oi_1 _23037_ (.Y(_06469_),
    .B1(net605),
    .B2(\top_ihp.oisc.regs[27][20] ),
    .A2(net451),
    .A1(\top_ihp.oisc.regs[7][20] ));
 sg13g2_a22oi_1 _23038_ (.Y(_06470_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][20] ),
    .A2(net332),
    .A1(\top_ihp.oisc.regs[3][20] ));
 sg13g2_nand4_1 _23039_ (.B(_06468_),
    .C(_06469_),
    .A(_06467_),
    .Y(_06471_),
    .D(_06470_));
 sg13g2_a22oi_1 _23040_ (.Y(_06472_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][20] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][20] ));
 sg13g2_a22oi_1 _23041_ (.Y(_06473_),
    .B1(_05504_),
    .B2(\top_ihp.oisc.regs[31][20] ),
    .A2(net175),
    .A1(\top_ihp.oisc.regs[13][20] ));
 sg13g2_mux2_1 _23042_ (.A0(\top_ihp.oisc.regs[29][20] ),
    .A1(\top_ihp.oisc.regs[25][20] ),
    .S(net598),
    .X(_06474_));
 sg13g2_nor2_1 _23043_ (.A(net681),
    .B(_05509_),
    .Y(_06475_));
 sg13g2_nand2_1 _23044_ (.Y(_06476_),
    .A(\top_ihp.oisc.regs[10][20] ),
    .B(net416));
 sg13g2_nand2_1 _23045_ (.Y(_06477_),
    .A(\top_ihp.oisc.regs[11][20] ),
    .B(net594));
 sg13g2_nand2_1 _23046_ (.Y(_06478_),
    .A(net607),
    .B(_05995_));
 sg13g2_a21oi_1 _23047_ (.A1(_06476_),
    .A2(_06477_),
    .Y(_06479_),
    .B1(_06478_));
 sg13g2_a21oi_1 _23048_ (.A1(_06474_),
    .A2(_06475_),
    .Y(_06480_),
    .B1(_06479_));
 sg13g2_nor2_1 _23049_ (.A(net676),
    .B(_05379_),
    .Y(_06481_));
 sg13g2_and3_1 _23050_ (.X(_06482_),
    .A(\top_ihp.oisc.regs[4][20] ),
    .B(_05847_),
    .C(_06481_));
 sg13g2_a221oi_1 _23051_ (.B2(\top_ihp.oisc.regs[1][20] ),
    .C1(_06482_),
    .B1(_05489_),
    .A1(\top_ihp.oisc.regs[19][20] ),
    .Y(_06483_),
    .A2(net445));
 sg13g2_nand4_1 _23052_ (.B(_06473_),
    .C(_06480_),
    .A(_06472_),
    .Y(_06484_),
    .D(_06483_));
 sg13g2_a22oi_1 _23053_ (.Y(_06485_),
    .B1(_06047_),
    .B2(\top_ihp.oisc.regs[49][20] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][20] ));
 sg13g2_a22oi_1 _23054_ (.Y(_06486_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][20] ),
    .A2(_05310_),
    .A1(\top_ihp.oisc.regs[60][20] ));
 sg13g2_a22oi_1 _23055_ (.Y(_06487_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][20] ),
    .A2(_05665_),
    .A1(\top_ihp.oisc.regs[54][20] ));
 sg13g2_a22oi_1 _23056_ (.Y(_06488_),
    .B1(net78),
    .B2(\top_ihp.oisc.regs[59][20] ),
    .A2(_05466_),
    .A1(\top_ihp.oisc.regs[62][20] ));
 sg13g2_nand4_1 _23057_ (.B(_06486_),
    .C(_06487_),
    .A(_06485_),
    .Y(_06489_),
    .D(_06488_));
 sg13g2_and2_1 _23058_ (.A(\top_ihp.oisc.regs[21][20] ),
    .B(net742),
    .X(_06490_));
 sg13g2_nor2_2 _23059_ (.A(net610),
    .B(_05426_),
    .Y(_06491_));
 sg13g2_a22oi_1 _23060_ (.Y(_06492_),
    .B1(_06490_),
    .B2(_06491_),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[8][20] ));
 sg13g2_a22oi_1 _23061_ (.Y(_06493_),
    .B1(_05828_),
    .B2(\top_ihp.oisc.regs[2][20] ),
    .A2(_05493_),
    .A1(\top_ihp.oisc.regs[26][20] ));
 sg13g2_mux2_1 _23062_ (.A0(\top_ihp.oisc.regs[14][20] ),
    .A1(\top_ihp.oisc.regs[6][20] ),
    .S(net681),
    .X(_06494_));
 sg13g2_nor2_1 _23063_ (.A(net594),
    .B(_05375_),
    .Y(_06495_));
 sg13g2_a22oi_1 _23064_ (.Y(_06496_),
    .B1(_06494_),
    .B2(_06495_),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][20] ));
 sg13g2_a22oi_1 _23065_ (.Y(_06497_),
    .B1(_05422_),
    .B2(\top_ihp.oisc.regs[18][20] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][20] ));
 sg13g2_and4_1 _23066_ (.A(_06492_),
    .B(_06493_),
    .C(_06496_),
    .D(_06497_),
    .X(_06498_));
 sg13g2_nand3_1 _23067_ (.B(net320),
    .C(net694),
    .A(\top_ihp.oisc.regs[23][20] ),
    .Y(_06499_));
 sg13g2_nand3_1 _23068_ (.B(net412),
    .C(net673),
    .A(\top_ihp.oisc.regs[16][20] ),
    .Y(_06500_));
 sg13g2_a21o_1 _23069_ (.A2(_06500_),
    .A1(_06499_),
    .B1(net415),
    .X(_06501_));
 sg13g2_a22oi_1 _23070_ (.Y(_06502_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][20] ),
    .A2(_05727_),
    .A1(\top_ihp.oisc.regs[12][20] ));
 sg13g2_a22oi_1 _23071_ (.Y(_06503_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][20] ),
    .A2(_05821_),
    .A1(\top_ihp.oisc.regs[28][20] ));
 sg13g2_nand4_1 _23072_ (.B(_06501_),
    .C(_06502_),
    .A(_06498_),
    .Y(_06504_),
    .D(_06503_));
 sg13g2_nor4_1 _23073_ (.A(_06471_),
    .B(_06484_),
    .C(_06489_),
    .D(_06504_),
    .Y(_06505_));
 sg13g2_buf_8 _23074_ (.A(net331),
    .X(_06506_));
 sg13g2_a21oi_1 _23075_ (.A1(_00261_),
    .A2(net150),
    .Y(_06507_),
    .B1(net34));
 sg13g2_a21oi_1 _23076_ (.A1(_08228_),
    .A2(net693),
    .Y(_06508_),
    .B1(_06507_));
 sg13g2_a21oi_1 _23077_ (.A1(_06466_),
    .A2(_06505_),
    .Y(_00432_),
    .B1(_06508_));
 sg13g2_nand2_1 _23078_ (.Y(_06509_),
    .A(\top_ihp.oisc.regs[51][21] ),
    .B(_05642_));
 sg13g2_a22oi_1 _23079_ (.Y(_06510_),
    .B1(_06114_),
    .B2(\top_ihp.oisc.regs[8][21] ),
    .A2(net154),
    .A1(\top_ihp.oisc.regs[47][21] ));
 sg13g2_nand2_1 _23080_ (.Y(_06511_),
    .A(_06509_),
    .B(_06510_));
 sg13g2_a22oi_1 _23081_ (.Y(_06512_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][21] ),
    .A2(_05539_),
    .A1(\top_ihp.oisc.regs[55][21] ));
 sg13g2_a22oi_1 _23082_ (.Y(_06513_),
    .B1(_05478_),
    .B2(\top_ihp.oisc.regs[43][21] ),
    .A2(_05465_),
    .A1(\top_ihp.oisc.regs[62][21] ));
 sg13g2_a22oi_1 _23083_ (.Y(_06514_),
    .B1(_05484_),
    .B2(\top_ihp.oisc.regs[42][21] ),
    .A2(_05337_),
    .A1(\top_ihp.oisc.regs[38][21] ));
 sg13g2_a22oi_1 _23084_ (.Y(_06515_),
    .B1(net435),
    .B2(\top_ihp.oisc.regs[40][21] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][21] ));
 sg13g2_and4_1 _23085_ (.A(_06512_),
    .B(_06513_),
    .C(_06514_),
    .D(_06515_),
    .X(_06516_));
 sg13g2_a22oi_1 _23086_ (.Y(_06517_),
    .B1(_05776_),
    .B2(\top_ihp.oisc.regs[57][21] ),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][21] ));
 sg13g2_nor4_2 _23087_ (.A(net613),
    .B(net678),
    .C(net671),
    .Y(_06518_),
    .D(_05335_));
 sg13g2_a22oi_1 _23088_ (.Y(_06519_),
    .B1(_06518_),
    .B2(\top_ihp.oisc.regs[52][21] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][21] ));
 sg13g2_a22oi_1 _23089_ (.Y(_06520_),
    .B1(_05900_),
    .B2(\top_ihp.oisc.regs[18][21] ),
    .A2(net696),
    .A1(\top_ihp.oisc.regs[30][21] ));
 sg13g2_nand2_1 _23090_ (.Y(_06521_),
    .A(\top_ihp.oisc.regs[50][21] ),
    .B(_05523_));
 sg13g2_o21ai_1 _23091_ (.B1(_06521_),
    .Y(_06522_),
    .A1(_05419_),
    .A2(_06520_));
 sg13g2_a221oi_1 _23092_ (.B2(\top_ihp.oisc.regs[56][21] ),
    .C1(_06522_),
    .B1(_05605_),
    .A1(\top_ihp.oisc.regs[35][21] ),
    .Y(_06523_),
    .A2(net433));
 sg13g2_nand4_1 _23093_ (.B(_06517_),
    .C(_06519_),
    .A(_06516_),
    .Y(_06524_),
    .D(_06523_));
 sg13g2_a22oi_1 _23094_ (.Y(_06525_),
    .B1(net302),
    .B2(\top_ihp.oisc.regs[32][21] ),
    .A2(_05311_),
    .A1(\top_ihp.oisc.regs[60][21] ));
 sg13g2_a22oi_1 _23095_ (.Y(_06526_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[33][21] ),
    .A2(_05661_),
    .A1(\top_ihp.oisc.regs[45][21] ));
 sg13g2_a22oi_1 _23096_ (.Y(_06527_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][21] ),
    .A2(_05762_),
    .A1(\top_ihp.oisc.regs[58][21] ));
 sg13g2_a22oi_1 _23097_ (.Y(_06528_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][21] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[63][21] ));
 sg13g2_nand4_1 _23098_ (.B(_06526_),
    .C(_06527_),
    .A(_06525_),
    .Y(_06529_),
    .D(_06528_));
 sg13g2_nor4_2 _23099_ (.A(net190),
    .B(_06511_),
    .C(_06524_),
    .Y(_06530_),
    .D(_06529_));
 sg13g2_a22oi_1 _23100_ (.Y(_06531_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][21] ),
    .A2(_05397_),
    .A1(\top_ihp.oisc.regs[12][21] ));
 sg13g2_a22oi_1 _23101_ (.Y(_06532_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][21] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[28][21] ));
 sg13g2_a22oi_1 _23102_ (.Y(_06533_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][21] ),
    .A2(_05327_),
    .A1(\top_ihp.oisc.regs[44][21] ));
 sg13g2_a22oi_1 _23103_ (.Y(_06534_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[25][21] ),
    .A2(net449),
    .A1(\top_ihp.oisc.regs[20][21] ));
 sg13g2_a22oi_1 _23104_ (.Y(_06535_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[15][21] ),
    .A2(_05685_),
    .A1(\top_ihp.oisc.regs[17][21] ));
 sg13g2_and2_1 _23105_ (.A(_06534_),
    .B(_06535_),
    .X(_06536_));
 sg13g2_nand4_1 _23106_ (.B(_06532_),
    .C(_06533_),
    .A(_06531_),
    .Y(_06537_),
    .D(_06536_));
 sg13g2_mux2_1 _23107_ (.A0(\top_ihp.oisc.regs[31][21] ),
    .A1(\top_ihp.oisc.regs[23][21] ),
    .S(_05696_),
    .X(_06538_));
 sg13g2_a22oi_1 _23108_ (.Y(_06539_),
    .B1(_06538_),
    .B2(_06215_),
    .A2(_05778_),
    .A1(\top_ihp.oisc.regs[54][21] ));
 sg13g2_a22oi_1 _23109_ (.Y(_06540_),
    .B1(net294),
    .B2(\top_ihp.oisc.regs[4][21] ),
    .A2(net332),
    .A1(\top_ihp.oisc.regs[3][21] ));
 sg13g2_nand2_1 _23110_ (.Y(_06541_),
    .A(\top_ihp.oisc.regs[13][21] ),
    .B(_05402_));
 sg13g2_nand4_1 _23111_ (.B(net594),
    .C(_05442_),
    .A(\top_ihp.oisc.regs[59][21] ),
    .Y(_06542_),
    .D(_06154_));
 sg13g2_nand2_1 _23112_ (.Y(_06543_),
    .A(_06541_),
    .B(_06542_));
 sg13g2_a221oi_1 _23113_ (.B2(\top_ihp.oisc.regs[21][21] ),
    .C1(_06543_),
    .B1(net444),
    .A1(\top_ihp.oisc.regs[27][21] ),
    .Y(_06544_),
    .A2(net603));
 sg13g2_a22oi_1 _23114_ (.Y(_06545_),
    .B1(net306),
    .B2(\top_ihp.oisc.regs[34][21] ),
    .A2(net155),
    .A1(\top_ihp.oisc.regs[39][21] ));
 sg13g2_nand4_1 _23115_ (.B(_06540_),
    .C(_06544_),
    .A(_06539_),
    .Y(_06546_),
    .D(_06545_));
 sg13g2_nand2_1 _23116_ (.Y(_06547_),
    .A(\top_ihp.oisc.regs[61][21] ),
    .B(net67));
 sg13g2_a22oi_1 _23117_ (.Y(_06548_),
    .B1(_05723_),
    .B2(\top_ihp.oisc.regs[9][21] ),
    .A2(net728),
    .A1(_08235_));
 sg13g2_a22oi_1 _23118_ (.Y(_06549_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[14][21] ),
    .A2(_05809_),
    .A1(\top_ihp.oisc.regs[5][21] ));
 sg13g2_a22oi_1 _23119_ (.Y(_06550_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[19][21] ),
    .A2(_05712_),
    .A1(\top_ihp.oisc.regs[16][21] ));
 sg13g2_nand4_1 _23120_ (.B(_06548_),
    .C(_06549_),
    .A(_06547_),
    .Y(_06551_),
    .D(_06550_));
 sg13g2_and4_1 _23121_ (.A(\top_ihp.oisc.regs[1][21] ),
    .B(_05609_),
    .C(net290),
    .D(_06014_),
    .X(_06552_));
 sg13g2_a21oi_1 _23122_ (.A1(\top_ihp.oisc.regs[7][21] ),
    .A2(_06256_),
    .Y(_06553_),
    .B1(_06552_));
 sg13g2_a22oi_1 _23123_ (.Y(_06554_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][21] ),
    .A2(net333),
    .A1(\top_ihp.oisc.regs[26][21] ));
 sg13g2_a22oi_1 _23124_ (.Y(_06555_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][21] ),
    .A2(net425),
    .A1(\top_ihp.oisc.regs[29][21] ));
 sg13g2_a22oi_1 _23125_ (.Y(_06556_),
    .B1(_05829_),
    .B2(\top_ihp.oisc.regs[2][21] ),
    .A2(_05876_),
    .A1(\top_ihp.oisc.regs[6][21] ));
 sg13g2_nand4_1 _23126_ (.B(_06554_),
    .C(_06555_),
    .A(_06553_),
    .Y(_06557_),
    .D(_06556_));
 sg13g2_nor4_1 _23127_ (.A(_06537_),
    .B(_06546_),
    .C(_06551_),
    .D(_06557_),
    .Y(_06558_));
 sg13g2_buf_1 _23128_ (.A(_05622_),
    .X(_06559_));
 sg13g2_a21oi_1 _23129_ (.A1(_00262_),
    .A2(net150),
    .Y(_06560_),
    .B1(net32));
 sg13g2_a21oi_1 _23130_ (.A1(_08235_),
    .A2(net693),
    .Y(_06561_),
    .B1(_06560_));
 sg13g2_a21oi_1 _23131_ (.A1(_06530_),
    .A2(_06558_),
    .Y(_00433_),
    .B1(_06561_));
 sg13g2_and2_1 _23132_ (.A(\top_ihp.oisc.regs[54][22] ),
    .B(net179),
    .X(_06562_));
 sg13g2_a221oi_1 _23133_ (.B2(\top_ihp.oisc.regs[52][22] ),
    .C1(_06562_),
    .B1(net311),
    .A1(\top_ihp.oisc.regs[36][22] ),
    .Y(_06563_),
    .A2(net156));
 sg13g2_a22oi_1 _23134_ (.Y(_06564_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][22] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][22] ));
 sg13g2_a22oi_1 _23135_ (.Y(_06565_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[47][22] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][22] ));
 sg13g2_a22oi_1 _23136_ (.Y(_06566_),
    .B1(net77),
    .B2(\top_ihp.oisc.regs[55][22] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][22] ));
 sg13g2_a22oi_1 _23137_ (.Y(_06567_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][22] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[58][22] ));
 sg13g2_nand4_1 _23138_ (.B(_06565_),
    .C(_06566_),
    .A(_06564_),
    .Y(_06568_),
    .D(_06567_));
 sg13g2_nand2_1 _23139_ (.Y(_06569_),
    .A(\top_ihp.oisc.regs[10][22] ),
    .B(_05728_));
 sg13g2_a22oi_1 _23140_ (.Y(_06570_),
    .B1(_05733_),
    .B2(\top_ihp.oisc.regs[14][22] ),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][22] ));
 sg13g2_a22oi_1 _23141_ (.Y(_06571_),
    .B1(_05817_),
    .B2(\top_ihp.oisc.regs[30][22] ),
    .A2(_05421_),
    .A1(\top_ihp.oisc.regs[18][22] ));
 sg13g2_a22oi_1 _23142_ (.Y(_06572_),
    .B1(_05493_),
    .B2(\top_ihp.oisc.regs[26][22] ),
    .A2(_05387_),
    .A1(\top_ihp.oisc.regs[6][22] ));
 sg13g2_nand4_1 _23143_ (.B(_06570_),
    .C(_06571_),
    .A(_06569_),
    .Y(_06573_),
    .D(_06572_));
 sg13g2_a22oi_1 _23144_ (.Y(_06574_),
    .B1(_05444_),
    .B2(\top_ihp.oisc.regs[27][22] ),
    .A2(_05402_),
    .A1(\top_ihp.oisc.regs[13][22] ));
 sg13g2_a22oi_1 _23145_ (.Y(_06575_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[15][22] ),
    .A2(_05450_),
    .A1(\top_ihp.oisc.regs[21][22] ));
 sg13g2_a22oi_1 _23146_ (.Y(_06576_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][22] ),
    .A2(_05455_),
    .A1(\top_ihp.oisc.regs[28][22] ));
 sg13g2_a22oi_1 _23147_ (.Y(_06577_),
    .B1(net611),
    .B2(\top_ihp.oisc.regs[31][22] ),
    .A2(_05395_),
    .A1(\top_ihp.oisc.regs[8][22] ));
 sg13g2_nand4_1 _23148_ (.B(_06575_),
    .C(_06576_),
    .A(_06574_),
    .Y(_06578_),
    .D(_06577_));
 sg13g2_mux2_1 _23149_ (.A0(\top_ihp.oisc.regs[3][22] ),
    .A1(\top_ihp.oisc.regs[2][22] ),
    .S(_05360_),
    .X(_06579_));
 sg13g2_a22oi_1 _23150_ (.Y(_06580_),
    .B1(_06579_),
    .B2(net595),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[11][22] ));
 sg13g2_nor2_1 _23151_ (.A(_05409_),
    .B(_06580_),
    .Y(_06581_));
 sg13g2_a22oi_1 _23152_ (.Y(_06582_),
    .B1(_05685_),
    .B2(\top_ihp.oisc.regs[17][22] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][22] ));
 sg13g2_a22oi_1 _23153_ (.Y(_06583_),
    .B1(_05725_),
    .B2(\top_ihp.oisc.regs[29][22] ),
    .A2(_05396_),
    .A1(\top_ihp.oisc.regs[12][22] ));
 sg13g2_a22oi_1 _23154_ (.Y(_06584_),
    .B1(_05436_),
    .B2(\top_ihp.oisc.regs[19][22] ),
    .A2(_05384_),
    .A1(\top_ihp.oisc.regs[7][22] ));
 sg13g2_a22oi_1 _23155_ (.Y(_06585_),
    .B1(_05507_),
    .B2(\top_ihp.oisc.regs[4][22] ),
    .A2(_05357_),
    .A1(\top_ihp.oisc.regs[16][22] ));
 sg13g2_nand4_1 _23156_ (.B(_06583_),
    .C(_06584_),
    .A(_06582_),
    .Y(_06586_),
    .D(_06585_));
 sg13g2_or4_2 _23157_ (.A(_06573_),
    .B(_06578_),
    .C(_06581_),
    .D(_06586_),
    .X(_06587_));
 sg13g2_a22oi_1 _23158_ (.Y(_06588_),
    .B1(_05593_),
    .B2(\top_ihp.oisc.regs[53][22] ),
    .A2(_05478_),
    .A1(\top_ihp.oisc.regs[43][22] ));
 sg13g2_a22oi_1 _23159_ (.Y(_06589_),
    .B1(_05605_),
    .B2(\top_ihp.oisc.regs[56][22] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[59][22] ));
 sg13g2_a22oi_1 _23160_ (.Y(_06590_),
    .B1(net324),
    .B2(\top_ihp.oisc.regs[63][22] ),
    .A2(_05523_),
    .A1(\top_ihp.oisc.regs[50][22] ));
 sg13g2_a22oi_1 _23161_ (.Y(_06591_),
    .B1(_05429_),
    .B2(\top_ihp.oisc.regs[32][22] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[44][22] ));
 sg13g2_nand4_1 _23162_ (.B(_06589_),
    .C(_06590_),
    .A(_06588_),
    .Y(_06592_),
    .D(_06591_));
 sg13g2_a22oi_1 _23163_ (.Y(_06593_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[49][22] ),
    .A2(_05465_),
    .A1(\top_ihp.oisc.regs[62][22] ));
 sg13g2_a22oi_1 _23164_ (.Y(_06594_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][22] ),
    .A2(net609),
    .A1(\top_ihp.oisc.regs[57][22] ));
 sg13g2_a22oi_1 _23165_ (.Y(_06595_),
    .B1(_05603_),
    .B2(\top_ihp.oisc.regs[46][22] ),
    .A2(_05484_),
    .A1(\top_ihp.oisc.regs[42][22] ));
 sg13g2_a22oi_1 _23166_ (.Y(_06596_),
    .B1(_05525_),
    .B2(\top_ihp.oisc.regs[45][22] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[40][22] ));
 sg13g2_nand4_1 _23167_ (.B(_06594_),
    .C(_06595_),
    .A(_06593_),
    .Y(_06597_),
    .D(_06596_));
 sg13g2_or2_1 _23168_ (.X(_06598_),
    .B(_06597_),
    .A(_06592_));
 sg13g2_a22oi_1 _23169_ (.Y(_06599_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[25][22] ),
    .A2(_05495_),
    .A1(\top_ihp.oisc.regs[23][22] ));
 sg13g2_nand3_1 _23170_ (.B(_06017_),
    .C(_06317_),
    .A(\top_ihp.oisc.regs[1][22] ),
    .Y(_06600_));
 sg13g2_nand2_2 _23171_ (.Y(_06601_),
    .A(_08391_),
    .B(net748));
 sg13g2_nand3_1 _23172_ (.B(net421),
    .C(_06056_),
    .A(\top_ihp.oisc.regs[22][22] ),
    .Y(_06602_));
 sg13g2_nand4_1 _23173_ (.B(_06600_),
    .C(_06601_),
    .A(_06599_),
    .Y(_06603_),
    .D(_06602_));
 sg13g2_a221oi_1 _23174_ (.B2(\top_ihp.oisc.regs[33][22] ),
    .C1(_06603_),
    .B1(_05633_),
    .A1(\top_ihp.oisc.regs[20][22] ),
    .Y(_06604_),
    .A2(net293));
 sg13g2_a22oi_1 _23175_ (.Y(_06605_),
    .B1(net174),
    .B2(\top_ihp.oisc.regs[39][22] ),
    .A2(net310),
    .A1(\top_ihp.oisc.regs[48][22] ));
 sg13g2_a22oi_1 _23176_ (.Y(_06606_),
    .B1(net307),
    .B2(\top_ihp.oisc.regs[34][22] ),
    .A2(net325),
    .A1(\top_ihp.oisc.regs[35][22] ));
 sg13g2_nand4_1 _23177_ (.B(_06604_),
    .C(_06605_),
    .A(_05918_),
    .Y(_06607_),
    .D(_06606_));
 sg13g2_nor4_1 _23178_ (.A(_06568_),
    .B(_06587_),
    .C(_06598_),
    .D(_06607_),
    .Y(_06608_));
 sg13g2_a21o_1 _23179_ (.A2(net159),
    .A1(_00263_),
    .B1(net33),
    .X(_06609_));
 sg13g2_a22oi_1 _23180_ (.Y(_00434_),
    .B1(_06609_),
    .B2(_06601_),
    .A2(_06608_),
    .A1(_06563_));
 sg13g2_a22oi_1 _23181_ (.Y(_06610_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][23] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][23] ));
 sg13g2_a22oi_1 _23182_ (.Y(_06611_),
    .B1(net600),
    .B2(\top_ihp.oisc.regs[12][23] ),
    .A2(net670),
    .A1(\top_ihp.oisc.regs[14][23] ));
 sg13g2_inv_1 _23183_ (.Y(_06612_),
    .A(_06611_));
 sg13g2_a22oi_1 _23184_ (.Y(_06613_),
    .B1(_05900_),
    .B2(\top_ihp.oisc.regs[17][23] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[21][23] ));
 sg13g2_nor2_1 _23185_ (.A(net734),
    .B(_06613_),
    .Y(_06614_));
 sg13g2_a221oi_1 _23186_ (.B2(_06612_),
    .C1(_06614_),
    .B1(net410),
    .A1(net1047),
    .Y(_06615_),
    .A2(net720));
 sg13g2_a22oi_1 _23187_ (.Y(_06616_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][23] ),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[1][23] ));
 sg13g2_a22oi_1 _23188_ (.Y(_06617_),
    .B1(net185),
    .B2(\top_ihp.oisc.regs[59][23] ),
    .A2(_05553_),
    .A1(\top_ihp.oisc.regs[39][23] ));
 sg13g2_a22oi_1 _23189_ (.Y(_06618_),
    .B1(_05588_),
    .B2(\top_ihp.oisc.regs[47][23] ),
    .A2(_05471_),
    .A1(\top_ihp.oisc.regs[37][23] ));
 sg13g2_and2_1 _23190_ (.A(_06617_),
    .B(_06618_),
    .X(_06619_));
 sg13g2_nand4_1 _23191_ (.B(_06615_),
    .C(_06616_),
    .A(_06610_),
    .Y(_06620_),
    .D(_06619_));
 sg13g2_nand2_1 _23192_ (.Y(_06621_),
    .A(\top_ihp.oisc.regs[5][23] ),
    .B(_05809_));
 sg13g2_a22oi_1 _23193_ (.Y(_06622_),
    .B1(net151),
    .B2(\top_ihp.oisc.regs[3][23] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[27][23] ));
 sg13g2_nand2_1 _23194_ (.Y(_06623_),
    .A(_06621_),
    .B(_06622_));
 sg13g2_a22oi_1 _23195_ (.Y(_06624_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[31][23] ),
    .A2(net283),
    .A1(\top_ihp.oisc.regs[23][23] ));
 sg13g2_nand3_1 _23196_ (.B(net291),
    .C(net697),
    .A(\top_ihp.oisc.regs[29][23] ),
    .Y(_06625_));
 sg13g2_nand3_1 _23197_ (.B(net598),
    .C(net695),
    .A(\top_ihp.oisc.regs[26][23] ),
    .Y(_06626_));
 sg13g2_nand2_1 _23198_ (.Y(_06627_),
    .A(_06625_),
    .B(_06626_));
 sg13g2_a22oi_1 _23199_ (.Y(_06628_),
    .B1(_06627_),
    .B2(net415),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][23] ));
 sg13g2_a22oi_1 _23200_ (.Y(_06629_),
    .B1(net294),
    .B2(\top_ihp.oisc.regs[4][23] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[19][23] ));
 sg13g2_a22oi_1 _23201_ (.Y(_06630_),
    .B1(net164),
    .B2(\top_ihp.oisc.regs[30][23] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][23] ));
 sg13g2_nand4_1 _23202_ (.B(_06628_),
    .C(_06629_),
    .A(_06624_),
    .Y(_06631_),
    .D(_06630_));
 sg13g2_a22oi_1 _23203_ (.Y(_06632_),
    .B1(_06158_),
    .B2(\top_ihp.oisc.regs[24][23] ),
    .A2(_05821_),
    .A1(\top_ihp.oisc.regs[28][23] ));
 sg13g2_nand2_1 _23204_ (.Y(_06633_),
    .A(\top_ihp.oisc.regs[22][23] ),
    .B(net152));
 sg13g2_a22oi_1 _23205_ (.Y(_06634_),
    .B1(_05422_),
    .B2(\top_ihp.oisc.regs[18][23] ),
    .A2(net411),
    .A1(\top_ihp.oisc.regs[8][23] ));
 sg13g2_a22oi_1 _23206_ (.Y(_06635_),
    .B1(_05403_),
    .B2(\top_ihp.oisc.regs[13][23] ),
    .A2(net449),
    .A1(\top_ihp.oisc.regs[20][23] ));
 sg13g2_a22oi_1 _23207_ (.Y(_06636_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[10][23] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[11][23] ));
 sg13g2_a22oi_1 _23208_ (.Y(_06637_),
    .B1(_05828_),
    .B2(\top_ihp.oisc.regs[2][23] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[9][23] ));
 sg13g2_and4_1 _23209_ (.A(_06634_),
    .B(_06635_),
    .C(_06636_),
    .D(_06637_),
    .X(_06638_));
 sg13g2_nand3_1 _23210_ (.B(_06633_),
    .C(_06638_),
    .A(_06632_),
    .Y(_06639_));
 sg13g2_nor4_1 _23211_ (.A(_06620_),
    .B(_06623_),
    .C(_06631_),
    .D(_06639_),
    .Y(_06640_));
 sg13g2_a22oi_1 _23212_ (.Y(_06641_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[42][23] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][23] ));
 sg13g2_a22oi_1 _23213_ (.Y(_06642_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[49][23] ),
    .A2(net302),
    .A1(\top_ihp.oisc.regs[32][23] ));
 sg13g2_a22oi_1 _23214_ (.Y(_06643_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][23] ),
    .A2(net310),
    .A1(\top_ihp.oisc.regs[48][23] ));
 sg13g2_a22oi_1 _23215_ (.Y(_06644_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][23] ),
    .A2(_05630_),
    .A1(\top_ihp.oisc.regs[61][23] ));
 sg13g2_nand4_1 _23216_ (.B(_06642_),
    .C(_06643_),
    .A(_06641_),
    .Y(_06645_),
    .D(_06644_));
 sg13g2_a22oi_1 _23217_ (.Y(_06646_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][23] ),
    .A2(net68),
    .A1(\top_ihp.oisc.regs[55][23] ));
 sg13g2_a22oi_1 _23218_ (.Y(_06647_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][23] ),
    .A2(_05776_),
    .A1(\top_ihp.oisc.regs[57][23] ));
 sg13g2_a22oi_1 _23219_ (.Y(_06648_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][23] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][23] ));
 sg13g2_a22oi_1 _23220_ (.Y(_06649_),
    .B1(net70),
    .B2(\top_ihp.oisc.regs[45][23] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][23] ));
 sg13g2_nand4_1 _23221_ (.B(_06647_),
    .C(_06648_),
    .A(_06646_),
    .Y(_06650_),
    .D(_06649_));
 sg13g2_o21ai_1 _23222_ (.B1(\top_ihp.oisc.regs[16][23] ),
    .Y(_06651_),
    .A1(net948),
    .A2(_05296_));
 sg13g2_nor2_1 _23223_ (.A(_05568_),
    .B(_06651_),
    .Y(_06652_));
 sg13g2_a22oi_1 _23224_ (.Y(_06653_),
    .B1(_06652_),
    .B2(_06260_),
    .A2(_06475_),
    .A1(\top_ihp.oisc.regs[25][23] ));
 sg13g2_nor2_2 _23225_ (.A(_05681_),
    .B(_06653_),
    .Y(_06654_));
 sg13g2_a221oi_1 _23226_ (.B2(\top_ihp.oisc.regs[41][23] ),
    .C1(_06654_),
    .B1(net323),
    .A1(\top_ihp.oisc.regs[56][23] ),
    .Y(_06655_),
    .A2(net301));
 sg13g2_a22oi_1 _23227_ (.Y(_06656_),
    .B1(net187),
    .B2(\top_ihp.oisc.regs[38][23] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][23] ));
 sg13g2_a22oi_1 _23228_ (.Y(_06657_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[53][23] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[40][23] ));
 sg13g2_a22oi_1 _23229_ (.Y(_06658_),
    .B1(net324),
    .B2(\top_ihp.oisc.regs[63][23] ),
    .A2(_05478_),
    .A1(\top_ihp.oisc.regs[43][23] ));
 sg13g2_a22oi_1 _23230_ (.Y(_06659_),
    .B1(net433),
    .B2(\top_ihp.oisc.regs[35][23] ),
    .A2(_05528_),
    .A1(\top_ihp.oisc.regs[33][23] ));
 sg13g2_and4_1 _23231_ (.A(_06656_),
    .B(_06657_),
    .C(_06658_),
    .D(_06659_),
    .X(_06660_));
 sg13g2_nand3_1 _23232_ (.B(_06655_),
    .C(_06660_),
    .A(_05918_),
    .Y(_06661_));
 sg13g2_nor3_1 _23233_ (.A(_06645_),
    .B(_06650_),
    .C(_06661_),
    .Y(_06662_));
 sg13g2_a21oi_1 _23234_ (.A1(_00069_),
    .A2(net150),
    .Y(_06663_),
    .B1(net32));
 sg13g2_a21oi_1 _23235_ (.A1(_08394_),
    .A2(net693),
    .Y(_06664_),
    .B1(_06663_));
 sg13g2_a21oi_1 _23236_ (.A1(_06640_),
    .A2(_06662_),
    .Y(_00435_),
    .B1(_06664_));
 sg13g2_nand2_1 _23237_ (.Y(_06665_),
    .A(_08380_),
    .B(net739));
 sg13g2_a21o_1 _23238_ (.A2(net158),
    .A1(_00070_),
    .B1(net33),
    .X(_06666_));
 sg13g2_a22oi_1 _23239_ (.Y(_06667_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][24] ),
    .A2(net314),
    .A1(\top_ihp.oisc.regs[9][24] ));
 sg13g2_a22oi_1 _23240_ (.Y(_06668_),
    .B1(net317),
    .B2(\top_ihp.oisc.regs[1][24] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[27][24] ));
 sg13g2_and2_1 _23241_ (.A(\top_ihp.oisc.regs[21][24] ),
    .B(net444),
    .X(_06669_));
 sg13g2_a221oi_1 _23242_ (.B2(\top_ihp.oisc.regs[61][24] ),
    .C1(_06669_),
    .B1(_05831_),
    .A1(\top_ihp.oisc.regs[20][24] ),
    .Y(_06670_),
    .A2(net449));
 sg13g2_a22oi_1 _23243_ (.Y(_06671_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][24] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][24] ));
 sg13g2_nand4_1 _23244_ (.B(_06668_),
    .C(_06670_),
    .A(_06667_),
    .Y(_06672_),
    .D(_06671_));
 sg13g2_a22oi_1 _23245_ (.Y(_06673_),
    .B1(_06143_),
    .B2(\top_ihp.oisc.regs[3][24] ),
    .A2(net600),
    .A1(\top_ihp.oisc.regs[5][24] ));
 sg13g2_o21ai_1 _23246_ (.B1(_06665_),
    .Y(_06674_),
    .A1(_05498_),
    .A2(_06673_));
 sg13g2_a221oi_1 _23247_ (.B2(\top_ihp.oisc.regs[2][24] ),
    .C1(_06674_),
    .B1(net295),
    .A1(\top_ihp.oisc.regs[42][24] ),
    .Y(_06675_),
    .A2(net334));
 sg13g2_and2_1 _23248_ (.A(\top_ihp.oisc.regs[23][24] ),
    .B(net694),
    .X(_06676_));
 sg13g2_and2_1 _23249_ (.A(\top_ihp.oisc.regs[26][24] ),
    .B(net695),
    .X(_06677_));
 sg13g2_a22oi_1 _23250_ (.Y(_06678_),
    .B1(net698),
    .B2(\top_ihp.oisc.regs[31][24] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[30][24] ));
 sg13g2_nor3_1 _23251_ (.A(net412),
    .B(net602),
    .C(_06678_),
    .Y(_06679_));
 sg13g2_a221oi_1 _23252_ (.B2(net699),
    .C1(_06679_),
    .B1(_06677_),
    .A1(net421),
    .Y(_06680_),
    .A2(_06676_));
 sg13g2_a22oi_1 _23253_ (.Y(_06681_),
    .B1(net429),
    .B2(\top_ihp.oisc.regs[8][24] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][24] ));
 sg13g2_nand3_1 _23254_ (.B(_06680_),
    .C(_06681_),
    .A(_06675_),
    .Y(_06682_));
 sg13g2_a22oi_1 _23255_ (.Y(_06683_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][24] ),
    .A2(_05712_),
    .A1(\top_ihp.oisc.regs[16][24] ));
 sg13g2_a22oi_1 _23256_ (.Y(_06684_),
    .B1(net296),
    .B2(\top_ihp.oisc.regs[28][24] ),
    .A2(_05717_),
    .A1(\top_ihp.oisc.regs[18][24] ));
 sg13g2_a22oi_1 _23257_ (.Y(_06685_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][24] ),
    .A2(_05859_),
    .A1(\top_ihp.oisc.regs[4][24] ));
 sg13g2_a22oi_1 _23258_ (.Y(_06686_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][24] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][24] ));
 sg13g2_nand4_1 _23259_ (.B(_06684_),
    .C(_06685_),
    .A(_06683_),
    .Y(_06687_),
    .D(_06686_));
 sg13g2_nor2_2 _23260_ (.A(_05317_),
    .B(net734),
    .Y(_06688_));
 sg13g2_a22oi_1 _23261_ (.Y(_06689_),
    .B1(_06688_),
    .B2(\top_ihp.oisc.regs[29][24] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[19][24] ));
 sg13g2_a22oi_1 _23262_ (.Y(_06690_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][24] ),
    .A2(net315),
    .A1(\top_ihp.oisc.regs[15][24] ));
 sg13g2_nand3_1 _23263_ (.B(net608),
    .C(net596),
    .A(\top_ihp.oisc.regs[10][24] ),
    .Y(_06691_));
 sg13g2_nand3_1 _23264_ (.B(net599),
    .C(net597),
    .A(\top_ihp.oisc.regs[6][24] ),
    .Y(_06692_));
 sg13g2_a21oi_1 _23265_ (.A1(_06691_),
    .A2(_06692_),
    .Y(_06693_),
    .B1(net414));
 sg13g2_a221oi_1 _23266_ (.B2(\top_ihp.oisc.regs[14][24] ),
    .C1(_06693_),
    .B1(net423),
    .A1(\top_ihp.oisc.regs[13][24] ),
    .Y(_06694_),
    .A2(net336));
 sg13g2_nand4_1 _23267_ (.B(_06689_),
    .C(_06690_),
    .A(_05918_),
    .Y(_06695_),
    .D(_06694_));
 sg13g2_nor4_1 _23268_ (.A(_06672_),
    .B(_06682_),
    .C(_06687_),
    .D(_06695_),
    .Y(_06696_));
 sg13g2_a22oi_1 _23269_ (.Y(_06697_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[63][24] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][24] ));
 sg13g2_a22oi_1 _23270_ (.Y(_06698_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][24] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][24] ));
 sg13g2_a22oi_1 _23271_ (.Y(_06699_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][24] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][24] ));
 sg13g2_a22oi_1 _23272_ (.Y(_06700_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[36][24] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][24] ));
 sg13g2_nand4_1 _23273_ (.B(_06698_),
    .C(_06699_),
    .A(_06697_),
    .Y(_06701_),
    .D(_06700_));
 sg13g2_a22oi_1 _23274_ (.Y(_06702_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][24] ),
    .A2(net68),
    .A1(\top_ihp.oisc.regs[55][24] ));
 sg13g2_a22oi_1 _23275_ (.Y(_06703_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][24] ),
    .A2(net70),
    .A1(\top_ihp.oisc.regs[45][24] ));
 sg13g2_nand2_1 _23276_ (.Y(_06704_),
    .A(_06702_),
    .B(_06703_));
 sg13g2_a22oi_1 _23277_ (.Y(_06705_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][24] ),
    .A2(net71),
    .A1(\top_ihp.oisc.regs[59][24] ));
 sg13g2_a22oi_1 _23278_ (.Y(_06706_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][24] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][24] ));
 sg13g2_a22oi_1 _23279_ (.Y(_06707_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][24] ),
    .A2(net422),
    .A1(\top_ihp.oisc.regs[57][24] ));
 sg13g2_nor4_2 _23280_ (.A(net594),
    .B(net678),
    .C(net671),
    .Y(_06708_),
    .D(net679));
 sg13g2_a22oi_1 _23281_ (.Y(_06709_),
    .B1(_06708_),
    .B2(\top_ihp.oisc.regs[56][24] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][24] ));
 sg13g2_nand4_1 _23282_ (.B(_06706_),
    .C(_06707_),
    .A(_06705_),
    .Y(_06710_),
    .D(_06709_));
 sg13g2_a22oi_1 _23283_ (.Y(_06711_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][24] ),
    .A2(net189),
    .A1(\top_ihp.oisc.regs[50][24] ));
 sg13g2_a22oi_1 _23284_ (.Y(_06712_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][24] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][24] ));
 sg13g2_a22oi_1 _23285_ (.Y(_06713_),
    .B1(net288),
    .B2(\top_ihp.oisc.regs[40][24] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][24] ));
 sg13g2_a22oi_1 _23286_ (.Y(_06714_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][24] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[33][24] ));
 sg13g2_nand4_1 _23287_ (.B(_06712_),
    .C(_06713_),
    .A(_06711_),
    .Y(_06715_),
    .D(_06714_));
 sg13g2_nor4_2 _23288_ (.A(_06701_),
    .B(_06704_),
    .C(_06710_),
    .Y(_06716_),
    .D(_06715_));
 sg13g2_a22oi_1 _23289_ (.Y(_00436_),
    .B1(_06696_),
    .B2(_06716_),
    .A2(_06666_),
    .A1(_06665_));
 sg13g2_nand2_1 _23290_ (.Y(_06717_),
    .A(_08384_),
    .B(net739));
 sg13g2_a21o_1 _23291_ (.A2(_05948_),
    .A1(_00071_),
    .B1(net33),
    .X(_06718_));
 sg13g2_nand2_1 _23292_ (.Y(_06719_),
    .A(\top_ihp.oisc.regs[45][25] ),
    .B(net70));
 sg13g2_a22oi_1 _23293_ (.Y(_06720_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][25] ),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][25] ));
 sg13g2_and2_1 _23294_ (.A(\top_ihp.oisc.regs[31][25] ),
    .B(_05503_),
    .X(_06721_));
 sg13g2_a221oi_1 _23295_ (.B2(\top_ihp.oisc.regs[3][25] ),
    .C1(_06721_),
    .B1(net332),
    .A1(\top_ihp.oisc.regs[38][25] ),
    .Y(_06722_),
    .A2(_05632_));
 sg13g2_a22oi_1 _23296_ (.Y(_06723_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][25] ),
    .A2(net609),
    .A1(\top_ihp.oisc.regs[57][25] ));
 sg13g2_nand4_1 _23297_ (.B(_06720_),
    .C(_06722_),
    .A(_06719_),
    .Y(_06724_),
    .D(_06723_));
 sg13g2_a22oi_1 _23298_ (.Y(_06725_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][25] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][25] ));
 sg13g2_a22oi_1 _23299_ (.Y(_06726_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][25] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][25] ));
 sg13g2_a22oi_1 _23300_ (.Y(_06727_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[63][25] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][25] ));
 sg13g2_a22oi_1 _23301_ (.Y(_06728_),
    .B1(net68),
    .B2(\top_ihp.oisc.regs[55][25] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][25] ));
 sg13g2_nand4_1 _23302_ (.B(_06726_),
    .C(_06727_),
    .A(_06725_),
    .Y(_06729_),
    .D(_06728_));
 sg13g2_a22oi_1 _23303_ (.Y(_06730_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][25] ),
    .A2(_06235_),
    .A1(\top_ihp.oisc.regs[39][25] ));
 sg13g2_a22oi_1 _23304_ (.Y(_06731_),
    .B1(_06518_),
    .B2(\top_ihp.oisc.regs[52][25] ),
    .A2(net184),
    .A1(\top_ihp.oisc.regs[51][25] ));
 sg13g2_a22oi_1 _23305_ (.Y(_06732_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[33][25] ),
    .A2(net179),
    .A1(\top_ihp.oisc.regs[54][25] ));
 sg13g2_a22oi_1 _23306_ (.Y(_06733_),
    .B1(_06047_),
    .B2(\top_ihp.oisc.regs[49][25] ),
    .A2(_05739_),
    .A1(\top_ihp.oisc.regs[37][25] ));
 sg13g2_nand4_1 _23307_ (.B(_06731_),
    .C(_06732_),
    .A(_06730_),
    .Y(_06734_),
    .D(_06733_));
 sg13g2_nor4_2 _23308_ (.A(net190),
    .B(_06724_),
    .C(_06729_),
    .Y(_06735_),
    .D(_06734_));
 sg13g2_a22oi_1 _23309_ (.Y(_06736_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][25] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][25] ));
 sg13g2_a22oi_1 _23310_ (.Y(_06737_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][25] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][25] ));
 sg13g2_a22oi_1 _23311_ (.Y(_06738_),
    .B1(net307),
    .B2(\top_ihp.oisc.regs[34][25] ),
    .A2(net433),
    .A1(\top_ihp.oisc.regs[35][25] ));
 sg13g2_a22oi_1 _23312_ (.Y(_06739_),
    .B1(net72),
    .B2(\top_ihp.oisc.regs[53][25] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][25] ));
 sg13g2_nand4_1 _23313_ (.B(_06737_),
    .C(_06738_),
    .A(_06736_),
    .Y(_06740_),
    .D(_06739_));
 sg13g2_a22oi_1 _23314_ (.Y(_06741_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][25] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][25] ));
 sg13g2_nand2_1 _23315_ (.Y(_06742_),
    .A(\top_ihp.oisc.regs[9][25] ),
    .B(net314));
 sg13g2_a22oi_1 _23316_ (.Y(_06743_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][25] ),
    .A2(net444),
    .A1(\top_ihp.oisc.regs[21][25] ));
 sg13g2_a22oi_1 _23317_ (.Y(_06744_),
    .B1(_05493_),
    .B2(\top_ihp.oisc.regs[26][25] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[28][25] ));
 sg13g2_a22oi_1 _23318_ (.Y(_06745_),
    .B1(net443),
    .B2(\top_ihp.oisc.regs[11][25] ),
    .A2(_05390_),
    .A1(\top_ihp.oisc.regs[20][25] ));
 sg13g2_a22oi_1 _23319_ (.Y(_06746_),
    .B1(net411),
    .B2(\top_ihp.oisc.regs[8][25] ),
    .A2(_05388_),
    .A1(\top_ihp.oisc.regs[6][25] ));
 sg13g2_nand3_1 _23320_ (.B(_05404_),
    .C(_05850_),
    .A(\top_ihp.oisc.regs[13][25] ),
    .Y(_06747_));
 sg13g2_nand3_1 _23321_ (.B(net682),
    .C(net670),
    .A(\top_ihp.oisc.regs[14][25] ),
    .Y(_06748_));
 sg13g2_nand2_1 _23322_ (.Y(_06749_),
    .A(_06747_),
    .B(_06748_));
 sg13g2_a22oi_1 _23323_ (.Y(_06750_),
    .B1(_06749_),
    .B2(net608),
    .A2(_05421_),
    .A1(\top_ihp.oisc.regs[18][25] ));
 sg13g2_and4_1 _23324_ (.A(_06744_),
    .B(_06745_),
    .C(_06746_),
    .D(_06750_),
    .X(_06751_));
 sg13g2_nand4_1 _23325_ (.B(_06742_),
    .C(_06743_),
    .A(_06741_),
    .Y(_06752_),
    .D(_06751_));
 sg13g2_a22oi_1 _23326_ (.Y(_06753_),
    .B1(_05710_),
    .B2(\top_ihp.oisc.regs[27][25] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][25] ));
 sg13g2_a22oi_1 _23327_ (.Y(_06754_),
    .B1(net294),
    .B2(\top_ihp.oisc.regs[4][25] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][25] ));
 sg13g2_a22oi_1 _23328_ (.Y(_06755_),
    .B1(_06308_),
    .B2(\top_ihp.oisc.regs[22][25] ),
    .A2(_05705_),
    .A1(\top_ihp.oisc.regs[1][25] ));
 sg13g2_a22oi_1 _23329_ (.Y(_06756_),
    .B1(_06688_),
    .B2(\top_ihp.oisc.regs[29][25] ),
    .A2(net164),
    .A1(\top_ihp.oisc.regs[30][25] ));
 sg13g2_nand4_1 _23330_ (.B(_06754_),
    .C(_06755_),
    .A(_06753_),
    .Y(_06757_),
    .D(_06756_));
 sg13g2_a22oi_1 _23331_ (.Y(_06758_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][25] ),
    .A2(net427),
    .A1(\top_ihp.oisc.regs[19][25] ));
 sg13g2_a22oi_1 _23332_ (.Y(_06759_),
    .B1(_06158_),
    .B2(\top_ihp.oisc.regs[24][25] ),
    .A2(net283),
    .A1(\top_ihp.oisc.regs[23][25] ));
 sg13g2_a22oi_1 _23333_ (.Y(_06760_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][25] ),
    .A2(net315),
    .A1(\top_ihp.oisc.regs[15][25] ));
 sg13g2_a22oi_1 _23334_ (.Y(_06761_),
    .B1(net697),
    .B2(\top_ihp.oisc.regs[17][25] ),
    .A2(net673),
    .A1(\top_ihp.oisc.regs[16][25] ));
 sg13g2_o21ai_1 _23335_ (.B1(_06717_),
    .Y(_06762_),
    .A1(net702),
    .A2(_06761_));
 sg13g2_a21oi_1 _23336_ (.A1(\top_ihp.oisc.regs[5][25] ),
    .A2(net297),
    .Y(_06763_),
    .B1(_06762_));
 sg13g2_nand4_1 _23337_ (.B(_06759_),
    .C(_06760_),
    .A(_06758_),
    .Y(_06764_),
    .D(_06763_));
 sg13g2_nor4_1 _23338_ (.A(_06740_),
    .B(_06752_),
    .C(_06757_),
    .D(_06764_),
    .Y(_06765_));
 sg13g2_a22oi_1 _23339_ (.Y(_00437_),
    .B1(_06735_),
    .B2(_06765_),
    .A2(_06718_),
    .A1(_06717_));
 sg13g2_a22oi_1 _23340_ (.Y(_06766_),
    .B1(_05829_),
    .B2(\top_ihp.oisc.regs[2][26] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][26] ));
 sg13g2_a22oi_1 _23341_ (.Y(_06767_),
    .B1(_05818_),
    .B2(\top_ihp.oisc.regs[30][26] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][26] ));
 sg13g2_nand2_1 _23342_ (.Y(_06768_),
    .A(\top_ihp.oisc.regs[10][26] ),
    .B(net416));
 sg13g2_nand2_1 _23343_ (.Y(_06769_),
    .A(\top_ihp.oisc.regs[11][26] ),
    .B(net594));
 sg13g2_a21oi_1 _23344_ (.A1(_06768_),
    .A2(_06769_),
    .Y(_06770_),
    .B1(_06478_));
 sg13g2_a21oi_1 _23345_ (.A1(\top_ihp.oisc.regs[19][26] ),
    .A2(_05437_),
    .Y(_06771_),
    .B1(_06770_));
 sg13g2_a22oi_1 _23346_ (.Y(_06772_),
    .B1(net151),
    .B2(\top_ihp.oisc.regs[3][26] ),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[1][26] ));
 sg13g2_nand4_1 _23347_ (.B(_06767_),
    .C(_06771_),
    .A(_06766_),
    .Y(_06773_),
    .D(_06772_));
 sg13g2_a22oi_1 _23348_ (.Y(_06774_),
    .B1(net314),
    .B2(\top_ihp.oisc.regs[9][26] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[8][26] ));
 sg13g2_a22oi_1 _23349_ (.Y(_06775_),
    .B1(_05720_),
    .B2(\top_ihp.oisc.regs[15][26] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[25][26] ));
 sg13g2_a22oi_1 _23350_ (.Y(_06776_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][26] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[28][26] ));
 sg13g2_mux2_1 _23351_ (.A0(\top_ihp.oisc.regs[5][26] ),
    .A1(\top_ihp.oisc.regs[4][26] ),
    .S(net416),
    .X(_06777_));
 sg13g2_a22oi_1 _23352_ (.Y(_06778_),
    .B1(_06777_),
    .B2(_06481_),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][26] ));
 sg13g2_nand4_1 _23353_ (.B(_06775_),
    .C(_06776_),
    .A(_06774_),
    .Y(_06779_),
    .D(_06778_));
 sg13g2_a22oi_1 _23354_ (.Y(_06780_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][26] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][26] ));
 sg13g2_and2_1 _23355_ (.A(\top_ihp.oisc.regs[14][26] ),
    .B(net423),
    .X(_06781_));
 sg13g2_a221oi_1 _23356_ (.B2(\top_ihp.oisc.regs[23][26] ),
    .C1(_06781_),
    .B1(_05496_),
    .A1(\top_ihp.oisc.regs[26][26] ),
    .Y(_06782_),
    .A2(net333));
 sg13g2_mux2_1 _23357_ (.A0(\top_ihp.oisc.regs[31][26] ),
    .A1(\top_ihp.oisc.regs[29][26] ),
    .S(net668),
    .X(_06783_));
 sg13g2_and2_1 _23358_ (.A(net669),
    .B(_05433_),
    .X(_06784_));
 sg13g2_nor2_2 _23359_ (.A(_05676_),
    .B(net734),
    .Y(_06785_));
 sg13g2_mux2_1 _23360_ (.A0(\top_ihp.oisc.regs[21][26] ),
    .A1(\top_ihp.oisc.regs[17][26] ),
    .S(net418),
    .X(_06786_));
 sg13g2_a22oi_1 _23361_ (.Y(_06787_),
    .B1(_06785_),
    .B2(_06786_),
    .A2(_06784_),
    .A1(_06783_));
 sg13g2_a22oi_1 _23362_ (.Y(_06788_),
    .B1(_05732_),
    .B2(\top_ihp.oisc.regs[13][26] ),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][26] ));
 sg13g2_nand4_1 _23363_ (.B(_06782_),
    .C(_06787_),
    .A(_06780_),
    .Y(_06789_),
    .D(_06788_));
 sg13g2_a22oi_1 _23364_ (.Y(_06790_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[54][26] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][26] ));
 sg13g2_a22oi_1 _23365_ (.Y(_06791_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][26] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][26] ));
 sg13g2_nand3_1 _23366_ (.B(_06790_),
    .C(_06791_),
    .A(_05918_),
    .Y(_06792_));
 sg13g2_nor4_2 _23367_ (.A(_06773_),
    .B(_06779_),
    .C(_06789_),
    .Y(_06793_),
    .D(_06792_));
 sg13g2_a22oi_1 _23368_ (.Y(_06794_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][26] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][26] ));
 sg13g2_a22oi_1 _23369_ (.Y(_06795_),
    .B1(_06035_),
    .B2(\top_ihp.oisc.regs[39][26] ),
    .A2(_05327_),
    .A1(\top_ihp.oisc.regs[44][26] ));
 sg13g2_a22oi_1 _23370_ (.Y(_06796_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][26] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][26] ));
 sg13g2_a22oi_1 _23371_ (.Y(_06797_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[58][26] ),
    .A2(net329),
    .A1(\top_ihp.oisc.regs[50][26] ));
 sg13g2_nand4_1 _23372_ (.B(_06795_),
    .C(_06796_),
    .A(_06794_),
    .Y(_06798_),
    .D(_06797_));
 sg13g2_a22oi_1 _23373_ (.Y(_06799_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][26] ),
    .A2(net433),
    .A1(\top_ihp.oisc.regs[35][26] ));
 sg13g2_a22oi_1 _23374_ (.Y(_06800_),
    .B1(_05637_),
    .B2(\top_ihp.oisc.regs[59][26] ),
    .A2(net324),
    .A1(\top_ihp.oisc.regs[63][26] ));
 sg13g2_a22oi_1 _23375_ (.Y(_06801_),
    .B1(net186),
    .B2(\top_ihp.oisc.regs[33][26] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][26] ));
 sg13g2_a22oi_1 _23376_ (.Y(_06802_),
    .B1(net326),
    .B2(\top_ihp.oisc.regs[51][26] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][26] ));
 sg13g2_nand4_1 _23377_ (.B(_06800_),
    .C(_06801_),
    .A(_06799_),
    .Y(_06803_),
    .D(_06802_));
 sg13g2_nand2_1 _23378_ (.Y(_06804_),
    .A(\top_ihp.oisc.regs[37][26] ),
    .B(net74));
 sg13g2_a22oi_1 _23379_ (.Y(_06805_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][26] ),
    .A2(net307),
    .A1(\top_ihp.oisc.regs[34][26] ));
 sg13g2_nand2_1 _23380_ (.Y(_06806_),
    .A(_06804_),
    .B(_06805_));
 sg13g2_mux2_1 _23381_ (.A0(\top_ihp.oisc.regs[24][26] ),
    .A1(\top_ihp.oisc.regs[16][26] ),
    .S(_06162_),
    .X(_06807_));
 sg13g2_a22oi_1 _23382_ (.Y(_06808_),
    .B1(_06807_),
    .B2(_06313_),
    .A2(_06334_),
    .A1(\top_ihp.oisc.regs[61][26] ));
 sg13g2_nand2_1 _23383_ (.Y(_06809_),
    .A(\top_ihp.oisc.regs[40][26] ),
    .B(_05279_));
 sg13g2_nand3_1 _23384_ (.B(_05319_),
    .C(_05548_),
    .A(\top_ihp.oisc.regs[57][26] ),
    .Y(_06810_));
 sg13g2_o21ai_1 _23385_ (.B1(_06810_),
    .Y(_06811_),
    .A1(net707),
    .A2(_06809_));
 sg13g2_nor2_1 _23386_ (.A(net671),
    .B(net679),
    .Y(_06812_));
 sg13g2_a22oi_1 _23387_ (.Y(_06813_),
    .B1(_06811_),
    .B2(_06812_),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][26] ));
 sg13g2_nand2_1 _23388_ (.Y(_06814_),
    .A(_08217_),
    .B(net748));
 sg13g2_nand3_1 _23389_ (.B(net597),
    .C(_06017_),
    .A(\top_ihp.oisc.regs[7][26] ),
    .Y(_06815_));
 sg13g2_nand3_1 _23390_ (.B(_05851_),
    .C(_06240_),
    .A(\top_ihp.oisc.regs[12][26] ),
    .Y(_06816_));
 sg13g2_nand3_1 _23391_ (.B(_06815_),
    .C(_06816_),
    .A(_06814_),
    .Y(_06817_));
 sg13g2_a21oi_1 _23392_ (.A1(\top_ihp.oisc.regs[53][26] ),
    .A2(net72),
    .Y(_06818_),
    .B1(_06817_));
 sg13g2_a22oi_1 _23393_ (.Y(_06819_),
    .B1(_05745_),
    .B2(\top_ihp.oisc.regs[56][26] ),
    .A2(_05652_),
    .A1(\top_ihp.oisc.regs[55][26] ));
 sg13g2_nand4_1 _23394_ (.B(_06813_),
    .C(_06818_),
    .A(_06808_),
    .Y(_06820_),
    .D(_06819_));
 sg13g2_nor4_2 _23395_ (.A(_06798_),
    .B(_06803_),
    .C(_06806_),
    .Y(_06821_),
    .D(_06820_));
 sg13g2_a21o_1 _23396_ (.A2(_05945_),
    .A1(_00072_),
    .B1(_05946_),
    .X(_06822_));
 sg13g2_a22oi_1 _23397_ (.Y(_00438_),
    .B1(_06822_),
    .B2(_06814_),
    .A2(_06821_),
    .A1(_06793_));
 sg13g2_a22oi_1 _23398_ (.Y(_06823_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][27] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][27] ));
 sg13g2_a22oi_1 _23399_ (.Y(_06824_),
    .B1(net181),
    .B2(\top_ihp.oisc.regs[47][27] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][27] ));
 sg13g2_a22oi_1 _23400_ (.Y(_06825_),
    .B1(net77),
    .B2(\top_ihp.oisc.regs[55][27] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][27] ));
 sg13g2_a22oi_1 _23401_ (.Y(_06826_),
    .B1(net325),
    .B2(\top_ihp.oisc.regs[35][27] ),
    .A2(net329),
    .A1(\top_ihp.oisc.regs[50][27] ));
 sg13g2_nand4_1 _23402_ (.B(_06824_),
    .C(_06825_),
    .A(_06823_),
    .Y(_06827_),
    .D(_06826_));
 sg13g2_a22oi_1 _23403_ (.Y(_06828_),
    .B1(net183),
    .B2(\top_ihp.oisc.regs[63][27] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][27] ));
 sg13g2_a22oi_1 _23404_ (.Y(_06829_),
    .B1(net174),
    .B2(\top_ihp.oisc.regs[39][27] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][27] ));
 sg13g2_a22oi_1 _23405_ (.Y(_06830_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][27] ),
    .A2(_05605_),
    .A1(\top_ihp.oisc.regs[56][27] ));
 sg13g2_a22oi_1 _23406_ (.Y(_06831_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][27] ),
    .A2(net609),
    .A1(\top_ihp.oisc.regs[57][27] ));
 sg13g2_nand4_1 _23407_ (.B(_06829_),
    .C(_06830_),
    .A(_06828_),
    .Y(_06832_),
    .D(_06831_));
 sg13g2_a22oi_1 _23408_ (.Y(_06833_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][27] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][27] ));
 sg13g2_a22oi_1 _23409_ (.Y(_06834_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][27] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[45][27] ));
 sg13g2_a22oi_1 _23410_ (.Y(_06835_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][27] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][27] ));
 sg13g2_a22oi_1 _23411_ (.Y(_06836_),
    .B1(net178),
    .B2(\top_ihp.oisc.regs[46][27] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[36][27] ));
 sg13g2_nand4_1 _23412_ (.B(_06834_),
    .C(_06835_),
    .A(_06833_),
    .Y(_06837_),
    .D(_06836_));
 sg13g2_nor4_2 _23413_ (.A(net190),
    .B(_06827_),
    .C(_06832_),
    .Y(_06838_),
    .D(_06837_));
 sg13g2_and4_1 _23414_ (.A(\top_ihp.oisc.regs[28][27] ),
    .B(net291),
    .C(net608),
    .D(net673),
    .X(_06839_));
 sg13g2_a221oi_1 _23415_ (.B2(\top_ihp.oisc.regs[19][27] ),
    .C1(_06839_),
    .B1(net445),
    .A1(_08450_),
    .Y(_06840_),
    .A2(_06312_));
 sg13g2_a22oi_1 _23416_ (.Y(_06841_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[9][27] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[8][27] ));
 sg13g2_a22oi_1 _23417_ (.Y(_06842_),
    .B1(_05818_),
    .B2(\top_ihp.oisc.regs[30][27] ),
    .A2(net283),
    .A1(\top_ihp.oisc.regs[23][27] ));
 sg13g2_a22oi_1 _23418_ (.Y(_06843_),
    .B1(net603),
    .B2(\top_ihp.oisc.regs[27][27] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[13][27] ));
 sg13g2_nand4_1 _23419_ (.B(_06841_),
    .C(_06842_),
    .A(_06840_),
    .Y(_06844_),
    .D(_06843_));
 sg13g2_a22oi_1 _23420_ (.Y(_06845_),
    .B1(_05730_),
    .B2(\top_ihp.oisc.regs[10][27] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[31][27] ));
 sg13g2_a22oi_1 _23421_ (.Y(_06846_),
    .B1(net152),
    .B2(\top_ihp.oisc.regs[22][27] ),
    .A2(_05501_),
    .A1(\top_ihp.oisc.regs[3][27] ));
 sg13g2_a22oi_1 _23422_ (.Y(_06847_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][27] ),
    .A2(_05717_),
    .A1(\top_ihp.oisc.regs[18][27] ));
 sg13g2_a22oi_1 _23423_ (.Y(_06848_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][27] ),
    .A2(net318),
    .A1(\top_ihp.oisc.regs[11][27] ));
 sg13g2_nand4_1 _23424_ (.B(_06846_),
    .C(_06847_),
    .A(_06845_),
    .Y(_06849_),
    .D(_06848_));
 sg13g2_mux2_1 _23425_ (.A0(\top_ihp.oisc.regs[7][27] ),
    .A1(\top_ihp.oisc.regs[6][27] ),
    .S(net682),
    .X(_06850_));
 sg13g2_a22oi_1 _23426_ (.Y(_06851_),
    .B1(_06850_),
    .B2(net606),
    .A2(net410),
    .A1(\top_ihp.oisc.regs[14][27] ));
 sg13g2_nor2_1 _23427_ (.A(_05375_),
    .B(_06851_),
    .Y(_06852_));
 sg13g2_a221oi_1 _23428_ (.B2(\top_ihp.oisc.regs[48][27] ),
    .C1(_06852_),
    .B1(_05796_),
    .A1(\top_ihp.oisc.regs[43][27] ),
    .Y(_06853_),
    .A2(_05479_));
 sg13g2_nand2_1 _23429_ (.Y(_06854_),
    .A(\top_ihp.oisc.regs[20][27] ),
    .B(net419));
 sg13g2_nand2_1 _23430_ (.Y(_06855_),
    .A(\top_ihp.oisc.regs[16][27] ),
    .B(net604));
 sg13g2_a21oi_1 _23431_ (.A1(_06854_),
    .A2(_06855_),
    .Y(_06856_),
    .B1(_05355_));
 sg13g2_nand3_1 _23432_ (.B(net419),
    .C(net697),
    .A(\top_ihp.oisc.regs[29][27] ),
    .Y(_06857_));
 sg13g2_nand3_1 _23433_ (.B(net604),
    .C(net721),
    .A(\top_ihp.oisc.regs[26][27] ),
    .Y(_06858_));
 sg13g2_a21oi_1 _23434_ (.A1(_06857_),
    .A2(_06858_),
    .Y(_06859_),
    .B1(net602));
 sg13g2_a21oi_1 _23435_ (.A1(net417),
    .A2(_06856_),
    .Y(_06860_),
    .B1(_06859_));
 sg13g2_mux2_1 _23436_ (.A0(\top_ihp.oisc.regs[21][27] ),
    .A1(\top_ihp.oisc.regs[17][27] ),
    .S(net418),
    .X(_06861_));
 sg13g2_a22oi_1 _23437_ (.Y(_06862_),
    .B1(_06785_),
    .B2(_06861_),
    .A2(_05719_),
    .A1(\top_ihp.oisc.regs[15][27] ));
 sg13g2_nand2_1 _23438_ (.Y(_06863_),
    .A(\top_ihp.oisc.regs[25][27] ),
    .B(net316));
 sg13g2_nand4_1 _23439_ (.B(_06860_),
    .C(_06862_),
    .A(_06853_),
    .Y(_06864_),
    .D(_06863_));
 sg13g2_a22oi_1 _23440_ (.Y(_06865_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][27] ),
    .A2(net67),
    .A1(\top_ihp.oisc.regs[61][27] ));
 sg13g2_a22oi_1 _23441_ (.Y(_06866_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[49][27] ),
    .A2(_05634_),
    .A1(\top_ihp.oisc.regs[33][27] ));
 sg13g2_a22oi_1 _23442_ (.Y(_06867_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[12][27] ),
    .A2(_06017_),
    .A1(\top_ihp.oisc.regs[5][27] ));
 sg13g2_inv_1 _23443_ (.Y(_06868_),
    .A(_06867_));
 sg13g2_nand2_1 _23444_ (.Y(_06869_),
    .A(net674),
    .B(_05916_));
 sg13g2_a22oi_1 _23445_ (.Y(_06870_),
    .B1(_05556_),
    .B2(\top_ihp.oisc.regs[1][27] ),
    .A2(_05462_),
    .A1(\top_ihp.oisc.regs[4][27] ));
 sg13g2_nor2_1 _23446_ (.A(_06869_),
    .B(_06870_),
    .Y(_06871_));
 sg13g2_a21oi_1 _23447_ (.A1(net600),
    .A2(_06868_),
    .Y(_06872_),
    .B1(_06871_));
 sg13g2_a22oi_1 _23448_ (.Y(_06873_),
    .B1(net74),
    .B2(\top_ihp.oisc.regs[37][27] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][27] ));
 sg13g2_nand4_1 _23449_ (.B(_06866_),
    .C(_06872_),
    .A(_06865_),
    .Y(_06874_),
    .D(_06873_));
 sg13g2_nor4_1 _23450_ (.A(_06844_),
    .B(_06849_),
    .C(_06864_),
    .D(_06874_),
    .Y(_06875_));
 sg13g2_a21oi_1 _23451_ (.A1(_00073_),
    .A2(net150),
    .Y(_06876_),
    .B1(net32));
 sg13g2_a21oi_1 _23452_ (.A1(net1046),
    .A2(net693),
    .Y(_06877_),
    .B1(_06876_));
 sg13g2_a21oi_1 _23453_ (.A1(_06838_),
    .A2(_06875_),
    .Y(_00439_),
    .B1(_06877_));
 sg13g2_nand2_1 _23454_ (.Y(_06878_),
    .A(\top_ihp.oisc.regs[61][28] ),
    .B(net67));
 sg13g2_a22oi_1 _23455_ (.Y(_06879_),
    .B1(net72),
    .B2(\top_ihp.oisc.regs[53][28] ),
    .A2(net308),
    .A1(\top_ihp.oisc.regs[40][28] ));
 sg13g2_a22oi_1 _23456_ (.Y(_06880_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[36][28] ),
    .A2(net185),
    .A1(\top_ihp.oisc.regs[59][28] ));
 sg13g2_a22oi_1 _23457_ (.Y(_06881_),
    .B1(net306),
    .B2(\top_ihp.oisc.regs[34][28] ),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][28] ));
 sg13g2_nand4_1 _23458_ (.B(_06879_),
    .C(_06880_),
    .A(_06878_),
    .Y(_06882_),
    .D(_06881_));
 sg13g2_a22oi_1 _23459_ (.Y(_06883_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][28] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][28] ));
 sg13g2_a22oi_1 _23460_ (.Y(_06884_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][28] ),
    .A2(net325),
    .A1(\top_ihp.oisc.regs[35][28] ));
 sg13g2_a22oi_1 _23461_ (.Y(_06885_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][28] ),
    .A2(_06035_),
    .A1(\top_ihp.oisc.regs[39][28] ));
 sg13g2_a22oi_1 _23462_ (.Y(_06886_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[63][28] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][28] ));
 sg13g2_nand4_1 _23463_ (.B(_06884_),
    .C(_06885_),
    .A(_06883_),
    .Y(_06887_),
    .D(_06886_));
 sg13g2_a22oi_1 _23464_ (.Y(_06888_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[58][28] ),
    .A2(net329),
    .A1(\top_ihp.oisc.regs[50][28] ));
 sg13g2_a22oi_1 _23465_ (.Y(_06889_),
    .B1(_06518_),
    .B2(\top_ihp.oisc.regs[52][28] ),
    .A2(_05795_),
    .A1(\top_ihp.oisc.regs[45][28] ));
 sg13g2_and2_1 _23466_ (.A(_06888_),
    .B(_06889_),
    .X(_06890_));
 sg13g2_nand2_1 _23467_ (.Y(_06891_),
    .A(\top_ihp.oisc.regs[51][28] ),
    .B(net184));
 sg13g2_nand2_1 _23468_ (.Y(_06892_),
    .A(\top_ihp.oisc.regs[38][28] ),
    .B(net157));
 sg13g2_a22oi_1 _23469_ (.Y(_06893_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][28] ),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][28] ));
 sg13g2_nand4_1 _23470_ (.B(_06891_),
    .C(_06892_),
    .A(_06890_),
    .Y(_06894_),
    .D(_06893_));
 sg13g2_nor4_2 _23471_ (.A(net158),
    .B(_06882_),
    .C(_06887_),
    .Y(_06895_),
    .D(_06894_));
 sg13g2_a22oi_1 _23472_ (.Y(_06896_),
    .B1(net279),
    .B2(\top_ihp.oisc.regs[42][28] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][28] ));
 sg13g2_a22oi_1 _23473_ (.Y(_06897_),
    .B1(net77),
    .B2(\top_ihp.oisc.regs[55][28] ),
    .A2(net328),
    .A1(\top_ihp.oisc.regs[33][28] ));
 sg13g2_a22oi_1 _23474_ (.Y(_06898_),
    .B1(_05605_),
    .B2(\top_ihp.oisc.regs[56][28] ),
    .A2(net440),
    .A1(\top_ihp.oisc.regs[43][28] ));
 sg13g2_a22oi_1 _23475_ (.Y(_06899_),
    .B1(net290),
    .B2(\top_ihp.oisc.regs[17][28] ),
    .A2(net696),
    .A1(\top_ihp.oisc.regs[29][28] ));
 sg13g2_inv_1 _23476_ (.Y(_06900_),
    .A(_06899_));
 sg13g2_a22oi_1 _23477_ (.Y(_06901_),
    .B1(_06900_),
    .B2(_05932_),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][28] ));
 sg13g2_nand4_1 _23478_ (.B(_06897_),
    .C(_06898_),
    .A(_06896_),
    .Y(_06902_),
    .D(_06901_));
 sg13g2_a22oi_1 _23479_ (.Y(_06903_),
    .B1(_05817_),
    .B2(\top_ihp.oisc.regs[30][28] ),
    .A2(_05421_),
    .A1(\top_ihp.oisc.regs[18][28] ));
 sg13g2_a22oi_1 _23480_ (.Y(_06904_),
    .B1(_05493_),
    .B2(\top_ihp.oisc.regs[26][28] ),
    .A2(_05454_),
    .A1(\top_ihp.oisc.regs[11][28] ));
 sg13g2_a22oi_1 _23481_ (.Y(_06905_),
    .B1(net411),
    .B2(\top_ihp.oisc.regs[8][28] ),
    .A2(_05389_),
    .A1(\top_ihp.oisc.regs[20][28] ));
 sg13g2_a22oi_1 _23482_ (.Y(_06906_),
    .B1(net611),
    .B2(\top_ihp.oisc.regs[31][28] ),
    .A2(_05488_),
    .A1(\top_ihp.oisc.regs[1][28] ));
 sg13g2_and4_1 _23483_ (.A(_06903_),
    .B(_06904_),
    .C(_06905_),
    .D(_06906_),
    .X(_06907_));
 sg13g2_a22oi_1 _23484_ (.Y(_06908_),
    .B1(net172),
    .B2(\top_ihp.oisc.regs[37][28] ),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][28] ));
 sg13g2_nand2_1 _23485_ (.Y(_06909_),
    .A(\top_ihp.oisc.regs[13][28] ),
    .B(_05732_));
 sg13g2_a22oi_1 _23486_ (.Y(_06910_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][28] ),
    .A2(net426),
    .A1(\top_ihp.oisc.regs[25][28] ));
 sg13g2_nand4_1 _23487_ (.B(_06908_),
    .C(_06909_),
    .A(_06907_),
    .Y(_06911_),
    .D(_06910_));
 sg13g2_mux2_1 _23488_ (.A0(\top_ihp.oisc.regs[15][28] ),
    .A1(\top_ihp.oisc.regs[14][28] ),
    .S(_05847_),
    .X(_06912_));
 sg13g2_a22oi_1 _23489_ (.Y(_06913_),
    .B1(_06912_),
    .B2(_05376_),
    .A2(net151),
    .A1(\top_ihp.oisc.regs[3][28] ));
 sg13g2_a22oi_1 _23490_ (.Y(_06914_),
    .B1(net296),
    .B2(\top_ihp.oisc.regs[28][28] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][28] ));
 sg13g2_a22oi_1 _23491_ (.Y(_06915_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][28] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[4][28] ));
 sg13g2_a22oi_1 _23492_ (.Y(_06916_),
    .B1(net605),
    .B2(\top_ihp.oisc.regs[27][28] ),
    .A2(net297),
    .A1(\top_ihp.oisc.regs[5][28] ));
 sg13g2_nand4_1 _23493_ (.B(_06914_),
    .C(_06915_),
    .A(_06913_),
    .Y(_06917_),
    .D(_06916_));
 sg13g2_and3_1 _23494_ (.X(_06918_),
    .A(\top_ihp.oisc.regs[12][28] ),
    .B(net669),
    .C(_05813_));
 sg13g2_a221oi_1 _23495_ (.B2(\top_ihp.oisc.regs[19][28] ),
    .C1(_06918_),
    .B1(net427),
    .A1(_08443_),
    .Y(_06919_),
    .A2(_06312_));
 sg13g2_a22oi_1 _23496_ (.Y(_06920_),
    .B1(_05451_),
    .B2(\top_ihp.oisc.regs[21][28] ),
    .A2(net314),
    .A1(\top_ihp.oisc.regs[9][28] ));
 sg13g2_a22oi_1 _23497_ (.Y(_06921_),
    .B1(_05730_),
    .B2(\top_ihp.oisc.regs[10][28] ),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][28] ));
 sg13g2_nand3_1 _23498_ (.B(net291),
    .C(net694),
    .A(\top_ihp.oisc.regs[23][28] ),
    .Y(_06922_));
 sg13g2_nand3_1 _23499_ (.B(net598),
    .C(net673),
    .A(\top_ihp.oisc.regs[16][28] ),
    .Y(_06923_));
 sg13g2_nand2_1 _23500_ (.Y(_06924_),
    .A(_06922_),
    .B(_06923_));
 sg13g2_a22oi_1 _23501_ (.Y(_06925_),
    .B1(_06924_),
    .B2(_05890_),
    .A2(net152),
    .A1(\top_ihp.oisc.regs[22][28] ));
 sg13g2_nand4_1 _23502_ (.B(_06920_),
    .C(_06921_),
    .A(_06919_),
    .Y(_06926_),
    .D(_06925_));
 sg13g2_nor4_1 _23503_ (.A(_06902_),
    .B(_06911_),
    .C(_06917_),
    .D(_06926_),
    .Y(_06927_));
 sg13g2_a21oi_1 _23504_ (.A1(_00074_),
    .A2(net150),
    .Y(_06928_),
    .B1(net32));
 sg13g2_a21oi_1 _23505_ (.A1(_08443_),
    .A2(net693),
    .Y(_06929_),
    .B1(_06928_));
 sg13g2_a21oi_1 _23506_ (.A1(_06895_),
    .A2(_06927_),
    .Y(_00440_),
    .B1(_06929_));
 sg13g2_a22oi_1 _23507_ (.Y(_06930_),
    .B1(net179),
    .B2(\top_ihp.oisc.regs[54][29] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][29] ));
 sg13g2_a22oi_1 _23508_ (.Y(_06931_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[50][29] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][29] ));
 sg13g2_a22oi_1 _23509_ (.Y(_06932_),
    .B1(net307),
    .B2(\top_ihp.oisc.regs[34][29] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[42][29] ));
 sg13g2_a22oi_1 _23510_ (.Y(_06933_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[46][29] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[40][29] ));
 sg13g2_nand4_1 _23511_ (.B(_06931_),
    .C(_06932_),
    .A(_06930_),
    .Y(_06934_),
    .D(_06933_));
 sg13g2_a22oi_1 _23512_ (.Y(_06935_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][29] ),
    .A2(net74),
    .A1(\top_ihp.oisc.regs[37][29] ));
 sg13g2_a22oi_1 _23513_ (.Y(_06936_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][29] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[63][29] ));
 sg13g2_a22oi_1 _23514_ (.Y(_06937_),
    .B1(net310),
    .B2(\top_ihp.oisc.regs[48][29] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][29] ));
 sg13g2_a22oi_1 _23515_ (.Y(_06938_),
    .B1(net302),
    .B2(\top_ihp.oisc.regs[32][29] ),
    .A2(_05767_),
    .A1(\top_ihp.oisc.regs[44][29] ));
 sg13g2_nand4_1 _23516_ (.B(_06936_),
    .C(_06937_),
    .A(_06935_),
    .Y(_06939_),
    .D(_06938_));
 sg13g2_nand2_1 _23517_ (.Y(_06940_),
    .A(\top_ihp.oisc.regs[57][29] ),
    .B(net432));
 sg13g2_a22oi_1 _23518_ (.Y(_06941_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[33][29] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][29] ));
 sg13g2_a22oi_1 _23519_ (.Y(_06942_),
    .B1(_06233_),
    .B2(\top_ihp.oisc.regs[45][29] ),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][29] ));
 sg13g2_a22oi_1 _23520_ (.Y(_06943_),
    .B1(_05745_),
    .B2(\top_ihp.oisc.regs[56][29] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[36][29] ));
 sg13g2_nand4_1 _23521_ (.B(_06941_),
    .C(_06942_),
    .A(_06940_),
    .Y(_06944_),
    .D(_06943_));
 sg13g2_nor4_2 _23522_ (.A(net158),
    .B(_06934_),
    .C(_06939_),
    .Y(_06945_),
    .D(_06944_));
 sg13g2_a22oi_1 _23523_ (.Y(_06946_),
    .B1(_05705_),
    .B2(\top_ihp.oisc.regs[1][29] ),
    .A2(_06256_),
    .A1(\top_ihp.oisc.regs[7][29] ));
 sg13g2_a22oi_1 _23524_ (.Y(_06947_),
    .B1(_05504_),
    .B2(\top_ihp.oisc.regs[31][29] ),
    .A2(_05820_),
    .A1(\top_ihp.oisc.regs[27][29] ));
 sg13g2_a22oi_1 _23525_ (.Y(_06948_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][29] ),
    .A2(net444),
    .A1(\top_ihp.oisc.regs[21][29] ));
 sg13g2_mux2_1 _23526_ (.A0(\top_ihp.oisc.regs[14][29] ),
    .A1(\top_ihp.oisc.regs[6][29] ),
    .S(_05889_),
    .X(_06949_));
 sg13g2_and2_1 _23527_ (.A(_05892_),
    .B(_05825_),
    .X(_06950_));
 sg13g2_a22oi_1 _23528_ (.Y(_06951_),
    .B1(_06949_),
    .B2(_06950_),
    .A2(_05415_),
    .A1(\top_ihp.oisc.regs[9][29] ));
 sg13g2_nand4_1 _23529_ (.B(_06947_),
    .C(_06948_),
    .A(_06946_),
    .Y(_06952_),
    .D(_06951_));
 sg13g2_and3_1 _23530_ (.X(_06953_),
    .A(\top_ihp.oisc.regs[11][29] ),
    .B(_05845_),
    .C(net596));
 sg13g2_a21oi_1 _23531_ (.A1(\top_ihp.oisc.regs[22][29] ),
    .A2(_06066_),
    .Y(_06954_),
    .B1(_06953_));
 sg13g2_a22oi_1 _23532_ (.Y(_06955_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][29] ),
    .A2(net445),
    .A1(\top_ihp.oisc.regs[19][29] ));
 sg13g2_a22oi_1 _23533_ (.Y(_06956_),
    .B1(_05727_),
    .B2(\top_ihp.oisc.regs[12][29] ),
    .A2(_05683_),
    .A1(\top_ihp.oisc.regs[8][29] ));
 sg13g2_a22oi_1 _23534_ (.Y(_06957_),
    .B1(net151),
    .B2(\top_ihp.oisc.regs[3][29] ),
    .A2(net720),
    .A1(net1045));
 sg13g2_nand4_1 _23535_ (.B(_06955_),
    .C(_06956_),
    .A(_06954_),
    .Y(_06958_),
    .D(_06957_));
 sg13g2_a22oi_1 _23536_ (.Y(_06959_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][29] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[39][29] ));
 sg13g2_a22oi_1 _23537_ (.Y(_06960_),
    .B1(_05630_),
    .B2(\top_ihp.oisc.regs[61][29] ),
    .A2(net77),
    .A1(\top_ihp.oisc.regs[55][29] ));
 sg13g2_a22oi_1 _23538_ (.Y(_06961_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][29] ),
    .A2(net173),
    .A1(\top_ihp.oisc.regs[53][29] ));
 sg13g2_a22oi_1 _23539_ (.Y(_06962_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][29] ),
    .A2(_05662_),
    .A1(\top_ihp.oisc.regs[58][29] ));
 sg13g2_nand4_1 _23540_ (.B(_06960_),
    .C(_06961_),
    .A(_06959_),
    .Y(_06963_),
    .D(_06962_));
 sg13g2_a22oi_1 _23541_ (.Y(_06964_),
    .B1(_05715_),
    .B2(\top_ihp.oisc.regs[25][29] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][29] ));
 sg13g2_a22oi_1 _23542_ (.Y(_06965_),
    .B1(_05720_),
    .B2(\top_ihp.oisc.regs[15][29] ),
    .A2(net293),
    .A1(\top_ihp.oisc.regs[20][29] ));
 sg13g2_nand2_1 _23543_ (.Y(_06966_),
    .A(\top_ihp.oisc.regs[13][29] ),
    .B(_05403_));
 sg13g2_nor2_1 _23544_ (.A(net434),
    .B(_05279_),
    .Y(_06967_));
 sg13g2_nand4_1 _23545_ (.B(net595),
    .C(_06967_),
    .A(\top_ihp.oisc.regs[51][29] ),
    .Y(_06968_),
    .D(_06154_));
 sg13g2_a22oi_1 _23546_ (.Y(_06969_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[10][29] ),
    .A2(_05456_),
    .A1(\top_ihp.oisc.regs[28][29] ));
 sg13g2_and3_1 _23547_ (.X(_06970_),
    .A(_06966_),
    .B(_06968_),
    .C(_06969_));
 sg13g2_a22oi_1 _23548_ (.Y(_06971_),
    .B1(_05691_),
    .B2(\top_ihp.oisc.regs[2][29] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][29] ));
 sg13g2_a22oi_1 _23549_ (.Y(_06972_),
    .B1(net425),
    .B2(\top_ihp.oisc.regs[29][29] ),
    .A2(_05421_),
    .A1(\top_ihp.oisc.regs[18][29] ));
 sg13g2_a22oi_1 _23550_ (.Y(_06973_),
    .B1(_05507_),
    .B2(\top_ihp.oisc.regs[4][29] ),
    .A2(_05493_),
    .A1(\top_ihp.oisc.regs[26][29] ));
 sg13g2_a22oi_1 _23551_ (.Y(_06974_),
    .B1(_05817_),
    .B2(\top_ihp.oisc.regs[30][29] ),
    .A2(_05496_),
    .A1(\top_ihp.oisc.regs[23][29] ));
 sg13g2_and4_1 _23552_ (.A(_06971_),
    .B(_06972_),
    .C(_06973_),
    .D(_06974_),
    .X(_06975_));
 sg13g2_nand4_1 _23553_ (.B(_06965_),
    .C(_06970_),
    .A(_06964_),
    .Y(_06976_),
    .D(_06975_));
 sg13g2_nor4_1 _23554_ (.A(_06952_),
    .B(_06958_),
    .C(_06963_),
    .D(_06976_),
    .Y(_06977_));
 sg13g2_a21oi_1 _23555_ (.A1(_00075_),
    .A2(net150),
    .Y(_06978_),
    .B1(net32));
 sg13g2_a21oi_1 _23556_ (.A1(_08557_),
    .A2(_06390_),
    .Y(_06979_),
    .B1(_06978_));
 sg13g2_a21oi_1 _23557_ (.A1(_06945_),
    .A2(_06977_),
    .Y(_00441_),
    .B1(_06979_));
 sg13g2_nand2_2 _23558_ (.Y(_06980_),
    .A(_08329_),
    .B(net748));
 sg13g2_a21o_1 _23559_ (.A2(_05948_),
    .A1(_00243_),
    .B1(net34),
    .X(_06981_));
 sg13g2_nand3_1 _23560_ (.B(_05462_),
    .C(net668),
    .A(\top_ihp.oisc.regs[4][2] ),
    .Y(_06982_));
 sg13g2_nand3_1 _23561_ (.B(net671),
    .C(_05556_),
    .A(\top_ihp.oisc.regs[3][2] ),
    .Y(_06983_));
 sg13g2_nand2_1 _23562_ (.Y(_06984_),
    .A(net602),
    .B(_05609_));
 sg13g2_a21oi_1 _23563_ (.A1(_06982_),
    .A2(_06983_),
    .Y(_06985_),
    .B1(_06984_));
 sg13g2_a221oi_1 _23564_ (.B2(\top_ihp.oisc.regs[50][2] ),
    .C1(_06985_),
    .B1(net189),
    .A1(\top_ihp.oisc.regs[40][2] ),
    .Y(_06986_),
    .A2(net288));
 sg13g2_inv_1 _23565_ (.Y(_06987_),
    .A(_06986_));
 sg13g2_a22oi_1 _23566_ (.Y(_06988_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][2] ),
    .A2(net70),
    .A1(\top_ihp.oisc.regs[45][2] ));
 sg13g2_a22oi_1 _23567_ (.Y(_06989_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][2] ),
    .A2(net179),
    .A1(\top_ihp.oisc.regs[54][2] ));
 sg13g2_a22oi_1 _23568_ (.Y(_06990_),
    .B1(net311),
    .B2(\top_ihp.oisc.regs[52][2] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][2] ));
 sg13g2_a22oi_1 _23569_ (.Y(_06991_),
    .B1(_05955_),
    .B2(\top_ihp.oisc.regs[56][2] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][2] ));
 sg13g2_nand4_1 _23570_ (.B(_06989_),
    .C(_06990_),
    .A(_06988_),
    .Y(_06992_),
    .D(_06991_));
 sg13g2_nor3_1 _23571_ (.A(net159),
    .B(_06987_),
    .C(_06992_),
    .Y(_06993_));
 sg13g2_and2_1 _23572_ (.A(\top_ihp.oisc.regs[59][2] ),
    .B(_06967_),
    .X(_06994_));
 sg13g2_nand2_1 _23573_ (.Y(_06995_),
    .A(\top_ihp.oisc.regs[10][2] ),
    .B(_05914_));
 sg13g2_nand2_1 _23574_ (.Y(_06996_),
    .A(\top_ihp.oisc.regs[11][2] ),
    .B(_06433_));
 sg13g2_a21oi_1 _23575_ (.A1(_06995_),
    .A2(_06996_),
    .Y(_06997_),
    .B1(_06478_));
 sg13g2_a221oi_1 _23576_ (.B2(_06994_),
    .C1(_06997_),
    .B1(_05463_),
    .A1(\top_ihp.oisc.regs[8][2] ),
    .Y(_06998_),
    .A2(net429));
 sg13g2_a22oi_1 _23577_ (.Y(_06999_),
    .B1(net698),
    .B2(\top_ihp.oisc.regs[19][2] ),
    .A2(net672),
    .A1(\top_ihp.oisc.regs[16][2] ));
 sg13g2_a221oi_1 _23578_ (.B2(\top_ihp.oisc.regs[25][2] ),
    .C1(net599),
    .B1(net722),
    .A1(\top_ihp.oisc.regs[27][2] ),
    .Y(_07000_),
    .A2(net698));
 sg13g2_a21oi_1 _23579_ (.A1(net602),
    .A2(_06999_),
    .Y(_07001_),
    .B1(_07000_));
 sg13g2_a22oi_1 _23580_ (.Y(_07002_),
    .B1(_07001_),
    .B2(net412),
    .A2(net317),
    .A1(\top_ihp.oisc.regs[1][2] ));
 sg13g2_nand3_1 _23581_ (.B(_05938_),
    .C(_05825_),
    .A(\top_ihp.oisc.regs[2][2] ),
    .Y(_07003_));
 sg13g2_mux2_1 _23582_ (.A0(\top_ihp.oisc.regs[23][2] ),
    .A1(\top_ihp.oisc.regs[21][2] ),
    .S(_05303_),
    .X(_07004_));
 sg13g2_nand3_1 _23583_ (.B(_05433_),
    .C(_07004_),
    .A(net419),
    .Y(_07005_));
 sg13g2_nand2_1 _23584_ (.Y(_07006_),
    .A(_07003_),
    .B(_07005_));
 sg13g2_a22oi_1 _23585_ (.Y(_07007_),
    .B1(_07006_),
    .B2(net417),
    .A2(_05494_),
    .A1(\top_ihp.oisc.regs[26][2] ));
 sg13g2_mux2_1 _23586_ (.A0(\top_ihp.oisc.regs[30][2] ),
    .A1(\top_ihp.oisc.regs[28][2] ),
    .S(net701),
    .X(_07008_));
 sg13g2_a22oi_1 _23587_ (.Y(_07009_),
    .B1(_06059_),
    .B2(_07008_),
    .A2(_05381_),
    .A1(\top_ihp.oisc.regs[5][2] ));
 sg13g2_nand3_1 _23588_ (.B(_06021_),
    .C(_06002_),
    .A(\top_ihp.oisc.regs[6][2] ),
    .Y(_07010_));
 sg13g2_nand3_1 _23589_ (.B(_05850_),
    .C(_05845_),
    .A(\top_ihp.oisc.regs[13][2] ),
    .Y(_07011_));
 sg13g2_nand4_1 _23590_ (.B(_07009_),
    .C(_07010_),
    .A(_06980_),
    .Y(_07012_),
    .D(_07011_));
 sg13g2_a22oi_1 _23591_ (.Y(_07013_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][2] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[31][2] ));
 sg13g2_a22oi_1 _23592_ (.Y(_07014_),
    .B1(_05579_),
    .B2(\top_ihp.oisc.regs[18][2] ),
    .A2(_05447_),
    .A1(\top_ihp.oisc.regs[17][2] ));
 sg13g2_or4_1 _23593_ (.A(net434),
    .B(_05566_),
    .C(_05351_),
    .D(_07014_),
    .X(_07015_));
 sg13g2_nand4_1 _23594_ (.B(_05319_),
    .C(net607),
    .A(\top_ihp.oisc.regs[15][2] ),
    .Y(_07016_),
    .D(_06021_));
 sg13g2_nand2_1 _23595_ (.Y(_07017_),
    .A(\top_ihp.oisc.regs[29][2] ),
    .B(_05724_));
 sg13g2_nand4_1 _23596_ (.B(_07015_),
    .C(_07016_),
    .A(_07013_),
    .Y(_07018_),
    .D(_07017_));
 sg13g2_nor2_1 _23597_ (.A(_07012_),
    .B(_07018_),
    .Y(_07019_));
 sg13g2_nand4_1 _23598_ (.B(_07002_),
    .C(_07007_),
    .A(_06998_),
    .Y(_07020_),
    .D(_07019_));
 sg13g2_a22oi_1 _23599_ (.Y(_07021_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][2] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[33][2] ));
 sg13g2_a22oi_1 _23600_ (.Y(_07022_),
    .B1(net174),
    .B2(\top_ihp.oisc.regs[39][2] ),
    .A2(net172),
    .A1(\top_ihp.oisc.regs[37][2] ));
 sg13g2_a22oi_1 _23601_ (.Y(_07023_),
    .B1(net72),
    .B2(\top_ihp.oisc.regs[53][2] ),
    .A2(net160),
    .A1(\top_ihp.oisc.regs[63][2] ));
 sg13g2_a22oi_1 _23602_ (.Y(_07024_),
    .B1(_05442_),
    .B2(\top_ihp.oisc.regs[24][2] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[20][2] ));
 sg13g2_inv_1 _23603_ (.Y(_07025_),
    .A(_07024_));
 sg13g2_a22oi_1 _23604_ (.Y(_07026_),
    .B1(_07025_),
    .B2(net673),
    .A2(_05765_),
    .A1(\top_ihp.oisc.regs[49][2] ));
 sg13g2_nand4_1 _23605_ (.B(_07022_),
    .C(_07023_),
    .A(_07021_),
    .Y(_07027_),
    .D(_07026_));
 sg13g2_a22oi_1 _23606_ (.Y(_07028_),
    .B1(_06240_),
    .B2(\top_ihp.oisc.regs[14][2] ),
    .A2(_06017_),
    .A1(\top_ihp.oisc.regs[7][2] ));
 sg13g2_inv_1 _23607_ (.Y(_07029_),
    .A(_07028_));
 sg13g2_a22oi_1 _23608_ (.Y(_07030_),
    .B1(_05556_),
    .B2(\top_ihp.oisc.regs[9][2] ),
    .A2(_05462_),
    .A1(\top_ihp.oisc.regs[12][2] ));
 sg13g2_nor3_1 _23609_ (.A(net602),
    .B(_05610_),
    .C(_07030_),
    .Y(_07031_));
 sg13g2_a21oi_2 _23610_ (.B1(_07031_),
    .Y(_07032_),
    .A2(_07029_),
    .A1(net597));
 sg13g2_a22oi_1 _23611_ (.Y(_07033_),
    .B1(_05659_),
    .B2(\top_ihp.oisc.regs[47][2] ),
    .A2(_06403_),
    .A1(\top_ihp.oisc.regs[62][2] ));
 sg13g2_a22oi_1 _23612_ (.Y(_07034_),
    .B1(net68),
    .B2(\top_ihp.oisc.regs[55][2] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][2] ));
 sg13g2_a22oi_1 _23613_ (.Y(_07035_),
    .B1(net67),
    .B2(\top_ihp.oisc.regs[61][2] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][2] ));
 sg13g2_nand4_1 _23614_ (.B(_07033_),
    .C(_07034_),
    .A(_07032_),
    .Y(_07036_),
    .D(_07035_));
 sg13g2_a22oi_1 _23615_ (.Y(_07037_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][2] ),
    .A2(net322),
    .A1(\top_ihp.oisc.regs[58][2] ));
 sg13g2_a22oi_1 _23616_ (.Y(_07038_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][2] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[42][2] ));
 sg13g2_a22oi_1 _23617_ (.Y(_07039_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][2] ),
    .A2(net178),
    .A1(\top_ihp.oisc.regs[46][2] ));
 sg13g2_a22oi_1 _23618_ (.Y(_07040_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][2] ),
    .A2(net302),
    .A1(\top_ihp.oisc.regs[32][2] ));
 sg13g2_nand4_1 _23619_ (.B(_07038_),
    .C(_07039_),
    .A(_07037_),
    .Y(_07041_),
    .D(_07040_));
 sg13g2_nor4_1 _23620_ (.A(_07020_),
    .B(_07027_),
    .C(_07036_),
    .D(_07041_),
    .Y(_07042_));
 sg13g2_a22oi_1 _23621_ (.Y(_00442_),
    .B1(_06993_),
    .B2(_07042_),
    .A2(_06981_),
    .A1(_06980_));
 sg13g2_a22oi_1 _23622_ (.Y(_07043_),
    .B1(_06138_),
    .B2(\top_ihp.oisc.regs[23][30] ),
    .A2(net605),
    .A1(\top_ihp.oisc.regs[27][30] ));
 sg13g2_a22oi_1 _23623_ (.Y(_07044_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[13][30] ),
    .A2(net297),
    .A1(\top_ihp.oisc.regs[5][30] ));
 sg13g2_a22oi_1 _23624_ (.Y(_07045_),
    .B1(_06354_),
    .B2(\top_ihp.oisc.regs[3][30] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][30] ));
 sg13g2_a22oi_1 _23625_ (.Y(_07046_),
    .B1(net286),
    .B2(\top_ihp.oisc.regs[22][30] ),
    .A2(_05876_),
    .A1(\top_ihp.oisc.regs[6][30] ));
 sg13g2_nand4_1 _23626_ (.B(_07044_),
    .C(_07045_),
    .A(_07043_),
    .Y(_07047_),
    .D(_07046_));
 sg13g2_a22oi_1 _23627_ (.Y(_07048_),
    .B1(_05884_),
    .B2(\top_ihp.oisc.regs[7][30] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][30] ));
 sg13g2_nand2_1 _23628_ (.Y(_07049_),
    .A(\top_ihp.oisc.regs[15][30] ),
    .B(_05700_));
 sg13g2_a22oi_1 _23629_ (.Y(_07050_),
    .B1(_05813_),
    .B2(\top_ihp.oisc.regs[12][30] ),
    .A2(net694),
    .A1(\top_ihp.oisc.regs[31][30] ));
 sg13g2_nand2_1 _23630_ (.Y(_07051_),
    .A(_07049_),
    .B(_07050_));
 sg13g2_a22oi_1 _23631_ (.Y(_07052_),
    .B1(net669),
    .B2(_07051_),
    .A2(net728),
    .A1(_08546_));
 sg13g2_a22oi_1 _23632_ (.Y(_07053_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][30] ),
    .A2(net318),
    .A1(\top_ihp.oisc.regs[11][30] ));
 sg13g2_nand3_1 _23633_ (.B(_07052_),
    .C(_07053_),
    .A(_07048_),
    .Y(_07054_));
 sg13g2_a22oi_1 _23634_ (.Y(_07055_),
    .B1(_05649_),
    .B2(\top_ihp.oisc.regs[63][30] ),
    .A2(_06276_),
    .A1(\top_ihp.oisc.regs[32][30] ));
 sg13g2_nand3_1 _23635_ (.B(_05914_),
    .C(_05407_),
    .A(\top_ihp.oisc.regs[14][30] ),
    .Y(_07056_));
 sg13g2_nand3_1 _23636_ (.B(net599),
    .C(net672),
    .A(\top_ihp.oisc.regs[20][30] ),
    .Y(_07057_));
 sg13g2_o21ai_1 _23637_ (.B1(_07057_),
    .Y(_07058_),
    .A1(_06162_),
    .A2(_07056_));
 sg13g2_nand3_1 _23638_ (.B(net291),
    .C(_06003_),
    .A(\top_ihp.oisc.regs[30][30] ),
    .Y(_07059_));
 sg13g2_nand3_1 _23639_ (.B(_05938_),
    .C(net668),
    .A(\top_ihp.oisc.regs[24][30] ),
    .Y(_07060_));
 sg13g2_nand2_1 _23640_ (.Y(_07061_),
    .A(_07059_),
    .B(_07060_));
 sg13g2_nor2_1 _23641_ (.A(_05832_),
    .B(_05568_),
    .Y(_07062_));
 sg13g2_a22oi_1 _23642_ (.Y(_07063_),
    .B1(_07061_),
    .B2(_07062_),
    .A2(_07058_),
    .A1(_05681_));
 sg13g2_a22oi_1 _23643_ (.Y(_07064_),
    .B1(_06708_),
    .B2(\top_ihp.oisc.regs[56][30] ),
    .A2(_05741_),
    .A1(\top_ihp.oisc.regs[52][30] ));
 sg13g2_a22oi_1 _23644_ (.Y(_07065_),
    .B1(net699),
    .B2(\top_ihp.oisc.regs[8][30] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[4][30] ));
 sg13g2_inv_1 _23645_ (.Y(_07066_),
    .A(_07065_));
 sg13g2_a22oi_1 _23646_ (.Y(_07067_),
    .B1(_05813_),
    .B2(_07066_),
    .A2(_05796_),
    .A1(\top_ihp.oisc.regs[48][30] ));
 sg13g2_nand4_1 _23647_ (.B(_07063_),
    .C(_07064_),
    .A(_07055_),
    .Y(_07068_),
    .D(_07067_));
 sg13g2_nand3_1 _23648_ (.B(_05674_),
    .C(net695),
    .A(\top_ihp.oisc.regs[26][30] ),
    .Y(_07069_));
 sg13g2_nand3_1 _23649_ (.B(_05696_),
    .C(net697),
    .A(\top_ihp.oisc.regs[17][30] ),
    .Y(_07070_));
 sg13g2_nand2_1 _23650_ (.Y(_07071_),
    .A(_07069_),
    .B(_07070_));
 sg13g2_mux2_1 _23651_ (.A0(\top_ihp.oisc.regs[29][30] ),
    .A1(\top_ihp.oisc.regs[21][30] ),
    .S(net595),
    .X(_07072_));
 sg13g2_a22oi_1 _23652_ (.Y(_07073_),
    .B1(_07072_),
    .B2(_05807_),
    .A2(_07071_),
    .A1(_06053_));
 sg13g2_a22oi_1 _23653_ (.Y(_07074_),
    .B1(_05709_),
    .B2(\top_ihp.oisc.regs[19][30] ),
    .A2(net176),
    .A1(\top_ihp.oisc.regs[18][30] ));
 sg13g2_nand3_1 _23654_ (.B(_05878_),
    .C(net672),
    .A(\top_ihp.oisc.regs[28][30] ),
    .Y(_07075_));
 sg13g2_nand3_1 _23655_ (.B(net604),
    .C(_05575_),
    .A(\top_ihp.oisc.regs[25][30] ),
    .Y(_07076_));
 sg13g2_nand2_1 _23656_ (.Y(_07077_),
    .A(_07075_),
    .B(_07076_));
 sg13g2_mux2_1 _23657_ (.A0(\top_ihp.oisc.regs[9][30] ),
    .A1(\top_ihp.oisc.regs[1][30] ),
    .S(net675),
    .X(_07078_));
 sg13g2_nand2_1 _23658_ (.Y(_07079_),
    .A(_06418_),
    .B(_07078_));
 sg13g2_nand4_1 _23659_ (.B(net599),
    .C(_05535_),
    .A(\top_ihp.oisc.regs[55][30] ),
    .Y(_07080_),
    .D(_06154_));
 sg13g2_nand2_1 _23660_ (.Y(_07081_),
    .A(_07079_),
    .B(_07080_));
 sg13g2_a221oi_1 _23661_ (.B2(net415),
    .C1(_07081_),
    .B1(_07077_),
    .A1(\top_ihp.oisc.regs[2][30] ),
    .Y(_07082_),
    .A2(net295));
 sg13g2_a22oi_1 _23662_ (.Y(_07083_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][30] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][30] ));
 sg13g2_nand4_1 _23663_ (.B(_07074_),
    .C(_07082_),
    .A(_07073_),
    .Y(_07084_),
    .D(_07083_));
 sg13g2_nor4_2 _23664_ (.A(_07047_),
    .B(_07054_),
    .C(_07068_),
    .Y(_07085_),
    .D(_07084_));
 sg13g2_a22oi_1 _23665_ (.Y(_07086_),
    .B1(_06233_),
    .B2(\top_ihp.oisc.regs[45][30] ),
    .A2(_05739_),
    .A1(\top_ihp.oisc.regs[37][30] ));
 sg13g2_a22oi_1 _23666_ (.Y(_07087_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][30] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][30] ));
 sg13g2_a22oi_1 _23667_ (.Y(_07088_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][30] ),
    .A2(net307),
    .A1(\top_ihp.oisc.regs[34][30] ));
 sg13g2_a22oi_1 _23668_ (.Y(_07089_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][30] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][30] ));
 sg13g2_nand4_1 _23669_ (.B(_07087_),
    .C(_07088_),
    .A(_07086_),
    .Y(_07090_),
    .D(_07089_));
 sg13g2_a22oi_1 _23670_ (.Y(_07091_),
    .B1(net288),
    .B2(\top_ihp.oisc.regs[40][30] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][30] ));
 sg13g2_a22oi_1 _23671_ (.Y(_07092_),
    .B1(net67),
    .B2(\top_ihp.oisc.regs[61][30] ),
    .A2(_06403_),
    .A1(\top_ihp.oisc.regs[62][30] ));
 sg13g2_a22oi_1 _23672_ (.Y(_07093_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][30] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][30] ));
 sg13g2_a22oi_1 _23673_ (.Y(_07094_),
    .B1(net154),
    .B2(\top_ihp.oisc.regs[47][30] ),
    .A2(net174),
    .A1(\top_ihp.oisc.regs[39][30] ));
 sg13g2_nand4_1 _23674_ (.B(_07092_),
    .C(_07093_),
    .A(_07091_),
    .Y(_07095_),
    .D(_07094_));
 sg13g2_a22oi_1 _23675_ (.Y(_07096_),
    .B1(net609),
    .B2(\top_ihp.oisc.regs[57][30] ),
    .A2(_05528_),
    .A1(\top_ihp.oisc.regs[33][30] ));
 sg13g2_inv_1 _23676_ (.Y(_07097_),
    .A(_07096_));
 sg13g2_a221oi_1 _23677_ (.B2(\top_ihp.oisc.regs[59][30] ),
    .C1(_07097_),
    .B1(_05637_),
    .A1(\top_ihp.oisc.regs[49][30] ),
    .Y(_07098_),
    .A2(net441));
 sg13g2_nand2_1 _23678_ (.Y(_07099_),
    .A(\top_ihp.oisc.regs[42][30] ),
    .B(net191));
 sg13g2_a22oi_1 _23679_ (.Y(_07100_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][30] ),
    .A2(net72),
    .A1(\top_ihp.oisc.regs[53][30] ));
 sg13g2_nand4_1 _23680_ (.B(_07098_),
    .C(_07099_),
    .A(_05918_),
    .Y(_07101_),
    .D(_07100_));
 sg13g2_nor3_1 _23681_ (.A(_07090_),
    .B(_07095_),
    .C(_07101_),
    .Y(_07102_));
 sg13g2_a21oi_1 _23682_ (.A1(_00076_),
    .A2(_06506_),
    .Y(_07103_),
    .B1(_06559_));
 sg13g2_a21oi_1 _23683_ (.A1(_08546_),
    .A2(net693),
    .Y(_07104_),
    .B1(_07103_));
 sg13g2_a21oi_1 _23684_ (.A1(_07085_),
    .A2(_07102_),
    .Y(_00443_),
    .B1(_07104_));
 sg13g2_nand2_1 _23685_ (.Y(_07105_),
    .A(\top_ihp.oisc.regs[35][31] ),
    .B(net300));
 sg13g2_a22oi_1 _23686_ (.Y(_07106_),
    .B1(_05646_),
    .B2(\top_ihp.oisc.regs[57][31] ),
    .A2(net302),
    .A1(\top_ihp.oisc.regs[32][31] ));
 sg13g2_nand2_1 _23687_ (.Y(_07107_),
    .A(_07105_),
    .B(_07106_));
 sg13g2_a22oi_1 _23688_ (.Y(_07108_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][31] ),
    .A2(net78),
    .A1(\top_ihp.oisc.regs[59][31] ));
 sg13g2_a22oi_1 _23689_ (.Y(_07109_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][31] ),
    .A2(net186),
    .A1(\top_ihp.oisc.regs[33][31] ));
 sg13g2_nand3_1 _23690_ (.B(net594),
    .C(_05900_),
    .A(\top_ihp.oisc.regs[3][31] ),
    .Y(_07110_));
 sg13g2_nand3_1 _23691_ (.B(net416),
    .C(net696),
    .A(\top_ihp.oisc.regs[14][31] ),
    .Y(_07111_));
 sg13g2_a21oi_1 _23692_ (.A1(_07110_),
    .A2(_07111_),
    .Y(_07112_),
    .B1(_05699_));
 sg13g2_a221oi_1 _23693_ (.B2(\top_ihp.oisc.regs[11][31] ),
    .C1(_07112_),
    .B1(net443),
    .A1(\top_ihp.oisc.regs[12][31] ),
    .Y(_07113_),
    .A2(net448));
 sg13g2_a22oi_1 _23694_ (.Y(_07114_),
    .B1(_05603_),
    .B2(\top_ihp.oisc.regs[46][31] ),
    .A2(_05516_),
    .A1(\top_ihp.oisc.regs[54][31] ));
 sg13g2_a22oi_1 _23695_ (.Y(_07115_),
    .B1(_05543_),
    .B2(\top_ihp.oisc.regs[61][31] ),
    .A2(_05326_),
    .A1(\top_ihp.oisc.regs[44][31] ));
 sg13g2_a22oi_1 _23696_ (.Y(_07116_),
    .B1(_05588_),
    .B2(\top_ihp.oisc.regs[47][31] ),
    .A2(_05519_),
    .A1(\top_ihp.oisc.regs[40][31] ));
 sg13g2_a22oi_1 _23697_ (.Y(_07117_),
    .B1(_05544_),
    .B2(\top_ihp.oisc.regs[58][31] ),
    .A2(_05471_),
    .A1(\top_ihp.oisc.regs[37][31] ));
 sg13g2_and4_1 _23698_ (.A(_07114_),
    .B(_07115_),
    .C(_07116_),
    .D(_07117_),
    .X(_07118_));
 sg13g2_nand4_1 _23699_ (.B(_07109_),
    .C(_07113_),
    .A(_07108_),
    .Y(_07119_),
    .D(_07118_));
 sg13g2_a22oi_1 _23700_ (.Y(_07120_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[50][31] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][31] ));
 sg13g2_a22oi_1 _23701_ (.Y(_07121_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][31] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][31] ));
 sg13g2_a22oi_1 _23702_ (.Y(_07122_),
    .B1(net68),
    .B2(\top_ihp.oisc.regs[55][31] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][31] ));
 sg13g2_a22oi_1 _23703_ (.Y(_07123_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][31] ),
    .A2(_05752_),
    .A1(\top_ihp.oisc.regs[34][31] ));
 sg13g2_nand4_1 _23704_ (.B(_07121_),
    .C(_07122_),
    .A(_07120_),
    .Y(_07124_),
    .D(_07123_));
 sg13g2_nor4_1 _23705_ (.A(net158),
    .B(_07107_),
    .C(_07119_),
    .D(_07124_),
    .Y(_07125_));
 sg13g2_a22oi_1 _23706_ (.Y(_07126_),
    .B1(net283),
    .B2(\top_ihp.oisc.regs[23][31] ),
    .A2(net281),
    .A1(\top_ihp.oisc.regs[7][31] ));
 sg13g2_a22oi_1 _23707_ (.Y(_07127_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][31] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[31][31] ));
 sg13g2_mux2_1 _23708_ (.A0(\top_ihp.oisc.regs[26][31] ),
    .A1(\top_ihp.oisc.regs[24][31] ),
    .S(_05530_),
    .X(_07128_));
 sg13g2_nand2_1 _23709_ (.Y(_07129_),
    .A(net724),
    .B(_07128_));
 sg13g2_nand3_1 _23710_ (.B(net594),
    .C(_05916_),
    .A(\top_ihp.oisc.regs[9][31] ),
    .Y(_07130_));
 sg13g2_a21oi_1 _23711_ (.A1(_07129_),
    .A2(_07130_),
    .Y(_07131_),
    .B1(_05508_));
 sg13g2_a221oi_1 _23712_ (.B2(\top_ihp.oisc.regs[13][31] ),
    .C1(_07131_),
    .B1(_06010_),
    .A1(\top_ihp.oisc.regs[2][31] ),
    .Y(_07132_),
    .A2(net295));
 sg13g2_nand3_1 _23713_ (.B(net434),
    .C(_05813_),
    .A(\top_ihp.oisc.regs[4][31] ),
    .Y(_07133_));
 sg13g2_nand3_1 _23714_ (.B(net610),
    .C(net698),
    .A(\top_ihp.oisc.regs[19][31] ),
    .Y(_07134_));
 sg13g2_a21oi_1 _23715_ (.A1(_07133_),
    .A2(_07134_),
    .Y(_07135_),
    .B1(net413));
 sg13g2_a221oi_1 _23716_ (.B2(\top_ihp.oisc.regs[18][31] ),
    .C1(_07135_),
    .B1(net335),
    .A1(\top_ihp.oisc.regs[5][31] ),
    .Y(_07136_),
    .A2(net297));
 sg13g2_nand4_1 _23717_ (.B(_07127_),
    .C(_07132_),
    .A(_07126_),
    .Y(_07137_),
    .D(_07136_));
 sg13g2_and3_1 _23718_ (.X(_07138_),
    .A(\top_ihp.oisc.regs[20][31] ),
    .B(_05799_),
    .C(_05802_));
 sg13g2_a221oi_1 _23719_ (.B2(\top_ihp.oisc.regs[27][31] ),
    .C1(_07138_),
    .B1(_05820_),
    .A1(_09673_),
    .Y(_07139_),
    .A2(net720));
 sg13g2_a22oi_1 _23720_ (.Y(_07140_),
    .B1(_06002_),
    .B2(\top_ihp.oisc.regs[6][31] ),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[15][31] ));
 sg13g2_nand2b_1 _23721_ (.Y(_07141_),
    .B(_06134_),
    .A_N(_07140_));
 sg13g2_a22oi_1 _23722_ (.Y(_07142_),
    .B1(_06066_),
    .B2(\top_ihp.oisc.regs[22][31] ),
    .A2(_05510_),
    .A1(\top_ihp.oisc.regs[25][31] ));
 sg13g2_a22oi_1 _23723_ (.Y(_07143_),
    .B1(net424),
    .B2(\top_ihp.oisc.regs[10][31] ),
    .A2(net439),
    .A1(\top_ihp.oisc.regs[1][31] ));
 sg13g2_nand4_1 _23724_ (.B(_07141_),
    .C(_07142_),
    .A(_07139_),
    .Y(_07144_),
    .D(_07143_));
 sg13g2_a22oi_1 _23725_ (.Y(_07145_),
    .B1(_05901_),
    .B2(\top_ihp.oisc.regs[16][31] ),
    .A2(_06119_),
    .A1(\top_ihp.oisc.regs[28][31] ));
 sg13g2_inv_1 _23726_ (.Y(_07146_),
    .A(_07145_));
 sg13g2_a22oi_1 _23727_ (.Y(_07147_),
    .B1(_05932_),
    .B2(\top_ihp.oisc.regs[29][31] ),
    .A2(net695),
    .A1(\top_ihp.oisc.regs[30][31] ));
 sg13g2_nand2_1 _23728_ (.Y(_07148_),
    .A(\top_ihp.oisc.regs[21][31] ),
    .B(_06785_));
 sg13g2_o21ai_1 _23729_ (.B1(_07148_),
    .Y(_07149_),
    .A1(_05832_),
    .A2(_07147_));
 sg13g2_a22oi_1 _23730_ (.Y(_07150_),
    .B1(_07149_),
    .B2(net320),
    .A2(_07146_),
    .A1(_05802_));
 sg13g2_a22oi_1 _23731_ (.Y(_07151_),
    .B1(_06047_),
    .B2(\top_ihp.oisc.regs[49][31] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[42][31] ));
 sg13g2_nand2_1 _23732_ (.Y(_07152_),
    .A(_07150_),
    .B(_07151_));
 sg13g2_a22oi_1 _23733_ (.Y(_07153_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][31] ),
    .A2(net183),
    .A1(\top_ihp.oisc.regs[63][31] ));
 sg13g2_a22oi_1 _23734_ (.Y(_07154_),
    .B1(_05957_),
    .B2(\top_ihp.oisc.regs[8][31] ),
    .A2(_05744_),
    .A1(\top_ihp.oisc.regs[48][31] ));
 sg13g2_a22oi_1 _23735_ (.Y(_07155_),
    .B1(net72),
    .B2(\top_ihp.oisc.regs[53][31] ),
    .A2(net180),
    .A1(\top_ihp.oisc.regs[45][31] ));
 sg13g2_a22oi_1 _23736_ (.Y(_07156_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][31] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][31] ));
 sg13g2_nand4_1 _23737_ (.B(_07154_),
    .C(_07155_),
    .A(_07153_),
    .Y(_07157_),
    .D(_07156_));
 sg13g2_nor4_1 _23738_ (.A(_07137_),
    .B(_07144_),
    .C(_07152_),
    .D(_07157_),
    .Y(_07158_));
 sg13g2_a21oi_1 _23739_ (.A1(_00077_),
    .A2(_06506_),
    .Y(_07159_),
    .B1(_06559_));
 sg13g2_a21oi_1 _23740_ (.A1(_09673_),
    .A2(_06390_),
    .Y(_07160_),
    .B1(_07159_));
 sg13g2_a21oi_1 _23741_ (.A1(_07125_),
    .A2(_07158_),
    .Y(_00444_),
    .B1(_07160_));
 sg13g2_a22oi_1 _23742_ (.Y(_07161_),
    .B1(net288),
    .B2(\top_ihp.oisc.regs[40][3] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][3] ));
 sg13g2_a22oi_1 _23743_ (.Y(_07162_),
    .B1(net151),
    .B2(\top_ihp.oisc.regs[3][3] ),
    .A2(net603),
    .A1(\top_ihp.oisc.regs[27][3] ));
 sg13g2_a22oi_1 _23744_ (.Y(_07163_),
    .B1(net175),
    .B2(\top_ihp.oisc.regs[13][3] ),
    .A2(net720),
    .A1(_08326_));
 sg13g2_a22oi_1 _23745_ (.Y(_07164_),
    .B1(_05741_),
    .B2(\top_ihp.oisc.regs[52][3] ),
    .A2(_05525_),
    .A1(\top_ihp.oisc.regs[45][3] ));
 sg13g2_a22oi_1 _23746_ (.Y(_07165_),
    .B1(_05543_),
    .B2(\top_ihp.oisc.regs[61][3] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][3] ));
 sg13g2_and2_1 _23747_ (.A(_07164_),
    .B(_07165_),
    .X(_07166_));
 sg13g2_nand4_1 _23748_ (.B(_07162_),
    .C(_07163_),
    .A(_07161_),
    .Y(_07167_),
    .D(_07166_));
 sg13g2_a22oi_1 _23749_ (.Y(_07168_),
    .B1(_05649_),
    .B2(\top_ihp.oisc.regs[63][3] ),
    .A2(_05634_),
    .A1(\top_ihp.oisc.regs[33][3] ));
 sg13g2_a22oi_1 _23750_ (.Y(_07169_),
    .B1(net300),
    .B2(\top_ihp.oisc.regs[35][3] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][3] ));
 sg13g2_a22oi_1 _23751_ (.Y(_07170_),
    .B1(net722),
    .B2(\top_ihp.oisc.regs[29][3] ),
    .A2(net672),
    .A1(\top_ihp.oisc.regs[28][3] ));
 sg13g2_nand2_1 _23752_ (.Y(_07171_),
    .A(\top_ihp.oisc.regs[24][3] ),
    .B(_06313_));
 sg13g2_o21ai_1 _23753_ (.B1(_07171_),
    .Y(_07172_),
    .A1(_06053_),
    .A2(_07170_));
 sg13g2_a22oi_1 _23754_ (.Y(_07173_),
    .B1(_07172_),
    .B2(net415),
    .A2(net306),
    .A1(\top_ihp.oisc.regs[34][3] ));
 sg13g2_a22oi_1 _23755_ (.Y(_07174_),
    .B1(net290),
    .B2(\top_ihp.oisc.regs[19][3] ),
    .A2(net696),
    .A1(\top_ihp.oisc.regs[31][3] ));
 sg13g2_inv_1 _23756_ (.Y(_07175_),
    .A(_07174_));
 sg13g2_a22oi_1 _23757_ (.Y(_07176_),
    .B1(_07175_),
    .B2(net694),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][3] ));
 sg13g2_nand4_1 _23758_ (.B(_07169_),
    .C(_07173_),
    .A(_07168_),
    .Y(_07177_),
    .D(_07176_));
 sg13g2_a22oi_1 _23759_ (.Y(_07178_),
    .B1(net314),
    .B2(\top_ihp.oisc.regs[9][3] ),
    .A2(_05861_),
    .A1(\top_ihp.oisc.regs[20][3] ));
 sg13g2_a22oi_1 _23760_ (.Y(_07179_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][3] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][3] ));
 sg13g2_a22oi_1 _23761_ (.Y(_07180_),
    .B1(net316),
    .B2(\top_ihp.oisc.regs[25][3] ),
    .A2(net297),
    .A1(\top_ihp.oisc.regs[5][3] ));
 sg13g2_a22oi_1 _23762_ (.Y(_07181_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[14][3] ),
    .A2(net295),
    .A1(\top_ihp.oisc.regs[2][3] ));
 sg13g2_nand4_1 _23763_ (.B(_07179_),
    .C(_07180_),
    .A(_07178_),
    .Y(_07182_),
    .D(_07181_));
 sg13g2_nand2_1 _23764_ (.Y(_07183_),
    .A(\top_ihp.oisc.regs[1][3] ),
    .B(net317));
 sg13g2_nand4_1 _23765_ (.B(net420),
    .C(net699),
    .A(\top_ihp.oisc.regs[58][3] ),
    .Y(_07184_),
    .D(_06154_));
 sg13g2_a22oi_1 _23766_ (.Y(_07185_),
    .B1(net429),
    .B2(\top_ihp.oisc.regs[8][3] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][3] ));
 sg13g2_mux2_1 _23767_ (.A0(\top_ihp.oisc.regs[30][3] ),
    .A1(\top_ihp.oisc.regs[22][3] ),
    .S(_05363_),
    .X(_07186_));
 sg13g2_a22oi_1 _23768_ (.Y(_07187_),
    .B1(_07186_),
    .B2(net320),
    .A2(net699),
    .A1(\top_ihp.oisc.regs[26][3] ));
 sg13g2_nand2b_1 _23769_ (.Y(_07188_),
    .B(net695),
    .A_N(_07187_));
 sg13g2_nand4_1 _23770_ (.B(_07184_),
    .C(_07185_),
    .A(_07183_),
    .Y(_07189_),
    .D(_07188_));
 sg13g2_nor4_1 _23771_ (.A(_07167_),
    .B(_07177_),
    .C(_07182_),
    .D(_07189_),
    .Y(_07190_));
 sg13g2_mux2_1 _23772_ (.A0(\top_ihp.oisc.regs[15][3] ),
    .A1(\top_ihp.oisc.regs[11][3] ),
    .S(net598),
    .X(_07191_));
 sg13g2_nand3_1 _23773_ (.B(_05700_),
    .C(_07191_),
    .A(net415),
    .Y(_07192_));
 sg13g2_nand3_1 _23774_ (.B(net291),
    .C(_06163_),
    .A(\top_ihp.oisc.regs[23][3] ),
    .Y(_07193_));
 sg13g2_nand3_1 _23775_ (.B(_05887_),
    .C(net697),
    .A(\top_ihp.oisc.regs[17][3] ),
    .Y(_07194_));
 sg13g2_a21o_1 _23776_ (.A2(_07194_),
    .A1(_07193_),
    .B1(_05931_),
    .X(_07195_));
 sg13g2_a22oi_1 _23777_ (.Y(_07196_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][3] ),
    .A2(net338),
    .A1(\top_ihp.oisc.regs[44][3] ));
 sg13g2_nand2_1 _23778_ (.Y(_07197_),
    .A(\top_ihp.oisc.regs[6][3] ),
    .B(_05825_));
 sg13g2_a22oi_1 _23779_ (.Y(_07198_),
    .B1(_05813_),
    .B2(\top_ihp.oisc.regs[4][3] ),
    .A2(_05574_),
    .A1(\top_ihp.oisc.regs[21][3] ));
 sg13g2_a21o_1 _23780_ (.A2(_07198_),
    .A1(_07197_),
    .B1(net610),
    .X(_07199_));
 sg13g2_nand3_1 _23781_ (.B(net604),
    .C(net721),
    .A(\top_ihp.oisc.regs[18][3] ),
    .Y(_07200_));
 sg13g2_a21oi_1 _23782_ (.A1(_07199_),
    .A2(_07200_),
    .Y(_07201_),
    .B1(_05998_));
 sg13g2_a221oi_1 _23783_ (.B2(\top_ihp.oisc.regs[46][3] ),
    .C1(_07201_),
    .B1(net169),
    .A1(\top_ihp.oisc.regs[62][3] ),
    .Y(_07202_),
    .A2(net193));
 sg13g2_nand4_1 _23784_ (.B(_07195_),
    .C(_07196_),
    .A(_07192_),
    .Y(_07203_),
    .D(_07202_));
 sg13g2_a22oi_1 _23785_ (.Y(_07204_),
    .B1(_06117_),
    .B2(\top_ihp.oisc.regs[47][3] ),
    .A2(_05784_),
    .A1(\top_ihp.oisc.regs[50][3] ));
 sg13g2_a22oi_1 _23786_ (.Y(_07205_),
    .B1(net323),
    .B2(\top_ihp.oisc.regs[41][3] ),
    .A2(_05590_),
    .A1(\top_ihp.oisc.regs[57][3] ));
 sg13g2_a22oi_1 _23787_ (.Y(_07206_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][3] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][3] ));
 sg13g2_a22oi_1 _23788_ (.Y(_07207_),
    .B1(_05779_),
    .B2(\top_ihp.oisc.regs[56][3] ),
    .A2(_05748_),
    .A1(\top_ihp.oisc.regs[53][3] ));
 sg13g2_nand4_1 _23789_ (.B(_07205_),
    .C(_07206_),
    .A(_07204_),
    .Y(_07208_),
    .D(_07207_));
 sg13g2_a22oi_1 _23790_ (.Y(_07209_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][3] ),
    .A2(_06287_),
    .A1(\top_ihp.oisc.regs[42][3] ));
 sg13g2_a22oi_1 _23791_ (.Y(_07210_),
    .B1(_06294_),
    .B2(\top_ihp.oisc.regs[55][3] ),
    .A2(net339),
    .A1(\top_ihp.oisc.regs[60][3] ));
 sg13g2_a22oi_1 _23792_ (.Y(_07211_),
    .B1(_05980_),
    .B2(\top_ihp.oisc.regs[59][3] ),
    .A2(_05778_),
    .A1(\top_ihp.oisc.regs[54][3] ));
 sg13g2_a22oi_1 _23793_ (.Y(_07212_),
    .B1(_05884_),
    .B2(\top_ihp.oisc.regs[7][3] ),
    .A2(_06276_),
    .A1(\top_ihp.oisc.regs[32][3] ));
 sg13g2_nand4_1 _23794_ (.B(_07210_),
    .C(_07211_),
    .A(_07209_),
    .Y(_07213_),
    .D(_07212_));
 sg13g2_nor4_1 _23795_ (.A(net158),
    .B(_07203_),
    .C(_07208_),
    .D(_07213_),
    .Y(_07214_));
 sg13g2_a21oi_1 _23796_ (.A1(_00244_),
    .A2(net150),
    .Y(_07215_),
    .B1(net32));
 sg13g2_a21oi_1 _23797_ (.A1(_08326_),
    .A2(net719),
    .Y(_07216_),
    .B1(_07215_));
 sg13g2_a21oi_1 _23798_ (.A1(_07190_),
    .A2(_07214_),
    .Y(_00445_),
    .B1(_07216_));
 sg13g2_a22oi_1 _23799_ (.Y(_07217_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][4] ),
    .A2(net171),
    .A1(\top_ihp.oisc.regs[44][4] ));
 sg13g2_a22oi_1 _23800_ (.Y(_07218_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][4] ),
    .A2(net430),
    .A1(\top_ihp.oisc.regs[58][4] ));
 sg13g2_a22oi_1 _23801_ (.Y(_07219_),
    .B1(net308),
    .B2(\top_ihp.oisc.regs[40][4] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][4] ));
 sg13g2_a22oi_1 _23802_ (.Y(_07220_),
    .B1(net161),
    .B2(\top_ihp.oisc.regs[36][4] ),
    .A2(net181),
    .A1(\top_ihp.oisc.regs[47][4] ));
 sg13g2_nand4_1 _23803_ (.B(_07218_),
    .C(_07219_),
    .A(_07217_),
    .Y(_07221_),
    .D(_07220_));
 sg13g2_a22oi_1 _23804_ (.Y(_07222_),
    .B1(net70),
    .B2(\top_ihp.oisc.regs[45][4] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][4] ));
 sg13g2_a22oi_1 _23805_ (.Y(_07223_),
    .B1(_05747_),
    .B2(\top_ihp.oisc.regs[39][4] ),
    .A2(net162),
    .A1(\top_ihp.oisc.regs[61][4] ));
 sg13g2_a22oi_1 _23806_ (.Y(_07224_),
    .B1(_06708_),
    .B2(\top_ihp.oisc.regs[56][4] ),
    .A2(net298),
    .A1(\top_ihp.oisc.regs[48][4] ));
 sg13g2_nand2_1 _23807_ (.Y(_07225_),
    .A(_05261_),
    .B(\top_ihp.oisc.regs[62][4] ));
 sg13g2_nand2_1 _23808_ (.Y(_07226_),
    .A(\top_ihp.oisc.regs[63][4] ),
    .B(_05319_));
 sg13g2_o21ai_1 _23809_ (.B1(_07226_),
    .Y(_07227_),
    .A1(_05319_),
    .A2(_07225_));
 sg13g2_nand2_1 _23810_ (.Y(_07228_),
    .A(_06154_),
    .B(_07227_));
 sg13g2_a22oi_1 _23811_ (.Y(_07229_),
    .B1(_05813_),
    .B2(\top_ihp.oisc.regs[12][4] ),
    .A2(net672),
    .A1(\top_ihp.oisc.regs[28][4] ));
 sg13g2_nand2_1 _23812_ (.Y(_07230_),
    .A(_07228_),
    .B(_07229_));
 sg13g2_a22oi_1 _23813_ (.Y(_07231_),
    .B1(_07230_),
    .B2(net669),
    .A2(net173),
    .A1(\top_ihp.oisc.regs[53][4] ));
 sg13g2_nand4_1 _23814_ (.B(_07223_),
    .C(_07224_),
    .A(_07222_),
    .Y(_07232_),
    .D(_07231_));
 sg13g2_a22oi_1 _23815_ (.Y(_07233_),
    .B1(net295),
    .B2(\top_ihp.oisc.regs[2][4] ),
    .A2(net611),
    .A1(\top_ihp.oisc.regs[31][4] ));
 sg13g2_nand3_1 _23816_ (.B(net676),
    .C(_05850_),
    .A(\top_ihp.oisc.regs[13][4] ),
    .Y(_07234_));
 sg13g2_nand3_1 _23817_ (.B(net675),
    .C(_06317_),
    .A(\top_ihp.oisc.regs[1][4] ),
    .Y(_07235_));
 sg13g2_nand2_1 _23818_ (.Y(_07236_),
    .A(_07234_),
    .B(_07235_));
 sg13g2_a22oi_1 _23819_ (.Y(_07237_),
    .B1(_07236_),
    .B2(net414),
    .A2(_05436_),
    .A1(\top_ihp.oisc.regs[19][4] ));
 sg13g2_a22oi_1 _23820_ (.Y(_07238_),
    .B1(_06688_),
    .B2(\top_ihp.oisc.regs[29][4] ),
    .A2(_05500_),
    .A1(\top_ihp.oisc.regs[3][4] ));
 sg13g2_nand2_1 _23821_ (.Y(_07239_),
    .A(\top_ihp.oisc.regs[10][4] ),
    .B(_05995_));
 sg13g2_nand3_1 _23822_ (.B(_05404_),
    .C(_06317_),
    .A(\top_ihp.oisc.regs[9][4] ),
    .Y(_07240_));
 sg13g2_o21ai_1 _23823_ (.B1(_07240_),
    .Y(_07241_),
    .A1(_06433_),
    .A2(_07239_));
 sg13g2_a22oi_1 _23824_ (.Y(_07242_),
    .B1(_07241_),
    .B2(_05674_),
    .A2(_05839_),
    .A1(\top_ihp.oisc.regs[22][4] ));
 sg13g2_and4_1 _23825_ (.A(_07233_),
    .B(_07237_),
    .C(_07238_),
    .D(_07242_),
    .X(_07243_));
 sg13g2_mux2_1 _23826_ (.A0(\top_ihp.oisc.regs[15][4] ),
    .A1(\top_ihp.oisc.regs[14][4] ),
    .S(_05279_),
    .X(_07244_));
 sg13g2_nand3_1 _23827_ (.B(net419),
    .C(_05825_),
    .A(\top_ihp.oisc.regs[6][4] ),
    .Y(_07245_));
 sg13g2_nand3_1 _23828_ (.B(net604),
    .C(_05934_),
    .A(\top_ihp.oisc.regs[16][4] ),
    .Y(_07246_));
 sg13g2_a21oi_1 _23829_ (.A1(_07245_),
    .A2(_07246_),
    .Y(_07247_),
    .B1(net413));
 sg13g2_a221oi_1 _23830_ (.B2(_07244_),
    .C1(_07247_),
    .B1(_05376_),
    .A1(_08338_),
    .Y(_07248_),
    .A2(net720));
 sg13g2_a22oi_1 _23831_ (.Y(_07249_),
    .B1(_05975_),
    .B2(\top_ihp.oisc.regs[43][4] ),
    .A2(net429),
    .A1(\top_ihp.oisc.regs[8][4] ));
 sg13g2_a22oi_1 _23832_ (.Y(_07250_),
    .B1(_05765_),
    .B2(\top_ihp.oisc.regs[49][4] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][4] ));
 sg13g2_nand4_1 _23833_ (.B(_07248_),
    .C(_07249_),
    .A(_07243_),
    .Y(_07251_),
    .D(_07250_));
 sg13g2_mux2_1 _23834_ (.A0(\top_ihp.oisc.regs[25][4] ),
    .A1(\top_ihp.oisc.regs[17][4] ),
    .S(net681),
    .X(_07252_));
 sg13g2_nand3_1 _23835_ (.B(net697),
    .C(_07252_),
    .A(net412),
    .Y(_07253_));
 sg13g2_nand4_1 _23836_ (.B(_05956_),
    .C(_05407_),
    .A(\top_ihp.oisc.regs[11][4] ),
    .Y(_07254_),
    .D(net699));
 sg13g2_a22oi_1 _23837_ (.Y(_07255_),
    .B1(_06083_),
    .B2(\top_ihp.oisc.regs[24][4] ),
    .A2(net335),
    .A1(\top_ihp.oisc.regs[18][4] ));
 sg13g2_nand3_1 _23838_ (.B(_05359_),
    .C(_05850_),
    .A(\top_ihp.oisc.regs[4][4] ),
    .Y(_07256_));
 sg13g2_nand3_1 _23839_ (.B(_05386_),
    .C(_06020_),
    .A(\top_ihp.oisc.regs[7][4] ),
    .Y(_07257_));
 sg13g2_nand2_1 _23840_ (.Y(_07258_),
    .A(_07256_),
    .B(_07257_));
 sg13g2_nand3_1 _23841_ (.B(net676),
    .C(_05582_),
    .A(\top_ihp.oisc.regs[30][4] ),
    .Y(_07259_));
 sg13g2_nand3_1 _23842_ (.B(net675),
    .C(_05440_),
    .A(\top_ihp.oisc.regs[23][4] ),
    .Y(_07260_));
 sg13g2_a21oi_1 _23843_ (.A1(_07259_),
    .A2(_07260_),
    .Y(_07261_),
    .B1(net610));
 sg13g2_a221oi_1 _23844_ (.B2(_05889_),
    .C1(_07261_),
    .B1(_07258_),
    .A1(\top_ihp.oisc.regs[5][4] ),
    .Y(_07262_),
    .A2(_05381_));
 sg13g2_nand4_1 _23845_ (.B(_07254_),
    .C(_07255_),
    .A(_07253_),
    .Y(_07263_),
    .D(_07262_));
 sg13g2_nor3_2 _23846_ (.A(_05342_),
    .B(net704),
    .C(_05530_),
    .Y(_07264_));
 sg13g2_a22oi_1 _23847_ (.Y(_07265_),
    .B1(_07264_),
    .B2(\top_ihp.oisc.regs[26][4] ),
    .A2(_06491_),
    .A1(\top_ihp.oisc.regs[20][4] ));
 sg13g2_nor2_1 _23848_ (.A(_05568_),
    .B(_07265_),
    .Y(_07266_));
 sg13g2_a22oi_1 _23849_ (.Y(_07267_),
    .B1(_07264_),
    .B2(\top_ihp.oisc.regs[27][4] ),
    .A2(_06491_),
    .A1(\top_ihp.oisc.regs[21][4] ));
 sg13g2_nor2b_1 _23850_ (.A(_07267_),
    .B_N(net742),
    .Y(_07268_));
 sg13g2_or3_1 _23851_ (.A(_07263_),
    .B(_07266_),
    .C(_07268_),
    .X(_07269_));
 sg13g2_nor4_1 _23852_ (.A(_07221_),
    .B(_07232_),
    .C(_07251_),
    .D(_07269_),
    .Y(_07270_));
 sg13g2_a22oi_1 _23853_ (.Y(_07271_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][4] ),
    .A2(net166),
    .A1(\top_ihp.oisc.regs[33][4] ));
 sg13g2_nand2_1 _23854_ (.Y(_07272_),
    .A(\top_ihp.oisc.regs[52][4] ),
    .B(net311));
 sg13g2_nand2_1 _23855_ (.Y(_07273_),
    .A(_07271_),
    .B(_07272_));
 sg13g2_a22oi_1 _23856_ (.Y(_07274_),
    .B1(net66),
    .B2(\top_ihp.oisc.regs[46][4] ),
    .A2(net68),
    .A1(\top_ihp.oisc.regs[55][4] ));
 sg13g2_a22oi_1 _23857_ (.Y(_07275_),
    .B1(_05600_),
    .B2(\top_ihp.oisc.regs[41][4] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[42][4] ));
 sg13g2_a22oi_1 _23858_ (.Y(_07276_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[50][4] ),
    .A2(net179),
    .A1(\top_ihp.oisc.regs[54][4] ));
 sg13g2_nor2_1 _23859_ (.A(net614),
    .B(net668),
    .Y(_07277_));
 sg13g2_a22oi_1 _23860_ (.Y(_07278_),
    .B1(_07277_),
    .B2(\top_ihp.oisc.regs[35][4] ),
    .A2(_06182_),
    .A1(\top_ihp.oisc.regs[32][4] ));
 sg13g2_nor3_1 _23861_ (.A(_05331_),
    .B(net702),
    .C(_07278_),
    .Y(_07279_));
 sg13g2_a21oi_1 _23862_ (.A1(\top_ihp.oisc.regs[57][4] ),
    .A2(net432),
    .Y(_07280_),
    .B1(_07279_));
 sg13g2_nand4_1 _23863_ (.B(_07275_),
    .C(_07276_),
    .A(_07274_),
    .Y(_07281_),
    .D(_07280_));
 sg13g2_nor3_1 _23864_ (.A(net159),
    .B(_07273_),
    .C(_07281_),
    .Y(_07282_));
 sg13g2_a21oi_1 _23865_ (.A1(_00245_),
    .A2(net150),
    .Y(_07283_),
    .B1(net32));
 sg13g2_a21oi_1 _23866_ (.A1(_08338_),
    .A2(net719),
    .Y(_07284_),
    .B1(_07283_));
 sg13g2_a21oi_1 _23867_ (.A1(_07270_),
    .A2(_07282_),
    .Y(_00446_),
    .B1(_07284_));
 sg13g2_a22oi_1 _23868_ (.Y(_07285_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][5] ),
    .A2(net309),
    .A1(\top_ihp.oisc.regs[56][5] ));
 sg13g2_a22oi_1 _23869_ (.Y(_07286_),
    .B1(net184),
    .B2(\top_ihp.oisc.regs[51][5] ),
    .A2(net191),
    .A1(\top_ihp.oisc.regs[42][5] ));
 sg13g2_a22oi_1 _23870_ (.Y(_07287_),
    .B1(net157),
    .B2(\top_ihp.oisc.regs[38][5] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][5] ));
 sg13g2_a22oi_1 _23871_ (.Y(_07288_),
    .B1(_05700_),
    .B2(\top_ihp.oisc.regs[7][5] ),
    .A2(net694),
    .A1(\top_ihp.oisc.regs[23][5] ));
 sg13g2_nor2_1 _23872_ (.A(_05335_),
    .B(_07288_),
    .Y(_07289_));
 sg13g2_a21oi_1 _23873_ (.A1(\top_ihp.oisc.regs[48][5] ),
    .A2(_06113_),
    .Y(_07290_),
    .B1(_07289_));
 sg13g2_nand4_1 _23874_ (.B(_07286_),
    .C(_07287_),
    .A(_07285_),
    .Y(_07291_),
    .D(_07290_));
 sg13g2_a22oi_1 _23875_ (.Y(_07292_),
    .B1(_06383_),
    .B2(\top_ihp.oisc.regs[46][5] ),
    .A2(net153),
    .A1(\top_ihp.oisc.regs[34][5] ));
 sg13g2_a22oi_1 _23876_ (.Y(_07293_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[50][5] ),
    .A2(_05666_),
    .A1(\top_ihp.oisc.regs[54][5] ));
 sg13g2_nand3_1 _23877_ (.B(_07292_),
    .C(_07293_),
    .A(_05918_),
    .Y(_07294_));
 sg13g2_nor2_1 _23878_ (.A(_07291_),
    .B(_07294_),
    .Y(_07295_));
 sg13g2_a22oi_1 _23879_ (.Y(_07296_),
    .B1(_05556_),
    .B2(\top_ihp.oisc.regs[1][5] ),
    .A2(_05462_),
    .A1(\top_ihp.oisc.regs[4][5] ));
 sg13g2_nor2_1 _23880_ (.A(_06869_),
    .B(_07296_),
    .Y(_07297_));
 sg13g2_a21oi_1 _23881_ (.A1(\top_ihp.oisc.regs[63][5] ),
    .A2(_05648_),
    .Y(_07298_),
    .B1(_07297_));
 sg13g2_a22oi_1 _23882_ (.Y(_07299_),
    .B1(_05442_),
    .B2(\top_ihp.oisc.regs[9][5] ),
    .A2(net421),
    .A1(\top_ihp.oisc.regs[5][5] ));
 sg13g2_inv_1 _23883_ (.Y(_07300_),
    .A(_07299_));
 sg13g2_a22oi_1 _23884_ (.Y(_07301_),
    .B1(_07300_),
    .B2(_05895_),
    .A2(_06047_),
    .A1(\top_ihp.oisc.regs[49][5] ));
 sg13g2_a22oi_1 _23885_ (.Y(_07302_),
    .B1(_05644_),
    .B2(\top_ihp.oisc.regs[35][5] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][5] ));
 sg13g2_a22oi_1 _23886_ (.Y(_07303_),
    .B1(_05748_),
    .B2(\top_ihp.oisc.regs[53][5] ),
    .A2(_05831_),
    .A1(\top_ihp.oisc.regs[61][5] ));
 sg13g2_nand4_1 _23887_ (.B(_07301_),
    .C(_07302_),
    .A(_07298_),
    .Y(_07304_),
    .D(_07303_));
 sg13g2_a22oi_1 _23888_ (.Y(_07305_),
    .B1(_06117_),
    .B2(\top_ihp.oisc.regs[47][5] ),
    .A2(net155),
    .A1(\top_ihp.oisc.regs[39][5] ));
 sg13g2_a22oi_1 _23889_ (.Y(_07306_),
    .B1(_05768_),
    .B2(\top_ihp.oisc.regs[36][5] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][5] ));
 sg13g2_a22oi_1 _23890_ (.Y(_07307_),
    .B1(net328),
    .B2(\top_ihp.oisc.regs[33][5] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][5] ));
 sg13g2_a22oi_1 _23891_ (.Y(_07308_),
    .B1(net430),
    .B2(\top_ihp.oisc.regs[58][5] ),
    .A2(net165),
    .A1(\top_ihp.oisc.regs[45][5] ));
 sg13g2_nand4_1 _23892_ (.B(_07306_),
    .C(_07307_),
    .A(_07305_),
    .Y(_07309_),
    .D(_07308_));
 sg13g2_mux2_1 _23893_ (.A0(\top_ihp.oisc.regs[11][5] ),
    .A1(\top_ihp.oisc.regs[3][5] ),
    .S(net704),
    .X(_07310_));
 sg13g2_nand2_1 _23894_ (.Y(_07311_),
    .A(net596),
    .B(_07310_));
 sg13g2_nand3_1 _23895_ (.B(_05548_),
    .C(_07264_),
    .A(\top_ihp.oisc.regs[59][5] ),
    .Y(_07312_));
 sg13g2_a21oi_1 _23896_ (.A1(_07311_),
    .A2(_07312_),
    .Y(_07313_),
    .B1(net420));
 sg13g2_mux2_1 _23897_ (.A0(\top_ihp.oisc.regs[14][5] ),
    .A1(\top_ihp.oisc.regs[10][5] ),
    .S(net677),
    .X(_07314_));
 sg13g2_and3_1 _23898_ (.X(_07315_),
    .A(net410),
    .B(_05407_),
    .C(_07314_));
 sg13g2_nand3_1 _23899_ (.B(net607),
    .C(net722),
    .A(\top_ihp.oisc.regs[25][5] ),
    .Y(_07316_));
 sg13g2_nand3_1 _23900_ (.B(net674),
    .C(_05871_),
    .A(\top_ihp.oisc.regs[19][5] ),
    .Y(_07317_));
 sg13g2_a21oi_1 _23901_ (.A1(_07316_),
    .A2(_07317_),
    .Y(_07318_),
    .B1(net320));
 sg13g2_nand3_1 _23902_ (.B(_05342_),
    .C(_05440_),
    .A(\top_ihp.oisc.regs[31][5] ),
    .Y(_07319_));
 sg13g2_nand3_1 _23903_ (.B(net677),
    .C(net721),
    .A(\top_ihp.oisc.regs[26][5] ),
    .Y(_07320_));
 sg13g2_a21oi_1 _23904_ (.A1(_07319_),
    .A2(_07320_),
    .Y(_07321_),
    .B1(_05678_));
 sg13g2_a21o_1 _23905_ (.A2(net335),
    .A1(\top_ihp.oisc.regs[18][5] ),
    .B1(_07321_),
    .X(_07322_));
 sg13g2_nor4_1 _23906_ (.A(_07313_),
    .B(_07315_),
    .C(_07318_),
    .D(_07322_),
    .Y(_07323_));
 sg13g2_a22oi_1 _23907_ (.Y(_07324_),
    .B1(net722),
    .B2(\top_ihp.oisc.regs[29][5] ),
    .A2(net721),
    .A1(\top_ihp.oisc.regs[30][5] ));
 sg13g2_nand2_1 _23908_ (.Y(_07325_),
    .A(_08341_),
    .B(_03714_));
 sg13g2_o21ai_1 _23909_ (.B1(_07325_),
    .Y(_07326_),
    .A1(_05317_),
    .A2(_07324_));
 sg13g2_a22oi_1 _23910_ (.Y(_07327_),
    .B1(_05575_),
    .B2(\top_ihp.oisc.regs[17][5] ),
    .A2(_05570_),
    .A1(\top_ihp.oisc.regs[16][5] ));
 sg13g2_nand3_1 _23911_ (.B(net421),
    .C(_05934_),
    .A(\top_ihp.oisc.regs[20][5] ),
    .Y(_07328_));
 sg13g2_o21ai_1 _23912_ (.B1(_07328_),
    .Y(_07329_),
    .A1(_05417_),
    .A2(_07327_));
 sg13g2_a22oi_1 _23913_ (.Y(_07330_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][5] ),
    .A2(_05444_),
    .A1(\top_ihp.oisc.regs[27][5] ));
 sg13g2_inv_1 _23914_ (.Y(_07331_),
    .A(_07330_));
 sg13g2_nor3_1 _23915_ (.A(_07326_),
    .B(_07329_),
    .C(_07331_),
    .Y(_07332_));
 sg13g2_a22oi_1 _23916_ (.Y(_07333_),
    .B1(_05814_),
    .B2(\top_ihp.oisc.regs[8][5] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[12][5] ));
 sg13g2_mux2_1 _23917_ (.A0(\top_ihp.oisc.regs[6][5] ),
    .A1(\top_ihp.oisc.regs[2][5] ),
    .S(net598),
    .X(_07334_));
 sg13g2_and2_1 _23918_ (.A(net595),
    .B(_05825_),
    .X(_07335_));
 sg13g2_a22oi_1 _23919_ (.Y(_07336_),
    .B1(_07334_),
    .B2(_07335_),
    .A2(_05863_),
    .A1(\top_ihp.oisc.regs[21][5] ));
 sg13g2_nand4_1 _23920_ (.B(_07332_),
    .C(_07333_),
    .A(_07323_),
    .Y(_07337_),
    .D(_07336_));
 sg13g2_a22oi_1 _23921_ (.Y(_07338_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][5] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][5] ));
 sg13g2_a22oi_1 _23922_ (.Y(_07339_),
    .B1(net288),
    .B2(\top_ihp.oisc.regs[40][5] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][5] ));
 sg13g2_a22oi_1 _23923_ (.Y(_07340_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][5] ),
    .A2(net75),
    .A1(\top_ihp.oisc.regs[62][5] ));
 sg13g2_a22oi_1 _23924_ (.Y(_07341_),
    .B1(_05895_),
    .B2(\top_ihp.oisc.regs[13][5] ),
    .A2(net672),
    .A1(\top_ihp.oisc.regs[28][5] ));
 sg13g2_nand2_1 _23925_ (.Y(_07342_),
    .A(\top_ihp.oisc.regs[24][5] ),
    .B(_06313_));
 sg13g2_o21ai_1 _23926_ (.B1(_07342_),
    .Y(_07343_),
    .A1(net412),
    .A2(_07341_));
 sg13g2_a22oi_1 _23927_ (.Y(_07344_),
    .B1(_07343_),
    .B2(net415),
    .A2(_05959_),
    .A1(\top_ihp.oisc.regs[15][5] ));
 sg13g2_nand4_1 _23928_ (.B(_07339_),
    .C(_07340_),
    .A(_07338_),
    .Y(_07345_),
    .D(_07344_));
 sg13g2_nor4_1 _23929_ (.A(_07304_),
    .B(_07309_),
    .C(_07337_),
    .D(_07345_),
    .Y(_07346_));
 sg13g2_a21o_1 _23930_ (.A2(_05945_),
    .A1(_00246_),
    .B1(net33),
    .X(_07347_));
 sg13g2_a22oi_1 _23931_ (.Y(_00447_),
    .B1(_07347_),
    .B2(_07325_),
    .A2(_07346_),
    .A1(_07295_));
 sg13g2_a22oi_1 _23932_ (.Y(_07348_),
    .B1(net317),
    .B2(\top_ihp.oisc.regs[1][6] ),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][6] ));
 sg13g2_a22oi_1 _23933_ (.Y(_07349_),
    .B1(net315),
    .B2(\top_ihp.oisc.regs[15][6] ),
    .A2(_06138_),
    .A1(\top_ihp.oisc.regs[23][6] ));
 sg13g2_and3_1 _23934_ (.X(_07350_),
    .A(\top_ihp.oisc.regs[33][6] ),
    .B(net414),
    .C(_06004_));
 sg13g2_nand3_1 _23935_ (.B(_06003_),
    .C(net724),
    .A(\top_ihp.oisc.regs[30][6] ),
    .Y(_07351_));
 sg13g2_nand3_1 _23936_ (.B(net668),
    .C(net742),
    .A(\top_ihp.oisc.regs[29][6] ),
    .Y(_07352_));
 sg13g2_nand2_1 _23937_ (.Y(_07353_),
    .A(_07351_),
    .B(_07352_));
 sg13g2_a22oi_1 _23938_ (.Y(_07354_),
    .B1(_07353_),
    .B2(_06119_),
    .A2(_07350_),
    .A1(_06429_));
 sg13g2_a22oi_1 _23939_ (.Y(_07355_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][6] ),
    .A2(net445),
    .A1(\top_ihp.oisc.regs[19][6] ));
 sg13g2_nand4_1 _23940_ (.B(_07349_),
    .C(_07354_),
    .A(_07348_),
    .Y(_07356_),
    .D(_07355_));
 sg13g2_a22oi_1 _23941_ (.Y(_07357_),
    .B1(net312),
    .B2(\top_ihp.oisc.regs[10][6] ),
    .A2(net437),
    .A1(\top_ihp.oisc.regs[31][6] ));
 sg13g2_a22oi_1 _23942_ (.Y(_07358_),
    .B1(net314),
    .B2(\top_ihp.oisc.regs[9][6] ),
    .A2(_05861_),
    .A1(\top_ihp.oisc.regs[20][6] ));
 sg13g2_and2_1 _23943_ (.A(\top_ihp.oisc.regs[27][6] ),
    .B(net742),
    .X(_07359_));
 sg13g2_a22oi_1 _23944_ (.Y(_07360_),
    .B1(_07264_),
    .B2(_07359_),
    .A2(net296),
    .A1(\top_ihp.oisc.regs[28][6] ));
 sg13g2_a22oi_1 _23945_ (.Y(_07361_),
    .B1(net600),
    .B2(\top_ihp.oisc.regs[12][6] ),
    .A2(net670),
    .A1(\top_ihp.oisc.regs[14][6] ));
 sg13g2_nor2b_1 _23946_ (.A(_07361_),
    .B_N(net410),
    .Y(_07362_));
 sg13g2_a221oi_1 _23947_ (.B2(\top_ihp.oisc.regs[3][6] ),
    .C1(_07362_),
    .B1(_05501_),
    .A1(_08345_),
    .Y(_07363_),
    .A2(_03715_));
 sg13g2_nand4_1 _23948_ (.B(_07358_),
    .C(_07360_),
    .A(_07357_),
    .Y(_07364_),
    .D(_07363_));
 sg13g2_a22oi_1 _23949_ (.Y(_07365_),
    .B1(net189),
    .B2(\top_ihp.oisc.regs[50][6] ),
    .A2(net74),
    .A1(\top_ihp.oisc.regs[37][6] ));
 sg13g2_a22oi_1 _23950_ (.Y(_07366_),
    .B1(net304),
    .B2(\top_ihp.oisc.regs[58][6] ),
    .A2(net279),
    .A1(\top_ihp.oisc.regs[42][6] ));
 sg13g2_a22oi_1 _23951_ (.Y(_07367_),
    .B1(net170),
    .B2(\top_ihp.oisc.regs[36][6] ),
    .A2(net77),
    .A1(\top_ihp.oisc.regs[55][6] ));
 sg13g2_a22oi_1 _23952_ (.Y(_07368_),
    .B1(_06002_),
    .B2(\top_ihp.oisc.regs[4][6] ),
    .A2(net601),
    .A1(\top_ihp.oisc.regs[13][6] ));
 sg13g2_inv_1 _23953_ (.Y(_07369_),
    .A(_07368_));
 sg13g2_a22oi_1 _23954_ (.Y(_07370_),
    .B1(_07369_),
    .B2(_05851_),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][6] ));
 sg13g2_nand4_1 _23955_ (.B(_07366_),
    .C(_07367_),
    .A(_07365_),
    .Y(_07371_),
    .D(_07370_));
 sg13g2_mux2_1 _23956_ (.A0(\top_ihp.oisc.regs[21][6] ),
    .A1(\top_ihp.oisc.regs[17][6] ),
    .S(net418),
    .X(_07372_));
 sg13g2_a22oi_1 _23957_ (.Y(_07373_),
    .B1(_07372_),
    .B2(_05890_),
    .A2(_05810_),
    .A1(\top_ihp.oisc.regs[25][6] ));
 sg13g2_mux2_1 _23958_ (.A0(\top_ihp.oisc.regs[22][6] ),
    .A1(\top_ihp.oisc.regs[18][6] ),
    .S(_05564_),
    .X(_07374_));
 sg13g2_a22oi_1 _23959_ (.Y(_07375_),
    .B1(_07374_),
    .B2(net595),
    .A2(net699),
    .A1(\top_ihp.oisc.regs[26][6] ));
 sg13g2_inv_1 _23960_ (.Y(_07376_),
    .A(_07375_));
 sg13g2_a22oi_1 _23961_ (.Y(_07377_),
    .B1(net451),
    .B2(\top_ihp.oisc.regs[7][6] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][6] ));
 sg13g2_mux2_1 _23962_ (.A0(\top_ihp.oisc.regs[24][6] ),
    .A1(\top_ihp.oisc.regs[16][6] ),
    .S(net675),
    .X(_07378_));
 sg13g2_nand4_1 _23963_ (.B(_06260_),
    .C(net724),
    .A(_05887_),
    .Y(_07379_),
    .D(_07378_));
 sg13g2_nor2_1 _23964_ (.A(net681),
    .B(_05331_),
    .Y(_07380_));
 sg13g2_nand4_1 _23965_ (.B(net598),
    .C(_06182_),
    .A(\top_ihp.oisc.regs[40][6] ),
    .Y(_07381_),
    .D(_07380_));
 sg13g2_nand3_1 _23966_ (.B(_07379_),
    .C(_07381_),
    .A(_07377_),
    .Y(_07382_));
 sg13g2_a21oi_1 _23967_ (.A1(net695),
    .A2(_07376_),
    .Y(_07383_),
    .B1(_07382_));
 sg13g2_o21ai_1 _23968_ (.B1(_07383_),
    .Y(_07384_),
    .A1(net734),
    .A2(_07373_));
 sg13g2_nor4_1 _23969_ (.A(_07356_),
    .B(_07364_),
    .C(_07371_),
    .D(_07384_),
    .Y(_07385_));
 sg13g2_a22oi_1 _23970_ (.Y(_07386_),
    .B1(_07277_),
    .B2(\top_ihp.oisc.regs[11][6] ),
    .A2(_06182_),
    .A1(\top_ihp.oisc.regs[8][6] ));
 sg13g2_nor3_1 _23971_ (.A(_05915_),
    .B(net679),
    .C(_07386_),
    .Y(_07387_));
 sg13g2_a21oi_1 _23972_ (.A1(\top_ihp.oisc.regs[46][6] ),
    .A2(net169),
    .Y(_07388_),
    .B1(_07387_));
 sg13g2_a22oi_1 _23973_ (.Y(_07389_),
    .B1(net180),
    .B2(\top_ihp.oisc.regs[45][6] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][6] ));
 sg13g2_a22oi_1 _23974_ (.Y(_07390_),
    .B1(net78),
    .B2(\top_ihp.oisc.regs[59][6] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][6] ));
 sg13g2_a22oi_1 _23975_ (.Y(_07391_),
    .B1(net422),
    .B2(\top_ihp.oisc.regs[57][6] ),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][6] ));
 sg13g2_nand4_1 _23976_ (.B(_07389_),
    .C(_07390_),
    .A(_07388_),
    .Y(_07392_),
    .D(_07391_));
 sg13g2_a22oi_1 _23977_ (.Y(_07393_),
    .B1(net307),
    .B2(\top_ihp.oisc.regs[34][6] ),
    .A2(_05645_),
    .A1(\top_ihp.oisc.regs[35][6] ));
 sg13g2_a22oi_1 _23978_ (.Y(_07394_),
    .B1(_05786_),
    .B2(\top_ihp.oisc.regs[53][6] ),
    .A2(net155),
    .A1(\top_ihp.oisc.regs[39][6] ));
 sg13g2_a22oi_1 _23979_ (.Y(_07395_),
    .B1(net75),
    .B2(\top_ihp.oisc.regs[62][6] ),
    .A2(net187),
    .A1(\top_ihp.oisc.regs[38][6] ));
 sg13g2_a22oi_1 _23980_ (.Y(_07396_),
    .B1(net431),
    .B2(\top_ihp.oisc.regs[41][6] ),
    .A2(_05532_),
    .A1(\top_ihp.oisc.regs[52][6] ));
 sg13g2_nand4_1 _23981_ (.B(_07394_),
    .C(_07395_),
    .A(_07393_),
    .Y(_07397_),
    .D(_07396_));
 sg13g2_a22oi_1 _23982_ (.Y(_07398_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][6] ),
    .A2(net183),
    .A1(\top_ihp.oisc.regs[63][6] ));
 sg13g2_a22oi_1 _23983_ (.Y(_07399_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][6] ),
    .A2(net305),
    .A1(\top_ihp.oisc.regs[51][6] ));
 sg13g2_a22oi_1 _23984_ (.Y(_07400_),
    .B1(net284),
    .B2(\top_ihp.oisc.regs[48][6] ),
    .A2(net188),
    .A1(\top_ihp.oisc.regs[61][6] ));
 sg13g2_a22oi_1 _23985_ (.Y(_07401_),
    .B1(_05328_),
    .B2(\top_ihp.oisc.regs[44][6] ),
    .A2(_06108_),
    .A1(\top_ihp.oisc.regs[60][6] ));
 sg13g2_nand4_1 _23986_ (.B(_07399_),
    .C(_07400_),
    .A(_07398_),
    .Y(_07402_),
    .D(_07401_));
 sg13g2_nor4_1 _23987_ (.A(net158),
    .B(_07392_),
    .C(_07397_),
    .D(_07402_),
    .Y(_07403_));
 sg13g2_a21oi_1 _23988_ (.A1(_00247_),
    .A2(net331),
    .Y(_07404_),
    .B1(net32));
 sg13g2_a21oi_1 _23989_ (.A1(_08345_),
    .A2(net719),
    .Y(_07405_),
    .B1(_07404_));
 sg13g2_a21oi_1 _23990_ (.A1(_07385_),
    .A2(_07403_),
    .Y(_00448_),
    .B1(_07405_));
 sg13g2_mux2_1 _23991_ (.A0(\top_ihp.oisc.regs[29][7] ),
    .A1(\top_ihp.oisc.regs[21][7] ),
    .S(net674),
    .X(_07406_));
 sg13g2_nand2_1 _23992_ (.Y(_07407_),
    .A(\top_ihp.oisc.regs[44][7] ),
    .B(net696));
 sg13g2_nand2_1 _23993_ (.Y(_07408_),
    .A(\top_ihp.oisc.regs[15][7] ),
    .B(_05719_));
 sg13g2_o21ai_1 _23994_ (.B1(_07408_),
    .Y(_07409_),
    .A1(_05325_),
    .A2(_07407_));
 sg13g2_a221oi_1 _23995_ (.B2(_07406_),
    .C1(_07409_),
    .B1(_05807_),
    .A1(\top_ihp.oisc.regs[8][7] ),
    .Y(_07410_),
    .A2(_05683_));
 sg13g2_a22oi_1 _23996_ (.Y(_07411_),
    .B1(net319),
    .B2(\top_ihp.oisc.regs[17][7] ),
    .A2(net447),
    .A1(\top_ihp.oisc.regs[9][7] ));
 sg13g2_a22oi_1 _23997_ (.Y(_07412_),
    .B1(_06308_),
    .B2(\top_ihp.oisc.regs[22][7] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[4][7] ));
 sg13g2_a22oi_1 _23998_ (.Y(_07413_),
    .B1(_05402_),
    .B2(\top_ihp.oisc.regs[13][7] ),
    .A2(_05396_),
    .A1(\top_ihp.oisc.regs[12][7] ));
 sg13g2_a22oi_1 _23999_ (.Y(_07414_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[25][7] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[6][7] ));
 sg13g2_a22oi_1 _24000_ (.Y(_07415_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][7] ),
    .A2(_05389_),
    .A1(\top_ihp.oisc.regs[20][7] ));
 sg13g2_nand3_1 _24001_ (.B(_05359_),
    .C(_05995_),
    .A(\top_ihp.oisc.regs[2][7] ),
    .Y(_07416_));
 sg13g2_nand3_1 _24002_ (.B(_05386_),
    .C(_06020_),
    .A(\top_ihp.oisc.regs[7][7] ),
    .Y(_07417_));
 sg13g2_nand2_1 _24003_ (.Y(_07418_),
    .A(_07416_),
    .B(_07417_));
 sg13g2_a22oi_1 _24004_ (.Y(_07419_),
    .B1(_07418_),
    .B2(net606),
    .A2(_05817_),
    .A1(\top_ihp.oisc.regs[30][7] ));
 sg13g2_and4_1 _24005_ (.A(_07413_),
    .B(_07414_),
    .C(_07415_),
    .D(_07419_),
    .X(_07420_));
 sg13g2_nand4_1 _24006_ (.B(_07411_),
    .C(_07412_),
    .A(_07410_),
    .Y(_07421_),
    .D(_07420_));
 sg13g2_a22oi_1 _24007_ (.Y(_07422_),
    .B1(_06354_),
    .B2(\top_ihp.oisc.regs[3][7] ),
    .A2(_05710_),
    .A1(\top_ihp.oisc.regs[27][7] ));
 sg13g2_a22oi_1 _24008_ (.Y(_07423_),
    .B1(net437),
    .B2(\top_ihp.oisc.regs[31][7] ),
    .A2(net296),
    .A1(\top_ihp.oisc.regs[28][7] ));
 sg13g2_mux2_1 _24009_ (.A0(\top_ihp.oisc.regs[5][7] ),
    .A1(\top_ihp.oisc.regs[1][7] ),
    .S(net677),
    .X(_07424_));
 sg13g2_nand3_1 _24010_ (.B(_05895_),
    .C(_07424_),
    .A(net599),
    .Y(_07425_));
 sg13g2_nand2_1 _24011_ (.Y(_07426_),
    .A(\top_ihp.oisc.regs[10][7] ),
    .B(_05728_));
 sg13g2_nand2_1 _24012_ (.Y(_07427_),
    .A(_07425_),
    .B(_07426_));
 sg13g2_a221oi_1 _24013_ (.B2(\top_ihp.oisc.regs[26][7] ),
    .C1(_07427_),
    .B1(net333),
    .A1(\top_ihp.oisc.regs[19][7] ),
    .Y(_07428_),
    .A2(_05437_));
 sg13g2_a22oi_1 _24014_ (.Y(_07429_),
    .B1(_05645_),
    .B2(\top_ihp.oisc.regs[35][7] ),
    .A2(net192),
    .A1(\top_ihp.oisc.regs[37][7] ));
 sg13g2_nand4_1 _24015_ (.B(_07423_),
    .C(_07428_),
    .A(_07422_),
    .Y(_07430_),
    .D(_07429_));
 sg13g2_a22oi_1 _24016_ (.Y(_07431_),
    .B1(net67),
    .B2(\top_ihp.oisc.regs[61][7] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][7] ));
 sg13g2_a22oi_1 _24017_ (.Y(_07432_),
    .B1(net305),
    .B2(\top_ihp.oisc.regs[51][7] ),
    .A2(net170),
    .A1(\top_ihp.oisc.regs[36][7] ));
 sg13g2_a22oi_1 _24018_ (.Y(_07433_),
    .B1(net169),
    .B2(\top_ihp.oisc.regs[46][7] ),
    .A2(net285),
    .A1(\top_ihp.oisc.regs[60][7] ));
 sg13g2_a22oi_1 _24019_ (.Y(_07434_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][7] ),
    .A2(net324),
    .A1(\top_ihp.oisc.regs[63][7] ));
 sg13g2_nand4_1 _24020_ (.B(_07432_),
    .C(_07433_),
    .A(_07431_),
    .Y(_07435_),
    .D(_07434_));
 sg13g2_a22oi_1 _24021_ (.Y(_07436_),
    .B1(net71),
    .B2(\top_ihp.oisc.regs[59][7] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][7] ));
 sg13g2_a22oi_1 _24022_ (.Y(_07437_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][7] ),
    .A2(net168),
    .A1(\top_ihp.oisc.regs[54][7] ));
 sg13g2_a22oi_1 _24023_ (.Y(_07438_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][7] ),
    .A2(net304),
    .A1(\top_ihp.oisc.regs[58][7] ));
 sg13g2_a22oi_1 _24024_ (.Y(_07439_),
    .B1(_05646_),
    .B2(\top_ihp.oisc.regs[57][7] ),
    .A2(net307),
    .A1(\top_ihp.oisc.regs[34][7] ));
 sg13g2_nand4_1 _24025_ (.B(_07437_),
    .C(_07438_),
    .A(_07436_),
    .Y(_07440_),
    .D(_07439_));
 sg13g2_nor4_1 _24026_ (.A(_07421_),
    .B(_07430_),
    .C(_07435_),
    .D(_07440_),
    .Y(_07441_));
 sg13g2_a22oi_1 _24027_ (.Y(_07442_),
    .B1(net166),
    .B2(\top_ihp.oisc.regs[33][7] ),
    .A2(net334),
    .A1(\top_ihp.oisc.regs[42][7] ));
 sg13g2_a22oi_1 _24028_ (.Y(_07443_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][7] ),
    .A2(net435),
    .A1(\top_ihp.oisc.regs[40][7] ));
 sg13g2_a22oi_1 _24029_ (.Y(_07444_),
    .B1(net173),
    .B2(\top_ihp.oisc.regs[53][7] ),
    .A2(_05795_),
    .A1(\top_ihp.oisc.regs[45][7] ));
 sg13g2_a22oi_1 _24030_ (.Y(_07445_),
    .B1(net75),
    .B2(\top_ihp.oisc.regs[62][7] ),
    .A2(net441),
    .A1(\top_ihp.oisc.regs[49][7] ));
 sg13g2_nand4_1 _24031_ (.B(_07443_),
    .C(_07444_),
    .A(_07442_),
    .Y(_07446_),
    .D(_07445_));
 sg13g2_nand2_1 _24032_ (.Y(_07447_),
    .A(\top_ihp.oisc.regs[48][7] ),
    .B(_06113_));
 sg13g2_a22oi_1 _24033_ (.Y(_07448_),
    .B1(net176),
    .B2(\top_ihp.oisc.regs[18][7] ),
    .A2(net728),
    .A1(_08314_));
 sg13g2_a22oi_1 _24034_ (.Y(_07449_),
    .B1(net318),
    .B2(\top_ihp.oisc.regs[11][7] ),
    .A2(net177),
    .A1(\top_ihp.oisc.regs[16][7] ));
 sg13g2_a22oi_1 _24035_ (.Y(_07450_),
    .B1(net282),
    .B2(\top_ihp.oisc.regs[24][7] ),
    .A2(net423),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_nand4_1 _24036_ (.B(_07448_),
    .C(_07449_),
    .A(_07447_),
    .Y(_07451_),
    .D(_07450_));
 sg13g2_a22oi_1 _24037_ (.Y(_07452_),
    .B1(_06235_),
    .B2(\top_ihp.oisc.regs[39][7] ),
    .A2(_05774_),
    .A1(\top_ihp.oisc.regs[32][7] ));
 sg13g2_a22oi_1 _24038_ (.Y(_07453_),
    .B1(net68),
    .B2(\top_ihp.oisc.regs[55][7] ),
    .A2(_05628_),
    .A1(\top_ihp.oisc.regs[50][7] ));
 sg13g2_nand2_1 _24039_ (.Y(_07454_),
    .A(_07452_),
    .B(_07453_));
 sg13g2_nor4_1 _24040_ (.A(_05616_),
    .B(_07446_),
    .C(_07451_),
    .D(_07454_),
    .Y(_07455_));
 sg13g2_a21oi_1 _24041_ (.A1(_00248_),
    .A2(net331),
    .Y(_07456_),
    .B1(_05622_));
 sg13g2_a21oi_1 _24042_ (.A1(_08314_),
    .A2(net719),
    .Y(_07457_),
    .B1(_07456_));
 sg13g2_a21oi_1 _24043_ (.A1(_07441_),
    .A2(_07455_),
    .Y(_00449_),
    .B1(_07457_));
 sg13g2_a22oi_1 _24044_ (.Y(_07458_),
    .B1(net74),
    .B2(\top_ihp.oisc.regs[37][8] ),
    .A2(net327),
    .A1(\top_ihp.oisc.regs[49][8] ));
 sg13g2_a22oi_1 _24045_ (.Y(_07459_),
    .B1(net325),
    .B2(\top_ihp.oisc.regs[35][8] ),
    .A2(_05633_),
    .A1(\top_ihp.oisc.regs[33][8] ));
 sg13g2_a22oi_1 _24046_ (.Y(_07460_),
    .B1(_05762_),
    .B2(\top_ihp.oisc.regs[58][8] ),
    .A2(net182),
    .A1(\top_ihp.oisc.regs[55][8] ));
 sg13g2_a22oi_1 _24047_ (.Y(_07461_),
    .B1(net167),
    .B2(\top_ihp.oisc.regs[50][8] ),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][8] ));
 sg13g2_nand4_1 _24048_ (.B(_07459_),
    .C(_07460_),
    .A(_07458_),
    .Y(_07462_),
    .D(_07461_));
 sg13g2_a22oi_1 _24049_ (.Y(_07463_),
    .B1(_05786_),
    .B2(\top_ihp.oisc.regs[53][8] ),
    .A2(net446),
    .A1(\top_ihp.oisc.regs[32][8] ));
 sg13g2_a22oi_1 _24050_ (.Y(_07464_),
    .B1(net301),
    .B2(\top_ihp.oisc.regs[56][8] ),
    .A2(net326),
    .A1(\top_ihp.oisc.regs[51][8] ));
 sg13g2_a22oi_1 _24051_ (.Y(_07465_),
    .B1(_05741_),
    .B2(\top_ihp.oisc.regs[52][8] ),
    .A2(net324),
    .A1(\top_ihp.oisc.regs[63][8] ));
 sg13g2_a22oi_1 _24052_ (.Y(_07466_),
    .B1(net290),
    .B2(\top_ihp.oisc.regs[18][8] ),
    .A2(net669),
    .A1(\top_ihp.oisc.regs[30][8] ));
 sg13g2_inv_1 _24053_ (.Y(_07467_),
    .A(_07466_));
 sg13g2_a22oi_1 _24054_ (.Y(_07468_),
    .B1(_06160_),
    .B2(_07467_),
    .A2(net452),
    .A1(\top_ihp.oisc.regs[60][8] ));
 sg13g2_nand4_1 _24055_ (.B(_07464_),
    .C(_07465_),
    .A(_07463_),
    .Y(_07469_),
    .D(_07468_));
 sg13g2_a22oi_1 _24056_ (.Y(_07470_),
    .B1(net439),
    .B2(\top_ihp.oisc.regs[1][8] ),
    .A2(_05436_),
    .A1(\top_ihp.oisc.regs[19][8] ));
 sg13g2_a22oi_1 _24057_ (.Y(_07471_),
    .B1(_06688_),
    .B2(\top_ihp.oisc.regs[29][8] ),
    .A2(net428),
    .A1(\top_ihp.oisc.regs[17][8] ));
 sg13g2_a22oi_1 _24058_ (.Y(_07472_),
    .B1(net426),
    .B2(\top_ihp.oisc.regs[25][8] ),
    .A2(net442),
    .A1(\top_ihp.oisc.regs[28][8] ));
 sg13g2_a22oi_1 _24059_ (.Y(_07473_),
    .B1(_05734_),
    .B2(\top_ihp.oisc.regs[14][8] ),
    .A2(_05450_),
    .A1(\top_ihp.oisc.regs[21][8] ));
 sg13g2_and4_1 _24060_ (.A(_07470_),
    .B(_07471_),
    .C(_07472_),
    .D(_07473_),
    .X(_07474_));
 sg13g2_nand2_1 _24061_ (.Y(_07475_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(_05688_));
 sg13g2_nand3_1 _24062_ (.B(net291),
    .C(_06163_),
    .A(\top_ihp.oisc.regs[31][8] ),
    .Y(_07476_));
 sg13g2_nand3_1 _24063_ (.B(net598),
    .C(_06160_),
    .A(\top_ihp.oisc.regs[26][8] ),
    .Y(_07477_));
 sg13g2_nand2_1 _24064_ (.Y(_07478_),
    .A(_07476_),
    .B(_07477_));
 sg13g2_a22oi_1 _24065_ (.Y(_07479_),
    .B1(_07478_),
    .B2(_05931_),
    .A2(net282),
    .A1(\top_ihp.oisc.regs[24][8] ));
 sg13g2_nand3_1 _24066_ (.B(_07475_),
    .C(_07479_),
    .A(_07474_),
    .Y(_07480_));
 sg13g2_a22oi_1 _24067_ (.Y(_07481_),
    .B1(net191),
    .B2(\top_ihp.oisc.regs[42][8] ),
    .A2(net195),
    .A1(\top_ihp.oisc.regs[44][8] ));
 sg13g2_a22oi_1 _24068_ (.Y(_07482_),
    .B1(net153),
    .B2(\top_ihp.oisc.regs[34][8] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][8] ));
 sg13g2_a22oi_1 _24069_ (.Y(_07483_),
    .B1(_05729_),
    .B2(\top_ihp.oisc.regs[10][8] ),
    .A2(net336),
    .A1(\top_ihp.oisc.regs[13][8] ));
 sg13g2_a22oi_1 _24070_ (.Y(_07484_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][8] ),
    .A2(_06070_),
    .A1(\top_ihp.oisc.regs[8][8] ));
 sg13g2_and2_1 _24071_ (.A(_07483_),
    .B(_07484_),
    .X(_07485_));
 sg13g2_nand2_1 _24072_ (.Y(_07486_),
    .A(\top_ihp.oisc.regs[16][8] ),
    .B(net672));
 sg13g2_nand2_1 _24073_ (.Y(_07487_),
    .A(_08350_),
    .B(net748));
 sg13g2_o21ai_1 _24074_ (.B1(_07487_),
    .Y(_07488_),
    .A1(net702),
    .A2(_07486_));
 sg13g2_a221oi_1 _24075_ (.B2(\top_ihp.oisc.regs[59][8] ),
    .C1(_07488_),
    .B1(net185),
    .A1(\top_ihp.oisc.regs[20][8] ),
    .Y(_07489_),
    .A2(net449));
 sg13g2_nand4_1 _24076_ (.B(_07482_),
    .C(_07485_),
    .A(_07481_),
    .Y(_07490_),
    .D(_07489_));
 sg13g2_nor4_1 _24077_ (.A(_07462_),
    .B(_07469_),
    .C(_07480_),
    .D(_07490_),
    .Y(_07491_));
 sg13g2_a22oi_1 _24078_ (.Y(_07492_),
    .B1(net76),
    .B2(\top_ihp.oisc.regs[47][8] ),
    .A2(net70),
    .A1(\top_ihp.oisc.regs[45][8] ));
 sg13g2_a22oi_1 _24079_ (.Y(_07493_),
    .B1(net303),
    .B2(\top_ihp.oisc.regs[41][8] ),
    .A2(net169),
    .A1(\top_ihp.oisc.regs[46][8] ));
 sg13g2_a22oi_1 _24080_ (.Y(_07494_),
    .B1(net67),
    .B2(\top_ihp.oisc.regs[61][8] ),
    .A2(net299),
    .A1(\top_ihp.oisc.regs[43][8] ));
 sg13g2_a22oi_1 _24081_ (.Y(_07495_),
    .B1(net156),
    .B2(\top_ihp.oisc.regs[36][8] ),
    .A2(net194),
    .A1(\top_ihp.oisc.regs[38][8] ));
 sg13g2_nand4_1 _24082_ (.B(_07493_),
    .C(_07494_),
    .A(_07492_),
    .Y(_07496_),
    .D(_07495_));
 sg13g2_a22oi_1 _24083_ (.Y(_07497_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][8] ),
    .A2(net288),
    .A1(\top_ihp.oisc.regs[40][8] ));
 sg13g2_a22oi_1 _24084_ (.Y(_07498_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][8] ),
    .A2(net284),
    .A1(\top_ihp.oisc.regs[48][8] ));
 sg13g2_nand2_1 _24085_ (.Y(_07499_),
    .A(_07497_),
    .B(_07498_));
 sg13g2_nand2_1 _24086_ (.Y(_07500_),
    .A(\top_ihp.oisc.regs[3][8] ),
    .B(net151));
 sg13g2_a22oi_1 _24087_ (.Y(_07501_),
    .B1(net163),
    .B2(\top_ihp.oisc.regs[2][8] ),
    .A2(net292),
    .A1(\top_ihp.oisc.regs[6][8] ));
 sg13g2_a22oi_1 _24088_ (.Y(_07502_),
    .B1(net447),
    .B2(\top_ihp.oisc.regs[9][8] ),
    .A2(net448),
    .A1(\top_ihp.oisc.regs[12][8] ));
 sg13g2_a22oi_1 _24089_ (.Y(_07503_),
    .B1(_05719_),
    .B2(\top_ihp.oisc.regs[15][8] ),
    .A2(_05444_),
    .A1(\top_ihp.oisc.regs[27][8] ));
 sg13g2_a22oi_1 _24090_ (.Y(_07504_),
    .B1(net451),
    .B2(\top_ihp.oisc.regs[7][8] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][8] ));
 sg13g2_a22oi_1 _24091_ (.Y(_07505_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][8] ),
    .A2(net436),
    .A1(\top_ihp.oisc.regs[4][8] ));
 sg13g2_and4_1 _24092_ (.A(_07502_),
    .B(_07503_),
    .C(_07504_),
    .D(_07505_),
    .X(_07506_));
 sg13g2_nand4_1 _24093_ (.B(_07500_),
    .C(_07501_),
    .A(_05918_),
    .Y(_07507_),
    .D(_07506_));
 sg13g2_nor3_1 _24094_ (.A(_07496_),
    .B(_07499_),
    .C(_07507_),
    .Y(_07508_));
 sg13g2_a21o_1 _24095_ (.A2(_05626_),
    .A1(_00249_),
    .B1(_05946_),
    .X(_07509_));
 sg13g2_a22oi_1 _24096_ (.Y(_00450_),
    .B1(_07509_),
    .B2(_07487_),
    .A2(_07508_),
    .A1(_07491_));
 sg13g2_a22oi_1 _24097_ (.Y(_07510_),
    .B1(_05655_),
    .B2(\top_ihp.oisc.regs[41][9] ),
    .A2(net280),
    .A1(\top_ihp.oisc.regs[32][9] ));
 sg13g2_a22oi_1 _24098_ (.Y(_07511_),
    .B1(net77),
    .B2(\top_ihp.oisc.regs[55][9] ),
    .A2(net321),
    .A1(\top_ihp.oisc.regs[54][9] ));
 sg13g2_a22oi_1 _24099_ (.Y(_07512_),
    .B1(net325),
    .B2(\top_ihp.oisc.regs[35][9] ),
    .A2(_05636_),
    .A1(\top_ihp.oisc.regs[59][9] ));
 sg13g2_a22oi_1 _24100_ (.Y(_07513_),
    .B1(net160),
    .B2(\top_ihp.oisc.regs[63][9] ),
    .A2(net328),
    .A1(\top_ihp.oisc.regs[33][9] ));
 sg13g2_nand4_1 _24101_ (.B(_07511_),
    .C(_07512_),
    .A(_07510_),
    .Y(_07514_),
    .D(_07513_));
 sg13g2_a22oi_1 _24102_ (.Y(_07515_),
    .B1(net289),
    .B2(\top_ihp.oisc.regs[52][9] ),
    .A2(_05771_),
    .A1(\top_ihp.oisc.regs[46][9] ));
 sg13g2_a22oi_1 _24103_ (.Y(_07516_),
    .B1(_05744_),
    .B2(\top_ihp.oisc.regs[48][9] ),
    .A2(_05485_),
    .A1(\top_ihp.oisc.regs[42][9] ));
 sg13g2_a22oi_1 _24104_ (.Y(_07517_),
    .B1(net188),
    .B2(\top_ihp.oisc.regs[61][9] ),
    .A2(net167),
    .A1(\top_ihp.oisc.regs[50][9] ));
 sg13g2_a22oi_1 _24105_ (.Y(_07518_),
    .B1(net410),
    .B2(\top_ihp.oisc.regs[10][9] ),
    .A2(_06017_),
    .A1(\top_ihp.oisc.regs[3][9] ));
 sg13g2_inv_1 _24106_ (.Y(_07519_),
    .A(_07518_));
 sg13g2_a22oi_1 _24107_ (.Y(_07520_),
    .B1(_07519_),
    .B2(net596),
    .A2(_05641_),
    .A1(\top_ihp.oisc.regs[51][9] ));
 sg13g2_nand4_1 _24108_ (.B(_07516_),
    .C(_07517_),
    .A(_07515_),
    .Y(_07521_),
    .D(_07520_));
 sg13g2_a22oi_1 _24109_ (.Y(_07522_),
    .B1(net438),
    .B2(\top_ihp.oisc.regs[23][9] ),
    .A2(_05488_),
    .A1(\top_ihp.oisc.regs[1][9] ));
 sg13g2_a22oi_1 _24110_ (.Y(_07523_),
    .B1(_05863_),
    .B2(\top_ihp.oisc.regs[21][9] ),
    .A2(_05414_),
    .A1(\top_ihp.oisc.regs[9][9] ));
 sg13g2_a22oi_1 _24111_ (.Y(_07524_),
    .B1(net442),
    .B2(\top_ihp.oisc.regs[28][9] ),
    .A2(net443),
    .A1(\top_ihp.oisc.regs[11][9] ));
 sg13g2_a22oi_1 _24112_ (.Y(_07525_),
    .B1(net335),
    .B2(\top_ihp.oisc.regs[18][9] ),
    .A2(_06070_),
    .A1(\top_ihp.oisc.regs[8][9] ));
 sg13g2_and4_1 _24113_ (.A(_07522_),
    .B(_07523_),
    .C(_07524_),
    .D(_07525_),
    .X(_07526_));
 sg13g2_nand3_1 _24114_ (.B(net291),
    .C(_05879_),
    .A(\top_ihp.oisc.regs[30][9] ),
    .Y(_07527_));
 sg13g2_nand3_1 _24115_ (.B(net418),
    .C(_06429_),
    .A(\top_ihp.oisc.regs[16][9] ),
    .Y(_07528_));
 sg13g2_a21o_1 _24116_ (.A2(_07528_),
    .A1(_07527_),
    .B1(_05568_),
    .X(_07529_));
 sg13g2_a22oi_1 _24117_ (.Y(_07530_),
    .B1(net427),
    .B2(\top_ihp.oisc.regs[19][9] ),
    .A2(net313),
    .A1(\top_ihp.oisc.regs[12][9] ));
 sg13g2_nand3_1 _24118_ (.B(net671),
    .C(net724),
    .A(\top_ihp.oisc.regs[26][9] ),
    .Y(_07531_));
 sg13g2_nand3_1 _24119_ (.B(net668),
    .C(net742),
    .A(\top_ihp.oisc.regs[25][9] ),
    .Y(_07532_));
 sg13g2_nand2_1 _24120_ (.Y(_07533_),
    .A(_07531_),
    .B(_07532_));
 sg13g2_a22oi_1 _24121_ (.Y(_07534_),
    .B1(_07533_),
    .B2(_05810_),
    .A2(_05859_),
    .A1(\top_ihp.oisc.regs[4][9] ));
 sg13g2_nand4_1 _24122_ (.B(_07529_),
    .C(_07530_),
    .A(_07526_),
    .Y(_07535_),
    .D(_07534_));
 sg13g2_a22oi_1 _24123_ (.Y(_07536_),
    .B1(_05736_),
    .B2(\top_ihp.oisc.regs[24][9] ),
    .A2(_05390_),
    .A1(\top_ihp.oisc.regs[20][9] ));
 sg13g2_a22oi_1 _24124_ (.Y(_07537_),
    .B1(net423),
    .B2(\top_ihp.oisc.regs[14][9] ),
    .A2(net425),
    .A1(\top_ihp.oisc.regs[29][9] ));
 sg13g2_a22oi_1 _24125_ (.Y(_07538_),
    .B1(_05839_),
    .B2(\top_ihp.oisc.regs[22][9] ),
    .A2(net450),
    .A1(\top_ihp.oisc.regs[6][9] ));
 sg13g2_a22oi_1 _24126_ (.Y(_07539_),
    .B1(_05691_),
    .B2(\top_ihp.oisc.regs[2][9] ),
    .A2(net337),
    .A1(\top_ihp.oisc.regs[5][9] ));
 sg13g2_and4_1 _24127_ (.A(_07536_),
    .B(_07537_),
    .C(_07538_),
    .D(_07539_),
    .X(_07540_));
 sg13g2_a22oi_1 _24128_ (.Y(_07541_),
    .B1(net309),
    .B2(\top_ihp.oisc.regs[56][9] ),
    .A2(_05640_),
    .A1(\top_ihp.oisc.regs[49][9] ));
 sg13g2_nand2_1 _24129_ (.Y(_07542_),
    .A(\top_ihp.oisc.regs[34][9] ),
    .B(_06148_));
 sg13g2_and3_1 _24130_ (.X(_07543_),
    .A(\top_ihp.oisc.regs[15][9] ),
    .B(net597),
    .C(net601));
 sg13g2_a221oi_1 _24131_ (.B2(\top_ihp.oisc.regs[7][9] ),
    .C1(_07543_),
    .B1(net281),
    .A1(_08353_),
    .Y(_07544_),
    .A2(net720));
 sg13g2_nand4_1 _24132_ (.B(_07541_),
    .C(_07542_),
    .A(_07540_),
    .Y(_07545_),
    .D(_07544_));
 sg13g2_nor4_1 _24133_ (.A(_07514_),
    .B(_07521_),
    .C(_07535_),
    .D(_07545_),
    .Y(_07546_));
 sg13g2_a22oi_1 _24134_ (.Y(_07547_),
    .B1(net69),
    .B2(\top_ihp.oisc.regs[39][9] ),
    .A2(net157),
    .A1(\top_ihp.oisc.regs[38][9] ));
 sg13g2_a22oi_1 _24135_ (.Y(_07548_),
    .B1(net70),
    .B2(\top_ihp.oisc.regs[45][9] ),
    .A2(net287),
    .A1(\top_ihp.oisc.regs[43][9] ));
 sg13g2_a22oi_1 _24136_ (.Y(_07549_),
    .B1(net432),
    .B2(\top_ihp.oisc.regs[57][9] ),
    .A2(_05311_),
    .A1(\top_ihp.oisc.regs[60][9] ));
 sg13g2_nand3_1 _24137_ (.B(net604),
    .C(net697),
    .A(\top_ihp.oisc.regs[17][9] ),
    .Y(_07550_));
 sg13g2_nand4_1 _24138_ (.B(_05956_),
    .C(net608),
    .A(\top_ihp.oisc.regs[13][9] ),
    .Y(_07551_),
    .D(net600));
 sg13g2_o21ai_1 _24139_ (.B1(_07551_),
    .Y(_07552_),
    .A1(net413),
    .A2(_07550_));
 sg13g2_a21oi_1 _24140_ (.A1(\top_ihp.oisc.regs[40][9] ),
    .A2(net288),
    .Y(_07553_),
    .B1(_07552_));
 sg13g2_nand4_1 _24141_ (.B(_07548_),
    .C(_07549_),
    .A(_07547_),
    .Y(_07554_),
    .D(_07553_));
 sg13g2_nand2_1 _24142_ (.Y(_07555_),
    .A(\top_ihp.oisc.regs[47][9] ),
    .B(net76));
 sg13g2_a22oi_1 _24143_ (.Y(_07556_),
    .B1(net73),
    .B2(\top_ihp.oisc.regs[53][9] ),
    .A2(net74),
    .A1(\top_ihp.oisc.regs[37][9] ));
 sg13g2_a22oi_1 _24144_ (.Y(_07557_),
    .B1(net322),
    .B2(\top_ihp.oisc.regs[58][9] ),
    .A2(net65),
    .A1(\top_ihp.oisc.regs[62][9] ));
 sg13g2_nand3_1 _24145_ (.B(net419),
    .C(net698),
    .A(\top_ihp.oisc.regs[31][9] ),
    .Y(_07558_));
 sg13g2_nand3_1 _24146_ (.B(net604),
    .C(net698),
    .A(\top_ihp.oisc.regs[27][9] ),
    .Y(_07559_));
 sg13g2_a21oi_2 _24147_ (.B1(net417),
    .Y(_07560_),
    .A2(_07559_),
    .A1(_07558_));
 sg13g2_a221oi_1 _24148_ (.B2(\top_ihp.oisc.regs[36][9] ),
    .C1(_07560_),
    .B1(net161),
    .A1(\top_ihp.oisc.regs[44][9] ),
    .Y(_07561_),
    .A2(net338));
 sg13g2_nand4_1 _24149_ (.B(_07556_),
    .C(_07557_),
    .A(_07555_),
    .Y(_07562_),
    .D(_07561_));
 sg13g2_nor3_1 _24150_ (.A(net159),
    .B(_07554_),
    .C(_07562_),
    .Y(_07563_));
 sg13g2_a21oi_1 _24151_ (.A1(_00250_),
    .A2(net331),
    .Y(_07564_),
    .B1(_05622_));
 sg13g2_a21oi_1 _24152_ (.A1(_08353_),
    .A2(net719),
    .Y(_07565_),
    .B1(_07564_));
 sg13g2_a21oi_1 _24153_ (.A1(_07546_),
    .A2(_07563_),
    .Y(_00451_),
    .B1(_07565_));
 sg13g2_nor3_1 _24154_ (.A(net1020),
    .B(_08989_),
    .C(\top_ihp.oisc.reg_rb[3] ),
    .Y(_07566_));
 sg13g2_buf_2 _24155_ (.A(_07566_),
    .X(_07567_));
 sg13g2_buf_1 _24156_ (.A(_07567_),
    .X(_07568_));
 sg13g2_buf_2 _24157_ (.A(_08997_),
    .X(_07569_));
 sg13g2_buf_1 _24158_ (.A(_07569_),
    .X(_07570_));
 sg13g2_buf_1 _24159_ (.A(net810),
    .X(_07571_));
 sg13g2_buf_1 _24160_ (.A(net776),
    .X(_07572_));
 sg13g2_mux2_1 _24161_ (.A0(\top_ihp.oisc.regs[5][0] ),
    .A1(\top_ihp.oisc.regs[1][0] ),
    .S(net758),
    .X(_07573_));
 sg13g2_nor2_1 _24162_ (.A(_08989_),
    .B(\top_ihp.oisc.reg_rb[3] ),
    .Y(_07574_));
 sg13g2_and2_1 _24163_ (.A(net1020),
    .B(_07574_),
    .X(_07575_));
 sg13g2_buf_2 _24164_ (.A(_07575_),
    .X(_07576_));
 sg13g2_buf_1 _24165_ (.A(_07576_),
    .X(_07577_));
 sg13g2_mux2_1 _24166_ (.A0(\top_ihp.oisc.regs[7][0] ),
    .A1(\top_ihp.oisc.regs[3][0] ),
    .S(net758),
    .X(_07578_));
 sg13g2_nor3_2 _24167_ (.A(\top_ihp.oisc.micro_op[11] ),
    .B(_08988_),
    .C(_08991_),
    .Y(_07579_));
 sg13g2_and2_1 _24168_ (.A(net1020),
    .B(_07579_),
    .X(_07580_));
 sg13g2_buf_1 _24169_ (.A(_07580_),
    .X(_07581_));
 sg13g2_buf_1 _24170_ (.A(net865),
    .X(_07582_));
 sg13g2_buf_1 _24171_ (.A(_07569_),
    .X(_07583_));
 sg13g2_mux2_1 _24172_ (.A0(\top_ihp.oisc.regs[6][0] ),
    .A1(\top_ihp.oisc.regs[2][0] ),
    .S(net808),
    .X(_07584_));
 sg13g2_nand2_1 _24173_ (.Y(_07585_),
    .A(net853),
    .B(_07584_));
 sg13g2_nand3_1 _24174_ (.B(\top_ihp.oisc.reg_rb[0] ),
    .C(\top_ihp.oisc.reg_rb[3] ),
    .A(net1020),
    .Y(_07586_));
 sg13g2_nor2_1 _24175_ (.A(_09141_),
    .B(_07586_),
    .Y(_07587_));
 sg13g2_buf_1 _24176_ (.A(_07587_),
    .X(_07588_));
 sg13g2_buf_1 _24177_ (.A(_07588_),
    .X(_07589_));
 sg13g2_buf_1 _24178_ (.A(net775),
    .X(_07590_));
 sg13g2_nand2_1 _24179_ (.Y(_07591_),
    .A(\top_ihp.oisc.regs[15][0] ),
    .B(net757));
 sg13g2_nor4_2 _24180_ (.A(\top_ihp.oisc.reg_rb[1] ),
    .B(\top_ihp.oisc.reg_rb[0] ),
    .C(\top_ihp.oisc.reg_rb[3] ),
    .Y(_07592_),
    .D(_08997_));
 sg13g2_buf_1 _24181_ (.A(_07592_),
    .X(_07593_));
 sg13g2_buf_1 _24182_ (.A(_07593_),
    .X(_07594_));
 sg13g2_nor4_2 _24183_ (.A(_08990_),
    .B(_08988_),
    .C(_08984_),
    .Y(_07595_),
    .D(_08991_));
 sg13g2_buf_2 _24184_ (.A(_07595_),
    .X(_07596_));
 sg13g2_and2_1 _24185_ (.A(net1041),
    .B(_07596_),
    .X(_07597_));
 sg13g2_buf_1 _24186_ (.A(_07597_),
    .X(_07598_));
 sg13g2_buf_1 _24187_ (.A(_07598_),
    .X(_07599_));
 sg13g2_nand2_1 _24188_ (.Y(_07600_),
    .A(\top_ihp.oisc.regs[12][0] ),
    .B(net838));
 sg13g2_nor2_2 _24189_ (.A(_08211_),
    .B(_08987_),
    .Y(_07601_));
 sg13g2_buf_1 _24190_ (.A(_07601_),
    .X(_07602_));
 sg13g2_and4_1 _24191_ (.A(\top_ihp.oisc.micro_op[11] ),
    .B(_09569_),
    .C(_08984_),
    .D(_08987_),
    .X(_07603_));
 sg13g2_buf_1 _24192_ (.A(_07603_),
    .X(_07604_));
 sg13g2_and2_1 _24193_ (.A(_09141_),
    .B(_07604_),
    .X(_07605_));
 sg13g2_buf_1 _24194_ (.A(_07605_),
    .X(_07606_));
 sg13g2_a22oi_1 _24195_ (.Y(_07607_),
    .B1(_07606_),
    .B2(\top_ihp.oisc.regs[10][0] ),
    .A2(net837),
    .A1(\top_ihp.oisc.regs[32][0] ));
 sg13g2_and2_1 _24196_ (.A(net1041),
    .B(_07604_),
    .X(_07608_));
 sg13g2_buf_2 _24197_ (.A(_07608_),
    .X(_07609_));
 sg13g2_nor2_1 _24198_ (.A(net1041),
    .B(net1020),
    .Y(_07610_));
 sg13g2_and2_1 _24199_ (.A(_07579_),
    .B(_07610_),
    .X(_07611_));
 sg13g2_buf_1 _24200_ (.A(_07611_),
    .X(_07612_));
 sg13g2_a22oi_1 _24201_ (.Y(_07613_),
    .B1(_07612_),
    .B2(\top_ihp.oisc.regs[0][0] ),
    .A2(_07609_),
    .A1(\top_ihp.oisc.regs[14][0] ));
 sg13g2_nand2_1 _24202_ (.Y(_07614_),
    .A(\top_ihp.oisc.reg_rb[0] ),
    .B(\top_ihp.oisc.reg_rb[3] ));
 sg13g2_nor2b_1 _24203_ (.A(_07614_),
    .B_N(_07610_),
    .Y(_07615_));
 sg13g2_buf_1 _24204_ (.A(_07615_),
    .X(_07616_));
 sg13g2_nor3_1 _24205_ (.A(_09141_),
    .B(net1020),
    .C(_07614_),
    .Y(_07617_));
 sg13g2_buf_1 _24206_ (.A(_07617_),
    .X(_07618_));
 sg13g2_a22oi_1 _24207_ (.Y(_07619_),
    .B1(_07618_),
    .B2(\top_ihp.oisc.regs[13][0] ),
    .A2(_07616_),
    .A1(\top_ihp.oisc.regs[9][0] ));
 sg13g2_nand4_1 _24208_ (.B(_07607_),
    .C(_07613_),
    .A(_07600_),
    .Y(_07620_),
    .D(_07619_));
 sg13g2_a21oi_1 _24209_ (.A1(\top_ihp.oisc.regs[4][0] ),
    .A2(net774),
    .Y(_07621_),
    .B1(_07620_));
 sg13g2_nor2_1 _24210_ (.A(net1041),
    .B(_07586_),
    .Y(_07622_));
 sg13g2_buf_1 _24211_ (.A(_07622_),
    .X(_07623_));
 sg13g2_buf_1 _24212_ (.A(_07623_),
    .X(_07624_));
 sg13g2_buf_1 _24213_ (.A(net773),
    .X(_07625_));
 sg13g2_and2_1 _24214_ (.A(_09141_),
    .B(_07596_),
    .X(_07626_));
 sg13g2_buf_1 _24215_ (.A(_07626_),
    .X(_07627_));
 sg13g2_buf_1 _24216_ (.A(net852),
    .X(_07628_));
 sg13g2_a22oi_1 _24217_ (.Y(_07629_),
    .B1(net836),
    .B2(\top_ihp.oisc.regs[8][0] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][0] ));
 sg13g2_nand4_1 _24218_ (.B(_07591_),
    .C(_07621_),
    .A(_07585_),
    .Y(_07630_),
    .D(_07629_));
 sg13g2_a221oi_1 _24219_ (.B2(_07578_),
    .C1(_07630_),
    .B1(net809),
    .A1(net839),
    .Y(_07631_),
    .A2(_07573_));
 sg13g2_nand2_1 _24220_ (.Y(_07632_),
    .A(net890),
    .B(_08991_));
 sg13g2_buf_4 _24221_ (.X(_07633_),
    .A(_07632_));
 sg13g2_o21ai_1 _24222_ (.B1(_07633_),
    .Y(_07634_),
    .A1(net982),
    .A2(net793));
 sg13g2_buf_1 _24223_ (.A(_07634_),
    .X(_07635_));
 sg13g2_buf_1 _24224_ (.A(net741),
    .X(_07636_));
 sg13g2_buf_1 _24225_ (.A(net719),
    .X(_07637_));
 sg13g2_nand2_1 _24226_ (.Y(_07638_),
    .A(_08320_),
    .B(net667));
 sg13g2_o21ai_1 _24227_ (.B1(_07638_),
    .Y(_00452_),
    .A1(_07631_),
    .A2(net733));
 sg13g2_buf_1 _24228_ (.A(_07569_),
    .X(_07639_));
 sg13g2_buf_1 _24229_ (.A(net807),
    .X(_07640_));
 sg13g2_mux2_1 _24230_ (.A0(\top_ihp.oisc.regs[7][10] ),
    .A1(\top_ihp.oisc.regs[3][10] ),
    .S(net772),
    .X(_07641_));
 sg13g2_buf_1 _24231_ (.A(net1041),
    .X(_07642_));
 sg13g2_buf_1 _24232_ (.A(net985),
    .X(_07643_));
 sg13g2_a22oi_1 _24233_ (.Y(_07644_),
    .B1(_07604_),
    .B2(\top_ihp.oisc.regs[10][10] ),
    .A2(_07596_),
    .A1(\top_ihp.oisc.regs[8][10] ));
 sg13g2_or2_1 _24234_ (.X(_07645_),
    .B(_07644_),
    .A(net935));
 sg13g2_buf_1 _24235_ (.A(_07616_),
    .X(_07646_));
 sg13g2_and2_1 _24236_ (.A(\top_ihp.oisc.regs[14][10] ),
    .B(_07609_),
    .X(_07647_));
 sg13g2_a221oi_1 _24237_ (.B2(\top_ihp.oisc.regs[9][10] ),
    .C1(_07647_),
    .B1(net771),
    .A1(\top_ihp.oisc.regs[32][10] ),
    .Y(_07648_),
    .A2(net837));
 sg13g2_buf_1 _24238_ (.A(_07618_),
    .X(_07649_));
 sg13g2_nand2_1 _24239_ (.Y(_07650_),
    .A(_07579_),
    .B(_07610_));
 sg13g2_buf_2 _24240_ (.A(_07650_),
    .X(_07651_));
 sg13g2_nor2_1 _24241_ (.A(_00251_),
    .B(_07651_),
    .Y(_07652_));
 sg13g2_a221oi_1 _24242_ (.B2(\top_ihp.oisc.regs[13][10] ),
    .C1(_07652_),
    .B1(net770),
    .A1(\top_ihp.oisc.regs[11][10] ),
    .Y(_07653_),
    .A2(net773));
 sg13g2_a22oi_1 _24243_ (.Y(_07654_),
    .B1(net775),
    .B2(\top_ihp.oisc.regs[15][10] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[12][10] ));
 sg13g2_nand4_1 _24244_ (.B(_07648_),
    .C(_07653_),
    .A(_07645_),
    .Y(_07655_),
    .D(_07654_));
 sg13g2_a21oi_1 _24245_ (.A1(net809),
    .A2(_07641_),
    .Y(_07656_),
    .B1(_07655_));
 sg13g2_buf_1 _24246_ (.A(_07593_),
    .X(_07657_));
 sg13g2_and2_1 _24247_ (.A(_07569_),
    .B(_07567_),
    .X(_07658_));
 sg13g2_buf_1 _24248_ (.A(_07658_),
    .X(_07659_));
 sg13g2_a22oi_1 _24249_ (.Y(_07660_),
    .B1(_07567_),
    .B2(\top_ihp.oisc.regs[5][10] ),
    .A2(net865),
    .A1(\top_ihp.oisc.regs[6][10] ));
 sg13g2_nand2_1 _24250_ (.Y(_07661_),
    .A(_08985_),
    .B(_07579_));
 sg13g2_buf_2 _24251_ (.A(_07661_),
    .X(_07662_));
 sg13g2_nor2_2 _24252_ (.A(_08999_),
    .B(_07662_),
    .Y(_07663_));
 sg13g2_nand2_1 _24253_ (.Y(_07664_),
    .A(\top_ihp.oisc.regs[2][10] ),
    .B(_07663_));
 sg13g2_o21ai_1 _24254_ (.B1(_07664_),
    .Y(_07665_),
    .A1(net772),
    .A2(_07660_));
 sg13g2_a221oi_1 _24255_ (.B2(\top_ihp.oisc.regs[1][10] ),
    .C1(_07665_),
    .B1(_07659_),
    .A1(\top_ihp.oisc.regs[4][10] ),
    .Y(_07666_),
    .A2(net769));
 sg13g2_a21oi_1 _24256_ (.A1(_07656_),
    .A2(_07666_),
    .Y(_07667_),
    .B1(net741));
 sg13g2_a21o_1 _24257_ (.A2(net667),
    .A1(_08263_),
    .B1(_07667_),
    .X(_00453_));
 sg13g2_nand2_1 _24258_ (.Y(_07668_),
    .A(\top_ihp.oisc.regs[2][11] ),
    .B(net772));
 sg13g2_nand2_1 _24259_ (.Y(_07669_),
    .A(\top_ihp.oisc.regs[6][11] ),
    .B(net794));
 sg13g2_a21oi_1 _24260_ (.A1(_07668_),
    .A2(_07669_),
    .Y(_07670_),
    .B1(_07662_));
 sg13g2_buf_1 _24261_ (.A(_07576_),
    .X(_07671_));
 sg13g2_a22oi_1 _24262_ (.Y(_07672_),
    .B1(net806),
    .B2(\top_ihp.oisc.regs[7][11] ),
    .A2(_07567_),
    .A1(\top_ihp.oisc.regs[5][11] ));
 sg13g2_buf_1 _24263_ (.A(_07602_),
    .X(_07673_));
 sg13g2_buf_1 _24264_ (.A(_07651_),
    .X(_07674_));
 sg13g2_nor2_1 _24265_ (.A(_00252_),
    .B(net851),
    .Y(_07675_));
 sg13g2_a221oi_1 _24266_ (.B2(\top_ihp.oisc.regs[13][11] ),
    .C1(_07675_),
    .B1(net770),
    .A1(\top_ihp.oisc.regs[32][11] ),
    .Y(_07676_),
    .A2(net805));
 sg13g2_o21ai_1 _24267_ (.B1(_07676_),
    .Y(_07677_),
    .A1(net758),
    .A2(_07672_));
 sg13g2_buf_1 _24268_ (.A(net773),
    .X(_07678_));
 sg13g2_nand2_1 _24269_ (.Y(_07679_),
    .A(\top_ihp.oisc.regs[11][11] ),
    .B(net755));
 sg13g2_buf_1 _24270_ (.A(_07616_),
    .X(_07680_));
 sg13g2_buf_1 _24271_ (.A(_07606_),
    .X(_07681_));
 sg13g2_buf_1 _24272_ (.A(net804),
    .X(_07682_));
 sg13g2_a22oi_1 _24273_ (.Y(_07683_),
    .B1(net767),
    .B2(\top_ihp.oisc.regs[10][11] ),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][11] ));
 sg13g2_buf_1 _24274_ (.A(net775),
    .X(_07684_));
 sg13g2_a22oi_1 _24275_ (.Y(_07685_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][11] ),
    .A2(net836),
    .A1(\top_ihp.oisc.regs[8][11] ));
 sg13g2_nand3_1 _24276_ (.B(_07683_),
    .C(_07685_),
    .A(_07679_),
    .Y(_07686_));
 sg13g2_nand2_1 _24277_ (.Y(_07687_),
    .A(_08985_),
    .B(_07574_));
 sg13g2_buf_2 _24278_ (.A(_07687_),
    .X(_07688_));
 sg13g2_nor2_2 _24279_ (.A(net830),
    .B(_07688_),
    .Y(_07689_));
 sg13g2_a22oi_1 _24280_ (.Y(_07690_),
    .B1(_07689_),
    .B2(\top_ihp.oisc.regs[3][11] ),
    .A2(net774),
    .A1(\top_ihp.oisc.regs[4][11] ));
 sg13g2_buf_1 _24281_ (.A(_07596_),
    .X(_07691_));
 sg13g2_buf_1 _24282_ (.A(_07604_),
    .X(_07692_));
 sg13g2_a22oi_1 _24283_ (.Y(_07693_),
    .B1(net850),
    .B2(\top_ihp.oisc.regs[14][11] ),
    .A2(net864),
    .A1(\top_ihp.oisc.regs[12][11] ));
 sg13g2_inv_1 _24284_ (.Y(_07694_),
    .A(_07693_));
 sg13g2_buf_1 _24285_ (.A(net935),
    .X(_07695_));
 sg13g2_a22oi_1 _24286_ (.Y(_07696_),
    .B1(_07694_),
    .B2(net893),
    .A2(_07659_),
    .A1(\top_ihp.oisc.regs[1][11] ));
 sg13g2_nand2_1 _24287_ (.Y(_07697_),
    .A(_07690_),
    .B(_07696_));
 sg13g2_nor4_1 _24288_ (.A(_07670_),
    .B(_07677_),
    .C(_07686_),
    .D(_07697_),
    .Y(_07698_));
 sg13g2_nand2_1 _24289_ (.Y(_07699_),
    .A(_08261_),
    .B(net667));
 sg13g2_o21ai_1 _24290_ (.B1(_07699_),
    .Y(_00454_),
    .A1(net733),
    .A2(_07698_));
 sg13g2_buf_1 _24291_ (.A(_07569_),
    .X(_07700_));
 sg13g2_mux2_1 _24292_ (.A0(\top_ihp.oisc.regs[7][12] ),
    .A1(\top_ihp.oisc.regs[3][12] ),
    .S(net803),
    .X(_07701_));
 sg13g2_mux2_1 _24293_ (.A0(\top_ihp.oisc.regs[6][12] ),
    .A1(\top_ihp.oisc.regs[2][12] ),
    .S(net808),
    .X(_07702_));
 sg13g2_a22oi_1 _24294_ (.Y(_07703_),
    .B1(_07702_),
    .B2(net853),
    .A2(_07701_),
    .A1(net809));
 sg13g2_buf_1 _24295_ (.A(_07569_),
    .X(_07704_));
 sg13g2_mux2_1 _24296_ (.A0(\top_ihp.oisc.regs[5][12] ),
    .A1(\top_ihp.oisc.regs[1][12] ),
    .S(net802),
    .X(_07705_));
 sg13g2_nand2_1 _24297_ (.Y(_07706_),
    .A(net839),
    .B(_07705_));
 sg13g2_a22oi_1 _24298_ (.Y(_07707_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][12] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][12] ));
 sg13g2_nor2_1 _24299_ (.A(_00253_),
    .B(net851),
    .Y(_07708_));
 sg13g2_a221oi_1 _24300_ (.B2(\top_ihp.oisc.regs[10][12] ),
    .C1(_07708_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][12] ),
    .Y(_07709_),
    .A2(net836));
 sg13g2_nand4_1 _24301_ (.B(_07706_),
    .C(_07707_),
    .A(_07703_),
    .Y(_07710_),
    .D(_07709_));
 sg13g2_nand2_1 _24302_ (.Y(_07711_),
    .A(\top_ihp.oisc.regs[4][12] ),
    .B(net769));
 sg13g2_buf_1 _24303_ (.A(_07596_),
    .X(_07712_));
 sg13g2_buf_1 _24304_ (.A(net850),
    .X(_07713_));
 sg13g2_a22oi_1 _24305_ (.Y(_07714_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][12] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[12][12] ));
 sg13g2_nand2b_1 _24306_ (.Y(_07715_),
    .B(net893),
    .A_N(_07714_));
 sg13g2_buf_1 _24307_ (.A(net771),
    .X(_07716_));
 sg13g2_nand2_1 _24308_ (.Y(_07717_),
    .A(\top_ihp.oisc.regs[9][12] ),
    .B(net753));
 sg13g2_buf_1 _24309_ (.A(net805),
    .X(_07718_));
 sg13g2_buf_1 _24310_ (.A(_07618_),
    .X(_07719_));
 sg13g2_buf_1 _24311_ (.A(net765),
    .X(_07720_));
 sg13g2_a22oi_1 _24312_ (.Y(_07721_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][12] ),
    .A2(net766),
    .A1(\top_ihp.oisc.regs[32][12] ));
 sg13g2_nand4_1 _24313_ (.B(_07715_),
    .C(_07717_),
    .A(_07711_),
    .Y(_07722_),
    .D(_07721_));
 sg13g2_nor2_1 _24314_ (.A(_07710_),
    .B(_07722_),
    .Y(_07723_));
 sg13g2_buf_1 _24315_ (.A(_03717_),
    .X(_07724_));
 sg13g2_nand2_1 _24316_ (.Y(_07725_),
    .A(_08253_),
    .B(_07724_));
 sg13g2_o21ai_1 _24317_ (.B1(_07725_),
    .Y(_00455_),
    .A1(net733),
    .A2(_07723_));
 sg13g2_buf_1 _24318_ (.A(_07612_),
    .X(_07726_));
 sg13g2_a22oi_1 _24319_ (.Y(_07727_),
    .B1(net771),
    .B2(\top_ihp.oisc.regs[9][13] ),
    .A2(net805),
    .A1(\top_ihp.oisc.regs[32][13] ));
 sg13g2_buf_1 _24320_ (.A(_07609_),
    .X(_07728_));
 sg13g2_a22oi_1 _24321_ (.Y(_07729_),
    .B1(net804),
    .B2(\top_ihp.oisc.regs[10][13] ),
    .A2(net801),
    .A1(\top_ihp.oisc.regs[14][13] ));
 sg13g2_a221oi_1 _24322_ (.B2(\top_ihp.oisc.regs[13][13] ),
    .C1(net849),
    .B1(net765),
    .A1(\top_ihp.oisc.regs[8][13] ),
    .Y(_07730_),
    .A2(net852));
 sg13g2_nand3_1 _24323_ (.B(_07729_),
    .C(_07730_),
    .A(_07727_),
    .Y(_07731_));
 sg13g2_a21oi_1 _24324_ (.A1(\top_ihp.oisc.regs[4][13] ),
    .A2(net769),
    .Y(_07732_),
    .B1(_07731_));
 sg13g2_buf_1 _24325_ (.A(_07567_),
    .X(_07733_));
 sg13g2_mux2_1 _24326_ (.A0(\top_ihp.oisc.regs[5][13] ),
    .A1(\top_ihp.oisc.regs[1][13] ),
    .S(_07583_),
    .X(_07734_));
 sg13g2_mux2_1 _24327_ (.A0(\top_ihp.oisc.regs[6][13] ),
    .A1(\top_ihp.oisc.regs[2][13] ),
    .S(net776),
    .X(_07735_));
 sg13g2_and2_1 _24328_ (.A(\top_ihp.oisc.regs[7][13] ),
    .B(_08998_),
    .X(_07736_));
 sg13g2_a21oi_1 _24329_ (.A1(\top_ihp.oisc.regs[3][13] ),
    .A2(net807),
    .Y(_07737_),
    .B1(_07736_));
 sg13g2_and2_1 _24330_ (.A(\top_ihp.oisc.regs[12][13] ),
    .B(_07598_),
    .X(_07738_));
 sg13g2_a221oi_1 _24331_ (.B2(\top_ihp.oisc.regs[15][13] ),
    .C1(_07738_),
    .B1(_07588_),
    .A1(\top_ihp.oisc.regs[11][13] ),
    .Y(_07739_),
    .A2(_07623_));
 sg13g2_o21ai_1 _24332_ (.B1(_07739_),
    .Y(_07740_),
    .A1(_07688_),
    .A2(_07737_));
 sg13g2_a221oi_1 _24333_ (.B2(net853),
    .C1(_07740_),
    .B1(_07735_),
    .A1(net834),
    .Y(_07741_),
    .A2(_07734_));
 sg13g2_a221oi_1 _24334_ (.B2(_07741_),
    .C1(net766),
    .B1(_07732_),
    .A1(_00254_),
    .Y(_07742_),
    .A2(net849));
 sg13g2_mux2_1 _24335_ (.A0(_07742_),
    .A1(_08251_),
    .S(_07637_),
    .X(_00456_));
 sg13g2_buf_1 _24336_ (.A(net719),
    .X(_07743_));
 sg13g2_and2_1 _24337_ (.A(\top_ihp.oisc.regs[2][14] ),
    .B(net776),
    .X(_07744_));
 sg13g2_a21oi_1 _24338_ (.A1(\top_ihp.oisc.regs[6][14] ),
    .A2(net794),
    .Y(_07745_),
    .B1(_07744_));
 sg13g2_mux2_1 _24339_ (.A0(\top_ihp.oisc.regs[7][14] ),
    .A1(\top_ihp.oisc.regs[3][14] ),
    .S(_07639_),
    .X(_07746_));
 sg13g2_mux2_1 _24340_ (.A0(\top_ihp.oisc.regs[5][14] ),
    .A1(\top_ihp.oisc.regs[1][14] ),
    .S(net803),
    .X(_07747_));
 sg13g2_a22oi_1 _24341_ (.Y(_07748_),
    .B1(_07747_),
    .B2(net834),
    .A2(_07746_),
    .A1(net806));
 sg13g2_o21ai_1 _24342_ (.B1(_07748_),
    .Y(_07749_),
    .A1(_07662_),
    .A2(_07745_));
 sg13g2_a22oi_1 _24343_ (.Y(_07750_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][14] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][14] ));
 sg13g2_mux2_1 _24344_ (.A0(\top_ihp.oisc.regs[8][14] ),
    .A1(\top_ihp.oisc.regs[12][14] ),
    .S(net935),
    .X(_07751_));
 sg13g2_a22oi_1 _24345_ (.Y(_07752_),
    .B1(_07751_),
    .B2(net863),
    .A2(net770),
    .A1(\top_ihp.oisc.regs[13][14] ));
 sg13g2_a22oi_1 _24346_ (.Y(_07753_),
    .B1(net801),
    .B2(\top_ihp.oisc.regs[14][14] ),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][14] ));
 sg13g2_buf_1 _24347_ (.A(_07651_),
    .X(_07754_));
 sg13g2_nand2_1 _24348_ (.Y(_07755_),
    .A(\top_ihp.oisc.regs[10][14] ),
    .B(_07681_));
 sg13g2_o21ai_1 _24349_ (.B1(_07755_),
    .Y(_07756_),
    .A1(_00255_),
    .A2(net848));
 sg13g2_a221oi_1 _24350_ (.B2(\top_ihp.oisc.regs[4][14] ),
    .C1(_07756_),
    .B1(_07594_),
    .A1(\top_ihp.oisc.regs[32][14] ),
    .Y(_07757_),
    .A2(net805));
 sg13g2_nand4_1 _24351_ (.B(_07752_),
    .C(_07753_),
    .A(_07750_),
    .Y(_07758_),
    .D(_07757_));
 sg13g2_o21ai_1 _24352_ (.B1(_07633_),
    .Y(_07759_),
    .A1(_07749_),
    .A2(_07758_));
 sg13g2_nand2_1 _24353_ (.Y(_07760_),
    .A(_08278_),
    .B(net666));
 sg13g2_o21ai_1 _24354_ (.B1(_07760_),
    .Y(_00457_),
    .A1(net665),
    .A2(_07759_));
 sg13g2_buf_1 _24355_ (.A(net865),
    .X(_07761_));
 sg13g2_mux2_1 _24356_ (.A0(\top_ihp.oisc.regs[6][15] ),
    .A1(\top_ihp.oisc.regs[2][15] ),
    .S(net807),
    .X(_07762_));
 sg13g2_nand2_1 _24357_ (.Y(_07763_),
    .A(net847),
    .B(_07762_));
 sg13g2_a22oi_1 _24358_ (.Y(_07764_),
    .B1(net836),
    .B2(\top_ihp.oisc.regs[8][15] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][15] ));
 sg13g2_nand2_1 _24359_ (.Y(_07765_),
    .A(\top_ihp.oisc.regs[12][15] ),
    .B(net838));
 sg13g2_mux2_1 _24360_ (.A0(\top_ihp.oisc.regs[7][15] ),
    .A1(\top_ihp.oisc.regs[3][15] ),
    .S(net810),
    .X(_07766_));
 sg13g2_buf_1 _24361_ (.A(_07569_),
    .X(_07767_));
 sg13g2_mux2_1 _24362_ (.A0(\top_ihp.oisc.regs[5][15] ),
    .A1(\top_ihp.oisc.regs[1][15] ),
    .S(net800),
    .X(_07768_));
 sg13g2_buf_1 _24363_ (.A(_07567_),
    .X(_07769_));
 sg13g2_a22oi_1 _24364_ (.Y(_07770_),
    .B1(_07768_),
    .B2(net833),
    .A2(_07766_),
    .A1(net806));
 sg13g2_nand4_1 _24365_ (.B(_07764_),
    .C(_07765_),
    .A(_07763_),
    .Y(_07771_),
    .D(_07770_));
 sg13g2_buf_1 _24366_ (.A(_07593_),
    .X(_07772_));
 sg13g2_nand2_1 _24367_ (.Y(_07773_),
    .A(\top_ihp.oisc.regs[4][15] ),
    .B(net764));
 sg13g2_nand2_1 _24368_ (.Y(_07774_),
    .A(\top_ihp.oisc.regs[32][15] ),
    .B(net766));
 sg13g2_mux2_1 _24369_ (.A0(\top_ihp.oisc.regs[10][15] ),
    .A1(\top_ihp.oisc.regs[14][15] ),
    .S(net985),
    .X(_07775_));
 sg13g2_nor2_1 _24370_ (.A(_00256_),
    .B(net848),
    .Y(_07776_));
 sg13g2_a221oi_1 _24371_ (.B2(_07775_),
    .C1(_07776_),
    .B1(_07713_),
    .A1(\top_ihp.oisc.regs[15][15] ),
    .Y(_07777_),
    .A2(net775));
 sg13g2_a22oi_1 _24372_ (.Y(_07778_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][15] ),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][15] ));
 sg13g2_nand4_1 _24373_ (.B(_07774_),
    .C(_07777_),
    .A(_07773_),
    .Y(_07779_),
    .D(_07778_));
 sg13g2_o21ai_1 _24374_ (.B1(_07633_),
    .Y(_07780_),
    .A1(_07771_),
    .A2(_07779_));
 sg13g2_nand2_1 _24375_ (.Y(_07781_),
    .A(_08279_),
    .B(net666));
 sg13g2_o21ai_1 _24376_ (.B1(_07781_),
    .Y(_00458_),
    .A1(net665),
    .A2(_07780_));
 sg13g2_mux2_1 _24377_ (.A0(\top_ihp.oisc.regs[7][16] ),
    .A1(\top_ihp.oisc.regs[3][16] ),
    .S(net803),
    .X(_07782_));
 sg13g2_mux2_1 _24378_ (.A0(\top_ihp.oisc.regs[6][16] ),
    .A1(\top_ihp.oisc.regs[2][16] ),
    .S(_07583_),
    .X(_07783_));
 sg13g2_a22oi_1 _24379_ (.Y(_07784_),
    .B1(_07783_),
    .B2(net853),
    .A2(_07782_),
    .A1(_07577_));
 sg13g2_mux2_1 _24380_ (.A0(\top_ihp.oisc.regs[5][16] ),
    .A1(\top_ihp.oisc.regs[1][16] ),
    .S(net802),
    .X(_07785_));
 sg13g2_nand2_1 _24381_ (.Y(_07786_),
    .A(_07568_),
    .B(_07785_));
 sg13g2_a22oi_1 _24382_ (.Y(_07787_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][16] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][16] ));
 sg13g2_nor2_1 _24383_ (.A(_00257_),
    .B(_07674_),
    .Y(_07788_));
 sg13g2_a221oi_1 _24384_ (.B2(\top_ihp.oisc.regs[10][16] ),
    .C1(_07788_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][16] ),
    .Y(_07789_),
    .A2(_07628_));
 sg13g2_nand4_1 _24385_ (.B(_07786_),
    .C(_07787_),
    .A(_07784_),
    .Y(_07790_),
    .D(_07789_));
 sg13g2_nand2_1 _24386_ (.Y(_07791_),
    .A(\top_ihp.oisc.regs[4][16] ),
    .B(net769));
 sg13g2_a22oi_1 _24387_ (.Y(_07792_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][16] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[12][16] ));
 sg13g2_nand2b_1 _24388_ (.Y(_07793_),
    .B(net893),
    .A_N(_07792_));
 sg13g2_nand2_1 _24389_ (.Y(_07794_),
    .A(\top_ihp.oisc.regs[9][16] ),
    .B(_07716_));
 sg13g2_buf_1 _24390_ (.A(net837),
    .X(_07795_));
 sg13g2_a22oi_1 _24391_ (.Y(_07796_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][16] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][16] ));
 sg13g2_nand4_1 _24392_ (.B(_07793_),
    .C(_07794_),
    .A(_07791_),
    .Y(_07797_),
    .D(_07796_));
 sg13g2_nor2_1 _24393_ (.A(_07790_),
    .B(_07797_),
    .Y(_07798_));
 sg13g2_nand2_1 _24394_ (.Y(_07799_),
    .A(_08272_),
    .B(net666));
 sg13g2_o21ai_1 _24395_ (.B1(_07799_),
    .Y(_00459_),
    .A1(net733),
    .A2(_07798_));
 sg13g2_mux2_1 _24396_ (.A0(\top_ihp.oisc.regs[7][17] ),
    .A1(\top_ihp.oisc.regs[3][17] ),
    .S(net803),
    .X(_07800_));
 sg13g2_mux2_1 _24397_ (.A0(\top_ihp.oisc.regs[6][17] ),
    .A1(\top_ihp.oisc.regs[2][17] ),
    .S(net808),
    .X(_07801_));
 sg13g2_a22oi_1 _24398_ (.Y(_07802_),
    .B1(_07801_),
    .B2(_07582_),
    .A2(_07800_),
    .A1(_07577_));
 sg13g2_mux2_1 _24399_ (.A0(\top_ihp.oisc.regs[5][17] ),
    .A1(\top_ihp.oisc.regs[1][17] ),
    .S(_07704_),
    .X(_07803_));
 sg13g2_nand2_1 _24400_ (.Y(_07804_),
    .A(_07568_),
    .B(_07803_));
 sg13g2_a22oi_1 _24401_ (.Y(_07805_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][17] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][17] ));
 sg13g2_nor2_1 _24402_ (.A(_00258_),
    .B(net851),
    .Y(_07806_));
 sg13g2_a221oi_1 _24403_ (.B2(\top_ihp.oisc.regs[10][17] ),
    .C1(_07806_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][17] ),
    .Y(_07807_),
    .A2(net836));
 sg13g2_nand4_1 _24404_ (.B(_07804_),
    .C(_07805_),
    .A(_07802_),
    .Y(_07808_),
    .D(_07807_));
 sg13g2_nand2_1 _24405_ (.Y(_07809_),
    .A(\top_ihp.oisc.regs[4][17] ),
    .B(_07657_));
 sg13g2_a22oi_1 _24406_ (.Y(_07810_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][17] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[12][17] ));
 sg13g2_nand2b_1 _24407_ (.Y(_07811_),
    .B(net893),
    .A_N(_07810_));
 sg13g2_nand2_1 _24408_ (.Y(_07812_),
    .A(\top_ihp.oisc.regs[9][17] ),
    .B(net753));
 sg13g2_a22oi_1 _24409_ (.Y(_07813_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][17] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][17] ));
 sg13g2_nand4_1 _24410_ (.B(_07811_),
    .C(_07812_),
    .A(_07809_),
    .Y(_07814_),
    .D(_07813_));
 sg13g2_nor2_1 _24411_ (.A(_07808_),
    .B(_07814_),
    .Y(_07815_));
 sg13g2_nand2_1 _24412_ (.Y(_07816_),
    .A(_08275_),
    .B(net666));
 sg13g2_o21ai_1 _24413_ (.B1(_07816_),
    .Y(_00460_),
    .A1(net733),
    .A2(_07815_));
 sg13g2_and2_1 _24414_ (.A(\top_ihp.oisc.regs[2][18] ),
    .B(net802),
    .X(_07817_));
 sg13g2_a21oi_1 _24415_ (.A1(\top_ihp.oisc.regs[6][18] ),
    .A2(\top_ihp.oisc.reg_rb[2] ),
    .Y(_07818_),
    .B1(_07817_));
 sg13g2_mux2_1 _24416_ (.A0(\top_ihp.oisc.regs[7][18] ),
    .A1(\top_ihp.oisc.regs[3][18] ),
    .S(net800),
    .X(_07819_));
 sg13g2_mux2_1 _24417_ (.A0(\top_ihp.oisc.regs[5][18] ),
    .A1(\top_ihp.oisc.regs[1][18] ),
    .S(net803),
    .X(_07820_));
 sg13g2_a22oi_1 _24418_ (.Y(_07821_),
    .B1(_07820_),
    .B2(net834),
    .A2(_07819_),
    .A1(net806));
 sg13g2_o21ai_1 _24419_ (.B1(_07821_),
    .Y(_07822_),
    .A1(_07662_),
    .A2(_07818_));
 sg13g2_a22oi_1 _24420_ (.Y(_07823_),
    .B1(_07684_),
    .B2(\top_ihp.oisc.regs[15][18] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][18] ));
 sg13g2_mux2_1 _24421_ (.A0(\top_ihp.oisc.regs[8][18] ),
    .A1(\top_ihp.oisc.regs[12][18] ),
    .S(net1041),
    .X(_07824_));
 sg13g2_a22oi_1 _24422_ (.Y(_07825_),
    .B1(_07824_),
    .B2(_07596_),
    .A2(_07616_),
    .A1(\top_ihp.oisc.regs[9][18] ));
 sg13g2_o21ai_1 _24423_ (.B1(_07825_),
    .Y(_07826_),
    .A1(_00259_),
    .A2(net848));
 sg13g2_a21oi_1 _24424_ (.A1(\top_ihp.oisc.regs[4][18] ),
    .A2(net774),
    .Y(_07827_),
    .B1(_07826_));
 sg13g2_a22oi_1 _24425_ (.Y(_07828_),
    .B1(_07682_),
    .B2(\top_ihp.oisc.regs[10][18] ),
    .A2(net801),
    .A1(\top_ihp.oisc.regs[14][18] ));
 sg13g2_a22oi_1 _24426_ (.Y(_07829_),
    .B1(net770),
    .B2(\top_ihp.oisc.regs[13][18] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][18] ));
 sg13g2_nand4_1 _24427_ (.B(_07827_),
    .C(_07828_),
    .A(_07823_),
    .Y(_07830_),
    .D(_07829_));
 sg13g2_o21ai_1 _24428_ (.B1(_07633_),
    .Y(_07831_),
    .A1(_07822_),
    .A2(_07830_));
 sg13g2_nand2_1 _24429_ (.Y(_07832_),
    .A(_08220_),
    .B(_07724_));
 sg13g2_o21ai_1 _24430_ (.B1(_07832_),
    .Y(_00461_),
    .A1(net665),
    .A2(_07831_));
 sg13g2_mux2_1 _24431_ (.A0(\top_ihp.oisc.regs[5][19] ),
    .A1(\top_ihp.oisc.regs[1][19] ),
    .S(net772),
    .X(_07833_));
 sg13g2_nand2_1 _24432_ (.Y(_07834_),
    .A(\top_ihp.oisc.regs[11][19] ),
    .B(net773));
 sg13g2_mux2_1 _24433_ (.A0(\top_ihp.oisc.regs[8][19] ),
    .A1(\top_ihp.oisc.regs[12][19] ),
    .S(net985),
    .X(_07835_));
 sg13g2_nand2_1 _24434_ (.Y(_07836_),
    .A(\top_ihp.oisc.regs[32][19] ),
    .B(net837));
 sg13g2_o21ai_1 _24435_ (.B1(_07836_),
    .Y(_07837_),
    .A1(_00260_),
    .A2(_07651_));
 sg13g2_a221oi_1 _24436_ (.B2(net864),
    .C1(_07837_),
    .B1(_07835_),
    .A1(\top_ihp.oisc.regs[13][19] ),
    .Y(_07838_),
    .A2(net765));
 sg13g2_mux2_1 _24437_ (.A0(\top_ihp.oisc.regs[10][19] ),
    .A1(\top_ihp.oisc.regs[14][19] ),
    .S(net985),
    .X(_07839_));
 sg13g2_a22oi_1 _24438_ (.Y(_07840_),
    .B1(net850),
    .B2(_07839_),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[9][19] ));
 sg13g2_nor2_2 _24439_ (.A(net810),
    .B(_07662_),
    .Y(_07841_));
 sg13g2_a22oi_1 _24440_ (.Y(_07842_),
    .B1(_07841_),
    .B2(\top_ihp.oisc.regs[6][19] ),
    .A2(net775),
    .A1(\top_ihp.oisc.regs[15][19] ));
 sg13g2_nand4_1 _24441_ (.B(_07838_),
    .C(_07840_),
    .A(_07834_),
    .Y(_07843_),
    .D(_07842_));
 sg13g2_a21oi_1 _24442_ (.A1(net839),
    .A2(_07833_),
    .Y(_07844_),
    .B1(_07843_));
 sg13g2_nand3_1 _24443_ (.B(net776),
    .C(net865),
    .A(\top_ihp.oisc.regs[2][19] ),
    .Y(_07845_));
 sg13g2_nand3_1 _24444_ (.B(net830),
    .C(_07576_),
    .A(\top_ihp.oisc.regs[7][19] ),
    .Y(_07846_));
 sg13g2_nand2_1 _24445_ (.Y(_07847_),
    .A(_07845_),
    .B(_07846_));
 sg13g2_a221oi_1 _24446_ (.B2(\top_ihp.oisc.regs[3][19] ),
    .C1(_07847_),
    .B1(_07689_),
    .A1(\top_ihp.oisc.regs[4][19] ),
    .Y(_07848_),
    .A2(net769));
 sg13g2_a21oi_1 _24447_ (.A1(_07844_),
    .A2(_07848_),
    .Y(_07849_),
    .B1(net741));
 sg13g2_a21o_1 _24448_ (.A2(_07637_),
    .A1(_08219_),
    .B1(_07849_),
    .X(_00462_));
 sg13g2_mux2_1 _24449_ (.A0(\top_ihp.oisc.regs[6][1] ),
    .A1(\top_ihp.oisc.regs[2][1] ),
    .S(net808),
    .X(_07850_));
 sg13g2_mux2_1 _24450_ (.A0(\top_ihp.oisc.regs[5][1] ),
    .A1(\top_ihp.oisc.regs[1][1] ),
    .S(net776),
    .X(_07851_));
 sg13g2_and2_1 _24451_ (.A(\top_ihp.oisc.regs[7][1] ),
    .B(net830),
    .X(_07852_));
 sg13g2_a21oi_1 _24452_ (.A1(\top_ihp.oisc.regs[3][1] ),
    .A2(net808),
    .Y(_07853_),
    .B1(_07852_));
 sg13g2_and2_1 _24453_ (.A(\top_ihp.oisc.regs[12][1] ),
    .B(_07598_),
    .X(_07854_));
 sg13g2_a221oi_1 _24454_ (.B2(\top_ihp.oisc.regs[15][1] ),
    .C1(_07854_),
    .B1(_07588_),
    .A1(\top_ihp.oisc.regs[8][1] ),
    .Y(_07855_),
    .A2(net852));
 sg13g2_o21ai_1 _24455_ (.B1(_07855_),
    .Y(_07856_),
    .A1(_07688_),
    .A2(_07853_));
 sg13g2_a221oi_1 _24456_ (.B2(net839),
    .C1(_07856_),
    .B1(_07851_),
    .A1(net853),
    .Y(_07857_),
    .A2(_07850_));
 sg13g2_a22oi_1 _24457_ (.Y(_07858_),
    .B1(net771),
    .B2(\top_ihp.oisc.regs[9][1] ),
    .A2(_07602_),
    .A1(\top_ihp.oisc.regs[32][1] ));
 sg13g2_a22oi_1 _24458_ (.Y(_07859_),
    .B1(net804),
    .B2(\top_ihp.oisc.regs[10][1] ),
    .A2(net801),
    .A1(\top_ihp.oisc.regs[14][1] ));
 sg13g2_a221oi_1 _24459_ (.B2(\top_ihp.oisc.regs[13][1] ),
    .C1(_07726_),
    .B1(net765),
    .A1(\top_ihp.oisc.regs[11][1] ),
    .Y(_07860_),
    .A2(_07623_));
 sg13g2_nand3_1 _24460_ (.B(_07859_),
    .C(_07860_),
    .A(_07858_),
    .Y(_07861_));
 sg13g2_a21oi_1 _24461_ (.A1(\top_ihp.oisc.regs[4][1] ),
    .A2(net769),
    .Y(_07862_),
    .B1(_07861_));
 sg13g2_a221oi_1 _24462_ (.B2(_07862_),
    .C1(net766),
    .B1(_07857_),
    .A1(_00242_),
    .Y(_07863_),
    .A2(net849));
 sg13g2_mux2_1 _24463_ (.A0(_07863_),
    .A1(_08319_),
    .S(net667),
    .X(_00463_));
 sg13g2_and2_1 _24464_ (.A(\top_ihp.oisc.regs[2][20] ),
    .B(net802),
    .X(_07864_));
 sg13g2_a21oi_1 _24465_ (.A1(\top_ihp.oisc.regs[6][20] ),
    .A2(net794),
    .Y(_07865_),
    .B1(_07864_));
 sg13g2_mux2_1 _24466_ (.A0(\top_ihp.oisc.regs[7][20] ),
    .A1(\top_ihp.oisc.regs[3][20] ),
    .S(net800),
    .X(_07866_));
 sg13g2_mux2_1 _24467_ (.A0(\top_ihp.oisc.regs[5][20] ),
    .A1(\top_ihp.oisc.regs[1][20] ),
    .S(_07700_),
    .X(_07867_));
 sg13g2_a22oi_1 _24468_ (.Y(_07868_),
    .B1(_07867_),
    .B2(net834),
    .A2(_07866_),
    .A1(net806));
 sg13g2_o21ai_1 _24469_ (.B1(_07868_),
    .Y(_07869_),
    .A1(_07662_),
    .A2(_07865_));
 sg13g2_nand2_1 _24470_ (.Y(_07870_),
    .A(\top_ihp.oisc.regs[4][20] ),
    .B(net764));
 sg13g2_nand2_1 _24471_ (.Y(_07871_),
    .A(\top_ihp.oisc.regs[9][20] ),
    .B(net753));
 sg13g2_mux2_1 _24472_ (.A0(\top_ihp.oisc.regs[8][20] ),
    .A1(\top_ihp.oisc.regs[12][20] ),
    .S(net935),
    .X(_07872_));
 sg13g2_a22oi_1 _24473_ (.Y(_07873_),
    .B1(_07712_),
    .B2(_07872_),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][20] ));
 sg13g2_mux2_1 _24474_ (.A0(\top_ihp.oisc.regs[10][20] ),
    .A1(\top_ihp.oisc.regs[14][20] ),
    .S(_08993_),
    .X(_07874_));
 sg13g2_a221oi_1 _24475_ (.B2(_07604_),
    .C1(_07612_),
    .B1(_07874_),
    .A1(\top_ihp.oisc.regs[13][20] ),
    .Y(_07875_),
    .A2(_07618_));
 sg13g2_inv_1 _24476_ (.Y(_07876_),
    .A(_07875_));
 sg13g2_a221oi_1 _24477_ (.B2(\top_ihp.oisc.regs[15][20] ),
    .C1(_07876_),
    .B1(net775),
    .A1(\top_ihp.oisc.regs[11][20] ),
    .Y(_07877_),
    .A2(_07624_));
 sg13g2_nand4_1 _24478_ (.B(_07871_),
    .C(_07873_),
    .A(_07870_),
    .Y(_07878_),
    .D(_07877_));
 sg13g2_a21oi_1 _24479_ (.A1(_00261_),
    .A2(net849),
    .Y(_07879_),
    .B1(net766));
 sg13g2_o21ai_1 _24480_ (.B1(_07879_),
    .Y(_07880_),
    .A1(_07869_),
    .A2(_07878_));
 sg13g2_nand2_1 _24481_ (.Y(_07881_),
    .A(_08227_),
    .B(net666));
 sg13g2_o21ai_1 _24482_ (.B1(_07881_),
    .Y(_00464_),
    .A1(net665),
    .A2(_07880_));
 sg13g2_a22oi_1 _24483_ (.Y(_07882_),
    .B1(_07733_),
    .B2(\top_ihp.oisc.regs[5][21] ),
    .A2(net847),
    .A1(\top_ihp.oisc.regs[6][21] ));
 sg13g2_nor2_1 _24484_ (.A(net758),
    .B(_07882_),
    .Y(_07883_));
 sg13g2_a22oi_1 _24485_ (.Y(_07884_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][21] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][21] ));
 sg13g2_nand2_1 _24486_ (.Y(_07885_),
    .A(\top_ihp.oisc.regs[10][21] ),
    .B(net804));
 sg13g2_o21ai_1 _24487_ (.B1(_07885_),
    .Y(_07886_),
    .A1(_00262_),
    .A2(net848));
 sg13g2_a221oi_1 _24488_ (.B2(\top_ihp.oisc.regs[1][21] ),
    .C1(_07886_),
    .B1(_07659_),
    .A1(\top_ihp.oisc.regs[32][21] ),
    .Y(_07887_),
    .A2(net805));
 sg13g2_a22oi_1 _24489_ (.Y(_07888_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][21] ),
    .A2(net801),
    .A1(\top_ihp.oisc.regs[14][21] ));
 sg13g2_mux2_1 _24490_ (.A0(\top_ihp.oisc.regs[8][21] ),
    .A1(\top_ihp.oisc.regs[12][21] ),
    .S(_07643_),
    .X(_07889_));
 sg13g2_a22oi_1 _24491_ (.Y(_07890_),
    .B1(_07889_),
    .B2(net863),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][21] ));
 sg13g2_nand4_1 _24492_ (.B(_07887_),
    .C(_07888_),
    .A(_07884_),
    .Y(_07891_),
    .D(_07890_));
 sg13g2_and2_1 _24493_ (.A(\top_ihp.oisc.regs[7][21] ),
    .B(_08999_),
    .X(_07892_));
 sg13g2_a21oi_1 _24494_ (.A1(\top_ihp.oisc.regs[3][21] ),
    .A2(net758),
    .Y(_07893_),
    .B1(_07892_));
 sg13g2_a22oi_1 _24495_ (.Y(_07894_),
    .B1(_07663_),
    .B2(\top_ihp.oisc.regs[2][21] ),
    .A2(net764),
    .A1(\top_ihp.oisc.regs[4][21] ));
 sg13g2_o21ai_1 _24496_ (.B1(_07894_),
    .Y(_07895_),
    .A1(_07688_),
    .A2(_07893_));
 sg13g2_nor3_1 _24497_ (.A(_07883_),
    .B(_07891_),
    .C(_07895_),
    .Y(_07896_));
 sg13g2_nand2_1 _24498_ (.Y(_07897_),
    .A(_08231_),
    .B(net666));
 sg13g2_o21ai_1 _24499_ (.B1(_07897_),
    .Y(_00465_),
    .A1(net733),
    .A2(_07896_));
 sg13g2_mux2_1 _24500_ (.A0(\top_ihp.oisc.regs[6][22] ),
    .A1(\top_ihp.oisc.regs[2][22] ),
    .S(net807),
    .X(_07898_));
 sg13g2_nand2_1 _24501_ (.Y(_07899_),
    .A(net847),
    .B(_07898_));
 sg13g2_a22oi_1 _24502_ (.Y(_07900_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][22] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][22] ));
 sg13g2_nand2_1 _24503_ (.Y(_07901_),
    .A(\top_ihp.oisc.regs[12][22] ),
    .B(net838));
 sg13g2_mux2_1 _24504_ (.A0(\top_ihp.oisc.regs[7][22] ),
    .A1(\top_ihp.oisc.regs[3][22] ),
    .S(net810),
    .X(_07902_));
 sg13g2_mux2_1 _24505_ (.A0(\top_ihp.oisc.regs[5][22] ),
    .A1(\top_ihp.oisc.regs[1][22] ),
    .S(net800),
    .X(_07903_));
 sg13g2_a22oi_1 _24506_ (.Y(_07904_),
    .B1(_07903_),
    .B2(net833),
    .A2(_07902_),
    .A1(net806));
 sg13g2_nand4_1 _24507_ (.B(_07900_),
    .C(_07901_),
    .A(_07899_),
    .Y(_07905_),
    .D(_07904_));
 sg13g2_nand2_1 _24508_ (.Y(_07906_),
    .A(\top_ihp.oisc.regs[8][22] ),
    .B(net836));
 sg13g2_mux2_1 _24509_ (.A0(\top_ihp.oisc.regs[10][22] ),
    .A1(\top_ihp.oisc.regs[14][22] ),
    .S(net935),
    .X(_07907_));
 sg13g2_a22oi_1 _24510_ (.Y(_07908_),
    .B1(net835),
    .B2(_07907_),
    .A2(net753),
    .A1(\top_ihp.oisc.regs[9][22] ));
 sg13g2_nand2_1 _24511_ (.Y(_07909_),
    .A(\top_ihp.oisc.regs[13][22] ),
    .B(_07719_));
 sg13g2_o21ai_1 _24512_ (.B1(_07909_),
    .Y(_07910_),
    .A1(_00263_),
    .A2(net848));
 sg13g2_a221oi_1 _24513_ (.B2(\top_ihp.oisc.regs[4][22] ),
    .C1(_07910_),
    .B1(net774),
    .A1(\top_ihp.oisc.regs[32][22] ),
    .Y(_07911_),
    .A2(net805));
 sg13g2_nand3_1 _24514_ (.B(_07908_),
    .C(_07911_),
    .A(_07906_),
    .Y(_07912_));
 sg13g2_o21ai_1 _24515_ (.B1(_07633_),
    .Y(_07913_),
    .A1(_07905_),
    .A2(_07912_));
 sg13g2_nand2_1 _24516_ (.Y(_07914_),
    .A(_08392_),
    .B(net666));
 sg13g2_o21ai_1 _24517_ (.B1(_07914_),
    .Y(_00466_),
    .A1(net665),
    .A2(_07913_));
 sg13g2_nand2_1 _24518_ (.Y(_07915_),
    .A(\top_ihp.oisc.regs[3][23] ),
    .B(_07640_));
 sg13g2_nand2_1 _24519_ (.Y(_07916_),
    .A(\top_ihp.oisc.regs[7][23] ),
    .B(net794));
 sg13g2_a21oi_1 _24520_ (.A1(_07915_),
    .A2(_07916_),
    .Y(_07917_),
    .B1(_07688_));
 sg13g2_a22oi_1 _24521_ (.Y(_07918_),
    .B1(net833),
    .B2(\top_ihp.oisc.regs[5][23] ),
    .A2(net865),
    .A1(\top_ihp.oisc.regs[6][23] ));
 sg13g2_nor2_1 _24522_ (.A(_00069_),
    .B(net851),
    .Y(_07919_));
 sg13g2_a221oi_1 _24523_ (.B2(\top_ihp.oisc.regs[13][23] ),
    .C1(_07919_),
    .B1(_07649_),
    .A1(\top_ihp.oisc.regs[9][23] ),
    .Y(_07920_),
    .A2(net768));
 sg13g2_o21ai_1 _24524_ (.B1(_07920_),
    .Y(_07921_),
    .A1(net758),
    .A2(_07918_));
 sg13g2_nand2_1 _24525_ (.Y(_07922_),
    .A(\top_ihp.oisc.regs[11][23] ),
    .B(net755));
 sg13g2_a22oi_1 _24526_ (.Y(_07923_),
    .B1(_07728_),
    .B2(\top_ihp.oisc.regs[14][23] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][23] ));
 sg13g2_a22oi_1 _24527_ (.Y(_07924_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][23] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[12][23] ));
 sg13g2_nand3_1 _24528_ (.B(_07923_),
    .C(_07924_),
    .A(_07922_),
    .Y(_07925_));
 sg13g2_a22oi_1 _24529_ (.Y(_07926_),
    .B1(net833),
    .B2(\top_ihp.oisc.regs[1][23] ),
    .A2(net847),
    .A1(\top_ihp.oisc.regs[2][23] ));
 sg13g2_a22oi_1 _24530_ (.Y(_07927_),
    .B1(net850),
    .B2(\top_ihp.oisc.regs[10][23] ),
    .A2(_07691_),
    .A1(\top_ihp.oisc.regs[8][23] ));
 sg13g2_nor2_1 _24531_ (.A(_07695_),
    .B(_07927_),
    .Y(_07928_));
 sg13g2_a21oi_1 _24532_ (.A1(\top_ihp.oisc.regs[4][23] ),
    .A2(net774),
    .Y(_07929_),
    .B1(_07928_));
 sg13g2_o21ai_1 _24533_ (.B1(_07929_),
    .Y(_07930_),
    .A1(net794),
    .A2(_07926_));
 sg13g2_nor4_1 _24534_ (.A(_07917_),
    .B(_07921_),
    .C(_07925_),
    .D(_07930_),
    .Y(_07931_));
 sg13g2_nand2_1 _24535_ (.Y(_07932_),
    .A(_08395_),
    .B(net666));
 sg13g2_o21ai_1 _24536_ (.B1(_07932_),
    .Y(_00467_),
    .A1(_07636_),
    .A2(_07931_));
 sg13g2_mux2_1 _24537_ (.A0(\top_ihp.oisc.regs[5][24] ),
    .A1(\top_ihp.oisc.regs[1][24] ),
    .S(net758),
    .X(_07933_));
 sg13g2_mux2_1 _24538_ (.A0(\top_ihp.oisc.regs[7][24] ),
    .A1(\top_ihp.oisc.regs[3][24] ),
    .S(net758),
    .X(_07934_));
 sg13g2_a22oi_1 _24539_ (.Y(_07935_),
    .B1(net850),
    .B2(\top_ihp.oisc.regs[14][24] ),
    .A2(_07596_),
    .A1(\top_ihp.oisc.regs[12][24] ));
 sg13g2_nor2_1 _24540_ (.A(_09141_),
    .B(_07935_),
    .Y(_07936_));
 sg13g2_a221oi_1 _24541_ (.B2(\top_ihp.oisc.regs[2][24] ),
    .C1(_07936_),
    .B1(_07663_),
    .A1(\top_ihp.oisc.regs[4][24] ),
    .Y(_07937_),
    .A2(net774));
 sg13g2_a22oi_1 _24542_ (.Y(_07938_),
    .B1(net765),
    .B2(\top_ihp.oisc.regs[13][24] ),
    .A2(_07616_),
    .A1(\top_ihp.oisc.regs[9][24] ));
 sg13g2_o21ai_1 _24543_ (.B1(_07938_),
    .Y(_07939_),
    .A1(_00070_),
    .A2(net851));
 sg13g2_a21oi_1 _24544_ (.A1(\top_ihp.oisc.regs[6][24] ),
    .A2(_07841_),
    .Y(_07940_),
    .B1(_07939_));
 sg13g2_and2_1 _24545_ (.A(\top_ihp.oisc.regs[10][24] ),
    .B(net804),
    .X(_07941_));
 sg13g2_a221oi_1 _24546_ (.B2(\top_ihp.oisc.regs[11][24] ),
    .C1(_07941_),
    .B1(net773),
    .A1(\top_ihp.oisc.regs[32][24] ),
    .Y(_07942_),
    .A2(net805));
 sg13g2_a22oi_1 _24547_ (.Y(_07943_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][24] ),
    .A2(net836),
    .A1(\top_ihp.oisc.regs[8][24] ));
 sg13g2_nand4_1 _24548_ (.B(_07940_),
    .C(_07942_),
    .A(_07937_),
    .Y(_07944_),
    .D(_07943_));
 sg13g2_a221oi_1 _24549_ (.B2(net809),
    .C1(_07944_),
    .B1(_07934_),
    .A1(net839),
    .Y(_07945_),
    .A2(_07933_));
 sg13g2_buf_1 _24550_ (.A(_03717_),
    .X(_07946_));
 sg13g2_nand2_1 _24551_ (.Y(_07947_),
    .A(_08379_),
    .B(net664));
 sg13g2_o21ai_1 _24552_ (.B1(_07947_),
    .Y(_00468_),
    .A1(net733),
    .A2(_07945_));
 sg13g2_nand2_1 _24553_ (.Y(_07948_),
    .A(\top_ihp.oisc.regs[3][25] ),
    .B(net772));
 sg13g2_nand2_1 _24554_ (.Y(_07949_),
    .A(\top_ihp.oisc.regs[7][25] ),
    .B(net794));
 sg13g2_a21oi_1 _24555_ (.A1(_07948_),
    .A2(_07949_),
    .Y(_07950_),
    .B1(_07688_));
 sg13g2_a22oi_1 _24556_ (.Y(_07951_),
    .B1(_07567_),
    .B2(\top_ihp.oisc.regs[5][25] ),
    .A2(_07581_),
    .A1(\top_ihp.oisc.regs[6][25] ));
 sg13g2_nor2_1 _24557_ (.A(_00071_),
    .B(net848),
    .Y(_07952_));
 sg13g2_a221oi_1 _24558_ (.B2(\top_ihp.oisc.regs[13][25] ),
    .C1(_07952_),
    .B1(net770),
    .A1(\top_ihp.oisc.regs[9][25] ),
    .Y(_07953_),
    .A2(_07680_));
 sg13g2_o21ai_1 _24559_ (.B1(_07953_),
    .Y(_07954_),
    .A1(_07572_),
    .A2(_07951_));
 sg13g2_nand2_1 _24560_ (.Y(_07955_),
    .A(\top_ihp.oisc.regs[11][25] ),
    .B(_07678_));
 sg13g2_a22oi_1 _24561_ (.Y(_07956_),
    .B1(net801),
    .B2(\top_ihp.oisc.regs[14][25] ),
    .A2(_07795_),
    .A1(\top_ihp.oisc.regs[32][25] ));
 sg13g2_a22oi_1 _24562_ (.Y(_07957_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][25] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[12][25] ));
 sg13g2_nand3_1 _24563_ (.B(_07956_),
    .C(_07957_),
    .A(_07955_),
    .Y(_07958_));
 sg13g2_a22oi_1 _24564_ (.Y(_07959_),
    .B1(net833),
    .B2(\top_ihp.oisc.regs[1][25] ),
    .A2(_07761_),
    .A1(\top_ihp.oisc.regs[2][25] ));
 sg13g2_a22oi_1 _24565_ (.Y(_07960_),
    .B1(_07692_),
    .B2(\top_ihp.oisc.regs[10][25] ),
    .A2(net864),
    .A1(\top_ihp.oisc.regs[8][25] ));
 sg13g2_nor2_1 _24566_ (.A(_07643_),
    .B(_07960_),
    .Y(_07961_));
 sg13g2_a21oi_1 _24567_ (.A1(\top_ihp.oisc.regs[4][25] ),
    .A2(net774),
    .Y(_07962_),
    .B1(_07961_));
 sg13g2_o21ai_1 _24568_ (.B1(_07962_),
    .Y(_07963_),
    .A1(net794),
    .A2(_07959_));
 sg13g2_nor4_1 _24569_ (.A(_07950_),
    .B(_07954_),
    .C(_07958_),
    .D(_07963_),
    .Y(_07964_));
 sg13g2_nand2_1 _24570_ (.Y(_07965_),
    .A(_08385_),
    .B(net664));
 sg13g2_o21ai_1 _24571_ (.B1(_07965_),
    .Y(_00469_),
    .A1(_07636_),
    .A2(_07964_));
 sg13g2_a221oi_1 _24572_ (.B2(\top_ihp.oisc.regs[14][26] ),
    .C1(net849),
    .B1(_07609_),
    .A1(\top_ihp.oisc.regs[8][26] ),
    .Y(_07966_),
    .A2(_07627_));
 sg13g2_a22oi_1 _24573_ (.Y(_07967_),
    .B1(_07646_),
    .B2(\top_ihp.oisc.regs[9][26] ),
    .A2(net837),
    .A1(\top_ihp.oisc.regs[32][26] ));
 sg13g2_a22oi_1 _24574_ (.Y(_07968_),
    .B1(net804),
    .B2(\top_ihp.oisc.regs[10][26] ),
    .A2(_07719_),
    .A1(\top_ihp.oisc.regs[13][26] ));
 sg13g2_nand3_1 _24575_ (.B(_07967_),
    .C(_07968_),
    .A(_07966_),
    .Y(_07969_));
 sg13g2_a21oi_1 _24576_ (.A1(\top_ihp.oisc.regs[4][26] ),
    .A2(net764),
    .Y(_07970_),
    .B1(_07969_));
 sg13g2_mux2_1 _24577_ (.A0(\top_ihp.oisc.regs[6][26] ),
    .A1(\top_ihp.oisc.regs[2][26] ),
    .S(net810),
    .X(_07971_));
 sg13g2_mux2_1 _24578_ (.A0(\top_ihp.oisc.regs[7][26] ),
    .A1(\top_ihp.oisc.regs[3][26] ),
    .S(net800),
    .X(_07972_));
 sg13g2_a22oi_1 _24579_ (.Y(_07973_),
    .B1(_07588_),
    .B2(\top_ihp.oisc.regs[15][26] ),
    .A2(_07623_),
    .A1(\top_ihp.oisc.regs[11][26] ));
 sg13g2_mux2_1 _24580_ (.A0(\top_ihp.oisc.regs[5][26] ),
    .A1(\top_ihp.oisc.regs[1][26] ),
    .S(_07569_),
    .X(_07974_));
 sg13g2_nand2_1 _24581_ (.Y(_07975_),
    .A(_07567_),
    .B(_07974_));
 sg13g2_nand2_1 _24582_ (.Y(_07976_),
    .A(\top_ihp.oisc.regs[12][26] ),
    .B(_07599_));
 sg13g2_nand3_1 _24583_ (.B(_07975_),
    .C(_07976_),
    .A(_07973_),
    .Y(_07977_));
 sg13g2_a221oi_1 _24584_ (.B2(_07671_),
    .C1(_07977_),
    .B1(_07972_),
    .A1(net847),
    .Y(_07978_),
    .A2(_07971_));
 sg13g2_a221oi_1 _24585_ (.B2(_07978_),
    .C1(net766),
    .B1(_07970_),
    .A1(_00072_),
    .Y(_07979_),
    .A2(net849));
 sg13g2_nor2_1 _24586_ (.A(net718),
    .B(_07979_),
    .Y(_07980_));
 sg13g2_a21oi_1 _24587_ (.A1(_08218_),
    .A2(net665),
    .Y(_00470_),
    .B1(_07980_));
 sg13g2_mux2_1 _24588_ (.A0(\top_ihp.oisc.regs[7][27] ),
    .A1(\top_ihp.oisc.regs[3][27] ),
    .S(net803),
    .X(_07981_));
 sg13g2_mux2_1 _24589_ (.A0(\top_ihp.oisc.regs[6][27] ),
    .A1(\top_ihp.oisc.regs[2][27] ),
    .S(net808),
    .X(_07982_));
 sg13g2_a22oi_1 _24590_ (.Y(_07983_),
    .B1(_07982_),
    .B2(net853),
    .A2(_07981_),
    .A1(net809));
 sg13g2_mux2_1 _24591_ (.A0(\top_ihp.oisc.regs[5][27] ),
    .A1(\top_ihp.oisc.regs[1][27] ),
    .S(net802),
    .X(_07984_));
 sg13g2_nand2_1 _24592_ (.Y(_07985_),
    .A(net834),
    .B(_07984_));
 sg13g2_a22oi_1 _24593_ (.Y(_07986_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][27] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][27] ));
 sg13g2_nor2_1 _24594_ (.A(_00073_),
    .B(net851),
    .Y(_07987_));
 sg13g2_a221oi_1 _24595_ (.B2(\top_ihp.oisc.regs[10][27] ),
    .C1(_07987_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][27] ),
    .Y(_07988_),
    .A2(net836));
 sg13g2_nand4_1 _24596_ (.B(_07985_),
    .C(_07986_),
    .A(_07983_),
    .Y(_07989_),
    .D(_07988_));
 sg13g2_nand2_1 _24597_ (.Y(_07990_),
    .A(\top_ihp.oisc.regs[4][27] ),
    .B(net764));
 sg13g2_a22oi_1 _24598_ (.Y(_07991_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][27] ),
    .A2(net863),
    .A1(\top_ihp.oisc.regs[12][27] ));
 sg13g2_nand2b_1 _24599_ (.Y(_07992_),
    .B(net893),
    .A_N(_07991_));
 sg13g2_nand2_1 _24600_ (.Y(_07993_),
    .A(\top_ihp.oisc.regs[9][27] ),
    .B(net753));
 sg13g2_a22oi_1 _24601_ (.Y(_07994_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][27] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][27] ));
 sg13g2_nand4_1 _24602_ (.B(_07992_),
    .C(_07993_),
    .A(_07990_),
    .Y(_07995_),
    .D(_07994_));
 sg13g2_nor2_1 _24603_ (.A(_07989_),
    .B(_07995_),
    .Y(_07996_));
 sg13g2_nand2_1 _24604_ (.Y(_07997_),
    .A(\top_ihp.oisc.op_b[27] ),
    .B(net664));
 sg13g2_o21ai_1 _24605_ (.B1(_07997_),
    .Y(_00471_),
    .A1(net733),
    .A2(_07996_));
 sg13g2_and2_1 _24606_ (.A(\top_ihp.oisc.regs[6][28] ),
    .B(net830),
    .X(_07998_));
 sg13g2_a21oi_1 _24607_ (.A1(\top_ihp.oisc.regs[2][28] ),
    .A2(net772),
    .Y(_07999_),
    .B1(_07998_));
 sg13g2_mux2_1 _24608_ (.A0(\top_ihp.oisc.regs[7][28] ),
    .A1(\top_ihp.oisc.regs[3][28] ),
    .S(net800),
    .X(_08000_));
 sg13g2_mux2_1 _24609_ (.A0(\top_ihp.oisc.regs[5][28] ),
    .A1(\top_ihp.oisc.regs[1][28] ),
    .S(net803),
    .X(_08001_));
 sg13g2_a22oi_1 _24610_ (.Y(_08002_),
    .B1(_08001_),
    .B2(net833),
    .A2(_08000_),
    .A1(net806));
 sg13g2_o21ai_1 _24611_ (.B1(_08002_),
    .Y(_08003_),
    .A1(_07662_),
    .A2(_07999_));
 sg13g2_a22oi_1 _24612_ (.Y(_08004_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][28] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][28] ));
 sg13g2_a22oi_1 _24613_ (.Y(_08005_),
    .B1(net765),
    .B2(\top_ihp.oisc.regs[13][28] ),
    .A2(_07609_),
    .A1(\top_ihp.oisc.regs[14][28] ));
 sg13g2_inv_1 _24614_ (.Y(_08006_),
    .A(_08005_));
 sg13g2_a221oi_1 _24615_ (.B2(\top_ihp.oisc.regs[10][28] ),
    .C1(_08006_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[4][28] ),
    .Y(_08007_),
    .A2(_07593_));
 sg13g2_mux2_1 _24616_ (.A0(\top_ihp.oisc.regs[8][28] ),
    .A1(\top_ihp.oisc.regs[12][28] ),
    .S(net935),
    .X(_08008_));
 sg13g2_a21oi_1 _24617_ (.A1(_07712_),
    .A2(_08008_),
    .Y(_08009_),
    .B1(_07726_));
 sg13g2_a22oi_1 _24618_ (.Y(_08010_),
    .B1(net753),
    .B2(\top_ihp.oisc.regs[9][28] ),
    .A2(net805),
    .A1(\top_ihp.oisc.regs[32][28] ));
 sg13g2_nand4_1 _24619_ (.B(_08007_),
    .C(_08009_),
    .A(_08004_),
    .Y(_08011_),
    .D(_08010_));
 sg13g2_a21oi_1 _24620_ (.A1(_00074_),
    .A2(net849),
    .Y(_08012_),
    .B1(net766));
 sg13g2_o21ai_1 _24621_ (.B1(_08012_),
    .Y(_08013_),
    .A1(_08003_),
    .A2(_08011_));
 sg13g2_nand2_1 _24622_ (.Y(_08014_),
    .A(_08444_),
    .B(_07946_));
 sg13g2_o21ai_1 _24623_ (.B1(_08014_),
    .Y(_00472_),
    .A1(net665),
    .A2(_08013_));
 sg13g2_and2_1 _24624_ (.A(\top_ihp.oisc.regs[2][29] ),
    .B(net802),
    .X(_08015_));
 sg13g2_a21oi_1 _24625_ (.A1(\top_ihp.oisc.regs[6][29] ),
    .A2(net794),
    .Y(_08016_),
    .B1(_08015_));
 sg13g2_mux2_1 _24626_ (.A0(\top_ihp.oisc.regs[7][29] ),
    .A1(\top_ihp.oisc.regs[3][29] ),
    .S(_07767_),
    .X(_08017_));
 sg13g2_mux2_1 _24627_ (.A0(\top_ihp.oisc.regs[5][29] ),
    .A1(\top_ihp.oisc.regs[1][29] ),
    .S(_07700_),
    .X(_08018_));
 sg13g2_a22oi_1 _24628_ (.Y(_08019_),
    .B1(_08018_),
    .B2(_07769_),
    .A2(_08017_),
    .A1(_07671_));
 sg13g2_o21ai_1 _24629_ (.B1(_08019_),
    .Y(_08020_),
    .A1(_07662_),
    .A2(_08016_));
 sg13g2_a22oi_1 _24630_ (.Y(_08021_),
    .B1(_07684_),
    .B2(\top_ihp.oisc.regs[15][29] ),
    .A2(_07625_),
    .A1(\top_ihp.oisc.regs[11][29] ));
 sg13g2_mux2_1 _24631_ (.A0(\top_ihp.oisc.regs[8][29] ),
    .A1(\top_ihp.oisc.regs[12][29] ),
    .S(net935),
    .X(_08022_));
 sg13g2_a22oi_1 _24632_ (.Y(_08023_),
    .B1(_08022_),
    .B2(net863),
    .A2(net770),
    .A1(\top_ihp.oisc.regs[13][29] ));
 sg13g2_a22oi_1 _24633_ (.Y(_08024_),
    .B1(_07728_),
    .B2(\top_ihp.oisc.regs[14][29] ),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][29] ));
 sg13g2_nand2_1 _24634_ (.Y(_08025_),
    .A(\top_ihp.oisc.regs[10][29] ),
    .B(net804));
 sg13g2_o21ai_1 _24635_ (.B1(_08025_),
    .Y(_08026_),
    .A1(_00075_),
    .A2(_07754_));
 sg13g2_a221oi_1 _24636_ (.B2(\top_ihp.oisc.regs[4][29] ),
    .C1(_08026_),
    .B1(_07593_),
    .A1(\top_ihp.oisc.regs[32][29] ),
    .Y(_08027_),
    .A2(_07673_));
 sg13g2_nand4_1 _24637_ (.B(_08023_),
    .C(_08024_),
    .A(_08021_),
    .Y(_08028_),
    .D(_08027_));
 sg13g2_o21ai_1 _24638_ (.B1(_07633_),
    .Y(_08029_),
    .A1(_08020_),
    .A2(_08028_));
 sg13g2_nand2_1 _24639_ (.Y(_08030_),
    .A(_08558_),
    .B(_07946_));
 sg13g2_o21ai_1 _24640_ (.B1(_08030_),
    .Y(_00473_),
    .A1(_07743_),
    .A2(_08029_));
 sg13g2_mux2_1 _24641_ (.A0(\top_ihp.oisc.regs[6][2] ),
    .A1(\top_ihp.oisc.regs[2][2] ),
    .S(net807),
    .X(_08031_));
 sg13g2_nand2_1 _24642_ (.Y(_08032_),
    .A(_07761_),
    .B(_08031_));
 sg13g2_a22oi_1 _24643_ (.Y(_08033_),
    .B1(_07628_),
    .B2(\top_ihp.oisc.regs[8][2] ),
    .A2(_07625_),
    .A1(\top_ihp.oisc.regs[11][2] ));
 sg13g2_nand2_1 _24644_ (.Y(_08034_),
    .A(\top_ihp.oisc.regs[12][2] ),
    .B(_07599_));
 sg13g2_mux2_1 _24645_ (.A0(\top_ihp.oisc.regs[7][2] ),
    .A1(\top_ihp.oisc.regs[3][2] ),
    .S(_07570_),
    .X(_08035_));
 sg13g2_mux2_1 _24646_ (.A0(\top_ihp.oisc.regs[5][2] ),
    .A1(\top_ihp.oisc.regs[1][2] ),
    .S(_07767_),
    .X(_08036_));
 sg13g2_a22oi_1 _24647_ (.Y(_08037_),
    .B1(_08036_),
    .B2(_07769_),
    .A2(_08035_),
    .A1(_07576_));
 sg13g2_nand4_1 _24648_ (.B(_08033_),
    .C(_08034_),
    .A(_08032_),
    .Y(_08038_),
    .D(_08037_));
 sg13g2_nand2_1 _24649_ (.Y(_08039_),
    .A(\top_ihp.oisc.regs[4][2] ),
    .B(_07772_));
 sg13g2_nand2_1 _24650_ (.Y(_08040_),
    .A(\top_ihp.oisc.regs[32][2] ),
    .B(_07718_));
 sg13g2_mux2_1 _24651_ (.A0(\top_ihp.oisc.regs[10][2] ),
    .A1(\top_ihp.oisc.regs[14][2] ),
    .S(net985),
    .X(_08041_));
 sg13g2_nor2_1 _24652_ (.A(_00243_),
    .B(net848),
    .Y(_08042_));
 sg13g2_a221oi_1 _24653_ (.B2(_08041_),
    .C1(_08042_),
    .B1(_07713_),
    .A1(\top_ihp.oisc.regs[15][2] ),
    .Y(_08043_),
    .A2(_07589_));
 sg13g2_a22oi_1 _24654_ (.Y(_08044_),
    .B1(_07649_),
    .B2(\top_ihp.oisc.regs[13][2] ),
    .A2(_07680_),
    .A1(\top_ihp.oisc.regs[9][2] ));
 sg13g2_nand4_1 _24655_ (.B(_08040_),
    .C(_08043_),
    .A(_08039_),
    .Y(_08045_),
    .D(_08044_));
 sg13g2_o21ai_1 _24656_ (.B1(_07633_),
    .Y(_08046_),
    .A1(_08038_),
    .A2(_08045_));
 sg13g2_nand2_1 _24657_ (.Y(_08047_),
    .A(_08330_),
    .B(net664));
 sg13g2_o21ai_1 _24658_ (.B1(_08047_),
    .Y(_00474_),
    .A1(_07743_),
    .A2(_08046_));
 sg13g2_mux2_1 _24659_ (.A0(\top_ihp.oisc.regs[6][30] ),
    .A1(\top_ihp.oisc.regs[2][30] ),
    .S(net810),
    .X(_08048_));
 sg13g2_mux2_1 _24660_ (.A0(\top_ihp.oisc.regs[5][30] ),
    .A1(\top_ihp.oisc.regs[1][30] ),
    .S(net800),
    .X(_08049_));
 sg13g2_and2_1 _24661_ (.A(\top_ihp.oisc.regs[7][30] ),
    .B(_08998_),
    .X(_08050_));
 sg13g2_a21oi_1 _24662_ (.A1(\top_ihp.oisc.regs[3][30] ),
    .A2(_07570_),
    .Y(_08051_),
    .B1(_08050_));
 sg13g2_and2_1 _24663_ (.A(\top_ihp.oisc.regs[12][30] ),
    .B(_07598_),
    .X(_08052_));
 sg13g2_a221oi_1 _24664_ (.B2(\top_ihp.oisc.regs[15][30] ),
    .C1(_08052_),
    .B1(_07588_),
    .A1(\top_ihp.oisc.regs[8][30] ),
    .Y(_08053_),
    .A2(net852));
 sg13g2_o21ai_1 _24665_ (.B1(_08053_),
    .Y(_08054_),
    .A1(_07688_),
    .A2(_08051_));
 sg13g2_a221oi_1 _24666_ (.B2(net833),
    .C1(_08054_),
    .B1(_08049_),
    .A1(net847),
    .Y(_08055_),
    .A2(_08048_));
 sg13g2_a22oi_1 _24667_ (.Y(_08056_),
    .B1(_07646_),
    .B2(\top_ihp.oisc.regs[9][30] ),
    .A2(net837),
    .A1(\top_ihp.oisc.regs[32][30] ));
 sg13g2_a22oi_1 _24668_ (.Y(_08057_),
    .B1(net804),
    .B2(\top_ihp.oisc.regs[10][30] ),
    .A2(_07609_),
    .A1(\top_ihp.oisc.regs[14][30] ));
 sg13g2_a221oi_1 _24669_ (.B2(\top_ihp.oisc.regs[13][30] ),
    .C1(_07612_),
    .B1(_07618_),
    .A1(\top_ihp.oisc.regs[11][30] ),
    .Y(_08058_),
    .A2(_07623_));
 sg13g2_nand3_1 _24670_ (.B(_08057_),
    .C(_08058_),
    .A(_08056_),
    .Y(_08059_));
 sg13g2_a21oi_1 _24671_ (.A1(\top_ihp.oisc.regs[4][30] ),
    .A2(_07594_),
    .Y(_08060_),
    .B1(_08059_));
 sg13g2_a221oi_1 _24672_ (.B2(_08060_),
    .C1(_07718_),
    .B1(_08055_),
    .A1(_00076_),
    .Y(_08061_),
    .A2(net849));
 sg13g2_nor2_1 _24673_ (.A(net718),
    .B(_08061_),
    .Y(_08062_));
 sg13g2_a21oi_1 _24674_ (.A1(_08549_),
    .A2(net665),
    .Y(_00475_),
    .B1(_08062_));
 sg13g2_mux2_1 _24675_ (.A0(\top_ihp.oisc.regs[7][31] ),
    .A1(\top_ihp.oisc.regs[3][31] ),
    .S(_07639_),
    .X(_08063_));
 sg13g2_nand2_1 _24676_ (.Y(_08064_),
    .A(\top_ihp.oisc.regs[2][31] ),
    .B(net803));
 sg13g2_o21ai_1 _24677_ (.B1(_08064_),
    .Y(_08065_),
    .A1(_03617_),
    .A2(net776));
 sg13g2_a22oi_1 _24678_ (.Y(_08066_),
    .B1(_08065_),
    .B2(_07582_),
    .A2(_08063_),
    .A1(net809));
 sg13g2_mux2_1 _24679_ (.A0(\top_ihp.oisc.regs[5][31] ),
    .A1(\top_ihp.oisc.regs[1][31] ),
    .S(_07704_),
    .X(_08067_));
 sg13g2_nand2_1 _24680_ (.Y(_08068_),
    .A(_07733_),
    .B(_08067_));
 sg13g2_a22oi_1 _24681_ (.Y(_08069_),
    .B1(_07590_),
    .B2(\top_ihp.oisc.regs[15][31] ),
    .A2(_07678_),
    .A1(\top_ihp.oisc.regs[11][31] ));
 sg13g2_nor2_1 _24682_ (.A(_00077_),
    .B(_07674_),
    .Y(_08070_));
 sg13g2_a221oi_1 _24683_ (.B2(\top_ihp.oisc.regs[10][31] ),
    .C1(_08070_),
    .B1(_07682_),
    .A1(\top_ihp.oisc.regs[8][31] ),
    .Y(_08071_),
    .A2(net852));
 sg13g2_nand4_1 _24684_ (.B(_08068_),
    .C(_08069_),
    .A(_08066_),
    .Y(_08072_),
    .D(_08071_));
 sg13g2_nand2_1 _24685_ (.Y(_08073_),
    .A(\top_ihp.oisc.regs[4][31] ),
    .B(_07772_));
 sg13g2_a22oi_1 _24686_ (.Y(_08074_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][31] ),
    .A2(_07691_),
    .A1(\top_ihp.oisc.regs[12][31] ));
 sg13g2_nand2b_1 _24687_ (.Y(_08075_),
    .B(_07695_),
    .A_N(_08074_));
 sg13g2_nand2_1 _24688_ (.Y(_08076_),
    .A(\top_ihp.oisc.regs[9][31] ),
    .B(_07716_));
 sg13g2_a22oi_1 _24689_ (.Y(_08077_),
    .B1(_07720_),
    .B2(\top_ihp.oisc.regs[13][31] ),
    .A2(_07795_),
    .A1(\top_ihp.oisc.regs[32][31] ));
 sg13g2_nand4_1 _24690_ (.B(_08075_),
    .C(_08076_),
    .A(_08073_),
    .Y(_08078_),
    .D(_08077_));
 sg13g2_nor2_1 _24691_ (.A(_08072_),
    .B(_08078_),
    .Y(_08079_));
 sg13g2_nand2_1 _24692_ (.Y(_08080_),
    .A(\top_ihp.oisc.op_b[31] ),
    .B(net664));
 sg13g2_o21ai_1 _24693_ (.B1(_08080_),
    .Y(_00476_),
    .A1(net741),
    .A2(_08079_));
 sg13g2_mux2_1 _24694_ (.A0(\top_ihp.oisc.regs[7][3] ),
    .A1(\top_ihp.oisc.regs[3][3] ),
    .S(net807),
    .X(_08081_));
 sg13g2_mux2_1 _24695_ (.A0(\top_ihp.oisc.regs[6][3] ),
    .A1(\top_ihp.oisc.regs[2][3] ),
    .S(net808),
    .X(_08082_));
 sg13g2_a22oi_1 _24696_ (.Y(_08083_),
    .B1(_08082_),
    .B2(net853),
    .A2(_08081_),
    .A1(net809));
 sg13g2_mux2_1 _24697_ (.A0(\top_ihp.oisc.regs[5][3] ),
    .A1(\top_ihp.oisc.regs[1][3] ),
    .S(net802),
    .X(_08084_));
 sg13g2_nand2_1 _24698_ (.Y(_08085_),
    .A(net834),
    .B(_08084_));
 sg13g2_a22oi_1 _24699_ (.Y(_08086_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][3] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][3] ));
 sg13g2_nor2_1 _24700_ (.A(_00244_),
    .B(net851),
    .Y(_08087_));
 sg13g2_a221oi_1 _24701_ (.B2(\top_ihp.oisc.regs[10][3] ),
    .C1(_08087_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][3] ),
    .Y(_08088_),
    .A2(net852));
 sg13g2_nand4_1 _24702_ (.B(_08085_),
    .C(_08086_),
    .A(_08083_),
    .Y(_08089_),
    .D(_08088_));
 sg13g2_nand2_1 _24703_ (.Y(_08090_),
    .A(\top_ihp.oisc.regs[4][3] ),
    .B(net764));
 sg13g2_a22oi_1 _24704_ (.Y(_08091_),
    .B1(net835),
    .B2(\top_ihp.oisc.regs[14][3] ),
    .A2(net864),
    .A1(\top_ihp.oisc.regs[12][3] ));
 sg13g2_nand2b_1 _24705_ (.Y(_08092_),
    .B(net893),
    .A_N(_08091_));
 sg13g2_nand2_1 _24706_ (.Y(_08093_),
    .A(\top_ihp.oisc.regs[9][3] ),
    .B(net753));
 sg13g2_a22oi_1 _24707_ (.Y(_08094_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][3] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][3] ));
 sg13g2_nand4_1 _24708_ (.B(_08092_),
    .C(_08093_),
    .A(_08090_),
    .Y(_08095_),
    .D(_08094_));
 sg13g2_nor2_1 _24709_ (.A(_08089_),
    .B(_08095_),
    .Y(_08096_));
 sg13g2_nand2_1 _24710_ (.Y(_08097_),
    .A(_08328_),
    .B(net664));
 sg13g2_o21ai_1 _24711_ (.B1(_08097_),
    .Y(_00477_),
    .A1(net741),
    .A2(_08096_));
 sg13g2_mux2_1 _24712_ (.A0(\top_ihp.oisc.regs[5][4] ),
    .A1(\top_ihp.oisc.regs[1][4] ),
    .S(net772),
    .X(_08098_));
 sg13g2_nand2_1 _24713_ (.Y(_08099_),
    .A(\top_ihp.oisc.regs[11][4] ),
    .B(net773));
 sg13g2_mux2_1 _24714_ (.A0(\top_ihp.oisc.regs[8][4] ),
    .A1(\top_ihp.oisc.regs[12][4] ),
    .S(net985),
    .X(_08100_));
 sg13g2_nand2_1 _24715_ (.Y(_08101_),
    .A(\top_ihp.oisc.regs[32][4] ),
    .B(net837));
 sg13g2_o21ai_1 _24716_ (.B1(_08101_),
    .Y(_08102_),
    .A1(_00245_),
    .A2(_07651_));
 sg13g2_a221oi_1 _24717_ (.B2(net864),
    .C1(_08102_),
    .B1(_08100_),
    .A1(\top_ihp.oisc.regs[13][4] ),
    .Y(_08103_),
    .A2(net765));
 sg13g2_mux2_1 _24718_ (.A0(\top_ihp.oisc.regs[10][4] ),
    .A1(\top_ihp.oisc.regs[14][4] ),
    .S(net985),
    .X(_08104_));
 sg13g2_a22oi_1 _24719_ (.Y(_08105_),
    .B1(net850),
    .B2(_08104_),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[9][4] ));
 sg13g2_a22oi_1 _24720_ (.Y(_08106_),
    .B1(_07841_),
    .B2(\top_ihp.oisc.regs[6][4] ),
    .A2(net775),
    .A1(\top_ihp.oisc.regs[15][4] ));
 sg13g2_nand4_1 _24721_ (.B(_08103_),
    .C(_08105_),
    .A(_08099_),
    .Y(_08107_),
    .D(_08106_));
 sg13g2_a21oi_1 _24722_ (.A1(net839),
    .A2(_08098_),
    .Y(_08108_),
    .B1(_08107_));
 sg13g2_nand3_1 _24723_ (.B(_07571_),
    .C(net865),
    .A(\top_ihp.oisc.regs[2][4] ),
    .Y(_08109_));
 sg13g2_nand3_1 _24724_ (.B(net830),
    .C(_07576_),
    .A(\top_ihp.oisc.regs[7][4] ),
    .Y(_08110_));
 sg13g2_nand2_1 _24725_ (.Y(_08111_),
    .A(_08109_),
    .B(_08110_));
 sg13g2_a221oi_1 _24726_ (.B2(\top_ihp.oisc.regs[3][4] ),
    .C1(_08111_),
    .B1(_07689_),
    .A1(\top_ihp.oisc.regs[4][4] ),
    .Y(_08112_),
    .A2(net769));
 sg13g2_a21oi_1 _24727_ (.A1(_08108_),
    .A2(_08112_),
    .Y(_08113_),
    .B1(net741));
 sg13g2_a21o_1 _24728_ (.A2(net667),
    .A1(_08339_),
    .B1(_08113_),
    .X(_00478_));
 sg13g2_mux2_1 _24729_ (.A0(\top_ihp.oisc.regs[7][5] ),
    .A1(\top_ihp.oisc.regs[3][5] ),
    .S(net807),
    .X(_08114_));
 sg13g2_mux2_1 _24730_ (.A0(\top_ihp.oisc.regs[6][5] ),
    .A1(\top_ihp.oisc.regs[2][5] ),
    .S(net808),
    .X(_08115_));
 sg13g2_a22oi_1 _24731_ (.Y(_08116_),
    .B1(_08115_),
    .B2(net853),
    .A2(_08114_),
    .A1(net806));
 sg13g2_mux2_1 _24732_ (.A0(\top_ihp.oisc.regs[5][5] ),
    .A1(\top_ihp.oisc.regs[1][5] ),
    .S(net802),
    .X(_08117_));
 sg13g2_nand2_1 _24733_ (.Y(_08118_),
    .A(net834),
    .B(_08117_));
 sg13g2_a22oi_1 _24734_ (.Y(_08119_),
    .B1(net757),
    .B2(\top_ihp.oisc.regs[15][5] ),
    .A2(net755),
    .A1(\top_ihp.oisc.regs[11][5] ));
 sg13g2_nor2_1 _24735_ (.A(_00246_),
    .B(net851),
    .Y(_08120_));
 sg13g2_a221oi_1 _24736_ (.B2(\top_ihp.oisc.regs[10][5] ),
    .C1(_08120_),
    .B1(net767),
    .A1(\top_ihp.oisc.regs[8][5] ),
    .Y(_08121_),
    .A2(net852));
 sg13g2_nand4_1 _24737_ (.B(_08118_),
    .C(_08119_),
    .A(_08116_),
    .Y(_08122_),
    .D(_08121_));
 sg13g2_nand2_1 _24738_ (.Y(_08123_),
    .A(\top_ihp.oisc.regs[4][5] ),
    .B(net764));
 sg13g2_a22oi_1 _24739_ (.Y(_08124_),
    .B1(net850),
    .B2(\top_ihp.oisc.regs[14][5] ),
    .A2(net864),
    .A1(\top_ihp.oisc.regs[12][5] ));
 sg13g2_nand2b_1 _24740_ (.Y(_08125_),
    .B(net893),
    .A_N(_08124_));
 sg13g2_nand2_1 _24741_ (.Y(_08126_),
    .A(\top_ihp.oisc.regs[9][5] ),
    .B(net753));
 sg13g2_a22oi_1 _24742_ (.Y(_08127_),
    .B1(net752),
    .B2(\top_ihp.oisc.regs[13][5] ),
    .A2(net799),
    .A1(\top_ihp.oisc.regs[32][5] ));
 sg13g2_nand4_1 _24743_ (.B(_08125_),
    .C(_08126_),
    .A(_08123_),
    .Y(_08128_),
    .D(_08127_));
 sg13g2_nor2_1 _24744_ (.A(_08122_),
    .B(_08128_),
    .Y(_08129_));
 sg13g2_nand2_1 _24745_ (.Y(_08130_),
    .A(_08342_),
    .B(net664));
 sg13g2_o21ai_1 _24746_ (.B1(_08130_),
    .Y(_00479_),
    .A1(net741),
    .A2(_08129_));
 sg13g2_mux2_1 _24747_ (.A0(\top_ihp.oisc.regs[6][6] ),
    .A1(\top_ihp.oisc.regs[2][6] ),
    .S(net807),
    .X(_08131_));
 sg13g2_nand2_1 _24748_ (.Y(_08132_),
    .A(net847),
    .B(_08131_));
 sg13g2_a22oi_1 _24749_ (.Y(_08133_),
    .B1(net754),
    .B2(\top_ihp.oisc.regs[15][6] ),
    .A2(net773),
    .A1(\top_ihp.oisc.regs[11][6] ));
 sg13g2_nand2_1 _24750_ (.Y(_08134_),
    .A(\top_ihp.oisc.regs[12][6] ),
    .B(net838));
 sg13g2_mux2_1 _24751_ (.A0(\top_ihp.oisc.regs[7][6] ),
    .A1(\top_ihp.oisc.regs[3][6] ),
    .S(net810),
    .X(_08135_));
 sg13g2_mux2_1 _24752_ (.A0(\top_ihp.oisc.regs[5][6] ),
    .A1(\top_ihp.oisc.regs[1][6] ),
    .S(net800),
    .X(_08136_));
 sg13g2_a22oi_1 _24753_ (.Y(_08137_),
    .B1(_08136_),
    .B2(net833),
    .A2(_08135_),
    .A1(_07576_));
 sg13g2_nand4_1 _24754_ (.B(_08133_),
    .C(_08134_),
    .A(_08132_),
    .Y(_08138_),
    .D(_08137_));
 sg13g2_nand2_1 _24755_ (.Y(_08139_),
    .A(\top_ihp.oisc.regs[4][6] ),
    .B(net764));
 sg13g2_nand2_1 _24756_ (.Y(_08140_),
    .A(\top_ihp.oisc.regs[32][6] ),
    .B(net766));
 sg13g2_mux2_1 _24757_ (.A0(\top_ihp.oisc.regs[10][6] ),
    .A1(\top_ihp.oisc.regs[14][6] ),
    .S(net985),
    .X(_08141_));
 sg13g2_nor2_1 _24758_ (.A(_00247_),
    .B(_07754_),
    .Y(_08142_));
 sg13g2_a221oi_1 _24759_ (.B2(_08141_),
    .C1(_08142_),
    .B1(net835),
    .A1(\top_ihp.oisc.regs[8][6] ),
    .Y(_08143_),
    .A2(net852));
 sg13g2_a22oi_1 _24760_ (.Y(_08144_),
    .B1(net770),
    .B2(\top_ihp.oisc.regs[13][6] ),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][6] ));
 sg13g2_nand4_1 _24761_ (.B(_08140_),
    .C(_08143_),
    .A(_08139_),
    .Y(_08145_),
    .D(_08144_));
 sg13g2_o21ai_1 _24762_ (.B1(_07633_),
    .Y(_08146_),
    .A1(_08138_),
    .A2(_08145_));
 sg13g2_nand2_1 _24763_ (.Y(_08147_),
    .A(_08366_),
    .B(net664));
 sg13g2_o21ai_1 _24764_ (.B1(_08147_),
    .Y(_00480_),
    .A1(net667),
    .A2(_08146_));
 sg13g2_a22oi_1 _24765_ (.Y(_08148_),
    .B1(net834),
    .B2(\top_ihp.oisc.regs[5][7] ),
    .A2(net847),
    .A1(\top_ihp.oisc.regs[6][7] ));
 sg13g2_nor2_1 _24766_ (.A(_07572_),
    .B(_08148_),
    .Y(_08149_));
 sg13g2_a22oi_1 _24767_ (.Y(_08150_),
    .B1(_07590_),
    .B2(\top_ihp.oisc.regs[15][7] ),
    .A2(net756),
    .A1(\top_ihp.oisc.regs[11][7] ));
 sg13g2_nand2_1 _24768_ (.Y(_08151_),
    .A(\top_ihp.oisc.regs[10][7] ),
    .B(_07681_));
 sg13g2_o21ai_1 _24769_ (.B1(_08151_),
    .Y(_08152_),
    .A1(_00248_),
    .A2(net848));
 sg13g2_a221oi_1 _24770_ (.B2(\top_ihp.oisc.regs[1][7] ),
    .C1(_08152_),
    .B1(_07659_),
    .A1(\top_ihp.oisc.regs[32][7] ),
    .Y(_08153_),
    .A2(_07673_));
 sg13g2_a22oi_1 _24771_ (.Y(_08154_),
    .B1(_07720_),
    .B2(\top_ihp.oisc.regs[13][7] ),
    .A2(net801),
    .A1(\top_ihp.oisc.regs[14][7] ));
 sg13g2_mux2_1 _24772_ (.A0(\top_ihp.oisc.regs[8][7] ),
    .A1(\top_ihp.oisc.regs[12][7] ),
    .S(net935),
    .X(_08155_));
 sg13g2_a22oi_1 _24773_ (.Y(_08156_),
    .B1(_08155_),
    .B2(net863),
    .A2(net768),
    .A1(\top_ihp.oisc.regs[9][7] ));
 sg13g2_nand4_1 _24774_ (.B(_08153_),
    .C(_08154_),
    .A(_08150_),
    .Y(_08157_),
    .D(_08156_));
 sg13g2_and2_1 _24775_ (.A(\top_ihp.oisc.regs[7][7] ),
    .B(net830),
    .X(_08158_));
 sg13g2_a21oi_1 _24776_ (.A1(\top_ihp.oisc.regs[3][7] ),
    .A2(net772),
    .Y(_08159_),
    .B1(_08158_));
 sg13g2_a22oi_1 _24777_ (.Y(_08160_),
    .B1(_07663_),
    .B2(\top_ihp.oisc.regs[2][7] ),
    .A2(net774),
    .A1(\top_ihp.oisc.regs[4][7] ));
 sg13g2_o21ai_1 _24778_ (.B1(_08160_),
    .Y(_08161_),
    .A1(_07688_),
    .A2(_08159_));
 sg13g2_nor3_1 _24779_ (.A(_08149_),
    .B(_08157_),
    .C(_08161_),
    .Y(_08162_));
 sg13g2_nand2_1 _24780_ (.Y(_08163_),
    .A(_08315_),
    .B(_03733_));
 sg13g2_o21ai_1 _24781_ (.B1(_08163_),
    .Y(_00481_),
    .A1(net741),
    .A2(_08162_));
 sg13g2_mux2_1 _24782_ (.A0(\top_ihp.oisc.regs[5][8] ),
    .A1(\top_ihp.oisc.regs[1][8] ),
    .S(_07640_),
    .X(_08164_));
 sg13g2_nand2_1 _24783_ (.Y(_08165_),
    .A(\top_ihp.oisc.regs[11][8] ),
    .B(_07624_));
 sg13g2_mux2_1 _24784_ (.A0(\top_ihp.oisc.regs[8][8] ),
    .A1(\top_ihp.oisc.regs[12][8] ),
    .S(_07642_),
    .X(_08166_));
 sg13g2_nand2_1 _24785_ (.Y(_08167_),
    .A(\top_ihp.oisc.regs[32][8] ),
    .B(_07601_));
 sg13g2_o21ai_1 _24786_ (.B1(_08167_),
    .Y(_08168_),
    .A1(_00249_),
    .A2(_07651_));
 sg13g2_a221oi_1 _24787_ (.B2(net864),
    .C1(_08168_),
    .B1(_08166_),
    .A1(\top_ihp.oisc.regs[13][8] ),
    .Y(_08169_),
    .A2(net765));
 sg13g2_mux2_1 _24788_ (.A0(\top_ihp.oisc.regs[10][8] ),
    .A1(\top_ihp.oisc.regs[14][8] ),
    .S(_07642_),
    .X(_08170_));
 sg13g2_a22oi_1 _24789_ (.Y(_08171_),
    .B1(_07692_),
    .B2(_08170_),
    .A2(net771),
    .A1(\top_ihp.oisc.regs[9][8] ));
 sg13g2_a22oi_1 _24790_ (.Y(_08172_),
    .B1(_07841_),
    .B2(\top_ihp.oisc.regs[6][8] ),
    .A2(_07589_),
    .A1(\top_ihp.oisc.regs[15][8] ));
 sg13g2_nand4_1 _24791_ (.B(_08169_),
    .C(_08171_),
    .A(_08165_),
    .Y(_08173_),
    .D(_08172_));
 sg13g2_a21oi_1 _24792_ (.A1(net839),
    .A2(_08164_),
    .Y(_08174_),
    .B1(_08173_));
 sg13g2_nand3_1 _24793_ (.B(net776),
    .C(net865),
    .A(\top_ihp.oisc.regs[2][8] ),
    .Y(_08175_));
 sg13g2_nand3_1 _24794_ (.B(net830),
    .C(_07576_),
    .A(\top_ihp.oisc.regs[7][8] ),
    .Y(_08176_));
 sg13g2_nand2_1 _24795_ (.Y(_08177_),
    .A(_08175_),
    .B(_08176_));
 sg13g2_a221oi_1 _24796_ (.B2(\top_ihp.oisc.regs[3][8] ),
    .C1(_08177_),
    .B1(_07689_),
    .A1(\top_ihp.oisc.regs[4][8] ),
    .Y(_08178_),
    .A2(_07657_));
 sg13g2_a21oi_1 _24797_ (.A1(_08174_),
    .A2(_08178_),
    .Y(_08179_),
    .B1(_07635_));
 sg13g2_a21o_1 _24798_ (.A2(net667),
    .A1(_08351_),
    .B1(_08179_),
    .X(_00482_));
 sg13g2_mux2_1 _24799_ (.A0(\top_ihp.oisc.regs[7][9] ),
    .A1(\top_ihp.oisc.regs[3][9] ),
    .S(net776),
    .X(_08180_));
 sg13g2_mux2_1 _24800_ (.A0(\top_ihp.oisc.regs[5][9] ),
    .A1(\top_ihp.oisc.regs[1][9] ),
    .S(_07571_),
    .X(_08181_));
 sg13g2_mux2_1 _24801_ (.A0(\top_ihp.oisc.regs[6][9] ),
    .A1(\top_ihp.oisc.regs[2][9] ),
    .S(net810),
    .X(_08182_));
 sg13g2_nand2_1 _24802_ (.Y(_08183_),
    .A(net865),
    .B(_08182_));
 sg13g2_nand2_1 _24803_ (.Y(_08184_),
    .A(\top_ihp.oisc.regs[11][9] ),
    .B(net773));
 sg13g2_a22oi_1 _24804_ (.Y(_08185_),
    .B1(net801),
    .B2(\top_ihp.oisc.regs[14][9] ),
    .A2(net837),
    .A1(\top_ihp.oisc.regs[32][9] ));
 sg13g2_a22oi_1 _24805_ (.Y(_08186_),
    .B1(net775),
    .B2(\top_ihp.oisc.regs[15][9] ),
    .A2(net838),
    .A1(\top_ihp.oisc.regs[12][9] ));
 sg13g2_nand4_1 _24806_ (.B(_08184_),
    .C(_08185_),
    .A(_08183_),
    .Y(_08187_),
    .D(_08186_));
 sg13g2_a221oi_1 _24807_ (.B2(net839),
    .C1(_08187_),
    .B1(_08181_),
    .A1(net809),
    .Y(_08188_),
    .A2(_08180_));
 sg13g2_a22oi_1 _24808_ (.Y(_08189_),
    .B1(net850),
    .B2(\top_ihp.oisc.regs[10][9] ),
    .A2(net864),
    .A1(\top_ihp.oisc.regs[8][9] ));
 sg13g2_nor2_1 _24809_ (.A(_00250_),
    .B(_07651_),
    .Y(_08190_));
 sg13g2_a221oi_1 _24810_ (.B2(\top_ihp.oisc.regs[13][9] ),
    .C1(_08190_),
    .B1(net770),
    .A1(\top_ihp.oisc.regs[9][9] ),
    .Y(_08191_),
    .A2(net771));
 sg13g2_o21ai_1 _24811_ (.B1(_08191_),
    .Y(_08192_),
    .A1(net893),
    .A2(_08189_));
 sg13g2_a21oi_1 _24812_ (.A1(\top_ihp.oisc.regs[4][9] ),
    .A2(net769),
    .Y(_08193_),
    .B1(_08192_));
 sg13g2_a21oi_1 _24813_ (.A1(_08188_),
    .A2(_08193_),
    .Y(_08194_),
    .B1(_07635_));
 sg13g2_a21o_1 _24814_ (.A2(net667),
    .A1(_08354_),
    .B1(_08194_),
    .X(_00483_));
 sg13g2_nor2_1 _24815_ (.A(_09852_),
    .B(_04746_),
    .Y(_00355_));
 sg13g2_mux4_1 _24816_ (.S0(_08818_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ),
    .S1(_08819_),
    .X(_08195_));
 sg13g2_mux4_1 _24817_ (.S0(_08818_),
    .A0(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ),
    .A1(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ),
    .A2(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ),
    .A3(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ),
    .S1(_08819_),
    .X(_08196_));
 sg13g2_mux2_1 _24818_ (.A0(_08195_),
    .A1(_08196_),
    .S(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ),
    .X(_08197_));
 sg13g2_nand2_1 _24819_ (.Y(_08198_),
    .A(_05101_),
    .B(_08815_));
 sg13g2_o21ai_1 _24820_ (.B1(_08198_),
    .Y(_00356_),
    .A1(_08853_),
    .A2(_08197_));
 sg13g2_nor2_1 _24821_ (.A(_04318_),
    .B(net2124),
    .Y(\top_ihp.ram_clk_o ));
 sg13g2_and2_1 _24822_ (.A(net895),
    .B(\top_ihp.wb_emem.cmd[63] ),
    .X(\top_ihp.ram_data_o ));
 sg13g2_nor2_1 _24823_ (.A(net2123),
    .B(\top_ihp.rom_cs_o ),
    .Y(\top_ihp.rom_clk_o ));
 sg13g2_and2_1 _24824_ (.A(_08589_),
    .B(\top_ihp.wb_dati_rom[7] ),
    .X(\top_ihp.rom_data_o ));
 sg13g2_and2_1 _24825_ (.A(net983),
    .B(\top_ihp.wb_dati_spi[31] ),
    .X(\top_ihp.spi_data_o ));
 sg13g2_inv_1 _14598__1 (.Y(net2007),
    .A(clknet_leaf_62_clk));
 sg13g2_buf_1 _24827_ (.A(net1422),
    .X(uio_oe[0]));
 sg13g2_buf_1 _24828_ (.A(net1423),
    .X(uio_oe[1]));
 sg13g2_buf_1 _24829_ (.A(net1424),
    .X(uio_oe[2]));
 sg13g2_buf_1 _24830_ (.A(net1425),
    .X(uio_oe[3]));
 sg13g2_buf_1 _24831_ (.A(net1426),
    .X(uio_oe[4]));
 sg13g2_buf_1 _24832_ (.A(net1427),
    .X(uio_oe[5]));
 sg13g2_buf_1 _24833_ (.A(net1428),
    .X(uio_oe[6]));
 sg13g2_buf_1 _24834_ (.A(net1429),
    .X(uio_oe[7]));
 sg13g2_buf_1 _24835_ (.A(\top_ihp.spi_data_o ),
    .X(net10));
 sg13g2_buf_1 _24836_ (.A(\top_ihp.spi_cs_o_1 ),
    .X(net11));
 sg13g2_buf_1 _24837_ (.A(\top_ihp.spi_cs_o_2 ),
    .X(net12));
 sg13g2_buf_1 _24838_ (.A(\top_ihp.spi_cs_o_3 ),
    .X(net13));
 sg13g2_buf_1 _24839_ (.A(\top_ihp.gpio_o_1 ),
    .X(net14));
 sg13g2_buf_1 _24840_ (.A(\top_ihp.gpio_o_2 ),
    .X(net15));
 sg13g2_buf_1 _24841_ (.A(\top_ihp.gpio_o_3 ),
    .X(net16));
 sg13g2_buf_1 _24842_ (.A(\top_ihp.gpio_o_4 ),
    .X(net17));
 sg13g2_buf_1 _24843_ (.A(\top_ihp.tx ),
    .X(net18));
 sg13g2_buf_1 _24844_ (.A(\top_ihp.rom_clk_o ),
    .X(net19));
 sg13g2_buf_1 _24845_ (.A(\top_ihp.rom_data_o ),
    .X(net20));
 sg13g2_buf_1 _24846_ (.A(\top_ihp.rom_cs_o ),
    .X(net21));
 sg13g2_buf_1 _24847_ (.A(\top_ihp.ram_clk_o ),
    .X(net22));
 sg13g2_buf_1 _24848_ (.A(\top_ihp.ram_data_o ),
    .X(net23));
 sg13g2_buf_1 _24849_ (.A(\top_ihp.ram_cs_o ),
    .X(net24));
 sg13g2_buf_1 _24850_ (.A(\top_ihp.spi_clk_o ),
    .X(net25));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1104),
    .D(_00357_),
    .Q_N(_13621_),
    .Q(\top_ihp.oisc.decoder.decoded[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_00358_),
    .Q_N(_13620_),
    .Q(\top_ihp.oisc.decoder.decoded[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1110),
    .D(_00359_),
    .Q_N(_13619_),
    .Q(\top_ihp.oisc.decoder.decoded[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1110),
    .D(_00360_),
    .Q_N(_13618_),
    .Q(\top_ihp.oisc.decoder.decoded[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1110),
    .D(_00361_),
    .Q_N(_13617_),
    .Q(\top_ihp.oisc.decoder.decoded[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1110),
    .D(_00362_),
    .Q_N(_13616_),
    .Q(\top_ihp.oisc.decoder.decoded[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1110),
    .D(_00363_),
    .Q_N(_00090_),
    .Q(\top_ihp.oisc.decoder.decoded[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1104),
    .D(_00364_),
    .Q_N(_13615_),
    .Q(\top_ihp.oisc.decoder.decoded[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1104),
    .D(_00365_),
    .Q_N(_13614_),
    .Q(\top_ihp.oisc.decoder.decoded[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1104),
    .D(_00366_),
    .Q_N(_13613_),
    .Q(\top_ihp.oisc.decoder.decoded[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1104),
    .D(_00367_),
    .Q_N(_13612_),
    .Q(\top_ihp.oisc.decoder.decoded[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1111),
    .D(_00368_),
    .Q_N(_13611_),
    .Q(\top_ihp.oisc.decoder.decoded[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1104),
    .D(_00369_),
    .Q_N(_13610_),
    .Q(\top_ihp.oisc.decoder.decoded[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.decoded[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1104),
    .D(_00370_),
    .Q_N(_13609_),
    .Q(\top_ihp.oisc.decoder.decoded[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1112),
    .D(_00371_),
    .Q_N(_13608_),
    .Q(\top_ihp.oisc.decoder.instruction[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1112),
    .D(_00372_),
    .Q_N(_13607_),
    .Q(\top_ihp.oisc.decoder.instruction[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1104),
    .D(_00373_),
    .Q_N(_13606_),
    .Q(\top_ihp.oisc.decoder.instruction[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1108),
    .D(_00374_),
    .Q_N(_13605_),
    .Q(\top_ihp.oisc.decoder.instruction[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1105),
    .D(_00375_),
    .Q_N(_00079_),
    .Q(\top_ihp.oisc.decoder.instruction[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1115),
    .D(_00241_),
    .Q_N(_13604_),
    .Q(\top_ihp.oisc.decoder.instruction[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1115),
    .D(_00376_),
    .Q_N(_00237_),
    .Q(\top_ihp.oisc.decoder.instruction[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1115),
    .D(_00377_),
    .Q_N(_00238_),
    .Q(\top_ihp.oisc.decoder.instruction[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1115),
    .D(_00378_),
    .Q_N(_00239_),
    .Q(\top_ihp.oisc.decoder.instruction[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1115),
    .D(_00379_),
    .Q_N(_00240_),
    .Q(\top_ihp.oisc.decoder.instruction[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1105),
    .D(_00380_),
    .Q_N(_13603_),
    .Q(\top_ihp.oisc.decoder.instruction[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1115),
    .D(_00381_),
    .Q_N(_00233_),
    .Q(\top_ihp.oisc.decoder.instruction[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1116),
    .D(_00382_),
    .Q_N(_00234_),
    .Q(\top_ihp.oisc.decoder.instruction[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1112),
    .D(_00383_),
    .Q_N(_00235_),
    .Q(\top_ihp.oisc.decoder.instruction[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1116),
    .D(_00384_),
    .Q_N(_00236_),
    .Q(\top_ihp.oisc.decoder.instruction[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1116),
    .D(_00385_),
    .Q_N(_13602_),
    .Q(\top_ihp.oisc.decoder.instruction[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1115),
    .D(_00386_),
    .Q_N(_13601_),
    .Q(\top_ihp.oisc.decoder.instruction[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net1108),
    .D(_00387_),
    .Q_N(_13600_),
    .Q(\top_ihp.oisc.decoder.instruction[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net1115),
    .D(_00388_),
    .Q_N(_13599_),
    .Q(\top_ihp.oisc.decoder.instruction[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1116),
    .D(_00389_),
    .Q_N(_13598_),
    .Q(\top_ihp.oisc.decoder.instruction[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1112),
    .D(_00390_),
    .Q_N(_13597_),
    .Q(\top_ihp.oisc.decoder.instruction[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1110),
    .D(_00391_),
    .Q_N(_13596_),
    .Q(\top_ihp.oisc.decoder.instruction[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1112),
    .D(_00392_),
    .Q_N(_13595_),
    .Q(\top_ihp.oisc.decoder.instruction[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1112),
    .D(_00393_),
    .Q_N(_13594_),
    .Q(\top_ihp.oisc.decoder.instruction[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.decoder.instruction[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1112),
    .D(_00394_),
    .Q_N(_13622_),
    .Q(\top_ihp.oisc.decoder.instruction[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net1430),
    .D(\top_ihp.oisc.wb_adr_o[0] ),
    .Q_N(_13623_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1431),
    .D(\top_ihp.oisc.wb_adr_o[1] ),
    .Q_N(_13593_),
    .Q(\top_ihp.oisc.mem_addr_lowbits[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1101),
    .D(_00395_),
    .Q_N(_13592_),
    .Q(\top_ihp.oisc.micro_op[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1138),
    .D(_00396_),
    .Q_N(_13591_),
    .Q(\top_ihp.oisc.micro_op[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1113),
    .D(_00397_),
    .Q_N(_13590_),
    .Q(\top_ihp.oisc.micro_op[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1102),
    .D(_00398_),
    .Q_N(_13589_),
    .Q(\top_ihp.oisc.micro_op[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1105),
    .D(_00399_),
    .Q_N(_13588_),
    .Q(\top_ihp.oisc.micro_op[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net1105),
    .D(_00400_),
    .Q_N(_13587_),
    .Q(\top_ihp.oisc.micro_op[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1102),
    .D(_00401_),
    .Q_N(_13586_),
    .Q(\top_ihp.oisc.micro_op[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1102),
    .D(_00402_),
    .Q_N(_13585_),
    .Q(\top_ihp.oisc.micro_op[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1103),
    .D(_00403_),
    .Q_N(_13584_),
    .Q(\top_ihp.oisc.micro_op[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1103),
    .D(_00404_),
    .Q_N(_13583_),
    .Q(\top_ihp.oisc.micro_op[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1101),
    .D(_00405_),
    .Q_N(_13582_),
    .Q(\top_ihp.oisc.micro_op[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1101),
    .D(_00406_),
    .Q_N(_13581_),
    .Q(\top_ihp.oisc.micro_op[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1113),
    .D(_00407_),
    .Q_N(_13580_),
    .Q(\top_ihp.oisc.micro_op[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_op[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1105),
    .D(_00408_),
    .Q_N(_13579_),
    .Q(\top_ihp.oisc.micro_op[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[0]$_DFFE_PP_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1432),
    .D(_00409_),
    .Q_N(_00218_),
    .Q(\top_ihp.oisc.micro_pc[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[1]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1433),
    .D(_00410_),
    .Q_N(_00219_),
    .Q(\top_ihp.oisc.micro_pc[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[2]$_DFFE_PP_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1434),
    .D(_00411_),
    .Q_N(_00217_),
    .Q(\top_ihp.oisc.micro_pc[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[3]$_DFFE_PP_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1435),
    .D(_00412_),
    .Q_N(_00216_),
    .Q(\top_ihp.oisc.micro_pc[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[4]$_DFFE_PP_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1436),
    .D(_00413_),
    .Q_N(_00215_),
    .Q(\top_ihp.oisc.micro_pc[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[5]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1437),
    .D(_00414_),
    .Q_N(_00214_),
    .Q(\top_ihp.oisc.micro_pc[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[6]$_DFFE_PP_  (.CLK(clknet_leaf_324_clk),
    .RESET_B(net1438),
    .D(_00415_),
    .Q_N(_00213_),
    .Q(\top_ihp.oisc.micro_pc[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_pc[7]$_DFFE_PP_  (.CLK(clknet_leaf_325_clk),
    .RESET_B(net1439),
    .D(_00416_),
    .Q_N(_00212_),
    .Q(\top_ihp.oisc.micro_pc[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[0]$_DFF_PN0_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1140),
    .D(\top_ihp.oisc.reg_rb[0] ),
    .Q_N(_13624_),
    .Q(\top_ihp.oisc.micro_res_addr[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[1]$_DFF_PN0_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1140),
    .D(\top_ihp.oisc.reg_rb[1] ),
    .Q_N(_13625_),
    .Q(\top_ihp.oisc.micro_res_addr[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[2]$_DFF_PN0_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1326),
    .D(\top_ihp.oisc.reg_rb[2] ),
    .Q_N(_13626_),
    .Q(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_res_addr[3]$_DFF_PN0_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1140),
    .D(\top_ihp.oisc.reg_rb[3] ),
    .Q_N(_13578_),
    .Q(\top_ihp.oisc.micro_res_addr[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1110),
    .D(_00417_),
    .Q_N(\top_ihp.oisc.micro_state[0] ),
    .Q(_13698_));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_323_clk),
    .RESET_B(net1113),
    .D(_00418_),
    .Q_N(_13577_),
    .Q(\top_ihp.oisc.micro_state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.micro_state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1110),
    .D(_00419_),
    .Q_N(_13576_),
    .Q(\top_ihp.oisc.micro_state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1326),
    .D(_00420_),
    .Q_N(_13575_),
    .Q(\top_ihp.oisc.op_a[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1326),
    .D(_00421_),
    .Q_N(_13574_),
    .Q(\top_ihp.oisc.op_a[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1158),
    .D(_00422_),
    .Q_N(_13573_),
    .Q(\top_ihp.oisc.op_a[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1330),
    .D(_00423_),
    .Q_N(_13572_),
    .Q(\top_ihp.oisc.op_a[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1314),
    .D(_00424_),
    .Q_N(_13571_),
    .Q(\top_ihp.oisc.op_a[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1236),
    .D(_00425_),
    .Q_N(_13570_),
    .Q(\top_ihp.oisc.op_a[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1314),
    .D(_00426_),
    .Q_N(_13569_),
    .Q(\top_ihp.oisc.op_a[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1349),
    .D(_00427_),
    .Q_N(_13568_),
    .Q(\top_ihp.oisc.op_a[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1355),
    .D(_00428_),
    .Q_N(_13567_),
    .Q(\top_ihp.oisc.op_a[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1354),
    .D(_00429_),
    .Q_N(_13566_),
    .Q(\top_ihp.oisc.op_a[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1313),
    .D(_00430_),
    .Q_N(_13565_),
    .Q(\top_ihp.oisc.op_a[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1331),
    .D(_00431_),
    .Q_N(_13564_),
    .Q(\top_ihp.oisc.op_a[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1133),
    .D(_00432_),
    .Q_N(_13563_),
    .Q(\top_ihp.oisc.op_a[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1358),
    .D(_00433_),
    .Q_N(_13562_),
    .Q(\top_ihp.oisc.op_a[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1172),
    .D(_00434_),
    .Q_N(_13561_),
    .Q(\top_ihp.oisc.op_a[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1355),
    .D(_00435_),
    .Q_N(_13560_),
    .Q(\top_ihp.oisc.op_a[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1326),
    .D(_00436_),
    .Q_N(_13559_),
    .Q(\top_ihp.oisc.op_a[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1354),
    .D(_00437_),
    .Q_N(_13558_),
    .Q(\top_ihp.oisc.op_a[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1320),
    .D(_00438_),
    .Q_N(_13557_),
    .Q(\top_ihp.oisc.op_a[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1330),
    .D(_00439_),
    .Q_N(_13556_),
    .Q(\top_ihp.oisc.op_a[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1333),
    .D(_00440_),
    .Q_N(_13555_),
    .Q(\top_ihp.oisc.op_a[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1358),
    .D(_00441_),
    .Q_N(_13554_),
    .Q(\top_ihp.oisc.op_a[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_00442_),
    .Q_N(_13553_),
    .Q(\top_ihp.oisc.op_a[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_00443_),
    .Q_N(_13552_),
    .Q(\top_ihp.oisc.op_a[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1352),
    .D(_00444_),
    .Q_N(_13551_),
    .Q(\top_ihp.oisc.op_a[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1328),
    .D(_00445_),
    .Q_N(_13550_),
    .Q(\top_ihp.oisc.op_a[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1286),
    .D(_00446_),
    .Q_N(_13549_),
    .Q(\top_ihp.oisc.op_a[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1287),
    .D(_00447_),
    .Q_N(_13548_),
    .Q(\top_ihp.oisc.op_a[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1326),
    .D(_00448_),
    .Q_N(_13547_),
    .Q(\top_ihp.oisc.op_a[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1331),
    .D(_00449_),
    .Q_N(_13546_),
    .Q(\top_ihp.oisc.op_a[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1209),
    .D(_00450_),
    .Q_N(_13545_),
    .Q(\top_ihp.oisc.op_a[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_a[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1268),
    .D(_00451_),
    .Q_N(_13544_),
    .Q(\top_ihp.oisc.op_a[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[0]$_DFFE_PN0N_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1292),
    .D(_00452_),
    .Q_N(_13543_),
    .Q(\top_ihp.oisc.op_b[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[10]$_DFFE_PN0N_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1292),
    .D(_00453_),
    .Q_N(_13542_),
    .Q(\top_ihp.oisc.op_b[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[11]$_DFFE_PN0N_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1292),
    .D(_00454_),
    .Q_N(_13541_),
    .Q(\top_ihp.oisc.op_b[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[12]$_DFFE_PN0N_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1315),
    .D(_00455_),
    .Q_N(_13540_),
    .Q(\top_ihp.oisc.op_b[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[13]$_DFFE_PN0N_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1315),
    .D(_00456_),
    .Q_N(_13539_),
    .Q(\top_ihp.oisc.op_b[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[14]$_DFFE_PN0N_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1312),
    .D(_00457_),
    .Q_N(_13538_),
    .Q(\top_ihp.oisc.op_b[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[15]$_DFFE_PN0N_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1312),
    .D(_00458_),
    .Q_N(_13537_),
    .Q(\top_ihp.oisc.op_b[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[16]$_DFFE_PN0N_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1316),
    .D(_00459_),
    .Q_N(_13536_),
    .Q(\top_ihp.oisc.op_b[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[17]$_DFFE_PN0N_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1316),
    .D(_00460_),
    .Q_N(_13535_),
    .Q(\top_ihp.oisc.op_b[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[18]$_DFFE_PN0N_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1320),
    .D(_00461_),
    .Q_N(_13534_),
    .Q(\top_ihp.oisc.op_b[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[19]$_DFFE_PN0N_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1315),
    .D(_00462_),
    .Q_N(_13533_),
    .Q(\top_ihp.oisc.op_b[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[1]$_DFFE_PN0N_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1331),
    .D(_00463_),
    .Q_N(_13532_),
    .Q(\top_ihp.oisc.op_b[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[20]$_DFFE_PN0N_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1307),
    .D(_00464_),
    .Q_N(_13531_),
    .Q(\top_ihp.oisc.op_b[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[21]$_DFFE_PN0N_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1320),
    .D(_00465_),
    .Q_N(_13530_),
    .Q(\top_ihp.oisc.op_b[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[22]$_DFFE_PN0N_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1318),
    .D(_00466_),
    .Q_N(_13529_),
    .Q(\top_ihp.oisc.op_b[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[23]$_DFFE_PN0N_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1320),
    .D(_00467_),
    .Q_N(_13528_),
    .Q(\top_ihp.oisc.op_b[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[24]$_DFFE_PN0N_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1320),
    .D(_00468_),
    .Q_N(_13527_),
    .Q(\top_ihp.oisc.op_b[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[25]$_DFFE_PN0N_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1320),
    .D(_00469_),
    .Q_N(_13526_),
    .Q(\top_ihp.oisc.op_b[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[26]$_DFFE_PN0N_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1172),
    .D(_00470_),
    .Q_N(_13525_),
    .Q(\top_ihp.oisc.op_b[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[27]$_DFFE_PN0N_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1292),
    .D(_00471_),
    .Q_N(_13524_),
    .Q(\top_ihp.oisc.op_b[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[28]$_DFFE_PN0N_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1314),
    .D(_00472_),
    .Q_N(_13523_),
    .Q(\top_ihp.oisc.op_b[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[29]$_DFFE_PN0N_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1314),
    .D(_00473_),
    .Q_N(_13522_),
    .Q(\top_ihp.oisc.op_b[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[2]$_DFFE_PN0N_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1313),
    .D(_00474_),
    .Q_N(_13521_),
    .Q(\top_ihp.oisc.op_b[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[30]$_DFFE_PN0N_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_00475_),
    .Q_N(_13520_),
    .Q(\top_ihp.oisc.op_b[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[31]$_DFFE_PN0N_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1315),
    .D(_00476_),
    .Q_N(_13519_),
    .Q(\top_ihp.oisc.op_b[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[3]$_DFFE_PN0N_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1287),
    .D(_00477_),
    .Q_N(_13518_),
    .Q(\top_ihp.oisc.op_b[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[4]$_DFFE_PN0N_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1330),
    .D(_00478_),
    .Q_N(_13517_),
    .Q(\top_ihp.oisc.op_b[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[5]$_DFFE_PN0N_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1292),
    .D(_00479_),
    .Q_N(_13516_),
    .Q(\top_ihp.oisc.op_b[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[6]$_DFFE_PN0N_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1293),
    .D(_00480_),
    .Q_N(_13515_),
    .Q(\top_ihp.oisc.op_b[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[7]$_DFFE_PN0N_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1348),
    .D(_00481_),
    .Q_N(_13514_),
    .Q(\top_ihp.oisc.op_b[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[8]$_DFFE_PN0N_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1293),
    .D(_00482_),
    .Q_N(_13513_),
    .Q(\top_ihp.oisc.op_b[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.op_b[9]$_DFFE_PN0N_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1330),
    .D(_00483_),
    .Q_N(_13512_),
    .Q(\top_ihp.oisc.op_b[9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1326),
    .D(_00484_),
    .Q_N(_13511_),
    .Q(\top_ihp.oisc.regs[0][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1325),
    .D(_00485_),
    .Q_N(_00251_),
    .Q(\top_ihp.oisc.regs[0][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1330),
    .D(_00486_),
    .Q_N(_00252_),
    .Q(\top_ihp.oisc.regs[0][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1330),
    .D(_00487_),
    .Q_N(_00253_),
    .Q(\top_ihp.oisc.regs[0][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1349),
    .D(_00488_),
    .Q_N(_00254_),
    .Q(\top_ihp.oisc.regs[0][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1349),
    .D(_00489_),
    .Q_N(_00255_),
    .Q(\top_ihp.oisc.regs[0][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1349),
    .D(_00490_),
    .Q_N(_00256_),
    .Q(\top_ihp.oisc.regs[0][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1350),
    .D(_00491_),
    .Q_N(_00257_),
    .Q(\top_ihp.oisc.regs[0][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1354),
    .D(_00492_),
    .Q_N(_00258_),
    .Q(\top_ihp.oisc.regs[0][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1354),
    .D(_00493_),
    .Q_N(_00259_),
    .Q(\top_ihp.oisc.regs[0][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1330),
    .D(_00494_),
    .Q_N(_00260_),
    .Q(\top_ihp.oisc.regs[0][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1331),
    .D(_00495_),
    .Q_N(_00242_),
    .Q(\top_ihp.oisc.regs[0][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1354),
    .D(_00496_),
    .Q_N(_00261_),
    .Q(\top_ihp.oisc.regs[0][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1357),
    .D(_00497_),
    .Q_N(_00262_),
    .Q(\top_ihp.oisc.regs[0][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1357),
    .D(_00498_),
    .Q_N(_00263_),
    .Q(\top_ihp.oisc.regs[0][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1357),
    .D(_00499_),
    .Q_N(_00069_),
    .Q(\top_ihp.oisc.regs[0][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1325),
    .D(_00500_),
    .Q_N(_00070_),
    .Q(\top_ihp.oisc.regs[0][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1354),
    .D(_00501_),
    .Q_N(_00071_),
    .Q(\top_ihp.oisc.regs[0][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1354),
    .D(_00502_),
    .Q_N(_00072_),
    .Q(\top_ihp.oisc.regs[0][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1330),
    .D(_00503_),
    .Q_N(_00073_),
    .Q(\top_ihp.oisc.regs[0][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1331),
    .D(_00504_),
    .Q_N(_00074_),
    .Q(\top_ihp.oisc.regs[0][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1350),
    .D(_00505_),
    .Q_N(_00075_),
    .Q(\top_ihp.oisc.regs[0][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1348),
    .D(_00506_),
    .Q_N(_00243_),
    .Q(\top_ihp.oisc.regs[0][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1349),
    .D(_00507_),
    .Q_N(_00076_),
    .Q(\top_ihp.oisc.regs[0][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1349),
    .D(_00508_),
    .Q_N(_00077_),
    .Q(\top_ihp.oisc.regs[0][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1325),
    .D(_00509_),
    .Q_N(_00244_),
    .Q(\top_ihp.oisc.regs[0][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1325),
    .D(_00510_),
    .Q_N(_00245_),
    .Q(\top_ihp.oisc.regs[0][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1328),
    .D(_00511_),
    .Q_N(_00246_),
    .Q(\top_ihp.oisc.regs[0][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1327),
    .D(_00512_),
    .Q_N(_00247_),
    .Q(\top_ihp.oisc.regs[0][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1349),
    .D(_00513_),
    .Q_N(_00248_),
    .Q(\top_ihp.oisc.regs[0][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1331),
    .D(_00514_),
    .Q_N(_00249_),
    .Q(\top_ihp.oisc.regs[0][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[0][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1327),
    .D(_00515_),
    .Q_N(_00250_),
    .Q(\top_ihp.oisc.regs[0][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1378),
    .D(_00516_),
    .Q_N(\top_ihp.oisc.regs[10][0] ),
    .Q(_00267_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1384),
    .D(_00517_),
    .Q_N(_13510_),
    .Q(\top_ihp.oisc.regs[10][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1389),
    .D(_00518_),
    .Q_N(_13509_),
    .Q(\top_ihp.oisc.regs[10][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1344),
    .D(_00519_),
    .Q_N(_13508_),
    .Q(\top_ihp.oisc.regs[10][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1405),
    .D(_00520_),
    .Q_N(_13507_),
    .Q(\top_ihp.oisc.regs[10][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1396),
    .D(_00521_),
    .Q_N(_13506_),
    .Q(\top_ihp.oisc.regs[10][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1396),
    .D(_00522_),
    .Q_N(_13505_),
    .Q(\top_ihp.oisc.regs[10][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1351),
    .D(_00523_),
    .Q_N(_13504_),
    .Q(\top_ihp.oisc.regs[10][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1367),
    .D(_00524_),
    .Q_N(_13503_),
    .Q(\top_ihp.oisc.regs[10][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1369),
    .D(_00525_),
    .Q_N(_13502_),
    .Q(\top_ihp.oisc.regs[10][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1342),
    .D(_00526_),
    .Q_N(_13501_),
    .Q(\top_ihp.oisc.regs[10][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1379),
    .D(_00527_),
    .Q_N(_13500_),
    .Q(\top_ihp.oisc.regs[10][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1395),
    .D(_00528_),
    .Q_N(_13499_),
    .Q(\top_ihp.oisc.regs[10][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1400),
    .D(_00529_),
    .Q_N(_13498_),
    .Q(\top_ihp.oisc.regs[10][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1411),
    .D(_00530_),
    .Q_N(_13497_),
    .Q(\top_ihp.oisc.regs[10][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1401),
    .D(_00531_),
    .Q_N(_13496_),
    .Q(\top_ihp.oisc.regs[10][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1339),
    .D(_00532_),
    .Q_N(_13495_),
    .Q(\top_ihp.oisc.regs[10][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1395),
    .D(_00533_),
    .Q_N(_13494_),
    .Q(\top_ihp.oisc.regs[10][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1396),
    .D(_00534_),
    .Q_N(_13493_),
    .Q(\top_ihp.oisc.regs[10][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1380),
    .D(_00535_),
    .Q_N(_13492_),
    .Q(\top_ihp.oisc.regs[10][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1390),
    .D(_00536_),
    .Q_N(_13491_),
    .Q(\top_ihp.oisc.regs[10][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1407),
    .D(_00537_),
    .Q_N(_13490_),
    .Q(\top_ihp.oisc.regs[10][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1395),
    .D(_00538_),
    .Q_N(_13489_),
    .Q(\top_ihp.oisc.regs[10][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1394),
    .D(_00539_),
    .Q_N(_13488_),
    .Q(\top_ihp.oisc.regs[10][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1361),
    .D(_00540_),
    .Q_N(_13487_),
    .Q(\top_ihp.oisc.regs[10][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1336),
    .D(_00541_),
    .Q_N(_13486_),
    .Q(\top_ihp.oisc.regs[10][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1374),
    .D(_00542_),
    .Q_N(_13485_),
    .Q(\top_ihp.oisc.regs[10][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1340),
    .D(_00543_),
    .Q_N(_13484_),
    .Q(\top_ihp.oisc.regs[10][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1383),
    .D(_00544_),
    .Q_N(_13483_),
    .Q(\top_ihp.oisc.regs[10][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1394),
    .D(_00545_),
    .Q_N(_13482_),
    .Q(\top_ihp.oisc.regs[10][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1405),
    .D(_00546_),
    .Q_N(_13481_),
    .Q(\top_ihp.oisc.regs[10][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[10][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1373),
    .D(_00547_),
    .Q_N(_13480_),
    .Q(\top_ihp.oisc.regs[10][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1376),
    .D(_00548_),
    .Q_N(\top_ihp.oisc.regs[11][0] ),
    .Q(_00268_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1384),
    .D(_00549_),
    .Q_N(_13479_),
    .Q(\top_ihp.oisc.regs[11][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1380),
    .D(_00550_),
    .Q_N(_13478_),
    .Q(\top_ihp.oisc.regs[11][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1344),
    .D(_00551_),
    .Q_N(_13477_),
    .Q(\top_ihp.oisc.regs[11][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_00552_),
    .Q_N(_13476_),
    .Q(\top_ihp.oisc.regs[11][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1401),
    .D(_00553_),
    .Q_N(_13475_),
    .Q(\top_ihp.oisc.regs[11][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1402),
    .D(_00554_),
    .Q_N(_13474_),
    .Q(\top_ihp.oisc.regs[11][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1367),
    .D(_00555_),
    .Q_N(_13473_),
    .Q(\top_ihp.oisc.regs[11][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1367),
    .D(_00556_),
    .Q_N(_13472_),
    .Q(\top_ihp.oisc.regs[11][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1400),
    .D(_00557_),
    .Q_N(_13471_),
    .Q(\top_ihp.oisc.regs[11][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1344),
    .D(_00558_),
    .Q_N(_13470_),
    .Q(\top_ihp.oisc.regs[11][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1345),
    .D(_00559_),
    .Q_N(\top_ihp.oisc.regs[11][1] ),
    .Q(_00269_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1396),
    .D(_00560_),
    .Q_N(_13469_),
    .Q(\top_ihp.oisc.regs[11][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1369),
    .D(_00561_),
    .Q_N(_13468_),
    .Q(\top_ihp.oisc.regs[11][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1401),
    .D(_00562_),
    .Q_N(_13467_),
    .Q(\top_ihp.oisc.regs[11][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1401),
    .D(_00563_),
    .Q_N(_13466_),
    .Q(\top_ihp.oisc.regs[11][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1339),
    .D(_00564_),
    .Q_N(_13465_),
    .Q(\top_ihp.oisc.regs[11][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1400),
    .D(_00565_),
    .Q_N(_13464_),
    .Q(\top_ihp.oisc.regs[11][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1395),
    .D(_00566_),
    .Q_N(_13463_),
    .Q(\top_ihp.oisc.regs[11][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1385),
    .D(_00567_),
    .Q_N(_13462_),
    .Q(\top_ihp.oisc.regs[11][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1380),
    .D(_00568_),
    .Q_N(_13461_),
    .Q(\top_ihp.oisc.regs[11][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1401),
    .D(_00569_),
    .Q_N(_13460_),
    .Q(\top_ihp.oisc.regs[11][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1394),
    .D(_00570_),
    .Q_N(\top_ihp.oisc.regs[11][2] ),
    .Q(_00270_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1363),
    .D(_00571_),
    .Q_N(_13459_),
    .Q(\top_ihp.oisc.regs[11][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1342),
    .D(_00572_),
    .Q_N(_13458_),
    .Q(\top_ihp.oisc.regs[11][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1336),
    .D(_00573_),
    .Q_N(\top_ihp.oisc.regs[11][3] ),
    .Q(_00271_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1372),
    .D(_00574_),
    .Q_N(\top_ihp.oisc.regs[11][4] ),
    .Q(_00272_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1336),
    .D(_00575_),
    .Q_N(_13457_),
    .Q(\top_ihp.oisc.regs[11][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1376),
    .D(_00576_),
    .Q_N(_13456_),
    .Q(\top_ihp.oisc.regs[11][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1345),
    .D(_00577_),
    .Q_N(_13455_),
    .Q(\top_ihp.oisc.regs[11][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1405),
    .D(_00578_),
    .Q_N(_13454_),
    .Q(\top_ihp.oisc.regs[11][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[11][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1385),
    .D(_00579_),
    .Q_N(_13453_),
    .Q(\top_ihp.oisc.regs[11][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][0]$_DFFE_PN1P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1376),
    .D(_00580_),
    .Q_N(\top_ihp.oisc.regs[12][0] ),
    .Q(_00273_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1375),
    .D(_00581_),
    .Q_N(\top_ihp.oisc.regs[12][10] ),
    .Q(_00274_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1378),
    .D(_00582_),
    .Q_N(\top_ihp.oisc.regs[12][11] ),
    .Q(_00275_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1332),
    .D(_00583_),
    .Q_N(\top_ihp.oisc.regs[12][12] ),
    .Q(_00276_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_00584_),
    .Q_N(\top_ihp.oisc.regs[12][13] ),
    .Q(_00277_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1402),
    .D(_00585_),
    .Q_N(\top_ihp.oisc.regs[12][14] ),
    .Q(_00278_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1399),
    .D(_00586_),
    .Q_N(\top_ihp.oisc.regs[12][15] ),
    .Q(_00279_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1333),
    .D(_00587_),
    .Q_N(\top_ihp.oisc.regs[12][16] ),
    .Q(_00280_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1367),
    .D(_00588_),
    .Q_N(\top_ihp.oisc.regs[12][17] ),
    .Q(_00281_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1368),
    .D(_00589_),
    .Q_N(\top_ihp.oisc.regs[12][18] ),
    .Q(_00282_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1344),
    .D(_00590_),
    .Q_N(\top_ihp.oisc.regs[12][19] ),
    .Q(_00283_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][1]$_DFFE_PN1P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1345),
    .D(_00591_),
    .Q_N(\top_ihp.oisc.regs[12][1] ),
    .Q(_00284_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1413),
    .D(_00592_),
    .Q_N(\top_ihp.oisc.regs[12][20] ),
    .Q(_00285_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1363),
    .D(_00593_),
    .Q_N(\top_ihp.oisc.regs[12][21] ),
    .Q(_00286_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1413),
    .D(_00594_),
    .Q_N(\top_ihp.oisc.regs[12][22] ),
    .Q(_00287_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1399),
    .D(_00595_),
    .Q_N(\top_ihp.oisc.regs[12][23] ),
    .Q(_00288_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1372),
    .D(_00596_),
    .Q_N(\top_ihp.oisc.regs[12][24] ),
    .Q(_00289_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1368),
    .D(_00597_),
    .Q_N(\top_ihp.oisc.regs[12][25] ),
    .Q(_00290_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1369),
    .D(_00598_),
    .Q_N(\top_ihp.oisc.regs[12][26] ),
    .Q(_00291_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1378),
    .D(_00599_),
    .Q_N(\top_ihp.oisc.regs[12][27] ),
    .Q(_00292_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1391),
    .D(_00600_),
    .Q_N(\top_ihp.oisc.regs[12][28] ),
    .Q(_00293_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1410),
    .D(_00601_),
    .Q_N(\top_ihp.oisc.regs[12][29] ),
    .Q(_00294_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1394),
    .D(_00602_),
    .Q_N(\top_ihp.oisc.regs[12][2] ),
    .Q(_00295_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1345),
    .D(_00603_),
    .Q_N(\top_ihp.oisc.regs[12][30] ),
    .Q(_00296_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1342),
    .D(_00604_),
    .Q_N(\top_ihp.oisc.regs[12][31] ),
    .Q(_00297_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1328),
    .D(_00605_),
    .Q_N(\top_ihp.oisc.regs[12][3] ),
    .Q(_00298_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1339),
    .D(_00606_),
    .Q_N(\top_ihp.oisc.regs[12][4] ),
    .Q(_00299_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1339),
    .D(_00607_),
    .Q_N(\top_ihp.oisc.regs[12][5] ),
    .Q(_00300_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1375),
    .D(_00608_),
    .Q_N(\top_ihp.oisc.regs[12][6] ),
    .Q(_00301_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1410),
    .D(_00609_),
    .Q_N(\top_ihp.oisc.regs[12][7] ),
    .Q(_00302_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1406),
    .D(_00610_),
    .Q_N(\top_ihp.oisc.regs[12][8] ),
    .Q(_00303_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[12][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1375),
    .D(_00611_),
    .Q_N(\top_ihp.oisc.regs[12][9] ),
    .Q(_00304_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1372),
    .D(_00612_),
    .Q_N(_13452_),
    .Q(\top_ihp.oisc.regs[13][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][10]$_DFFE_PN1P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1375),
    .D(_00613_),
    .Q_N(\top_ihp.oisc.regs[13][10] ),
    .Q(_00305_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1344),
    .D(_00614_),
    .Q_N(\top_ihp.oisc.regs[13][11] ),
    .Q(_00306_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][12]$_DFFE_PN1P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1332),
    .D(_00615_),
    .Q_N(\top_ihp.oisc.regs[13][12] ),
    .Q(_00307_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][13]$_DFFE_PN1P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_00616_),
    .Q_N(\top_ihp.oisc.regs[13][13] ),
    .Q(_00308_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][14]$_DFFE_PN1P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1402),
    .D(_00617_),
    .Q_N(\top_ihp.oisc.regs[13][14] ),
    .Q(_00309_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1399),
    .D(_00618_),
    .Q_N(\top_ihp.oisc.regs[13][15] ),
    .Q(_00310_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][16]$_DFFE_PN1P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1352),
    .D(_00619_),
    .Q_N(\top_ihp.oisc.regs[13][16] ),
    .Q(_00311_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][17]$_DFFE_PN1P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1366),
    .D(_00620_),
    .Q_N(\top_ihp.oisc.regs[13][17] ),
    .Q(_00312_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][18]$_DFFE_PN1P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1368),
    .D(_00621_),
    .Q_N(\top_ihp.oisc.regs[13][18] ),
    .Q(_00313_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][19]$_DFFE_PN1P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1344),
    .D(_00622_),
    .Q_N(\top_ihp.oisc.regs[13][19] ),
    .Q(_00314_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1344),
    .D(_00623_),
    .Q_N(_13451_),
    .Q(\top_ihp.oisc.regs[13][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][20]$_DFFE_PN1P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1413),
    .D(_00624_),
    .Q_N(\top_ihp.oisc.regs[13][20] ),
    .Q(_00315_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][21]$_DFFE_PN1P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1363),
    .D(_00625_),
    .Q_N(\top_ihp.oisc.regs[13][21] ),
    .Q(_00316_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][22]$_DFFE_PN1P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1413),
    .D(_00626_),
    .Q_N(\top_ihp.oisc.regs[13][22] ),
    .Q(_00317_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][23]$_DFFE_PN1P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1413),
    .D(_00627_),
    .Q_N(\top_ihp.oisc.regs[13][23] ),
    .Q(_00318_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][24]$_DFFE_PN1P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1372),
    .D(_00628_),
    .Q_N(\top_ihp.oisc.regs[13][24] ),
    .Q(_00319_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][25]$_DFFE_PN1P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1361),
    .D(_00629_),
    .Q_N(\top_ihp.oisc.regs[13][25] ),
    .Q(_00320_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][26]$_DFFE_PN1P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1411),
    .D(_00630_),
    .Q_N(\top_ihp.oisc.regs[13][26] ),
    .Q(_00321_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1385),
    .D(_00631_),
    .Q_N(\top_ihp.oisc.regs[13][27] ),
    .Q(_00322_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][28]$_DFFE_PN1P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1391),
    .D(_00632_),
    .Q_N(\top_ihp.oisc.regs[13][28] ),
    .Q(_00323_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][29]$_DFFE_PN1P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1410),
    .D(_00633_),
    .Q_N(\top_ihp.oisc.regs[13][29] ),
    .Q(_00324_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][2]$_DFFE_PN1P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1397),
    .D(_00634_),
    .Q_N(\top_ihp.oisc.regs[13][2] ),
    .Q(_00325_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1363),
    .D(_00635_),
    .Q_N(\top_ihp.oisc.regs[13][30] ),
    .Q(_00326_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1352),
    .D(_00636_),
    .Q_N(\top_ihp.oisc.regs[13][31] ),
    .Q(_00327_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][3]$_DFFE_PN1P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1328),
    .D(_00637_),
    .Q_N(\top_ihp.oisc.regs[13][3] ),
    .Q(_00328_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][4]$_DFFE_PN1P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1373),
    .D(_00638_),
    .Q_N(\top_ihp.oisc.regs[13][4] ),
    .Q(_00329_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][5]$_DFFE_PN1P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1328),
    .D(_00639_),
    .Q_N(\top_ihp.oisc.regs[13][5] ),
    .Q(_00330_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][6]$_DFFE_PN1P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1338),
    .D(_00640_),
    .Q_N(\top_ihp.oisc.regs[13][6] ),
    .Q(_00331_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][7]$_DFFE_PN1P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1406),
    .D(_00641_),
    .Q_N(\top_ihp.oisc.regs[13][7] ),
    .Q(_00332_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][8]$_DFFE_PN1P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1405),
    .D(_00642_),
    .Q_N(\top_ihp.oisc.regs[13][8] ),
    .Q(_00333_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[13][9]$_DFFE_PN1P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1373),
    .D(_00643_),
    .Q_N(\top_ihp.oisc.regs[13][9] ),
    .Q(_00334_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1374),
    .D(_00644_),
    .Q_N(_13450_),
    .Q(\top_ihp.oisc.regs[14][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1384),
    .D(_00645_),
    .Q_N(_13449_),
    .Q(\top_ihp.oisc.regs[14][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1342),
    .D(_00646_),
    .Q_N(_13448_),
    .Q(\top_ihp.oisc.regs[14][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1341),
    .D(_00647_),
    .Q_N(_13447_),
    .Q(\top_ihp.oisc.regs[14][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1361),
    .D(_00648_),
    .Q_N(_13446_),
    .Q(\top_ihp.oisc.regs[14][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1396),
    .D(_00649_),
    .Q_N(_13445_),
    .Q(\top_ihp.oisc.regs[14][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1351),
    .D(_00650_),
    .Q_N(_13444_),
    .Q(\top_ihp.oisc.regs[14][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1353),
    .D(_00651_),
    .Q_N(_13443_),
    .Q(\top_ihp.oisc.regs[14][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1362),
    .D(_00652_),
    .Q_N(_13442_),
    .Q(\top_ihp.oisc.regs[14][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1364),
    .D(_00653_),
    .Q_N(_13441_),
    .Q(\top_ihp.oisc.regs[14][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1342),
    .D(_00654_),
    .Q_N(_13440_),
    .Q(\top_ihp.oisc.regs[14][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1379),
    .D(_00655_),
    .Q_N(_13439_),
    .Q(\top_ihp.oisc.regs[14][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1396),
    .D(_00656_),
    .Q_N(_13438_),
    .Q(\top_ihp.oisc.regs[14][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1400),
    .D(_00657_),
    .Q_N(_13437_),
    .Q(\top_ihp.oisc.regs[14][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1407),
    .D(_00658_),
    .Q_N(_13436_),
    .Q(\top_ihp.oisc.regs[14][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1400),
    .D(_00659_),
    .Q_N(_13435_),
    .Q(\top_ihp.oisc.regs[14][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1372),
    .D(_00660_),
    .Q_N(_13434_),
    .Q(\top_ihp.oisc.regs[14][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1341),
    .D(_00661_),
    .Q_N(_13433_),
    .Q(\top_ihp.oisc.regs[14][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1407),
    .D(_00662_),
    .Q_N(_13432_),
    .Q(\top_ihp.oisc.regs[14][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1379),
    .D(_00663_),
    .Q_N(_13431_),
    .Q(\top_ihp.oisc.regs[14][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1390),
    .D(_00664_),
    .Q_N(_13430_),
    .Q(\top_ihp.oisc.regs[14][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1407),
    .D(_00665_),
    .Q_N(_13429_),
    .Q(\top_ihp.oisc.regs[14][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1395),
    .D(_00666_),
    .Q_N(_13428_),
    .Q(\top_ihp.oisc.regs[14][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1379),
    .D(_00667_),
    .Q_N(_13427_),
    .Q(\top_ihp.oisc.regs[14][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1361),
    .D(_00668_),
    .Q_N(_13426_),
    .Q(\top_ihp.oisc.regs[14][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1336),
    .D(_00669_),
    .Q_N(_13425_),
    .Q(\top_ihp.oisc.regs[14][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1373),
    .D(_00670_),
    .Q_N(_13424_),
    .Q(\top_ihp.oisc.regs[14][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1340),
    .D(_00671_),
    .Q_N(_13423_),
    .Q(\top_ihp.oisc.regs[14][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1385),
    .D(_00672_),
    .Q_N(_13422_),
    .Q(\top_ihp.oisc.regs[14][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1379),
    .D(_00673_),
    .Q_N(_13421_),
    .Q(\top_ihp.oisc.regs[14][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1405),
    .D(_00674_),
    .Q_N(_13420_),
    .Q(\top_ihp.oisc.regs[14][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[14][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1384),
    .D(_00675_),
    .Q_N(_13419_),
    .Q(\top_ihp.oisc.regs[14][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1374),
    .D(_00676_),
    .Q_N(_13418_),
    .Q(\top_ihp.oisc.regs[15][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1384),
    .D(_00677_),
    .Q_N(_13417_),
    .Q(\top_ihp.oisc.regs[15][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1380),
    .D(_00678_),
    .Q_N(_13416_),
    .Q(\top_ihp.oisc.regs[15][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1341),
    .D(_00679_),
    .Q_N(_13415_),
    .Q(\top_ihp.oisc.regs[15][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1353),
    .D(_00680_),
    .Q_N(_13414_),
    .Q(\top_ihp.oisc.regs[15][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1402),
    .D(_00681_),
    .Q_N(_13413_),
    .Q(\top_ihp.oisc.regs[15][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1395),
    .D(_00682_),
    .Q_N(_13412_),
    .Q(\top_ihp.oisc.regs[15][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1366),
    .D(_00683_),
    .Q_N(_13411_),
    .Q(\top_ihp.oisc.regs[15][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1366),
    .D(_00684_),
    .Q_N(_13410_),
    .Q(\top_ihp.oisc.regs[15][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1400),
    .D(_00685_),
    .Q_N(_13409_),
    .Q(\top_ihp.oisc.regs[15][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1346),
    .D(_00686_),
    .Q_N(_13408_),
    .Q(\top_ihp.oisc.regs[15][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1379),
    .D(_00687_),
    .Q_N(_13407_),
    .Q(\top_ihp.oisc.regs[15][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1403),
    .D(_00688_),
    .Q_N(_13406_),
    .Q(\top_ihp.oisc.regs[15][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1399),
    .D(_00689_),
    .Q_N(_13405_),
    .Q(\top_ihp.oisc.regs[15][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1411),
    .D(_00690_),
    .Q_N(_13404_),
    .Q(\top_ihp.oisc.regs[15][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1399),
    .D(_00691_),
    .Q_N(_13403_),
    .Q(\top_ihp.oisc.regs[15][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1372),
    .D(_00692_),
    .Q_N(_13402_),
    .Q(\top_ihp.oisc.regs[15][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1368),
    .D(_00693_),
    .Q_N(_13401_),
    .Q(\top_ihp.oisc.regs[15][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1411),
    .D(_00694_),
    .Q_N(_13400_),
    .Q(\top_ihp.oisc.regs[15][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1389),
    .D(_00695_),
    .Q_N(_13399_),
    .Q(\top_ihp.oisc.regs[15][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1390),
    .D(_00696_),
    .Q_N(_13398_),
    .Q(\top_ihp.oisc.regs[15][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1411),
    .D(_00697_),
    .Q_N(_13397_),
    .Q(\top_ihp.oisc.regs[15][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1394),
    .D(_00698_),
    .Q_N(_13396_),
    .Q(\top_ihp.oisc.regs[15][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1345),
    .D(_00699_),
    .Q_N(_13395_),
    .Q(\top_ihp.oisc.regs[15][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1342),
    .D(_00700_),
    .Q_N(_13394_),
    .Q(\top_ihp.oisc.regs[15][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1336),
    .D(_00701_),
    .Q_N(_13393_),
    .Q(\top_ihp.oisc.regs[15][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1373),
    .D(_00702_),
    .Q_N(_13392_),
    .Q(\top_ihp.oisc.regs[15][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1336),
    .D(_00703_),
    .Q_N(_13391_),
    .Q(\top_ihp.oisc.regs[15][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1385),
    .D(_00704_),
    .Q_N(_13390_),
    .Q(\top_ihp.oisc.regs[15][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1346),
    .D(_00705_),
    .Q_N(_13389_),
    .Q(\top_ihp.oisc.regs[15][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1390),
    .D(_00706_),
    .Q_N(_13388_),
    .Q(\top_ihp.oisc.regs[15][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[15][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1373),
    .D(_00707_),
    .Q_N(_13387_),
    .Q(\top_ihp.oisc.regs[15][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][0]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1440),
    .D(_00708_),
    .Q_N(_13386_),
    .Q(\top_ihp.oisc.regs[16][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][10]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1441),
    .D(_00709_),
    .Q_N(_13385_),
    .Q(\top_ihp.oisc.regs[16][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1442),
    .D(_00710_),
    .Q_N(_13384_),
    .Q(\top_ihp.oisc.regs[16][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][12]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1443),
    .D(_00711_),
    .Q_N(_13383_),
    .Q(\top_ihp.oisc.regs[16][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1444),
    .D(_00712_),
    .Q_N(_13382_),
    .Q(\top_ihp.oisc.regs[16][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][14]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1445),
    .D(_00713_),
    .Q_N(_13381_),
    .Q(\top_ihp.oisc.regs[16][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][15]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1446),
    .D(_00714_),
    .Q_N(_13380_),
    .Q(\top_ihp.oisc.regs[16][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][16]$_DFFE_PP_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1447),
    .D(_00715_),
    .Q_N(_13379_),
    .Q(\top_ihp.oisc.regs[16][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][17]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1448),
    .D(_00716_),
    .Q_N(_13378_),
    .Q(\top_ihp.oisc.regs[16][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][18]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1449),
    .D(_00717_),
    .Q_N(_13377_),
    .Q(\top_ihp.oisc.regs[16][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][19]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1450),
    .D(_00718_),
    .Q_N(_13376_),
    .Q(\top_ihp.oisc.regs[16][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][1]$_DFFE_PP_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1451),
    .D(_00719_),
    .Q_N(_13375_),
    .Q(\top_ihp.oisc.regs[16][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][20]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1452),
    .D(_00720_),
    .Q_N(_13374_),
    .Q(\top_ihp.oisc.regs[16][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][21]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1453),
    .D(_00721_),
    .Q_N(_13373_),
    .Q(\top_ihp.oisc.regs[16][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][22]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1454),
    .D(_00722_),
    .Q_N(_13372_),
    .Q(\top_ihp.oisc.regs[16][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][23]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1455),
    .D(_00723_),
    .Q_N(_13371_),
    .Q(\top_ihp.oisc.regs[16][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][24]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1456),
    .D(_00724_),
    .Q_N(_13370_),
    .Q(\top_ihp.oisc.regs[16][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][25]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1457),
    .D(_00725_),
    .Q_N(_13369_),
    .Q(\top_ihp.oisc.regs[16][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][26]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1458),
    .D(_00726_),
    .Q_N(_13368_),
    .Q(\top_ihp.oisc.regs[16][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][27]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1459),
    .D(_00727_),
    .Q_N(_13367_),
    .Q(\top_ihp.oisc.regs[16][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][28]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1460),
    .D(_00728_),
    .Q_N(_13366_),
    .Q(\top_ihp.oisc.regs[16][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][29]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1461),
    .D(_00729_),
    .Q_N(_13365_),
    .Q(\top_ihp.oisc.regs[16][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1462),
    .D(_00730_),
    .Q_N(_13364_),
    .Q(\top_ihp.oisc.regs[16][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][30]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1463),
    .D(_00731_),
    .Q_N(_13363_),
    .Q(\top_ihp.oisc.regs[16][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][31]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1464),
    .D(_00732_),
    .Q_N(_13362_),
    .Q(\top_ihp.oisc.regs[16][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1465),
    .D(_00733_),
    .Q_N(_13361_),
    .Q(\top_ihp.oisc.regs[16][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][4]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1466),
    .D(_00734_),
    .Q_N(_13360_),
    .Q(\top_ihp.oisc.regs[16][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][5]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1467),
    .D(_00735_),
    .Q_N(_13359_),
    .Q(\top_ihp.oisc.regs[16][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1468),
    .D(_00736_),
    .Q_N(_13358_),
    .Q(\top_ihp.oisc.regs[16][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][7]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1469),
    .D(_00737_),
    .Q_N(_13357_),
    .Q(\top_ihp.oisc.regs[16][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][8]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1470),
    .D(_00738_),
    .Q_N(_13356_),
    .Q(\top_ihp.oisc.regs[16][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[16][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1471),
    .D(_00739_),
    .Q_N(_13355_),
    .Q(\top_ihp.oisc.regs[16][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1472),
    .D(_00740_),
    .Q_N(_13354_),
    .Q(\top_ihp.oisc.regs[17][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][10]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1473),
    .D(_00741_),
    .Q_N(_13353_),
    .Q(\top_ihp.oisc.regs[17][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][11]$_DFFE_PP_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1474),
    .D(_00742_),
    .Q_N(_13352_),
    .Q(\top_ihp.oisc.regs[17][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1475),
    .D(_00743_),
    .Q_N(_13351_),
    .Q(\top_ihp.oisc.regs[17][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][13]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1476),
    .D(_00744_),
    .Q_N(_13350_),
    .Q(\top_ihp.oisc.regs[17][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1477),
    .D(_00745_),
    .Q_N(_13349_),
    .Q(\top_ihp.oisc.regs[17][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][15]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1478),
    .D(_00746_),
    .Q_N(_13348_),
    .Q(\top_ihp.oisc.regs[17][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][16]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1479),
    .D(_00747_),
    .Q_N(_13347_),
    .Q(\top_ihp.oisc.regs[17][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][17]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1480),
    .D(_00748_),
    .Q_N(_13346_),
    .Q(\top_ihp.oisc.regs[17][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][18]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1481),
    .D(_00749_),
    .Q_N(_13345_),
    .Q(\top_ihp.oisc.regs[17][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][19]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1482),
    .D(_00750_),
    .Q_N(_13344_),
    .Q(\top_ihp.oisc.regs[17][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1483),
    .D(_00751_),
    .Q_N(_13343_),
    .Q(\top_ihp.oisc.regs[17][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][20]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1484),
    .D(_00752_),
    .Q_N(_13342_),
    .Q(\top_ihp.oisc.regs[17][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][21]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1485),
    .D(_00753_),
    .Q_N(_13341_),
    .Q(\top_ihp.oisc.regs[17][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][22]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1486),
    .D(_00754_),
    .Q_N(_13340_),
    .Q(\top_ihp.oisc.regs[17][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][23]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1487),
    .D(_00755_),
    .Q_N(_13339_),
    .Q(\top_ihp.oisc.regs[17][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][24]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1488),
    .D(_00756_),
    .Q_N(_13338_),
    .Q(\top_ihp.oisc.regs[17][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][25]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1489),
    .D(_00757_),
    .Q_N(_13337_),
    .Q(\top_ihp.oisc.regs[17][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][26]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1490),
    .D(_00758_),
    .Q_N(_13336_),
    .Q(\top_ihp.oisc.regs[17][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][27]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1491),
    .D(_00759_),
    .Q_N(_13335_),
    .Q(\top_ihp.oisc.regs[17][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][28]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1492),
    .D(_00760_),
    .Q_N(_13334_),
    .Q(\top_ihp.oisc.regs[17][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][29]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1493),
    .D(_00761_),
    .Q_N(_13333_),
    .Q(\top_ihp.oisc.regs[17][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1494),
    .D(_00762_),
    .Q_N(_13332_),
    .Q(\top_ihp.oisc.regs[17][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][30]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1495),
    .D(_00763_),
    .Q_N(_13331_),
    .Q(\top_ihp.oisc.regs[17][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][31]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1496),
    .D(_00764_),
    .Q_N(_13330_),
    .Q(\top_ihp.oisc.regs[17][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][3]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1497),
    .D(_00765_),
    .Q_N(_13329_),
    .Q(\top_ihp.oisc.regs[17][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1498),
    .D(_00766_),
    .Q_N(_13328_),
    .Q(\top_ihp.oisc.regs[17][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][5]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1499),
    .D(_00767_),
    .Q_N(_13327_),
    .Q(\top_ihp.oisc.regs[17][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][6]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1500),
    .D(_00768_),
    .Q_N(_13326_),
    .Q(\top_ihp.oisc.regs[17][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1501),
    .D(_00769_),
    .Q_N(_13325_),
    .Q(\top_ihp.oisc.regs[17][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1502),
    .D(_00770_),
    .Q_N(_13324_),
    .Q(\top_ihp.oisc.regs[17][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[17][9]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1503),
    .D(_00771_),
    .Q_N(_13323_),
    .Q(\top_ihp.oisc.regs[17][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][0]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1504),
    .D(_00772_),
    .Q_N(_13322_),
    .Q(\top_ihp.oisc.regs[18][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][10]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1505),
    .D(_00773_),
    .Q_N(_13321_),
    .Q(\top_ihp.oisc.regs[18][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1506),
    .D(_00774_),
    .Q_N(_13320_),
    .Q(\top_ihp.oisc.regs[18][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][12]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1507),
    .D(_00775_),
    .Q_N(_13319_),
    .Q(\top_ihp.oisc.regs[18][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][13]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1508),
    .D(_00776_),
    .Q_N(_13318_),
    .Q(\top_ihp.oisc.regs[18][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][14]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1509),
    .D(_00777_),
    .Q_N(_13317_),
    .Q(\top_ihp.oisc.regs[18][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][15]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1510),
    .D(_00778_),
    .Q_N(_13316_),
    .Q(\top_ihp.oisc.regs[18][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][16]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1511),
    .D(_00779_),
    .Q_N(_13315_),
    .Q(\top_ihp.oisc.regs[18][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][17]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1512),
    .D(_00780_),
    .Q_N(_13314_),
    .Q(\top_ihp.oisc.regs[18][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1513),
    .D(_00781_),
    .Q_N(_13313_),
    .Q(\top_ihp.oisc.regs[18][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][19]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1514),
    .D(_00782_),
    .Q_N(_13312_),
    .Q(\top_ihp.oisc.regs[18][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1515),
    .D(_00783_),
    .Q_N(_13311_),
    .Q(\top_ihp.oisc.regs[18][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][20]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1516),
    .D(_00784_),
    .Q_N(_13310_),
    .Q(\top_ihp.oisc.regs[18][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][21]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1517),
    .D(_00785_),
    .Q_N(_13309_),
    .Q(\top_ihp.oisc.regs[18][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1518),
    .D(_00786_),
    .Q_N(_13308_),
    .Q(\top_ihp.oisc.regs[18][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][23]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1519),
    .D(_00787_),
    .Q_N(_13307_),
    .Q(\top_ihp.oisc.regs[18][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][24]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1520),
    .D(_00788_),
    .Q_N(_13306_),
    .Q(\top_ihp.oisc.regs[18][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][25]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1521),
    .D(_00789_),
    .Q_N(_13305_),
    .Q(\top_ihp.oisc.regs[18][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][26]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1522),
    .D(_00790_),
    .Q_N(_13304_),
    .Q(\top_ihp.oisc.regs[18][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][27]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1523),
    .D(_00791_),
    .Q_N(_13303_),
    .Q(\top_ihp.oisc.regs[18][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1524),
    .D(_00792_),
    .Q_N(_13302_),
    .Q(\top_ihp.oisc.regs[18][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][29]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1525),
    .D(_00793_),
    .Q_N(_13301_),
    .Q(\top_ihp.oisc.regs[18][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][2]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1526),
    .D(_00794_),
    .Q_N(_13300_),
    .Q(\top_ihp.oisc.regs[18][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][30]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1527),
    .D(_00795_),
    .Q_N(_13299_),
    .Q(\top_ihp.oisc.regs[18][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][31]$_DFFE_PP_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1528),
    .D(_00796_),
    .Q_N(_13298_),
    .Q(\top_ihp.oisc.regs[18][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1529),
    .D(_00797_),
    .Q_N(_13297_),
    .Q(\top_ihp.oisc.regs[18][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][4]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1530),
    .D(_00798_),
    .Q_N(_13296_),
    .Q(\top_ihp.oisc.regs[18][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][5]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1531),
    .D(_00799_),
    .Q_N(_13295_),
    .Q(\top_ihp.oisc.regs[18][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][6]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1532),
    .D(_00800_),
    .Q_N(_13294_),
    .Q(\top_ihp.oisc.regs[18][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][7]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1533),
    .D(_00801_),
    .Q_N(_13293_),
    .Q(\top_ihp.oisc.regs[18][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][8]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1534),
    .D(_00802_),
    .Q_N(_13292_),
    .Q(\top_ihp.oisc.regs[18][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[18][9]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1535),
    .D(_00803_),
    .Q_N(_13291_),
    .Q(\top_ihp.oisc.regs[18][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][0]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1536),
    .D(_00804_),
    .Q_N(_13290_),
    .Q(\top_ihp.oisc.regs[19][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][10]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1537),
    .D(_00805_),
    .Q_N(_13289_),
    .Q(\top_ihp.oisc.regs[19][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1538),
    .D(_00806_),
    .Q_N(_13288_),
    .Q(\top_ihp.oisc.regs[19][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1539),
    .D(_00807_),
    .Q_N(_13287_),
    .Q(\top_ihp.oisc.regs[19][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][13]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1540),
    .D(_00808_),
    .Q_N(_13286_),
    .Q(\top_ihp.oisc.regs[19][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1541),
    .D(_00809_),
    .Q_N(_13285_),
    .Q(\top_ihp.oisc.regs[19][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][15]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1542),
    .D(_00810_),
    .Q_N(_13284_),
    .Q(\top_ihp.oisc.regs[19][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][16]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1543),
    .D(_00811_),
    .Q_N(_13283_),
    .Q(\top_ihp.oisc.regs[19][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][17]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1544),
    .D(_00812_),
    .Q_N(_13282_),
    .Q(\top_ihp.oisc.regs[19][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][18]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1545),
    .D(_00813_),
    .Q_N(_13281_),
    .Q(\top_ihp.oisc.regs[19][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][19]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1546),
    .D(_00814_),
    .Q_N(_13280_),
    .Q(\top_ihp.oisc.regs[19][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][1]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1547),
    .D(_00815_),
    .Q_N(_13279_),
    .Q(\top_ihp.oisc.regs[19][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1548),
    .D(_00816_),
    .Q_N(_13278_),
    .Q(\top_ihp.oisc.regs[19][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][21]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1549),
    .D(_00817_),
    .Q_N(_13277_),
    .Q(\top_ihp.oisc.regs[19][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][22]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1550),
    .D(_00818_),
    .Q_N(_13276_),
    .Q(\top_ihp.oisc.regs[19][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][23]$_DFFE_PP_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1551),
    .D(_00819_),
    .Q_N(_13275_),
    .Q(\top_ihp.oisc.regs[19][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][24]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1552),
    .D(_00820_),
    .Q_N(_13274_),
    .Q(\top_ihp.oisc.regs[19][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][25]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1553),
    .D(_00821_),
    .Q_N(_13273_),
    .Q(\top_ihp.oisc.regs[19][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][26]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1554),
    .D(_00822_),
    .Q_N(_13272_),
    .Q(\top_ihp.oisc.regs[19][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][27]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1555),
    .D(_00823_),
    .Q_N(_13271_),
    .Q(\top_ihp.oisc.regs[19][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][28]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1556),
    .D(_00824_),
    .Q_N(_13270_),
    .Q(\top_ihp.oisc.regs[19][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][29]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1557),
    .D(_00825_),
    .Q_N(_13269_),
    .Q(\top_ihp.oisc.regs[19][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][2]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1558),
    .D(_00826_),
    .Q_N(_13268_),
    .Q(\top_ihp.oisc.regs[19][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][30]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1559),
    .D(_00827_),
    .Q_N(_13267_),
    .Q(\top_ihp.oisc.regs[19][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][31]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1560),
    .D(_00828_),
    .Q_N(_13266_),
    .Q(\top_ihp.oisc.regs[19][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][3]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1561),
    .D(_00829_),
    .Q_N(_13265_),
    .Q(\top_ihp.oisc.regs[19][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1562),
    .D(_00830_),
    .Q_N(_13264_),
    .Q(\top_ihp.oisc.regs[19][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][5]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1563),
    .D(_00831_),
    .Q_N(_13263_),
    .Q(\top_ihp.oisc.regs[19][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][6]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1564),
    .D(_00832_),
    .Q_N(_13262_),
    .Q(\top_ihp.oisc.regs[19][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][7]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1565),
    .D(_00833_),
    .Q_N(_13261_),
    .Q(\top_ihp.oisc.regs[19][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1566),
    .D(_00834_),
    .Q_N(_13260_),
    .Q(\top_ihp.oisc.regs[19][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[19][9]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1567),
    .D(_00835_),
    .Q_N(_13259_),
    .Q(\top_ihp.oisc.regs[19][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1387),
    .D(_00836_),
    .Q_N(_13258_),
    .Q(\top_ihp.oisc.regs[1][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1387),
    .D(_00837_),
    .Q_N(_13257_),
    .Q(\top_ihp.oisc.regs[1][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1391),
    .D(_00838_),
    .Q_N(_13256_),
    .Q(\top_ihp.oisc.regs[1][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1342),
    .D(_00839_),
    .Q_N(_13255_),
    .Q(\top_ihp.oisc.regs[1][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_00840_),
    .Q_N(_13254_),
    .Q(\top_ihp.oisc.regs[1][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1366),
    .D(_00841_),
    .Q_N(_13253_),
    .Q(\top_ihp.oisc.regs[1][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1402),
    .D(_00842_),
    .Q_N(_13252_),
    .Q(\top_ihp.oisc.regs[1][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1367),
    .D(_00843_),
    .Q_N(_13251_),
    .Q(\top_ihp.oisc.regs[1][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1366),
    .D(_00844_),
    .Q_N(_13250_),
    .Q(\top_ihp.oisc.regs[1][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1367),
    .D(_00845_),
    .Q_N(_13249_),
    .Q(\top_ihp.oisc.regs[1][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1341),
    .D(_00846_),
    .Q_N(_13248_),
    .Q(\top_ihp.oisc.regs[1][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1378),
    .D(_00847_),
    .Q_N(_13247_),
    .Q(\top_ihp.oisc.regs[1][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1402),
    .D(_00848_),
    .Q_N(_13246_),
    .Q(\top_ihp.oisc.regs[1][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1366),
    .D(_00849_),
    .Q_N(_13245_),
    .Q(\top_ihp.oisc.regs[1][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1401),
    .D(_00850_),
    .Q_N(_13244_),
    .Q(\top_ihp.oisc.regs[1][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1404),
    .D(_00851_),
    .Q_N(_13243_),
    .Q(\top_ihp.oisc.regs[1][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1339),
    .D(_00852_),
    .Q_N(_13242_),
    .Q(\top_ihp.oisc.regs[1][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1399),
    .D(_00853_),
    .Q_N(_13241_),
    .Q(\top_ihp.oisc.regs[1][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_139_clk),
    .RESET_B(net1368),
    .D(_00854_),
    .Q_N(_13240_),
    .Q(\top_ihp.oisc.regs[1][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1338),
    .D(_00855_),
    .Q_N(_13239_),
    .Q(\top_ihp.oisc.regs[1][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1391),
    .D(_00856_),
    .Q_N(_13238_),
    .Q(\top_ihp.oisc.regs[1][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_143_clk),
    .RESET_B(net1401),
    .D(_00857_),
    .Q_N(_13237_),
    .Q(\top_ihp.oisc.regs[1][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1397),
    .D(_00858_),
    .Q_N(_13236_),
    .Q(\top_ihp.oisc.regs[1][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][30]$_DFFE_PN1P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1345),
    .D(_00859_),
    .Q_N(\top_ihp.oisc.regs[1][30] ),
    .Q(_00335_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1361),
    .D(_00860_),
    .Q_N(_13235_),
    .Q(\top_ihp.oisc.regs[1][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1337),
    .D(_00861_),
    .Q_N(_13234_),
    .Q(\top_ihp.oisc.regs[1][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1391),
    .D(_00862_),
    .Q_N(_13233_),
    .Q(\top_ihp.oisc.regs[1][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1338),
    .D(_00863_),
    .Q_N(_13232_),
    .Q(\top_ihp.oisc.regs[1][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1389),
    .D(_00864_),
    .Q_N(_13231_),
    .Q(\top_ihp.oisc.regs[1][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1394),
    .D(_00865_),
    .Q_N(_13230_),
    .Q(\top_ihp.oisc.regs[1][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1397),
    .D(_00866_),
    .Q_N(_13229_),
    .Q(\top_ihp.oisc.regs[1][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[1][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1387),
    .D(_00867_),
    .Q_N(_13228_),
    .Q(\top_ihp.oisc.regs[1][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][0]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1568),
    .D(_00868_),
    .Q_N(_13227_),
    .Q(\top_ihp.oisc.regs[20][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][10]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1569),
    .D(_00869_),
    .Q_N(_13226_),
    .Q(\top_ihp.oisc.regs[20][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][11]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1570),
    .D(_00870_),
    .Q_N(_13225_),
    .Q(\top_ihp.oisc.regs[20][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][12]$_DFFE_PP_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1571),
    .D(_00871_),
    .Q_N(_13224_),
    .Q(\top_ihp.oisc.regs[20][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][13]$_DFFE_PP_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1572),
    .D(_00872_),
    .Q_N(_13223_),
    .Q(\top_ihp.oisc.regs[20][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1573),
    .D(_00873_),
    .Q_N(_13222_),
    .Q(\top_ihp.oisc.regs[20][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][15]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1574),
    .D(_00874_),
    .Q_N(_13221_),
    .Q(\top_ihp.oisc.regs[20][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][16]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1575),
    .D(_00875_),
    .Q_N(_13220_),
    .Q(\top_ihp.oisc.regs[20][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][17]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1576),
    .D(_00876_),
    .Q_N(_13219_),
    .Q(\top_ihp.oisc.regs[20][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][18]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1577),
    .D(_00877_),
    .Q_N(_13218_),
    .Q(\top_ihp.oisc.regs[20][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][19]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1578),
    .D(_00878_),
    .Q_N(_13217_),
    .Q(\top_ihp.oisc.regs[20][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][1]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1579),
    .D(_00879_),
    .Q_N(_13216_),
    .Q(\top_ihp.oisc.regs[20][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][20]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1580),
    .D(_00880_),
    .Q_N(_13215_),
    .Q(\top_ihp.oisc.regs[20][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][21]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1581),
    .D(_00881_),
    .Q_N(_13214_),
    .Q(\top_ihp.oisc.regs[20][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][22]$_DFFE_PP_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1582),
    .D(_00882_),
    .Q_N(_13213_),
    .Q(\top_ihp.oisc.regs[20][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][23]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1583),
    .D(_00883_),
    .Q_N(_13212_),
    .Q(\top_ihp.oisc.regs[20][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][24]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1584),
    .D(_00884_),
    .Q_N(_13211_),
    .Q(\top_ihp.oisc.regs[20][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][25]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1585),
    .D(_00885_),
    .Q_N(_13210_),
    .Q(\top_ihp.oisc.regs[20][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][26]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1586),
    .D(_00886_),
    .Q_N(_13209_),
    .Q(\top_ihp.oisc.regs[20][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][27]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1587),
    .D(_00887_),
    .Q_N(_13208_),
    .Q(\top_ihp.oisc.regs[20][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][28]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1588),
    .D(_00888_),
    .Q_N(_13207_),
    .Q(\top_ihp.oisc.regs[20][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][29]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1589),
    .D(_00889_),
    .Q_N(_13206_),
    .Q(\top_ihp.oisc.regs[20][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][2]$_DFFE_PP_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1590),
    .D(_00890_),
    .Q_N(_13205_),
    .Q(\top_ihp.oisc.regs[20][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][30]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1591),
    .D(_00891_),
    .Q_N(_13204_),
    .Q(\top_ihp.oisc.regs[20][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][31]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1592),
    .D(_00892_),
    .Q_N(_13203_),
    .Q(\top_ihp.oisc.regs[20][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][3]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1593),
    .D(_00893_),
    .Q_N(_13202_),
    .Q(\top_ihp.oisc.regs[20][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][4]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1594),
    .D(_00894_),
    .Q_N(_13201_),
    .Q(\top_ihp.oisc.regs[20][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][5]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1595),
    .D(_00895_),
    .Q_N(_13200_),
    .Q(\top_ihp.oisc.regs[20][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][6]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1596),
    .D(_00896_),
    .Q_N(_13199_),
    .Q(\top_ihp.oisc.regs[20][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][7]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1597),
    .D(_00897_),
    .Q_N(_13198_),
    .Q(\top_ihp.oisc.regs[20][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][8]$_DFFE_PP_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1598),
    .D(_00898_),
    .Q_N(_13197_),
    .Q(\top_ihp.oisc.regs[20][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[20][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1599),
    .D(_00899_),
    .Q_N(_13196_),
    .Q(\top_ihp.oisc.regs[20][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][0]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1600),
    .D(_00900_),
    .Q_N(_13195_),
    .Q(\top_ihp.oisc.regs[21][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][10]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1601),
    .D(_00901_),
    .Q_N(_13194_),
    .Q(\top_ihp.oisc.regs[21][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][11]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1602),
    .D(_00902_),
    .Q_N(_13193_),
    .Q(\top_ihp.oisc.regs[21][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][12]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1603),
    .D(_00903_),
    .Q_N(_13192_),
    .Q(\top_ihp.oisc.regs[21][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][13]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1604),
    .D(_00904_),
    .Q_N(_13191_),
    .Q(\top_ihp.oisc.regs[21][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1605),
    .D(_00905_),
    .Q_N(_13190_),
    .Q(\top_ihp.oisc.regs[21][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][15]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1606),
    .D(_00906_),
    .Q_N(_13189_),
    .Q(\top_ihp.oisc.regs[21][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][16]$_DFFE_PP_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1607),
    .D(_00907_),
    .Q_N(_13188_),
    .Q(\top_ihp.oisc.regs[21][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][17]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1608),
    .D(_00908_),
    .Q_N(_13187_),
    .Q(\top_ihp.oisc.regs[21][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][18]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1609),
    .D(_00909_),
    .Q_N(_13186_),
    .Q(\top_ihp.oisc.regs[21][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][19]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1610),
    .D(_00910_),
    .Q_N(_13185_),
    .Q(\top_ihp.oisc.regs[21][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1611),
    .D(_00911_),
    .Q_N(_13184_),
    .Q(\top_ihp.oisc.regs[21][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][20]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1612),
    .D(_00912_),
    .Q_N(_13183_),
    .Q(\top_ihp.oisc.regs[21][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][21]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1613),
    .D(_00913_),
    .Q_N(_13182_),
    .Q(\top_ihp.oisc.regs[21][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1614),
    .D(_00914_),
    .Q_N(_13181_),
    .Q(\top_ihp.oisc.regs[21][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][23]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1615),
    .D(_00915_),
    .Q_N(_13180_),
    .Q(\top_ihp.oisc.regs[21][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][24]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1616),
    .D(_00916_),
    .Q_N(_13179_),
    .Q(\top_ihp.oisc.regs[21][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][25]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1617),
    .D(_00917_),
    .Q_N(_13178_),
    .Q(\top_ihp.oisc.regs[21][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][26]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1618),
    .D(_00918_),
    .Q_N(_13177_),
    .Q(\top_ihp.oisc.regs[21][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][27]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1619),
    .D(_00919_),
    .Q_N(_13176_),
    .Q(\top_ihp.oisc.regs[21][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][28]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1620),
    .D(_00920_),
    .Q_N(_13175_),
    .Q(\top_ihp.oisc.regs[21][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][29]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1621),
    .D(_00921_),
    .Q_N(_13174_),
    .Q(\top_ihp.oisc.regs[21][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][2]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1622),
    .D(_00922_),
    .Q_N(_13173_),
    .Q(\top_ihp.oisc.regs[21][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][30]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1623),
    .D(_00923_),
    .Q_N(_13172_),
    .Q(\top_ihp.oisc.regs[21][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][31]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1624),
    .D(_00924_),
    .Q_N(_13171_),
    .Q(\top_ihp.oisc.regs[21][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1625),
    .D(_00925_),
    .Q_N(_13170_),
    .Q(\top_ihp.oisc.regs[21][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1626),
    .D(_00926_),
    .Q_N(_13169_),
    .Q(\top_ihp.oisc.regs[21][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][5]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1627),
    .D(_00927_),
    .Q_N(_13168_),
    .Q(\top_ihp.oisc.regs[21][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][6]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1628),
    .D(_00928_),
    .Q_N(_13167_),
    .Q(\top_ihp.oisc.regs[21][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][7]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1629),
    .D(_00929_),
    .Q_N(_13166_),
    .Q(\top_ihp.oisc.regs[21][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1630),
    .D(_00930_),
    .Q_N(_13165_),
    .Q(\top_ihp.oisc.regs[21][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[21][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1631),
    .D(_00931_),
    .Q_N(_13164_),
    .Q(\top_ihp.oisc.regs[21][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1632),
    .D(_00932_),
    .Q_N(_13163_),
    .Q(\top_ihp.oisc.regs[22][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1633),
    .D(_00933_),
    .Q_N(_13162_),
    .Q(\top_ihp.oisc.regs[22][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1634),
    .D(_00934_),
    .Q_N(_13161_),
    .Q(\top_ihp.oisc.regs[22][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][12]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1635),
    .D(_00935_),
    .Q_N(_13160_),
    .Q(\top_ihp.oisc.regs[22][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][13]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1636),
    .D(_00936_),
    .Q_N(_13159_),
    .Q(\top_ihp.oisc.regs[22][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][14]$_DFFE_PP_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1637),
    .D(_00937_),
    .Q_N(_13158_),
    .Q(\top_ihp.oisc.regs[22][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][15]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1638),
    .D(_00938_),
    .Q_N(_13157_),
    .Q(\top_ihp.oisc.regs[22][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][16]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1639),
    .D(_00939_),
    .Q_N(_13156_),
    .Q(\top_ihp.oisc.regs[22][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][17]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1640),
    .D(_00940_),
    .Q_N(_13155_),
    .Q(\top_ihp.oisc.regs[22][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][18]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1641),
    .D(_00941_),
    .Q_N(_13154_),
    .Q(\top_ihp.oisc.regs[22][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][19]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1642),
    .D(_00942_),
    .Q_N(_13153_),
    .Q(\top_ihp.oisc.regs[22][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1643),
    .D(_00943_),
    .Q_N(_13152_),
    .Q(\top_ihp.oisc.regs[22][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][20]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1644),
    .D(_00944_),
    .Q_N(_13151_),
    .Q(\top_ihp.oisc.regs[22][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][21]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1645),
    .D(_00945_),
    .Q_N(_13150_),
    .Q(\top_ihp.oisc.regs[22][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][22]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1646),
    .D(_00946_),
    .Q_N(_13149_),
    .Q(\top_ihp.oisc.regs[22][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][23]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1647),
    .D(_00947_),
    .Q_N(_13148_),
    .Q(\top_ihp.oisc.regs[22][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][24]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1648),
    .D(_00948_),
    .Q_N(_13147_),
    .Q(\top_ihp.oisc.regs[22][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][25]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1649),
    .D(_00949_),
    .Q_N(_13146_),
    .Q(\top_ihp.oisc.regs[22][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1650),
    .D(_00950_),
    .Q_N(_13145_),
    .Q(\top_ihp.oisc.regs[22][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][27]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1651),
    .D(_00951_),
    .Q_N(_13144_),
    .Q(\top_ihp.oisc.regs[22][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][28]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1652),
    .D(_00952_),
    .Q_N(_13143_),
    .Q(\top_ihp.oisc.regs[22][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][29]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1653),
    .D(_00953_),
    .Q_N(_13142_),
    .Q(\top_ihp.oisc.regs[22][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1654),
    .D(_00954_),
    .Q_N(_13141_),
    .Q(\top_ihp.oisc.regs[22][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][30]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1655),
    .D(_00955_),
    .Q_N(_13140_),
    .Q(\top_ihp.oisc.regs[22][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][31]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1656),
    .D(_00956_),
    .Q_N(_13139_),
    .Q(\top_ihp.oisc.regs[22][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][3]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1657),
    .D(_00957_),
    .Q_N(_13138_),
    .Q(\top_ihp.oisc.regs[22][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1658),
    .D(_00958_),
    .Q_N(_13137_),
    .Q(\top_ihp.oisc.regs[22][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1659),
    .D(_00959_),
    .Q_N(_13136_),
    .Q(\top_ihp.oisc.regs[22][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][6]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1660),
    .D(_00960_),
    .Q_N(_13135_),
    .Q(\top_ihp.oisc.regs[22][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1661),
    .D(_00961_),
    .Q_N(_13134_),
    .Q(\top_ihp.oisc.regs[22][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1662),
    .D(_00962_),
    .Q_N(_13133_),
    .Q(\top_ihp.oisc.regs[22][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[22][9]$_DFFE_PP_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1663),
    .D(_00963_),
    .Q_N(_13132_),
    .Q(\top_ihp.oisc.regs[22][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][0]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1664),
    .D(_00964_),
    .Q_N(_13131_),
    .Q(\top_ihp.oisc.regs[23][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1665),
    .D(_00965_),
    .Q_N(_13130_),
    .Q(\top_ihp.oisc.regs[23][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][11]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1666),
    .D(_00966_),
    .Q_N(_13129_),
    .Q(\top_ihp.oisc.regs[23][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][12]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1667),
    .D(_00967_),
    .Q_N(_13128_),
    .Q(\top_ihp.oisc.regs[23][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][13]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1668),
    .D(_00968_),
    .Q_N(_13127_),
    .Q(\top_ihp.oisc.regs[23][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][14]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1669),
    .D(_00969_),
    .Q_N(_13126_),
    .Q(\top_ihp.oisc.regs[23][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][15]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1670),
    .D(_00970_),
    .Q_N(_13125_),
    .Q(\top_ihp.oisc.regs[23][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][16]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1671),
    .D(_00971_),
    .Q_N(_13124_),
    .Q(\top_ihp.oisc.regs[23][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][17]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1672),
    .D(_00972_),
    .Q_N(_13123_),
    .Q(\top_ihp.oisc.regs[23][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][18]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1673),
    .D(_00973_),
    .Q_N(_13122_),
    .Q(\top_ihp.oisc.regs[23][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][19]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1674),
    .D(_00974_),
    .Q_N(_13121_),
    .Q(\top_ihp.oisc.regs[23][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][1]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1675),
    .D(_00975_),
    .Q_N(_13120_),
    .Q(\top_ihp.oisc.regs[23][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][20]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1676),
    .D(_00976_),
    .Q_N(_13119_),
    .Q(\top_ihp.oisc.regs[23][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][21]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1677),
    .D(_00977_),
    .Q_N(_13118_),
    .Q(\top_ihp.oisc.regs[23][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][22]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1678),
    .D(_00978_),
    .Q_N(_13117_),
    .Q(\top_ihp.oisc.regs[23][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][23]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1679),
    .D(_00979_),
    .Q_N(_13116_),
    .Q(\top_ihp.oisc.regs[23][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][24]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1680),
    .D(_00980_),
    .Q_N(_13115_),
    .Q(\top_ihp.oisc.regs[23][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][25]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1681),
    .D(_00981_),
    .Q_N(_13114_),
    .Q(\top_ihp.oisc.regs[23][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][26]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1682),
    .D(_00982_),
    .Q_N(_13113_),
    .Q(\top_ihp.oisc.regs[23][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][27]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1683),
    .D(_00983_),
    .Q_N(_13112_),
    .Q(\top_ihp.oisc.regs[23][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][28]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1684),
    .D(_00984_),
    .Q_N(_13111_),
    .Q(\top_ihp.oisc.regs[23][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][29]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1685),
    .D(_00985_),
    .Q_N(_13110_),
    .Q(\top_ihp.oisc.regs[23][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][2]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1686),
    .D(_00986_),
    .Q_N(_13109_),
    .Q(\top_ihp.oisc.regs[23][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][30]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1687),
    .D(_00987_),
    .Q_N(_13108_),
    .Q(\top_ihp.oisc.regs[23][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][31]$_DFFE_PP_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1688),
    .D(_00988_),
    .Q_N(_13107_),
    .Q(\top_ihp.oisc.regs[23][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][3]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1689),
    .D(_00989_),
    .Q_N(_13106_),
    .Q(\top_ihp.oisc.regs[23][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][4]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1690),
    .D(_00990_),
    .Q_N(_13105_),
    .Q(\top_ihp.oisc.regs[23][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][5]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1691),
    .D(_00991_),
    .Q_N(_13104_),
    .Q(\top_ihp.oisc.regs[23][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][6]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1692),
    .D(_00992_),
    .Q_N(_13103_),
    .Q(\top_ihp.oisc.regs[23][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][7]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1693),
    .D(_00993_),
    .Q_N(_13102_),
    .Q(\top_ihp.oisc.regs[23][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1694),
    .D(_00994_),
    .Q_N(_13101_),
    .Q(\top_ihp.oisc.regs[23][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[23][9]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1695),
    .D(_00995_),
    .Q_N(_13100_),
    .Q(\top_ihp.oisc.regs[23][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][0]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1696),
    .D(_00996_),
    .Q_N(_13099_),
    .Q(\top_ihp.oisc.regs[24][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][10]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1697),
    .D(_00997_),
    .Q_N(_13098_),
    .Q(\top_ihp.oisc.regs[24][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][11]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1698),
    .D(_00998_),
    .Q_N(_13097_),
    .Q(\top_ihp.oisc.regs[24][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][12]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1699),
    .D(_00999_),
    .Q_N(_13096_),
    .Q(\top_ihp.oisc.regs[24][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][13]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1700),
    .D(_01000_),
    .Q_N(_13095_),
    .Q(\top_ihp.oisc.regs[24][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][14]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1701),
    .D(_01001_),
    .Q_N(_13094_),
    .Q(\top_ihp.oisc.regs[24][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][15]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1702),
    .D(_01002_),
    .Q_N(_13093_),
    .Q(\top_ihp.oisc.regs[24][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][16]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1703),
    .D(_01003_),
    .Q_N(_13092_),
    .Q(\top_ihp.oisc.regs[24][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][17]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1704),
    .D(_01004_),
    .Q_N(_13091_),
    .Q(\top_ihp.oisc.regs[24][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][18]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1705),
    .D(_01005_),
    .Q_N(_13090_),
    .Q(\top_ihp.oisc.regs[24][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][19]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1706),
    .D(_01006_),
    .Q_N(_13089_),
    .Q(\top_ihp.oisc.regs[24][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][1]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1707),
    .D(_01007_),
    .Q_N(_13088_),
    .Q(\top_ihp.oisc.regs[24][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1708),
    .D(_01008_),
    .Q_N(_13087_),
    .Q(\top_ihp.oisc.regs[24][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][21]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1709),
    .D(_01009_),
    .Q_N(_13086_),
    .Q(\top_ihp.oisc.regs[24][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1710),
    .D(_01010_),
    .Q_N(_13085_),
    .Q(\top_ihp.oisc.regs[24][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][23]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1711),
    .D(_01011_),
    .Q_N(_13084_),
    .Q(\top_ihp.oisc.regs[24][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][24]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1712),
    .D(_01012_),
    .Q_N(_13083_),
    .Q(\top_ihp.oisc.regs[24][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][25]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1713),
    .D(_01013_),
    .Q_N(_13082_),
    .Q(\top_ihp.oisc.regs[24][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][26]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1714),
    .D(_01014_),
    .Q_N(_13081_),
    .Q(\top_ihp.oisc.regs[24][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][27]$_DFFE_PP_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1715),
    .D(_01015_),
    .Q_N(_13080_),
    .Q(\top_ihp.oisc.regs[24][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][28]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1716),
    .D(_01016_),
    .Q_N(_13079_),
    .Q(\top_ihp.oisc.regs[24][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][29]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1717),
    .D(_01017_),
    .Q_N(_13078_),
    .Q(\top_ihp.oisc.regs[24][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][2]$_DFFE_PP_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1718),
    .D(_01018_),
    .Q_N(_13077_),
    .Q(\top_ihp.oisc.regs[24][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][30]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1719),
    .D(_01019_),
    .Q_N(_13076_),
    .Q(\top_ihp.oisc.regs[24][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][31]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1720),
    .D(_01020_),
    .Q_N(_13075_),
    .Q(\top_ihp.oisc.regs[24][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][3]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1721),
    .D(_01021_),
    .Q_N(_13074_),
    .Q(\top_ihp.oisc.regs[24][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][4]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1722),
    .D(_01022_),
    .Q_N(_13073_),
    .Q(\top_ihp.oisc.regs[24][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][5]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1723),
    .D(_01023_),
    .Q_N(_13072_),
    .Q(\top_ihp.oisc.regs[24][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][6]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1724),
    .D(_01024_),
    .Q_N(_13071_),
    .Q(\top_ihp.oisc.regs[24][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][7]$_DFFE_PP_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1725),
    .D(_01025_),
    .Q_N(_13070_),
    .Q(\top_ihp.oisc.regs[24][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][8]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1726),
    .D(_01026_),
    .Q_N(_13069_),
    .Q(\top_ihp.oisc.regs[24][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[24][9]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1727),
    .D(_01027_),
    .Q_N(_13068_),
    .Q(\top_ihp.oisc.regs[24][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][0]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1728),
    .D(_01028_),
    .Q_N(_13067_),
    .Q(\top_ihp.oisc.regs[25][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][10]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1729),
    .D(_01029_),
    .Q_N(_13066_),
    .Q(\top_ihp.oisc.regs[25][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][11]$_DFFE_PP_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1730),
    .D(_01030_),
    .Q_N(_13065_),
    .Q(\top_ihp.oisc.regs[25][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][12]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1731),
    .D(_01031_),
    .Q_N(_13064_),
    .Q(\top_ihp.oisc.regs[25][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1732),
    .D(_01032_),
    .Q_N(_13063_),
    .Q(\top_ihp.oisc.regs[25][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][14]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1733),
    .D(_01033_),
    .Q_N(_13062_),
    .Q(\top_ihp.oisc.regs[25][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][15]$_DFFE_PP_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1734),
    .D(_01034_),
    .Q_N(_13061_),
    .Q(\top_ihp.oisc.regs[25][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][16]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1735),
    .D(_01035_),
    .Q_N(_13060_),
    .Q(\top_ihp.oisc.regs[25][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][17]$_DFFE_PP_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1736),
    .D(_01036_),
    .Q_N(_13059_),
    .Q(\top_ihp.oisc.regs[25][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][18]$_DFFE_PP_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1737),
    .D(_01037_),
    .Q_N(_13058_),
    .Q(\top_ihp.oisc.regs[25][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][19]$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1738),
    .D(_01038_),
    .Q_N(_13057_),
    .Q(\top_ihp.oisc.regs[25][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1739),
    .D(_01039_),
    .Q_N(_13056_),
    .Q(\top_ihp.oisc.regs[25][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][20]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1740),
    .D(_01040_),
    .Q_N(_13055_),
    .Q(\top_ihp.oisc.regs[25][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][21]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1741),
    .D(_01041_),
    .Q_N(_13054_),
    .Q(\top_ihp.oisc.regs[25][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][22]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1742),
    .D(_01042_),
    .Q_N(_13053_),
    .Q(\top_ihp.oisc.regs[25][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][23]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1743),
    .D(_01043_),
    .Q_N(_13052_),
    .Q(\top_ihp.oisc.regs[25][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][24]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1744),
    .D(_01044_),
    .Q_N(_13051_),
    .Q(\top_ihp.oisc.regs[25][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][25]$_DFFE_PP_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1745),
    .D(_01045_),
    .Q_N(_13050_),
    .Q(\top_ihp.oisc.regs[25][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][26]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1746),
    .D(_01046_),
    .Q_N(_13049_),
    .Q(\top_ihp.oisc.regs[25][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][27]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1747),
    .D(_01047_),
    .Q_N(_13048_),
    .Q(\top_ihp.oisc.regs[25][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][28]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1748),
    .D(_01048_),
    .Q_N(_13047_),
    .Q(\top_ihp.oisc.regs[25][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][29]$_DFFE_PP_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1749),
    .D(_01049_),
    .Q_N(_13046_),
    .Q(\top_ihp.oisc.regs[25][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][2]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1750),
    .D(_01050_),
    .Q_N(_13045_),
    .Q(\top_ihp.oisc.regs[25][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][30]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1751),
    .D(_01051_),
    .Q_N(_13044_),
    .Q(\top_ihp.oisc.regs[25][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][31]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1752),
    .D(_01052_),
    .Q_N(_13043_),
    .Q(\top_ihp.oisc.regs[25][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][3]$_DFFE_PP_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1753),
    .D(_01053_),
    .Q_N(_13042_),
    .Q(\top_ihp.oisc.regs[25][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][4]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1754),
    .D(_01054_),
    .Q_N(_13041_),
    .Q(\top_ihp.oisc.regs[25][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][5]$_DFFE_PP_  (.CLK(clknet_leaf_234_clk),
    .RESET_B(net1755),
    .D(_01055_),
    .Q_N(_13040_),
    .Q(\top_ihp.oisc.regs[25][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][6]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1756),
    .D(_01056_),
    .Q_N(_13039_),
    .Q(\top_ihp.oisc.regs[25][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][7]$_DFFE_PP_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1757),
    .D(_01057_),
    .Q_N(_13038_),
    .Q(\top_ihp.oisc.regs[25][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1758),
    .D(_01058_),
    .Q_N(_13037_),
    .Q(\top_ihp.oisc.regs[25][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[25][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1759),
    .D(_01059_),
    .Q_N(_13036_),
    .Q(\top_ihp.oisc.regs[25][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][0]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1760),
    .D(_01060_),
    .Q_N(_13035_),
    .Q(\top_ihp.oisc.regs[26][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][10]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1761),
    .D(_01061_),
    .Q_N(_13034_),
    .Q(\top_ihp.oisc.regs[26][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1762),
    .D(_01062_),
    .Q_N(_13033_),
    .Q(\top_ihp.oisc.regs[26][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][12]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1763),
    .D(_01063_),
    .Q_N(_13032_),
    .Q(\top_ihp.oisc.regs[26][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][13]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1764),
    .D(_01064_),
    .Q_N(_13031_),
    .Q(\top_ihp.oisc.regs[26][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][14]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1765),
    .D(_01065_),
    .Q_N(_13030_),
    .Q(\top_ihp.oisc.regs[26][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1766),
    .D(_01066_),
    .Q_N(_13029_),
    .Q(\top_ihp.oisc.regs[26][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][16]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1767),
    .D(_01067_),
    .Q_N(_13028_),
    .Q(\top_ihp.oisc.regs[26][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][17]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1768),
    .D(_01068_),
    .Q_N(_13027_),
    .Q(\top_ihp.oisc.regs[26][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][18]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1769),
    .D(_01069_),
    .Q_N(_13026_),
    .Q(\top_ihp.oisc.regs[26][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][19]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1770),
    .D(_01070_),
    .Q_N(_13025_),
    .Q(\top_ihp.oisc.regs[26][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1771),
    .D(_01071_),
    .Q_N(_13024_),
    .Q(\top_ihp.oisc.regs[26][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][20]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1772),
    .D(_01072_),
    .Q_N(_13023_),
    .Q(\top_ihp.oisc.regs[26][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][21]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1773),
    .D(_01073_),
    .Q_N(_13022_),
    .Q(\top_ihp.oisc.regs[26][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][22]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1774),
    .D(_01074_),
    .Q_N(_13021_),
    .Q(\top_ihp.oisc.regs[26][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][23]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1775),
    .D(_01075_),
    .Q_N(_13020_),
    .Q(\top_ihp.oisc.regs[26][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][24]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1776),
    .D(_01076_),
    .Q_N(_13019_),
    .Q(\top_ihp.oisc.regs[26][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1777),
    .D(_01077_),
    .Q_N(_13018_),
    .Q(\top_ihp.oisc.regs[26][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][26]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1778),
    .D(_01078_),
    .Q_N(_13017_),
    .Q(\top_ihp.oisc.regs[26][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][27]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1779),
    .D(_01079_),
    .Q_N(_13016_),
    .Q(\top_ihp.oisc.regs[26][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][28]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1780),
    .D(_01080_),
    .Q_N(_13015_),
    .Q(\top_ihp.oisc.regs[26][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][29]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1781),
    .D(_01081_),
    .Q_N(_13014_),
    .Q(\top_ihp.oisc.regs[26][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][2]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1782),
    .D(_01082_),
    .Q_N(_13013_),
    .Q(\top_ihp.oisc.regs[26][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][30]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1783),
    .D(_01083_),
    .Q_N(_13012_),
    .Q(\top_ihp.oisc.regs[26][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][31]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1784),
    .D(_01084_),
    .Q_N(_13011_),
    .Q(\top_ihp.oisc.regs[26][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][3]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1785),
    .D(_01085_),
    .Q_N(_13010_),
    .Q(\top_ihp.oisc.regs[26][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][4]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1786),
    .D(_01086_),
    .Q_N(_13009_),
    .Q(\top_ihp.oisc.regs[26][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][5]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1787),
    .D(_01087_),
    .Q_N(_13008_),
    .Q(\top_ihp.oisc.regs[26][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][6]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1788),
    .D(_01088_),
    .Q_N(_13007_),
    .Q(\top_ihp.oisc.regs[26][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][7]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1789),
    .D(_01089_),
    .Q_N(_13006_),
    .Q(\top_ihp.oisc.regs[26][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1790),
    .D(_01090_),
    .Q_N(_13005_),
    .Q(\top_ihp.oisc.regs[26][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[26][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1791),
    .D(_01091_),
    .Q_N(_13004_),
    .Q(\top_ihp.oisc.regs[26][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][0]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1792),
    .D(_01092_),
    .Q_N(_13003_),
    .Q(\top_ihp.oisc.regs[27][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][10]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1793),
    .D(_01093_),
    .Q_N(_13002_),
    .Q(\top_ihp.oisc.regs[27][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][11]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1794),
    .D(_01094_),
    .Q_N(_13001_),
    .Q(\top_ihp.oisc.regs[27][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][12]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1795),
    .D(_01095_),
    .Q_N(_13000_),
    .Q(\top_ihp.oisc.regs[27][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][13]$_DFFE_PP_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1796),
    .D(_01096_),
    .Q_N(_12999_),
    .Q(\top_ihp.oisc.regs[27][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][14]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1797),
    .D(_01097_),
    .Q_N(_12998_),
    .Q(\top_ihp.oisc.regs[27][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][15]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1798),
    .D(_01098_),
    .Q_N(_12997_),
    .Q(\top_ihp.oisc.regs[27][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][16]$_DFFE_PP_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1799),
    .D(_01099_),
    .Q_N(_12996_),
    .Q(\top_ihp.oisc.regs[27][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1800),
    .D(_01100_),
    .Q_N(_12995_),
    .Q(\top_ihp.oisc.regs[27][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][18]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1801),
    .D(_01101_),
    .Q_N(_12994_),
    .Q(\top_ihp.oisc.regs[27][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][19]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1802),
    .D(_01102_),
    .Q_N(_12993_),
    .Q(\top_ihp.oisc.regs[27][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][1]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1803),
    .D(_01103_),
    .Q_N(_12992_),
    .Q(\top_ihp.oisc.regs[27][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][20]$_DFFE_PP_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1804),
    .D(_01104_),
    .Q_N(_12991_),
    .Q(\top_ihp.oisc.regs[27][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][21]$_DFFE_PP_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1805),
    .D(_01105_),
    .Q_N(_12990_),
    .Q(\top_ihp.oisc.regs[27][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][22]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1806),
    .D(_01106_),
    .Q_N(_12989_),
    .Q(\top_ihp.oisc.regs[27][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][23]$_DFFE_PP_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1807),
    .D(_01107_),
    .Q_N(_12988_),
    .Q(\top_ihp.oisc.regs[27][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][24]$_DFFE_PP_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1808),
    .D(_01108_),
    .Q_N(_12987_),
    .Q(\top_ihp.oisc.regs[27][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][25]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1809),
    .D(_01109_),
    .Q_N(_12986_),
    .Q(\top_ihp.oisc.regs[27][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][26]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1810),
    .D(_01110_),
    .Q_N(_12985_),
    .Q(\top_ihp.oisc.regs[27][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][27]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1811),
    .D(_01111_),
    .Q_N(_12984_),
    .Q(\top_ihp.oisc.regs[27][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][28]$_DFFE_PP_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1812),
    .D(_01112_),
    .Q_N(_12983_),
    .Q(\top_ihp.oisc.regs[27][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1813),
    .D(_01113_),
    .Q_N(_12982_),
    .Q(\top_ihp.oisc.regs[27][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][2]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1814),
    .D(_01114_),
    .Q_N(_12981_),
    .Q(\top_ihp.oisc.regs[27][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][30]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1815),
    .D(_01115_),
    .Q_N(_12980_),
    .Q(\top_ihp.oisc.regs[27][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][31]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1816),
    .D(_01116_),
    .Q_N(_12979_),
    .Q(\top_ihp.oisc.regs[27][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][3]$_DFFE_PP_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1817),
    .D(_01117_),
    .Q_N(_12978_),
    .Q(\top_ihp.oisc.regs[27][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][4]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1818),
    .D(_01118_),
    .Q_N(_12977_),
    .Q(\top_ihp.oisc.regs[27][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][5]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1819),
    .D(_01119_),
    .Q_N(_12976_),
    .Q(\top_ihp.oisc.regs[27][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][6]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1820),
    .D(_01120_),
    .Q_N(_12975_),
    .Q(\top_ihp.oisc.regs[27][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][7]$_DFFE_PP_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1821),
    .D(_01121_),
    .Q_N(_12974_),
    .Q(\top_ihp.oisc.regs[27][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][8]$_DFFE_PP_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1822),
    .D(_01122_),
    .Q_N(_12973_),
    .Q(\top_ihp.oisc.regs[27][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[27][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1823),
    .D(_01123_),
    .Q_N(_12972_),
    .Q(\top_ihp.oisc.regs[27][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][0]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1824),
    .D(_01124_),
    .Q_N(_12971_),
    .Q(\top_ihp.oisc.regs[28][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][10]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1825),
    .D(_01125_),
    .Q_N(_12970_),
    .Q(\top_ihp.oisc.regs[28][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][11]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1826),
    .D(_01126_),
    .Q_N(_12969_),
    .Q(\top_ihp.oisc.regs[28][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][12]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1827),
    .D(_01127_),
    .Q_N(_12968_),
    .Q(\top_ihp.oisc.regs[28][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][13]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1828),
    .D(_01128_),
    .Q_N(_12967_),
    .Q(\top_ihp.oisc.regs[28][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][14]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1829),
    .D(_01129_),
    .Q_N(_12966_),
    .Q(\top_ihp.oisc.regs[28][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][15]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1830),
    .D(_01130_),
    .Q_N(_12965_),
    .Q(\top_ihp.oisc.regs[28][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][16]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1831),
    .D(_01131_),
    .Q_N(_12964_),
    .Q(\top_ihp.oisc.regs[28][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][17]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1832),
    .D(_01132_),
    .Q_N(_12963_),
    .Q(\top_ihp.oisc.regs[28][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][18]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1833),
    .D(_01133_),
    .Q_N(_12962_),
    .Q(\top_ihp.oisc.regs[28][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][19]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1834),
    .D(_01134_),
    .Q_N(_12961_),
    .Q(\top_ihp.oisc.regs[28][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][1]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1835),
    .D(_01135_),
    .Q_N(_12960_),
    .Q(\top_ihp.oisc.regs[28][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][20]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1836),
    .D(_01136_),
    .Q_N(_12959_),
    .Q(\top_ihp.oisc.regs[28][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][21]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1837),
    .D(_01137_),
    .Q_N(_12958_),
    .Q(\top_ihp.oisc.regs[28][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][22]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1838),
    .D(_01138_),
    .Q_N(_12957_),
    .Q(\top_ihp.oisc.regs[28][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][23]$_DFFE_PP_  (.CLK(clknet_leaf_152_clk),
    .RESET_B(net1839),
    .D(_01139_),
    .Q_N(_12956_),
    .Q(\top_ihp.oisc.regs[28][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][24]$_DFFE_PP_  (.CLK(clknet_leaf_238_clk),
    .RESET_B(net1840),
    .D(_01140_),
    .Q_N(_12955_),
    .Q(\top_ihp.oisc.regs[28][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1841),
    .D(_01141_),
    .Q_N(_12954_),
    .Q(\top_ihp.oisc.regs[28][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][26]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1842),
    .D(_01142_),
    .Q_N(_12953_),
    .Q(\top_ihp.oisc.regs[28][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][27]$_DFFE_PP_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1843),
    .D(_01143_),
    .Q_N(_12952_),
    .Q(\top_ihp.oisc.regs[28][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][28]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1844),
    .D(_01144_),
    .Q_N(_12951_),
    .Q(\top_ihp.oisc.regs[28][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][29]$_DFFE_PP_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1845),
    .D(_01145_),
    .Q_N(_12950_),
    .Q(\top_ihp.oisc.regs[28][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][2]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1846),
    .D(_01146_),
    .Q_N(_12949_),
    .Q(\top_ihp.oisc.regs[28][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][30]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1847),
    .D(_01147_),
    .Q_N(_12948_),
    .Q(\top_ihp.oisc.regs[28][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][31]$_DFFE_PP_  (.CLK(clknet_leaf_241_clk),
    .RESET_B(net1848),
    .D(_01148_),
    .Q_N(_12947_),
    .Q(\top_ihp.oisc.regs[28][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][3]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1849),
    .D(_01149_),
    .Q_N(_12946_),
    .Q(\top_ihp.oisc.regs[28][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][4]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1850),
    .D(_01150_),
    .Q_N(_12945_),
    .Q(\top_ihp.oisc.regs[28][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][5]$_DFFE_PP_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1851),
    .D(_01151_),
    .Q_N(_12944_),
    .Q(\top_ihp.oisc.regs[28][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][6]$_DFFE_PP_  (.CLK(clknet_leaf_237_clk),
    .RESET_B(net1852),
    .D(_01152_),
    .Q_N(_12943_),
    .Q(\top_ihp.oisc.regs[28][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][7]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1853),
    .D(_01153_),
    .Q_N(_12942_),
    .Q(\top_ihp.oisc.regs[28][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][8]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1854),
    .D(_01154_),
    .Q_N(_12941_),
    .Q(\top_ihp.oisc.regs[28][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[28][9]$_DFFE_PP_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1855),
    .D(_01155_),
    .Q_N(_12940_),
    .Q(\top_ihp.oisc.regs[28][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1856),
    .D(_01156_),
    .Q_N(_12939_),
    .Q(\top_ihp.oisc.regs[29][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][10]$_DFFE_PP_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1857),
    .D(_01157_),
    .Q_N(_12938_),
    .Q(\top_ihp.oisc.regs[29][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][11]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1858),
    .D(_01158_),
    .Q_N(_12937_),
    .Q(\top_ihp.oisc.regs[29][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][12]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1859),
    .D(_01159_),
    .Q_N(_12936_),
    .Q(\top_ihp.oisc.regs[29][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][13]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1860),
    .D(_01160_),
    .Q_N(_12935_),
    .Q(\top_ihp.oisc.regs[29][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][14]$_DFFE_PP_  (.CLK(clknet_leaf_216_clk),
    .RESET_B(net1861),
    .D(_01161_),
    .Q_N(_12934_),
    .Q(\top_ihp.oisc.regs[29][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][15]$_DFFE_PP_  (.CLK(clknet_leaf_149_clk),
    .RESET_B(net1862),
    .D(_01162_),
    .Q_N(_12933_),
    .Q(\top_ihp.oisc.regs[29][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][16]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1863),
    .D(_01163_),
    .Q_N(_12932_),
    .Q(\top_ihp.oisc.regs[29][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][17]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1864),
    .D(_01164_),
    .Q_N(_12931_),
    .Q(\top_ihp.oisc.regs[29][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][18]$_DFFE_PP_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1865),
    .D(_01165_),
    .Q_N(_12930_),
    .Q(\top_ihp.oisc.regs[29][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][19]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1866),
    .D(_01166_),
    .Q_N(_12929_),
    .Q(\top_ihp.oisc.regs[29][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][1]$_DFFE_PP_  (.CLK(clknet_leaf_219_clk),
    .RESET_B(net1867),
    .D(_01167_),
    .Q_N(_12928_),
    .Q(\top_ihp.oisc.regs[29][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][20]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1868),
    .D(_01168_),
    .Q_N(_12927_),
    .Q(\top_ihp.oisc.regs[29][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][21]$_DFFE_PP_  (.CLK(clknet_leaf_163_clk),
    .RESET_B(net1869),
    .D(_01169_),
    .Q_N(_12926_),
    .Q(\top_ihp.oisc.regs[29][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][22]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1870),
    .D(_01170_),
    .Q_N(_12925_),
    .Q(\top_ihp.oisc.regs[29][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][23]$_DFFE_PP_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1871),
    .D(_01171_),
    .Q_N(_12924_),
    .Q(\top_ihp.oisc.regs[29][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][24]$_DFFE_PP_  (.CLK(clknet_leaf_242_clk),
    .RESET_B(net1872),
    .D(_01172_),
    .Q_N(_12923_),
    .Q(\top_ihp.oisc.regs[29][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][25]$_DFFE_PP_  (.CLK(clknet_leaf_157_clk),
    .RESET_B(net1873),
    .D(_01173_),
    .Q_N(_12922_),
    .Q(\top_ihp.oisc.regs[29][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][26]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1874),
    .D(_01174_),
    .Q_N(_12921_),
    .Q(\top_ihp.oisc.regs[29][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][27]$_DFFE_PP_  (.CLK(clknet_leaf_235_clk),
    .RESET_B(net1875),
    .D(_01175_),
    .Q_N(_12920_),
    .Q(\top_ihp.oisc.regs[29][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][28]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1876),
    .D(_01176_),
    .Q_N(_12919_),
    .Q(\top_ihp.oisc.regs[29][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][29]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1877),
    .D(_01177_),
    .Q_N(_12918_),
    .Q(\top_ihp.oisc.regs[29][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1878),
    .D(_01178_),
    .Q_N(_12917_),
    .Q(\top_ihp.oisc.regs[29][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][30]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1879),
    .D(_01179_),
    .Q_N(_12916_),
    .Q(\top_ihp.oisc.regs[29][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][31]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1880),
    .D(_01180_),
    .Q_N(_12915_),
    .Q(\top_ihp.oisc.regs[29][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][3]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1881),
    .D(_01181_),
    .Q_N(_12914_),
    .Q(\top_ihp.oisc.regs[29][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][4]$_DFFE_PP_  (.CLK(clknet_leaf_214_clk),
    .RESET_B(net1882),
    .D(_01182_),
    .Q_N(_12913_),
    .Q(\top_ihp.oisc.regs[29][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1883),
    .D(_01183_),
    .Q_N(_12912_),
    .Q(\top_ihp.oisc.regs[29][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][6]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1884),
    .D(_01184_),
    .Q_N(_12911_),
    .Q(\top_ihp.oisc.regs[29][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][7]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1885),
    .D(_01185_),
    .Q_N(_12910_),
    .Q(\top_ihp.oisc.regs[29][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][8]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1886),
    .D(_01186_),
    .Q_N(_12909_),
    .Q(\top_ihp.oisc.regs[29][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[29][9]$_DFFE_PP_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1887),
    .D(_01187_),
    .Q_N(_12908_),
    .Q(\top_ihp.oisc.regs[29][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1374),
    .D(_01188_),
    .Q_N(_12907_),
    .Q(\top_ihp.oisc.regs[2][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1383),
    .D(_01189_),
    .Q_N(_12906_),
    .Q(\top_ihp.oisc.regs[2][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1380),
    .D(_01190_),
    .Q_N(_12905_),
    .Q(\top_ihp.oisc.regs[2][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1342),
    .D(_01191_),
    .Q_N(_12904_),
    .Q(\top_ihp.oisc.regs[2][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1405),
    .D(_01192_),
    .Q_N(_12903_),
    .Q(\top_ihp.oisc.regs[2][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1397),
    .D(_01193_),
    .Q_N(_12902_),
    .Q(\top_ihp.oisc.regs[2][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1396),
    .D(_01194_),
    .Q_N(_12901_),
    .Q(\top_ihp.oisc.regs[2][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1362),
    .D(_01195_),
    .Q_N(_12900_),
    .Q(\top_ihp.oisc.regs[2][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1362),
    .D(_01196_),
    .Q_N(_12899_),
    .Q(\top_ihp.oisc.regs[2][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_189_clk),
    .RESET_B(net1398),
    .D(_01197_),
    .Q_N(_12898_),
    .Q(\top_ihp.oisc.regs[2][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1343),
    .D(_01198_),
    .Q_N(_12897_),
    .Q(\top_ihp.oisc.regs[2][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1382),
    .D(_01199_),
    .Q_N(_12896_),
    .Q(\top_ihp.oisc.regs[2][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1412),
    .D(_01200_),
    .Q_N(_12895_),
    .Q(\top_ihp.oisc.regs[2][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1399),
    .D(_01201_),
    .Q_N(_12894_),
    .Q(\top_ihp.oisc.regs[2][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1403),
    .D(_01202_),
    .Q_N(_12893_),
    .Q(\top_ihp.oisc.regs[2][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1403),
    .D(_01203_),
    .Q_N(_12892_),
    .Q(\top_ihp.oisc.regs[2][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1340),
    .D(_01204_),
    .Q_N(_12891_),
    .Q(\top_ihp.oisc.regs[2][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_145_clk),
    .RESET_B(net1399),
    .D(_01205_),
    .Q_N(_12890_),
    .Q(\top_ihp.oisc.regs[2][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1412),
    .D(_01206_),
    .Q_N(_12889_),
    .Q(\top_ihp.oisc.regs[2][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1381),
    .D(_01207_),
    .Q_N(_12888_),
    .Q(\top_ihp.oisc.regs[2][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1381),
    .D(_01208_),
    .Q_N(_12887_),
    .Q(\top_ihp.oisc.regs[2][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1396),
    .D(_01209_),
    .Q_N(_12886_),
    .Q(\top_ihp.oisc.regs[2][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1405),
    .D(_01210_),
    .Q_N(_12885_),
    .Q(\top_ihp.oisc.regs[2][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1394),
    .D(_01211_),
    .Q_N(_12884_),
    .Q(\top_ihp.oisc.regs[2][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1361),
    .D(_01212_),
    .Q_N(_12883_),
    .Q(\top_ihp.oisc.regs[2][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1336),
    .D(_01213_),
    .Q_N(_12882_),
    .Q(\top_ihp.oisc.regs[2][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_243_clk),
    .RESET_B(net1387),
    .D(_01214_),
    .Q_N(_12881_),
    .Q(\top_ihp.oisc.regs[2][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1339),
    .D(_01215_),
    .Q_N(_12880_),
    .Q(\top_ihp.oisc.regs[2][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1385),
    .D(_01216_),
    .Q_N(_12879_),
    .Q(\top_ihp.oisc.regs[2][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1394),
    .D(_01217_),
    .Q_N(_12878_),
    .Q(\top_ihp.oisc.regs[2][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1381),
    .D(_01218_),
    .Q_N(_12877_),
    .Q(\top_ihp.oisc.regs[2][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[2][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1387),
    .D(_01219_),
    .Q_N(_12876_),
    .Q(\top_ihp.oisc.regs[2][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][0]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1888),
    .D(_01220_),
    .Q_N(_12875_),
    .Q(\top_ihp.oisc.regs[30][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][10]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1889),
    .D(_01221_),
    .Q_N(_12874_),
    .Q(\top_ihp.oisc.regs[30][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][11]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1890),
    .D(_01222_),
    .Q_N(_12873_),
    .Q(\top_ihp.oisc.regs[30][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][12]$_DFFE_PP_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net1891),
    .D(_01223_),
    .Q_N(_12872_),
    .Q(\top_ihp.oisc.regs[30][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][13]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1892),
    .D(_01224_),
    .Q_N(_12871_),
    .Q(\top_ihp.oisc.regs[30][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][14]$_DFFE_PP_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1893),
    .D(_01225_),
    .Q_N(_12870_),
    .Q(\top_ihp.oisc.regs[30][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][15]$_DFFE_PP_  (.CLK(clknet_leaf_171_clk),
    .RESET_B(net1894),
    .D(_01226_),
    .Q_N(_12869_),
    .Q(\top_ihp.oisc.regs[30][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][16]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1895),
    .D(_01227_),
    .Q_N(_12868_),
    .Q(\top_ihp.oisc.regs[30][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][17]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1896),
    .D(_01228_),
    .Q_N(_12867_),
    .Q(\top_ihp.oisc.regs[30][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1897),
    .D(_01229_),
    .Q_N(_12866_),
    .Q(\top_ihp.oisc.regs[30][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][19]$_DFFE_PP_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1898),
    .D(_01230_),
    .Q_N(_12865_),
    .Q(\top_ihp.oisc.regs[30][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1899),
    .D(_01231_),
    .Q_N(_12864_),
    .Q(\top_ihp.oisc.regs[30][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][20]$_DFFE_PP_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1900),
    .D(_01232_),
    .Q_N(_12863_),
    .Q(\top_ihp.oisc.regs[30][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][21]$_DFFE_PP_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1901),
    .D(_01233_),
    .Q_N(_12862_),
    .Q(\top_ihp.oisc.regs[30][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1902),
    .D(_01234_),
    .Q_N(_12861_),
    .Q(\top_ihp.oisc.regs[30][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][23]$_DFFE_PP_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1903),
    .D(_01235_),
    .Q_N(_12860_),
    .Q(\top_ihp.oisc.regs[30][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][24]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1904),
    .D(_01236_),
    .Q_N(_12859_),
    .Q(\top_ihp.oisc.regs[30][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][25]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1905),
    .D(_01237_),
    .Q_N(_12858_),
    .Q(\top_ihp.oisc.regs[30][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][26]$_DFFE_PP_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1906),
    .D(_01238_),
    .Q_N(_12857_),
    .Q(\top_ihp.oisc.regs[30][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][27]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1907),
    .D(_01239_),
    .Q_N(_12856_),
    .Q(\top_ihp.oisc.regs[30][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][28]$_DFFE_PP_  (.CLK(clknet_leaf_175_clk),
    .RESET_B(net1908),
    .D(_01240_),
    .Q_N(_12855_),
    .Q(\top_ihp.oisc.regs[30][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][29]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1909),
    .D(_01241_),
    .Q_N(_12854_),
    .Q(\top_ihp.oisc.regs[30][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][2]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1910),
    .D(_01242_),
    .Q_N(_12853_),
    .Q(\top_ihp.oisc.regs[30][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][30]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1911),
    .D(_01243_),
    .Q_N(_12852_),
    .Q(\top_ihp.oisc.regs[30][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][31]$_DFFE_PP_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1912),
    .D(_01244_),
    .Q_N(_12851_),
    .Q(\top_ihp.oisc.regs[30][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][3]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1913),
    .D(_01245_),
    .Q_N(_12850_),
    .Q(\top_ihp.oisc.regs[30][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][4]$_DFFE_PP_  (.CLK(clknet_leaf_220_clk),
    .RESET_B(net1914),
    .D(_01246_),
    .Q_N(_12849_),
    .Q(\top_ihp.oisc.regs[30][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][5]$_DFFE_PP_  (.CLK(clknet_leaf_236_clk),
    .RESET_B(net1915),
    .D(_01247_),
    .Q_N(_12848_),
    .Q(\top_ihp.oisc.regs[30][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][6]$_DFFE_PP_  (.CLK(clknet_leaf_224_clk),
    .RESET_B(net1916),
    .D(_01248_),
    .Q_N(_12847_),
    .Q(\top_ihp.oisc.regs[30][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][7]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1917),
    .D(_01249_),
    .Q_N(_12846_),
    .Q(\top_ihp.oisc.regs[30][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][8]$_DFFE_PP_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1918),
    .D(_01250_),
    .Q_N(_12845_),
    .Q(\top_ihp.oisc.regs[30][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[30][9]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1919),
    .D(_01251_),
    .Q_N(_12844_),
    .Q(\top_ihp.oisc.regs[30][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][0]$_DFFE_PP_  (.CLK(clknet_leaf_232_clk),
    .RESET_B(net1920),
    .D(_01252_),
    .Q_N(_12843_),
    .Q(\top_ihp.oisc.regs[31][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][10]$_DFFE_PP_  (.CLK(clknet_leaf_233_clk),
    .RESET_B(net1921),
    .D(_01253_),
    .Q_N(_12842_),
    .Q(\top_ihp.oisc.regs[31][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][11]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1922),
    .D(_01254_),
    .Q_N(_12841_),
    .Q(\top_ihp.oisc.regs[31][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][12]$_DFFE_PP_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1923),
    .D(_01255_),
    .Q_N(_12840_),
    .Q(\top_ihp.oisc.regs[31][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][13]$_DFFE_PP_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1924),
    .D(_01256_),
    .Q_N(_12839_),
    .Q(\top_ihp.oisc.regs[31][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][14]$_DFFE_PP_  (.CLK(clknet_leaf_170_clk),
    .RESET_B(net1925),
    .D(_01257_),
    .Q_N(_12838_),
    .Q(\top_ihp.oisc.regs[31][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][15]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1926),
    .D(_01258_),
    .Q_N(_12837_),
    .Q(\top_ihp.oisc.regs[31][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][16]$_DFFE_PP_  (.CLK(clknet_leaf_174_clk),
    .RESET_B(net1927),
    .D(_01259_),
    .Q_N(_12836_),
    .Q(\top_ihp.oisc.regs[31][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][17]$_DFFE_PP_  (.CLK(clknet_leaf_154_clk),
    .RESET_B(net1928),
    .D(_01260_),
    .Q_N(_12835_),
    .Q(\top_ihp.oisc.regs[31][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][18]$_DFFE_PP_  (.CLK(clknet_leaf_158_clk),
    .RESET_B(net1929),
    .D(_01261_),
    .Q_N(_12834_),
    .Q(\top_ihp.oisc.regs[31][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][19]$_DFFE_PP_  (.CLK(clknet_leaf_240_clk),
    .RESET_B(net1930),
    .D(_01262_),
    .Q_N(_12833_),
    .Q(\top_ihp.oisc.regs[31][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][1]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1931),
    .D(_01263_),
    .Q_N(_12832_),
    .Q(\top_ihp.oisc.regs[31][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][20]$_DFFE_PP_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1932),
    .D(_01264_),
    .Q_N(_12831_),
    .Q(\top_ihp.oisc.regs[31][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][21]$_DFFE_PP_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1933),
    .D(_01265_),
    .Q_N(_12830_),
    .Q(\top_ihp.oisc.regs[31][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][22]$_DFFE_PP_  (.CLK(clknet_leaf_162_clk),
    .RESET_B(net1934),
    .D(_01266_),
    .Q_N(_12829_),
    .Q(\top_ihp.oisc.regs[31][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][23]$_DFFE_PP_  (.CLK(clknet_leaf_153_clk),
    .RESET_B(net1935),
    .D(_01267_),
    .Q_N(_12828_),
    .Q(\top_ihp.oisc.regs[31][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][24]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1936),
    .D(_01268_),
    .Q_N(_12827_),
    .Q(\top_ihp.oisc.regs[31][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][25]$_DFFE_PP_  (.CLK(clknet_leaf_151_clk),
    .RESET_B(net1937),
    .D(_01269_),
    .Q_N(_12826_),
    .Q(\top_ihp.oisc.regs[31][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][26]$_DFFE_PP_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1938),
    .D(_01270_),
    .Q_N(_12825_),
    .Q(\top_ihp.oisc.regs[31][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][27]$_DFFE_PP_  (.CLK(clknet_leaf_225_clk),
    .RESET_B(net1939),
    .D(_01271_),
    .Q_N(_12824_),
    .Q(\top_ihp.oisc.regs[31][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][28]$_DFFE_PP_  (.CLK(clknet_leaf_215_clk),
    .RESET_B(net1940),
    .D(_01272_),
    .Q_N(_12823_),
    .Q(\top_ihp.oisc.regs[31][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][29]$_DFFE_PP_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1941),
    .D(_01273_),
    .Q_N(_12822_),
    .Q(\top_ihp.oisc.regs[31][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][2]$_DFFE_PP_  (.CLK(clknet_leaf_180_clk),
    .RESET_B(net1942),
    .D(_01274_),
    .Q_N(_12821_),
    .Q(\top_ihp.oisc.regs[31][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][30]$_DFFE_PP_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1943),
    .D(_01275_),
    .Q_N(_12820_),
    .Q(\top_ihp.oisc.regs[31][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][31]$_DFFE_PP_  (.CLK(clknet_leaf_181_clk),
    .RESET_B(net1944),
    .D(_01276_),
    .Q_N(_12819_),
    .Q(\top_ihp.oisc.regs[31][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][3]$_DFFE_PP_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1945),
    .D(_01277_),
    .Q_N(_12818_),
    .Q(\top_ihp.oisc.regs[31][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][4]$_DFFE_PP_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1946),
    .D(_01278_),
    .Q_N(_12817_),
    .Q(\top_ihp.oisc.regs[31][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][5]$_DFFE_PP_  (.CLK(clknet_leaf_218_clk),
    .RESET_B(net1947),
    .D(_01279_),
    .Q_N(_12816_),
    .Q(\top_ihp.oisc.regs[31][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][6]$_DFFE_PP_  (.CLK(clknet_leaf_231_clk),
    .RESET_B(net1948),
    .D(_01280_),
    .Q_N(_12815_),
    .Q(\top_ihp.oisc.regs[31][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][7]$_DFFE_PP_  (.CLK(clknet_leaf_176_clk),
    .RESET_B(net1949),
    .D(_01281_),
    .Q_N(_12814_),
    .Q(\top_ihp.oisc.regs[31][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][8]$_DFFE_PP_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1950),
    .D(_01282_),
    .Q_N(_12813_),
    .Q(\top_ihp.oisc.regs[31][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[31][9]$_DFFE_PP_  (.CLK(clknet_leaf_239_clk),
    .RESET_B(net1951),
    .D(_01283_),
    .Q_N(_12812_),
    .Q(\top_ihp.oisc.regs[31][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][0]$_DFFE_PP_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1952),
    .D(_01284_),
    .Q_N(_12811_),
    .Q(\top_ihp.oisc.regs[32][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][10]$_DFFE_PP_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1953),
    .D(_01285_),
    .Q_N(_12810_),
    .Q(\top_ihp.oisc.regs[32][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][11]$_DFFE_PP_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1954),
    .D(_01286_),
    .Q_N(_12809_),
    .Q(\top_ihp.oisc.regs[32][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][12]$_DFFE_PP_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1955),
    .D(_01287_),
    .Q_N(_12808_),
    .Q(\top_ihp.oisc.regs[32][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][13]$_DFFE_PP_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1956),
    .D(_01288_),
    .Q_N(_12807_),
    .Q(\top_ihp.oisc.regs[32][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][14]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1957),
    .D(_01289_),
    .Q_N(_12806_),
    .Q(\top_ihp.oisc.regs[32][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][15]$_DFFE_PP_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1958),
    .D(_01290_),
    .Q_N(_12805_),
    .Q(\top_ihp.oisc.regs[32][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][16]$_DFFE_PP_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1959),
    .D(_01291_),
    .Q_N(_12804_),
    .Q(\top_ihp.oisc.regs[32][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][17]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1960),
    .D(_01292_),
    .Q_N(_12803_),
    .Q(\top_ihp.oisc.regs[32][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][18]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1961),
    .D(_01293_),
    .Q_N(_12802_),
    .Q(\top_ihp.oisc.regs[32][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][19]$_DFFE_PP_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1962),
    .D(_01294_),
    .Q_N(_12801_),
    .Q(\top_ihp.oisc.regs[32][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][1]$_DFFE_PP_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1963),
    .D(_01295_),
    .Q_N(_12800_),
    .Q(\top_ihp.oisc.regs[32][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][20]$_DFFE_PP_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1964),
    .D(_01296_),
    .Q_N(_12799_),
    .Q(\top_ihp.oisc.regs[32][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][21]$_DFFE_PP_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1965),
    .D(_01297_),
    .Q_N(_12798_),
    .Q(\top_ihp.oisc.regs[32][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][22]$_DFFE_PP_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1966),
    .D(_01298_),
    .Q_N(_12797_),
    .Q(\top_ihp.oisc.regs[32][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][23]$_DFFE_PP_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1967),
    .D(_01299_),
    .Q_N(_12796_),
    .Q(\top_ihp.oisc.regs[32][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][24]$_DFFE_PP_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1968),
    .D(_01300_),
    .Q_N(_12795_),
    .Q(\top_ihp.oisc.regs[32][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][25]$_DFFE_PP_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1969),
    .D(_01301_),
    .Q_N(_12794_),
    .Q(\top_ihp.oisc.regs[32][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][26]$_DFFE_PP_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1970),
    .D(_01302_),
    .Q_N(_12793_),
    .Q(\top_ihp.oisc.regs[32][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][27]$_DFFE_PP_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1971),
    .D(_01303_),
    .Q_N(_12792_),
    .Q(\top_ihp.oisc.regs[32][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][28]$_DFFE_PP_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1972),
    .D(_01304_),
    .Q_N(_12791_),
    .Q(\top_ihp.oisc.regs[32][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][29]$_DFFE_PP_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1973),
    .D(_01305_),
    .Q_N(_12790_),
    .Q(\top_ihp.oisc.regs[32][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][2]$_DFFE_PP_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1974),
    .D(_01306_),
    .Q_N(_12789_),
    .Q(\top_ihp.oisc.regs[32][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][30]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1975),
    .D(_01307_),
    .Q_N(_12788_),
    .Q(\top_ihp.oisc.regs[32][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][31]$_DFFE_PP_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1976),
    .D(_01308_),
    .Q_N(_12787_),
    .Q(\top_ihp.oisc.regs[32][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][3]$_DFFE_PP_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1977),
    .D(_01309_),
    .Q_N(_12786_),
    .Q(\top_ihp.oisc.regs[32][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][4]$_DFFE_PP_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1978),
    .D(_01310_),
    .Q_N(_12785_),
    .Q(\top_ihp.oisc.regs[32][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][5]$_DFFE_PP_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1979),
    .D(_01311_),
    .Q_N(_12784_),
    .Q(\top_ihp.oisc.regs[32][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][6]$_DFFE_PP_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1980),
    .D(_01312_),
    .Q_N(_12783_),
    .Q(\top_ihp.oisc.regs[32][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][7]$_DFFE_PP_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1981),
    .D(_01313_),
    .Q_N(_12782_),
    .Q(\top_ihp.oisc.regs[32][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][8]$_DFFE_PP_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1982),
    .D(_01314_),
    .Q_N(_12781_),
    .Q(\top_ihp.oisc.regs[32][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[32][9]$_DFFE_PP_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1983),
    .D(_01315_),
    .Q_N(_12780_),
    .Q(\top_ihp.oisc.regs[32][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1289),
    .D(_01316_),
    .Q_N(_12779_),
    .Q(\top_ihp.oisc.regs[33][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1151),
    .D(_01317_),
    .Q_N(_12778_),
    .Q(\top_ihp.oisc.regs[33][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1221),
    .D(_01318_),
    .Q_N(_12777_),
    .Q(\top_ihp.oisc.regs[33][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1225),
    .D(_01319_),
    .Q_N(_12776_),
    .Q(\top_ihp.oisc.regs[33][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1298),
    .D(_01320_),
    .Q_N(_12775_),
    .Q(\top_ihp.oisc.regs[33][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1299),
    .D(_01321_),
    .Q_N(_12774_),
    .Q(\top_ihp.oisc.regs[33][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1297),
    .D(_01322_),
    .Q_N(_12773_),
    .Q(\top_ihp.oisc.regs[33][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1299),
    .D(_01323_),
    .Q_N(_12772_),
    .Q(\top_ihp.oisc.regs[33][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_01324_),
    .Q_N(_12771_),
    .Q(\top_ihp.oisc.regs[33][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1295),
    .D(_01325_),
    .Q_N(_12770_),
    .Q(\top_ihp.oisc.regs[33][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1272),
    .D(_01326_),
    .Q_N(_12769_),
    .Q(\top_ihp.oisc.regs[33][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1209),
    .D(_01327_),
    .Q_N(_12768_),
    .Q(\top_ihp.oisc.regs[33][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1236),
    .D(_01328_),
    .Q_N(_12767_),
    .Q(\top_ihp.oisc.regs[33][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1236),
    .D(_01329_),
    .Q_N(_12766_),
    .Q(\top_ihp.oisc.regs[33][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1237),
    .D(_01330_),
    .Q_N(_12765_),
    .Q(\top_ihp.oisc.regs[33][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1177),
    .D(_01331_),
    .Q_N(_12764_),
    .Q(\top_ihp.oisc.regs[33][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1142),
    .D(_01332_),
    .Q_N(_12763_),
    .Q(\top_ihp.oisc.regs[33][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_01333_),
    .Q_N(_12762_),
    .Q(\top_ihp.oisc.regs[33][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1177),
    .D(_01334_),
    .Q_N(_12761_),
    .Q(\top_ihp.oisc.regs[33][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1284),
    .D(_01335_),
    .Q_N(_12760_),
    .Q(\top_ihp.oisc.regs[33][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1229),
    .D(_01336_),
    .Q_N(_12759_),
    .Q(\top_ihp.oisc.regs[33][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1168),
    .D(_01337_),
    .Q_N(_12758_),
    .Q(\top_ihp.oisc.regs[33][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1186),
    .D(_01338_),
    .Q_N(_12757_),
    .Q(\top_ihp.oisc.regs[33][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1185),
    .D(_01339_),
    .Q_N(_12756_),
    .Q(\top_ihp.oisc.regs[33][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1234),
    .D(_01340_),
    .Q_N(_12755_),
    .Q(\top_ihp.oisc.regs[33][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1283),
    .D(_01341_),
    .Q_N(_12754_),
    .Q(\top_ihp.oisc.regs[33][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1151),
    .D(_01342_),
    .Q_N(_12753_),
    .Q(\top_ihp.oisc.regs[33][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1266),
    .D(_01343_),
    .Q_N(_12752_),
    .Q(\top_ihp.oisc.regs[33][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1287),
    .D(_01344_),
    .Q_N(_12751_),
    .Q(\top_ihp.oisc.regs[33][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1160),
    .D(_01345_),
    .Q_N(_12750_),
    .Q(\top_ihp.oisc.regs[33][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1206),
    .D(_01346_),
    .Q_N(_12749_),
    .Q(\top_ihp.oisc.regs[33][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[33][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1214),
    .D(_01347_),
    .Q_N(_12748_),
    .Q(\top_ihp.oisc.regs[33][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1292),
    .D(_01348_),
    .Q_N(_12747_),
    .Q(\top_ihp.oisc.regs[34][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1151),
    .D(_01349_),
    .Q_N(_12746_),
    .Q(\top_ihp.oisc.regs[34][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1221),
    .D(_01350_),
    .Q_N(_12745_),
    .Q(\top_ihp.oisc.regs[34][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1225),
    .D(_01351_),
    .Q_N(_12744_),
    .Q(\top_ihp.oisc.regs[34][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1313),
    .D(_01352_),
    .Q_N(_12743_),
    .Q(\top_ihp.oisc.regs[34][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1300),
    .D(_01353_),
    .Q_N(_12742_),
    .Q(\top_ihp.oisc.regs[34][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][15]$_DFFE_PN1P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1297),
    .D(_01354_),
    .Q_N(\top_ihp.oisc.regs[34][15] ),
    .Q(_00336_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1312),
    .D(_01355_),
    .Q_N(_12741_),
    .Q(\top_ihp.oisc.regs[34][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1296),
    .D(_01356_),
    .Q_N(_12740_),
    .Q(\top_ihp.oisc.regs[34][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1295),
    .D(_01357_),
    .Q_N(_12739_),
    .Q(\top_ihp.oisc.regs[34][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1291),
    .D(_01358_),
    .Q_N(_12738_),
    .Q(\top_ihp.oisc.regs[34][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1208),
    .D(_01359_),
    .Q_N(_12737_),
    .Q(\top_ihp.oisc.regs[34][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1244),
    .D(_01360_),
    .Q_N(_12736_),
    .Q(\top_ihp.oisc.regs[34][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1245),
    .D(_01361_),
    .Q_N(_12735_),
    .Q(\top_ihp.oisc.regs[34][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1177),
    .D(_01362_),
    .Q_N(_12734_),
    .Q(\top_ihp.oisc.regs[34][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1178),
    .D(_01363_),
    .Q_N(_12733_),
    .Q(\top_ihp.oisc.regs[34][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1142),
    .D(_01364_),
    .Q_N(_12732_),
    .Q(\top_ihp.oisc.regs[34][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1180),
    .D(_01365_),
    .Q_N(_12731_),
    .Q(\top_ihp.oisc.regs[34][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1172),
    .D(_01366_),
    .Q_N(_12730_),
    .Q(\top_ihp.oisc.regs[34][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][27]$_DFFE_PN1P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1147),
    .D(_01367_),
    .Q_N(\top_ihp.oisc.regs[34][27] ),
    .Q(_00337_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1236),
    .D(_01368_),
    .Q_N(_12729_),
    .Q(\top_ihp.oisc.regs[34][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1168),
    .D(_01369_),
    .Q_N(_12728_),
    .Q(\top_ihp.oisc.regs[34][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1166),
    .D(_01370_),
    .Q_N(_12727_),
    .Q(\top_ihp.oisc.regs[34][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1166),
    .D(_01371_),
    .Q_N(_12726_),
    .Q(\top_ihp.oisc.regs[34][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1234),
    .D(_01372_),
    .Q_N(_12725_),
    .Q(\top_ihp.oisc.regs[34][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1286),
    .D(_01373_),
    .Q_N(_12724_),
    .Q(\top_ihp.oisc.regs[34][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1152),
    .D(_01374_),
    .Q_N(_12723_),
    .Q(\top_ihp.oisc.regs[34][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1217),
    .D(_01375_),
    .Q_N(_12722_),
    .Q(\top_ihp.oisc.regs[34][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1200),
    .D(_01376_),
    .Q_N(_12721_),
    .Q(\top_ihp.oisc.regs[34][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1185),
    .D(_01377_),
    .Q_N(_12720_),
    .Q(\top_ihp.oisc.regs[34][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1149),
    .D(_01378_),
    .Q_N(_12719_),
    .Q(\top_ihp.oisc.regs[34][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[34][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1268),
    .D(_01379_),
    .Q_N(_12718_),
    .Q(\top_ihp.oisc.regs[34][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1313),
    .D(_01380_),
    .Q_N(_12717_),
    .Q(\top_ihp.oisc.regs[35][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1156),
    .D(_01381_),
    .Q_N(_12716_),
    .Q(\top_ihp.oisc.regs[35][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][11]$_DFFE_PN1P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1208),
    .D(_01382_),
    .Q_N(\top_ihp.oisc.regs[35][11] ),
    .Q(_00338_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1225),
    .D(_01383_),
    .Q_N(_12715_),
    .Q(\top_ihp.oisc.regs[35][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1251),
    .D(_01384_),
    .Q_N(_12714_),
    .Q(\top_ihp.oisc.regs[35][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1318),
    .D(_01385_),
    .Q_N(_12713_),
    .Q(\top_ihp.oisc.regs[35][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1317),
    .D(_01386_),
    .Q_N(_12712_),
    .Q(\top_ihp.oisc.regs[35][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1317),
    .D(_01387_),
    .Q_N(_12711_),
    .Q(\top_ihp.oisc.regs[35][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1257),
    .D(_01388_),
    .Q_N(_12710_),
    .Q(\top_ihp.oisc.regs[35][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1305),
    .D(_01389_),
    .Q_N(_12709_),
    .Q(\top_ihp.oisc.regs[35][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_200_clk),
    .RESET_B(net1333),
    .D(_01390_),
    .Q_N(_12708_),
    .Q(\top_ihp.oisc.regs[35][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1225),
    .D(_01391_),
    .Q_N(_12707_),
    .Q(\top_ihp.oisc.regs[35][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1255),
    .D(_01392_),
    .Q_N(_12706_),
    .Q(\top_ihp.oisc.regs[35][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1248),
    .D(_01393_),
    .Q_N(_12705_),
    .Q(\top_ihp.oisc.regs[35][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1172),
    .D(_01394_),
    .Q_N(_12704_),
    .Q(\top_ihp.oisc.regs[35][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1172),
    .D(_01395_),
    .Q_N(_12703_),
    .Q(\top_ihp.oisc.regs[35][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1144),
    .D(_01396_),
    .Q_N(_12702_),
    .Q(\top_ihp.oisc.regs[35][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1177),
    .D(_01397_),
    .Q_N(_12701_),
    .Q(\top_ihp.oisc.regs[35][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1174),
    .D(_01398_),
    .Q_N(_12700_),
    .Q(\top_ihp.oisc.regs[35][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1147),
    .D(_01399_),
    .Q_N(_12699_),
    .Q(\top_ihp.oisc.regs[35][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1163),
    .D(_01400_),
    .Q_N(_12698_),
    .Q(\top_ihp.oisc.regs[35][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1172),
    .D(_01401_),
    .Q_N(_12697_),
    .Q(\top_ihp.oisc.regs[35][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1231),
    .D(_01402_),
    .Q_N(_12696_),
    .Q(\top_ihp.oisc.regs[35][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1229),
    .D(_01403_),
    .Q_N(_12695_),
    .Q(\top_ihp.oisc.regs[35][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][31]$_DFFE_PN1P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1234),
    .D(_01404_),
    .Q_N(\top_ihp.oisc.regs[35][31] ),
    .Q(_00339_));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1283),
    .D(_01405_),
    .Q_N(_12694_),
    .Q(\top_ihp.oisc.regs[35][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1329),
    .D(_01406_),
    .Q_N(_12693_),
    .Q(\top_ihp.oisc.regs[35][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1287),
    .D(_01407_),
    .Q_N(_12692_),
    .Q(\top_ihp.oisc.regs[35][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1200),
    .D(_01408_),
    .Q_N(_12691_),
    .Q(\top_ihp.oisc.regs[35][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1229),
    .D(_01409_),
    .Q_N(_12690_),
    .Q(\top_ihp.oisc.regs[35][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1206),
    .D(_01410_),
    .Q_N(_12689_),
    .Q(\top_ihp.oisc.regs[35][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[35][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1200),
    .D(_01411_),
    .Q_N(_12688_),
    .Q(\top_ihp.oisc.regs[35][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1289),
    .D(_01412_),
    .Q_N(_12687_),
    .Q(\top_ihp.oisc.regs[36][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1328),
    .D(_01413_),
    .Q_N(_12686_),
    .Q(\top_ihp.oisc.regs[36][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1221),
    .D(_01414_),
    .Q_N(_12685_),
    .Q(\top_ihp.oisc.regs[36][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1226),
    .D(_01415_),
    .Q_N(_12684_),
    .Q(\top_ihp.oisc.regs[36][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1295),
    .D(_01416_),
    .Q_N(_12683_),
    .Q(\top_ihp.oisc.regs[36][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1304),
    .D(_01417_),
    .Q_N(_12682_),
    .Q(\top_ihp.oisc.regs[36][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1297),
    .D(_01418_),
    .Q_N(_12681_),
    .Q(\top_ihp.oisc.regs[36][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1304),
    .D(_01419_),
    .Q_N(_12680_),
    .Q(\top_ihp.oisc.regs[36][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1262),
    .D(_01420_),
    .Q_N(_12679_),
    .Q(\top_ihp.oisc.regs[36][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1304),
    .D(_01421_),
    .Q_N(_12678_),
    .Q(\top_ihp.oisc.regs[36][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1272),
    .D(_01422_),
    .Q_N(_12677_),
    .Q(\top_ihp.oisc.regs[36][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1222),
    .D(_01423_),
    .Q_N(_12676_),
    .Q(\top_ihp.oisc.regs[36][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1244),
    .D(_01424_),
    .Q_N(_12675_),
    .Q(\top_ihp.oisc.regs[36][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1241),
    .D(_01425_),
    .Q_N(_12674_),
    .Q(\top_ihp.oisc.regs[36][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1179),
    .D(_01426_),
    .Q_N(_12673_),
    .Q(\top_ihp.oisc.regs[36][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(_01427_),
    .Q_N(_12672_),
    .Q(\top_ihp.oisc.regs[36][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1142),
    .D(_01428_),
    .Q_N(_12671_),
    .Q(\top_ihp.oisc.regs[36][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1240),
    .D(_01429_),
    .Q_N(_12670_),
    .Q(\top_ihp.oisc.regs[36][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1193),
    .D(_01430_),
    .Q_N(_12669_),
    .Q(\top_ihp.oisc.regs[36][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1147),
    .D(_01431_),
    .Q_N(_12668_),
    .Q(\top_ihp.oisc.regs[36][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1187),
    .D(_01432_),
    .Q_N(_12667_),
    .Q(\top_ihp.oisc.regs[36][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1179),
    .D(_01433_),
    .Q_N(_12666_),
    .Q(\top_ihp.oisc.regs[36][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1168),
    .D(_01434_),
    .Q_N(_12665_),
    .Q(\top_ihp.oisc.regs[36][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1166),
    .D(_01435_),
    .Q_N(_12664_),
    .Q(\top_ihp.oisc.regs[36][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1230),
    .D(_01436_),
    .Q_N(_12663_),
    .Q(\top_ihp.oisc.regs[36][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1283),
    .D(_01437_),
    .Q_N(_12662_),
    .Q(\top_ihp.oisc.regs[36][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1154),
    .D(_01438_),
    .Q_N(_12661_),
    .Q(\top_ihp.oisc.regs[36][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1267),
    .D(_01439_),
    .Q_N(_12660_),
    .Q(\top_ihp.oisc.regs[36][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1201),
    .D(_01440_),
    .Q_N(_12659_),
    .Q(\top_ihp.oisc.regs[36][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1158),
    .D(_01441_),
    .Q_N(_12658_),
    .Q(\top_ihp.oisc.regs[36][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1147),
    .D(_01442_),
    .Q_N(_12657_),
    .Q(\top_ihp.oisc.regs[36][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[36][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1212),
    .D(_01443_),
    .Q_N(_12656_),
    .Q(\top_ihp.oisc.regs[36][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1287),
    .D(_01444_),
    .Q_N(_12655_),
    .Q(\top_ihp.oisc.regs[37][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1154),
    .D(_01445_),
    .Q_N(_12654_),
    .Q(\top_ihp.oisc.regs[37][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1222),
    .D(_01446_),
    .Q_N(_12653_),
    .Q(\top_ihp.oisc.regs[37][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1225),
    .D(_01447_),
    .Q_N(_12652_),
    .Q(\top_ihp.oisc.regs[37][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1313),
    .D(_01448_),
    .Q_N(_12651_),
    .Q(\top_ihp.oisc.regs[37][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1307),
    .D(_01449_),
    .Q_N(_12650_),
    .Q(\top_ihp.oisc.regs[37][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1276),
    .D(_01450_),
    .Q_N(_12649_),
    .Q(\top_ihp.oisc.regs[37][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1312),
    .D(_01451_),
    .Q_N(_12648_),
    .Q(\top_ihp.oisc.regs[37][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1259),
    .D(_01452_),
    .Q_N(_12647_),
    .Q(\top_ihp.oisc.regs[37][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1318),
    .D(_01453_),
    .Q_N(_12646_),
    .Q(\top_ihp.oisc.regs[37][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1284),
    .D(_01454_),
    .Q_N(_12645_),
    .Q(\top_ihp.oisc.regs[37][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1222),
    .D(_01455_),
    .Q_N(_12644_),
    .Q(\top_ihp.oisc.regs[37][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1243),
    .D(_01456_),
    .Q_N(_12643_),
    .Q(\top_ihp.oisc.regs[37][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1243),
    .D(_01457_),
    .Q_N(_12642_),
    .Q(\top_ihp.oisc.regs[37][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1190),
    .D(_01458_),
    .Q_N(_12641_),
    .Q(\top_ihp.oisc.regs[37][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1244),
    .D(_01459_),
    .Q_N(_12640_),
    .Q(\top_ihp.oisc.regs[37][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1154),
    .D(_01460_),
    .Q_N(_12639_),
    .Q(\top_ihp.oisc.regs[37][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(_01461_),
    .Q_N(_12638_),
    .Q(\top_ihp.oisc.regs[37][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1190),
    .D(_01462_),
    .Q_N(_12637_),
    .Q(\top_ihp.oisc.regs[37][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1218),
    .D(_01463_),
    .Q_N(_12636_),
    .Q(\top_ihp.oisc.regs[37][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1185),
    .D(_01464_),
    .Q_N(_12635_),
    .Q(\top_ihp.oisc.regs[37][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1179),
    .D(_01465_),
    .Q_N(_12634_),
    .Q(\top_ihp.oisc.regs[37][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1186),
    .D(_01466_),
    .Q_N(_12633_),
    .Q(\top_ihp.oisc.regs[37][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1167),
    .D(_01467_),
    .Q_N(_12632_),
    .Q(\top_ihp.oisc.regs[37][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1234),
    .D(_01468_),
    .Q_N(_12631_),
    .Q(\top_ihp.oisc.regs[37][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1283),
    .D(_01469_),
    .Q_N(_12630_),
    .Q(\top_ihp.oisc.regs[37][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1198),
    .D(_01470_),
    .Q_N(_12629_),
    .Q(\top_ihp.oisc.regs[37][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1286),
    .D(_01471_),
    .Q_N(_12628_),
    .Q(\top_ihp.oisc.regs[37][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1201),
    .D(_01472_),
    .Q_N(_12627_),
    .Q(\top_ihp.oisc.regs[37][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1230),
    .D(_01473_),
    .Q_N(_12626_),
    .Q(\top_ihp.oisc.regs[37][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1209),
    .D(_01474_),
    .Q_N(_12625_),
    .Q(\top_ihp.oisc.regs[37][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[37][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1212),
    .D(_01475_),
    .Q_N(_12624_),
    .Q(\top_ihp.oisc.regs[37][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1272),
    .D(_01476_),
    .Q_N(_12623_),
    .Q(\top_ihp.oisc.regs[38][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1151),
    .D(_01477_),
    .Q_N(_12622_),
    .Q(\top_ihp.oisc.regs[38][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1224),
    .D(_01478_),
    .Q_N(_12621_),
    .Q(\top_ihp.oisc.regs[38][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1275),
    .D(_01479_),
    .Q_N(_12620_),
    .Q(\top_ihp.oisc.regs[38][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1252),
    .D(_01480_),
    .Q_N(_12619_),
    .Q(\top_ihp.oisc.regs[38][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1307),
    .D(_01481_),
    .Q_N(_12618_),
    .Q(\top_ihp.oisc.regs[38][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1298),
    .D(_01482_),
    .Q_N(_12617_),
    .Q(\top_ihp.oisc.regs[38][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1299),
    .D(_01483_),
    .Q_N(_12616_),
    .Q(\top_ihp.oisc.regs[38][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1259),
    .D(_01484_),
    .Q_N(_12615_),
    .Q(\top_ihp.oisc.regs[38][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1307),
    .D(_01485_),
    .Q_N(_12614_),
    .Q(\top_ihp.oisc.regs[38][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1280),
    .D(_01486_),
    .Q_N(_12613_),
    .Q(\top_ihp.oisc.regs[38][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1208),
    .D(_01487_),
    .Q_N(_12612_),
    .Q(\top_ihp.oisc.regs[38][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1244),
    .D(_01488_),
    .Q_N(_12611_),
    .Q(\top_ihp.oisc.regs[38][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1243),
    .D(_01489_),
    .Q_N(_12610_),
    .Q(\top_ihp.oisc.regs[38][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1191),
    .D(_01490_),
    .Q_N(_12609_),
    .Q(\top_ihp.oisc.regs[38][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1193),
    .D(_01491_),
    .Q_N(_12608_),
    .Q(\top_ihp.oisc.regs[38][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1142),
    .D(_01492_),
    .Q_N(_12607_),
    .Q(\top_ihp.oisc.regs[38][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1256),
    .D(_01493_),
    .Q_N(_12606_),
    .Q(\top_ihp.oisc.regs[38][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1189),
    .D(_01494_),
    .Q_N(_12605_),
    .Q(\top_ihp.oisc.regs[38][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1158),
    .D(_01495_),
    .Q_N(_12604_),
    .Q(\top_ihp.oisc.regs[38][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1162),
    .D(_01496_),
    .Q_N(_12603_),
    .Q(\top_ihp.oisc.regs[38][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1168),
    .D(_01497_),
    .Q_N(_12602_),
    .Q(\top_ihp.oisc.regs[38][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1167),
    .D(_01498_),
    .Q_N(_12601_),
    .Q(\top_ihp.oisc.regs[38][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1297),
    .D(_01499_),
    .Q_N(_12600_),
    .Q(\top_ihp.oisc.regs[38][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1248),
    .D(_01500_),
    .Q_N(_12599_),
    .Q(\top_ihp.oisc.regs[38][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1283),
    .D(_01501_),
    .Q_N(_12598_),
    .Q(\top_ihp.oisc.regs[38][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1285),
    .D(_01502_),
    .Q_N(_12597_),
    .Q(\top_ihp.oisc.regs[38][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1217),
    .D(_01503_),
    .Q_N(_12596_),
    .Q(\top_ihp.oisc.regs[38][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1200),
    .D(_01504_),
    .Q_N(_12595_),
    .Q(\top_ihp.oisc.regs[38][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1161),
    .D(_01505_),
    .Q_N(_12594_),
    .Q(\top_ihp.oisc.regs[38][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1147),
    .D(_01506_),
    .Q_N(_12593_),
    .Q(\top_ihp.oisc.regs[38][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[38][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1214),
    .D(_01507_),
    .Q_N(_12592_),
    .Q(\top_ihp.oisc.regs[38][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1289),
    .D(_01508_),
    .Q_N(_12591_),
    .Q(\top_ihp.oisc.regs[39][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1154),
    .D(_01509_),
    .Q_N(_12590_),
    .Q(\top_ihp.oisc.regs[39][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1276),
    .D(_01510_),
    .Q_N(_12589_),
    .Q(\top_ihp.oisc.regs[39][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1224),
    .D(_01511_),
    .Q_N(_12588_),
    .Q(\top_ihp.oisc.regs[39][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1252),
    .D(_01512_),
    .Q_N(_12587_),
    .Q(\top_ihp.oisc.regs[39][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1259),
    .D(_01513_),
    .Q_N(_12586_),
    .Q(\top_ihp.oisc.regs[39][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1252),
    .D(_01514_),
    .Q_N(_12585_),
    .Q(\top_ihp.oisc.regs[39][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1295),
    .D(_01515_),
    .Q_N(_12584_),
    .Q(\top_ihp.oisc.regs[39][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1259),
    .D(_01516_),
    .Q_N(_12583_),
    .Q(\top_ihp.oisc.regs[39][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1303),
    .D(_01517_),
    .Q_N(_12582_),
    .Q(\top_ihp.oisc.regs[39][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1280),
    .D(_01518_),
    .Q_N(_12581_),
    .Q(\top_ihp.oisc.regs[39][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1222),
    .D(_01519_),
    .Q_N(_12580_),
    .Q(\top_ihp.oisc.regs[39][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1255),
    .D(_01520_),
    .Q_N(_12579_),
    .Q(\top_ihp.oisc.regs[39][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1241),
    .D(_01521_),
    .Q_N(_12578_),
    .Q(\top_ihp.oisc.regs[39][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1186),
    .D(_01522_),
    .Q_N(_12577_),
    .Q(\top_ihp.oisc.regs[39][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1241),
    .D(_01523_),
    .Q_N(_12576_),
    .Q(\top_ihp.oisc.regs[39][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1154),
    .D(_01524_),
    .Q_N(_12575_),
    .Q(\top_ihp.oisc.regs[39][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1239),
    .D(_01525_),
    .Q_N(_12574_),
    .Q(\top_ihp.oisc.regs[39][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1240),
    .D(_01526_),
    .Q_N(_12573_),
    .Q(\top_ihp.oisc.regs[39][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1156),
    .D(_01527_),
    .Q_N(_12572_),
    .Q(\top_ihp.oisc.regs[39][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1231),
    .D(_01528_),
    .Q_N(_12571_),
    .Q(\top_ihp.oisc.regs[39][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1189),
    .D(_01529_),
    .Q_N(_12570_),
    .Q(\top_ihp.oisc.regs[39][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1186),
    .D(_01530_),
    .Q_N(_12569_),
    .Q(\top_ihp.oisc.regs[39][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1182),
    .D(_01531_),
    .Q_N(_12568_),
    .Q(\top_ihp.oisc.regs[39][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1229),
    .D(_01532_),
    .Q_N(_12567_),
    .Q(\top_ihp.oisc.regs[39][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1266),
    .D(_01533_),
    .Q_N(_12566_),
    .Q(\top_ihp.oisc.regs[39][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1270),
    .D(_01534_),
    .Q_N(_12565_),
    .Q(\top_ihp.oisc.regs[39][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1267),
    .D(_01535_),
    .Q_N(_12564_),
    .Q(\top_ihp.oisc.regs[39][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1203),
    .D(_01536_),
    .Q_N(_12563_),
    .Q(\top_ihp.oisc.regs[39][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1276),
    .D(_01537_),
    .Q_N(_12562_),
    .Q(\top_ihp.oisc.regs[39][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1163),
    .D(_01538_),
    .Q_N(_12561_),
    .Q(\top_ihp.oisc.regs[39][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[39][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1214),
    .D(_01539_),
    .Q_N(_12560_),
    .Q(\top_ihp.oisc.regs[39][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1388),
    .D(_01540_),
    .Q_N(_12559_),
    .Q(\top_ihp.oisc.regs[3][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1383),
    .D(_01541_),
    .Q_N(_12558_),
    .Q(\top_ihp.oisc.regs[3][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_226_clk),
    .RESET_B(net1391),
    .D(_01542_),
    .Q_N(_12557_),
    .Q(\top_ihp.oisc.regs[3][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1341),
    .D(_01543_),
    .Q_N(_12556_),
    .Q(\top_ihp.oisc.regs[3][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1350),
    .D(_01544_),
    .Q_N(_12555_),
    .Q(\top_ihp.oisc.regs[3][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1350),
    .D(_01545_),
    .Q_N(_12554_),
    .Q(\top_ihp.oisc.regs[3][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1359),
    .D(_01546_),
    .Q_N(_12553_),
    .Q(\top_ihp.oisc.regs[3][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1356),
    .D(_01547_),
    .Q_N(_12552_),
    .Q(\top_ihp.oisc.regs[3][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1356),
    .D(_01548_),
    .Q_N(_12551_),
    .Q(\top_ihp.oisc.regs[3][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1356),
    .D(_01549_),
    .Q_N(_12550_),
    .Q(\top_ihp.oisc.regs[3][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1344),
    .D(_01550_),
    .Q_N(_12549_),
    .Q(\top_ihp.oisc.regs[3][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1378),
    .D(_01551_),
    .Q_N(_12548_),
    .Q(\top_ihp.oisc.regs[3][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1356),
    .D(_01552_),
    .Q_N(_12547_),
    .Q(\top_ihp.oisc.regs[3][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1355),
    .D(_01553_),
    .Q_N(_12546_),
    .Q(\top_ihp.oisc.regs[3][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1356),
    .D(_01554_),
    .Q_N(_12545_),
    .Q(\top_ihp.oisc.regs[3][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_135_clk),
    .RESET_B(net1355),
    .D(_01555_),
    .Q_N(_12544_),
    .Q(\top_ihp.oisc.regs[3][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1340),
    .D(_01556_),
    .Q_N(_12543_),
    .Q(\top_ihp.oisc.regs[3][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1355),
    .D(_01557_),
    .Q_N(_12542_),
    .Q(\top_ihp.oisc.regs[3][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1355),
    .D(_01558_),
    .Q_N(_12541_),
    .Q(\top_ihp.oisc.regs[3][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1380),
    .D(_01559_),
    .Q_N(_12540_),
    .Q(\top_ihp.oisc.regs[3][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1389),
    .D(_01560_),
    .Q_N(_12539_),
    .Q(\top_ihp.oisc.regs[3][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1354),
    .D(_01561_),
    .Q_N(_12538_),
    .Q(\top_ihp.oisc.regs[3][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1348),
    .D(_01562_),
    .Q_N(_12537_),
    .Q(\top_ihp.oisc.regs[3][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1348),
    .D(_01563_),
    .Q_N(_12536_),
    .Q(\top_ihp.oisc.regs[3][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1348),
    .D(_01564_),
    .Q_N(_12535_),
    .Q(\top_ihp.oisc.regs[3][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1337),
    .D(_01565_),
    .Q_N(_12534_),
    .Q(\top_ihp.oisc.regs[3][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1391),
    .D(_01566_),
    .Q_N(_12533_),
    .Q(\top_ihp.oisc.regs[3][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1338),
    .D(_01567_),
    .Q_N(_12532_),
    .Q(\top_ihp.oisc.regs[3][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1385),
    .D(_01568_),
    .Q_N(_12531_),
    .Q(\top_ihp.oisc.regs[3][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1348),
    .D(_01569_),
    .Q_N(_12530_),
    .Q(\top_ihp.oisc.regs[3][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1331),
    .D(_01570_),
    .Q_N(_12529_),
    .Q(\top_ihp.oisc.regs[3][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[3][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_251_clk),
    .RESET_B(net1373),
    .D(_01571_),
    .Q_N(_12528_),
    .Q(\top_ihp.oisc.regs[3][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1279),
    .D(_01572_),
    .Q_N(_12527_),
    .Q(\top_ihp.oisc.regs[40][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1151),
    .D(_01573_),
    .Q_N(_12526_),
    .Q(\top_ihp.oisc.regs[40][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1275),
    .D(_01574_),
    .Q_N(_12525_),
    .Q(\top_ihp.oisc.regs[40][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1278),
    .D(_01575_),
    .Q_N(_12524_),
    .Q(\top_ihp.oisc.regs[40][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1251),
    .D(_01576_),
    .Q_N(_12523_),
    .Q(\top_ihp.oisc.regs[40][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1299),
    .D(_01577_),
    .Q_N(_12522_),
    .Q(\top_ihp.oisc.regs[40][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1276),
    .D(_01578_),
    .Q_N(_12521_),
    .Q(\top_ihp.oisc.regs[40][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1299),
    .D(_01579_),
    .Q_N(_12520_),
    .Q(\top_ihp.oisc.regs[40][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1259),
    .D(_01580_),
    .Q_N(_12519_),
    .Q(\top_ihp.oisc.regs[40][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1303),
    .D(_01581_),
    .Q_N(_12518_),
    .Q(\top_ihp.oisc.regs[40][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1268),
    .D(_01582_),
    .Q_N(_12517_),
    .Q(\top_ihp.oisc.regs[40][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1203),
    .D(_01583_),
    .Q_N(_12516_),
    .Q(\top_ihp.oisc.regs[40][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1243),
    .D(_01584_),
    .Q_N(_12515_),
    .Q(\top_ihp.oisc.regs[40][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1239),
    .D(_01585_),
    .Q_N(_12514_),
    .Q(\top_ihp.oisc.regs[40][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_01586_),
    .Q_N(_12513_),
    .Q(\top_ihp.oisc.regs[40][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1195),
    .D(_01587_),
    .Q_N(_12512_),
    .Q(\top_ihp.oisc.regs[40][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1144),
    .D(_01588_),
    .Q_N(_12511_),
    .Q(\top_ihp.oisc.regs[40][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1195),
    .D(_01589_),
    .Q_N(_12510_),
    .Q(\top_ihp.oisc.regs[40][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1298),
    .D(_01590_),
    .Q_N(_12509_),
    .Q(\top_ihp.oisc.regs[40][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1144),
    .D(_01591_),
    .Q_N(_12508_),
    .Q(\top_ihp.oisc.regs[40][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1156),
    .D(_01592_),
    .Q_N(_12507_),
    .Q(\top_ihp.oisc.regs[40][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1186),
    .D(_01593_),
    .Q_N(_12506_),
    .Q(\top_ihp.oisc.regs[40][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1187),
    .D(_01594_),
    .Q_N(_12505_),
    .Q(\top_ihp.oisc.regs[40][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1159),
    .D(_01595_),
    .Q_N(_12504_),
    .Q(\top_ihp.oisc.regs[40][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1206),
    .D(_01596_),
    .Q_N(_12503_),
    .Q(\top_ihp.oisc.regs[40][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1267),
    .D(_01597_),
    .Q_N(_12502_),
    .Q(\top_ihp.oisc.regs[40][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1198),
    .D(_01598_),
    .Q_N(_12501_),
    .Q(\top_ihp.oisc.regs[40][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1198),
    .D(_01599_),
    .Q_N(_12500_),
    .Q(\top_ihp.oisc.regs[40][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1269),
    .D(_01600_),
    .Q_N(_12499_),
    .Q(\top_ihp.oisc.regs[40][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1160),
    .D(_01601_),
    .Q_N(_12498_),
    .Q(\top_ihp.oisc.regs[40][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1163),
    .D(_01602_),
    .Q_N(_12497_),
    .Q(\top_ihp.oisc.regs[40][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[40][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1217),
    .D(_01603_),
    .Q_N(_12496_),
    .Q(\top_ihp.oisc.regs[40][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1279),
    .D(_01604_),
    .Q_N(_12495_),
    .Q(\top_ihp.oisc.regs[41][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1153),
    .D(_01605_),
    .Q_N(_12494_),
    .Q(\top_ihp.oisc.regs[41][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1224),
    .D(_01606_),
    .Q_N(_12493_),
    .Q(\top_ihp.oisc.regs[41][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1275),
    .D(_01607_),
    .Q_N(_12492_),
    .Q(\top_ihp.oisc.regs[41][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1251),
    .D(_01608_),
    .Q_N(_12491_),
    .Q(\top_ihp.oisc.regs[41][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1305),
    .D(_01609_),
    .Q_N(_12490_),
    .Q(\top_ihp.oisc.regs[41][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1297),
    .D(_01610_),
    .Q_N(_12489_),
    .Q(\top_ihp.oisc.regs[41][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1304),
    .D(_01611_),
    .Q_N(_12488_),
    .Q(\top_ihp.oisc.regs[41][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1261),
    .D(_01612_),
    .Q_N(_12487_),
    .Q(\top_ihp.oisc.regs[41][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1261),
    .D(_01613_),
    .Q_N(_12486_),
    .Q(\top_ihp.oisc.regs[41][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1280),
    .D(_01614_),
    .Q_N(_12485_),
    .Q(\top_ihp.oisc.regs[41][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1209),
    .D(_01615_),
    .Q_N(_12484_),
    .Q(\top_ihp.oisc.regs[41][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1244),
    .D(_01616_),
    .Q_N(_12483_),
    .Q(\top_ihp.oisc.regs[41][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1244),
    .D(_01617_),
    .Q_N(_12482_),
    .Q(\top_ihp.oisc.regs[41][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1240),
    .D(_01618_),
    .Q_N(_12481_),
    .Q(\top_ihp.oisc.regs[41][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(_01619_),
    .Q_N(_12480_),
    .Q(\top_ihp.oisc.regs[41][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1155),
    .D(_01620_),
    .Q_N(_12479_),
    .Q(\top_ihp.oisc.regs[41][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1191),
    .D(_01621_),
    .Q_N(_12478_),
    .Q(\top_ihp.oisc.regs[41][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1190),
    .D(_01622_),
    .Q_N(_12477_),
    .Q(\top_ihp.oisc.regs[41][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1153),
    .D(_01623_),
    .Q_N(_12476_),
    .Q(\top_ihp.oisc.regs[41][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1231),
    .D(_01624_),
    .Q_N(_12475_),
    .Q(\top_ihp.oisc.regs[41][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1190),
    .D(_01625_),
    .Q_N(_12474_),
    .Q(\top_ihp.oisc.regs[41][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1183),
    .D(_01626_),
    .Q_N(_12473_),
    .Q(\top_ihp.oisc.regs[41][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1182),
    .D(_01627_),
    .Q_N(_12472_),
    .Q(\top_ihp.oisc.regs[41][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1234),
    .D(_01628_),
    .Q_N(_12471_),
    .Q(\top_ihp.oisc.regs[41][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1270),
    .D(_01629_),
    .Q_N(_12470_),
    .Q(\top_ihp.oisc.regs[41][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1151),
    .D(_01630_),
    .Q_N(_12469_),
    .Q(\top_ihp.oisc.regs[41][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1199),
    .D(_01631_),
    .Q_N(_12468_),
    .Q(\top_ihp.oisc.regs[41][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1203),
    .D(_01632_),
    .Q_N(_12467_),
    .Q(\top_ihp.oisc.regs[41][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1206),
    .D(_01633_),
    .Q_N(_12466_),
    .Q(\top_ihp.oisc.regs[41][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1158),
    .D(_01634_),
    .Q_N(_12465_),
    .Q(\top_ihp.oisc.regs[41][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[41][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1215),
    .D(_01635_),
    .Q_N(_12464_),
    .Q(\top_ihp.oisc.regs[41][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1287),
    .D(_01636_),
    .Q_N(_12463_),
    .Q(\top_ihp.oisc.regs[42][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1153),
    .D(_01637_),
    .Q_N(_12462_),
    .Q(\top_ihp.oisc.regs[42][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1223),
    .D(_01638_),
    .Q_N(_12461_),
    .Q(\top_ihp.oisc.regs[42][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1276),
    .D(_01639_),
    .Q_N(_12460_),
    .Q(\top_ihp.oisc.regs[42][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1295),
    .D(_01640_),
    .Q_N(_12459_),
    .Q(\top_ihp.oisc.regs[42][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_01641_),
    .Q_N(_12458_),
    .Q(\top_ihp.oisc.regs[42][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1297),
    .D(_01642_),
    .Q_N(_12457_),
    .Q(\top_ihp.oisc.regs[42][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1296),
    .D(_01643_),
    .Q_N(_12456_),
    .Q(\top_ihp.oisc.regs[42][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1255),
    .D(_01644_),
    .Q_N(_12455_),
    .Q(\top_ihp.oisc.regs[42][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1259),
    .D(_01645_),
    .Q_N(_12454_),
    .Q(\top_ihp.oisc.regs[42][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1276),
    .D(_01646_),
    .Q_N(_12453_),
    .Q(\top_ihp.oisc.regs[42][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1208),
    .D(_01647_),
    .Q_N(_12452_),
    .Q(\top_ihp.oisc.regs[42][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1243),
    .D(_01648_),
    .Q_N(_12451_),
    .Q(\top_ihp.oisc.regs[42][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1246),
    .D(_01649_),
    .Q_N(_12450_),
    .Q(\top_ihp.oisc.regs[42][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1231),
    .D(_01650_),
    .Q_N(_12449_),
    .Q(\top_ihp.oisc.regs[42][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1195),
    .D(_01651_),
    .Q_N(_12448_),
    .Q(\top_ihp.oisc.regs[42][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1325),
    .D(_01652_),
    .Q_N(_12447_),
    .Q(\top_ihp.oisc.regs[42][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1189),
    .D(_01653_),
    .Q_N(_12446_),
    .Q(\top_ihp.oisc.regs[42][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1195),
    .D(_01654_),
    .Q_N(_12445_),
    .Q(\top_ihp.oisc.regs[42][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1158),
    .D(_01655_),
    .Q_N(_12444_),
    .Q(\top_ihp.oisc.regs[42][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1207),
    .D(_01656_),
    .Q_N(_12443_),
    .Q(\top_ihp.oisc.regs[42][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1183),
    .D(_01657_),
    .Q_N(_12442_),
    .Q(\top_ihp.oisc.regs[42][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1182),
    .D(_01658_),
    .Q_N(_12441_),
    .Q(\top_ihp.oisc.regs[42][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1182),
    .D(_01659_),
    .Q_N(_12440_),
    .Q(\top_ihp.oisc.regs[42][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1250),
    .D(_01660_),
    .Q_N(_12439_),
    .Q(\top_ihp.oisc.regs[42][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1266),
    .D(_01661_),
    .Q_N(_12438_),
    .Q(\top_ihp.oisc.regs[42][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1151),
    .D(_01662_),
    .Q_N(_12437_),
    .Q(\top_ihp.oisc.regs[42][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1213),
    .D(_01663_),
    .Q_N(_12436_),
    .Q(\top_ihp.oisc.regs[42][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1201),
    .D(_01664_),
    .Q_N(_12435_),
    .Q(\top_ihp.oisc.regs[42][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1160),
    .D(_01665_),
    .Q_N(_12434_),
    .Q(\top_ihp.oisc.regs[42][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1159),
    .D(_01666_),
    .Q_N(_12433_),
    .Q(\top_ihp.oisc.regs[42][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[42][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1266),
    .D(_01667_),
    .Q_N(_12432_),
    .Q(\top_ihp.oisc.regs[42][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1284),
    .D(_01668_),
    .Q_N(_12431_),
    .Q(\top_ihp.oisc.regs[43][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1144),
    .D(_01669_),
    .Q_N(_12430_),
    .Q(\top_ihp.oisc.regs[43][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1207),
    .D(_01670_),
    .Q_N(_12429_),
    .Q(\top_ihp.oisc.regs[43][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1219),
    .D(_01671_),
    .Q_N(_12428_),
    .Q(\top_ihp.oisc.regs[43][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1253),
    .D(_01672_),
    .Q_N(_12427_),
    .Q(\top_ihp.oisc.regs[43][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1305),
    .D(_01673_),
    .Q_N(_12426_),
    .Q(\top_ihp.oisc.regs[43][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1261),
    .D(_01674_),
    .Q_N(_12425_),
    .Q(\top_ihp.oisc.regs[43][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1305),
    .D(_01675_),
    .Q_N(_12424_),
    .Q(\top_ihp.oisc.regs[43][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1255),
    .D(_01676_),
    .Q_N(_12423_),
    .Q(\top_ihp.oisc.regs[43][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1259),
    .D(_01677_),
    .Q_N(_12422_),
    .Q(\top_ihp.oisc.regs[43][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1268),
    .D(_01678_),
    .Q_N(_12421_),
    .Q(\top_ihp.oisc.regs[43][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1215),
    .D(_01679_),
    .Q_N(_12420_),
    .Q(\top_ihp.oisc.regs[43][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1245),
    .D(_01680_),
    .Q_N(_12419_),
    .Q(\top_ihp.oisc.regs[43][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1245),
    .D(_01681_),
    .Q_N(_12418_),
    .Q(\top_ihp.oisc.regs[43][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1239),
    .D(_01682_),
    .Q_N(_12417_),
    .Q(\top_ihp.oisc.regs[43][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1194),
    .D(_01683_),
    .Q_N(_12416_),
    .Q(\top_ihp.oisc.regs[43][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1142),
    .D(_01684_),
    .Q_N(_12415_),
    .Q(\top_ihp.oisc.regs[43][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1179),
    .D(_01685_),
    .Q_N(_12414_),
    .Q(\top_ihp.oisc.regs[43][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(_01686_),
    .Q_N(_12413_),
    .Q(\top_ihp.oisc.regs[43][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1288),
    .D(_01687_),
    .Q_N(_12412_),
    .Q(\top_ihp.oisc.regs[43][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1200),
    .D(_01688_),
    .Q_N(_12411_),
    .Q(\top_ihp.oisc.regs[43][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1169),
    .D(_01689_),
    .Q_N(_12410_),
    .Q(\top_ihp.oisc.regs[43][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1168),
    .D(_01690_),
    .Q_N(_12409_),
    .Q(\top_ihp.oisc.regs[43][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1167),
    .D(_01691_),
    .Q_N(_12408_),
    .Q(\top_ihp.oisc.regs[43][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1185),
    .D(_01692_),
    .Q_N(_12407_),
    .Q(\top_ihp.oisc.regs[43][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1267),
    .D(_01693_),
    .Q_N(_12406_),
    .Q(\top_ihp.oisc.regs[43][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1286),
    .D(_01694_),
    .Q_N(_12405_),
    .Q(\top_ihp.oisc.regs[43][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1199),
    .D(_01695_),
    .Q_N(_12404_),
    .Q(\top_ihp.oisc.regs[43][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1268),
    .D(_01696_),
    .Q_N(_12403_),
    .Q(\top_ihp.oisc.regs[43][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1163),
    .D(_01697_),
    .Q_N(_12402_),
    .Q(\top_ihp.oisc.regs[43][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1147),
    .D(_01698_),
    .Q_N(_12401_),
    .Q(\top_ihp.oisc.regs[43][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[43][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1203),
    .D(_01699_),
    .Q_N(_12400_),
    .Q(\top_ihp.oisc.regs[43][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1272),
    .D(_01700_),
    .Q_N(_12399_),
    .Q(\top_ihp.oisc.regs[44][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1140),
    .D(_01701_),
    .Q_N(_12398_),
    .Q(\top_ihp.oisc.regs[44][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1221),
    .D(_01702_),
    .Q_N(_12397_),
    .Q(\top_ihp.oisc.regs[44][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1224),
    .D(_01703_),
    .Q_N(_12396_),
    .Q(\top_ihp.oisc.regs[44][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1253),
    .D(_01704_),
    .Q_N(_12395_),
    .Q(\top_ihp.oisc.regs[44][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1260),
    .D(_01705_),
    .Q_N(_12394_),
    .Q(\top_ihp.oisc.regs[44][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1317),
    .D(_01706_),
    .Q_N(_12393_),
    .Q(\top_ihp.oisc.regs[44][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1309),
    .D(_01707_),
    .Q_N(_12392_),
    .Q(\top_ihp.oisc.regs[44][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1255),
    .D(_01708_),
    .Q_N(_12391_),
    .Q(\top_ihp.oisc.regs[44][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1261),
    .D(_01709_),
    .Q_N(_12390_),
    .Q(\top_ihp.oisc.regs[44][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1280),
    .D(_01710_),
    .Q_N(_12389_),
    .Q(\top_ihp.oisc.regs[44][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1203),
    .D(_01711_),
    .Q_N(_12388_),
    .Q(\top_ihp.oisc.regs[44][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1244),
    .D(_01712_),
    .Q_N(_12387_),
    .Q(\top_ihp.oisc.regs[44][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1245),
    .D(_01713_),
    .Q_N(_12386_),
    .Q(\top_ihp.oisc.regs[44][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1317),
    .D(_01714_),
    .Q_N(_12385_),
    .Q(\top_ihp.oisc.regs[44][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1240),
    .D(_01715_),
    .Q_N(_12384_),
    .Q(\top_ihp.oisc.regs[44][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1142),
    .D(_01716_),
    .Q_N(_12383_),
    .Q(\top_ihp.oisc.regs[44][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1240),
    .D(_01717_),
    .Q_N(_12382_),
    .Q(\top_ihp.oisc.regs[44][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1240),
    .D(_01718_),
    .Q_N(_12381_),
    .Q(\top_ihp.oisc.regs[44][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1218),
    .D(_01719_),
    .Q_N(_12380_),
    .Q(\top_ihp.oisc.regs[44][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1162),
    .D(_01720_),
    .Q_N(_12379_),
    .Q(\top_ihp.oisc.regs[44][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1231),
    .D(_01721_),
    .Q_N(_12378_),
    .Q(\top_ihp.oisc.regs[44][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1169),
    .D(_01722_),
    .Q_N(_12377_),
    .Q(\top_ihp.oisc.regs[44][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1159),
    .D(_01723_),
    .Q_N(_12376_),
    .Q(\top_ihp.oisc.regs[44][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1226),
    .D(_01724_),
    .Q_N(_12375_),
    .Q(\top_ihp.oisc.regs[44][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1270),
    .D(_01725_),
    .Q_N(_12374_),
    .Q(\top_ihp.oisc.regs[44][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1198),
    .D(_01726_),
    .Q_N(_12373_),
    .Q(\top_ihp.oisc.regs[44][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1217),
    .D(_01727_),
    .Q_N(_12372_),
    .Q(\top_ihp.oisc.regs[44][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1212),
    .D(_01728_),
    .Q_N(_12371_),
    .Q(\top_ihp.oisc.regs[44][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1253),
    .D(_01729_),
    .Q_N(_12370_),
    .Q(\top_ihp.oisc.regs[44][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1159),
    .D(_01730_),
    .Q_N(_12369_),
    .Q(\top_ihp.oisc.regs[44][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[44][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1213),
    .D(_01731_),
    .Q_N(_12368_),
    .Q(\top_ihp.oisc.regs[44][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1289),
    .D(_01732_),
    .Q_N(_12367_),
    .Q(\top_ihp.oisc.regs[45][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1140),
    .D(_01733_),
    .Q_N(_12366_),
    .Q(\top_ihp.oisc.regs[45][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1275),
    .D(_01734_),
    .Q_N(_12365_),
    .Q(\top_ihp.oisc.regs[45][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1278),
    .D(_01735_),
    .Q_N(_12364_),
    .Q(\top_ihp.oisc.regs[45][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1250),
    .D(_01736_),
    .Q_N(_12363_),
    .Q(\top_ihp.oisc.regs[45][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1303),
    .D(_01737_),
    .Q_N(_12362_),
    .Q(\top_ihp.oisc.regs[45][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1251),
    .D(_01738_),
    .Q_N(_12361_),
    .Q(\top_ihp.oisc.regs[45][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1303),
    .D(_01739_),
    .Q_N(_12360_),
    .Q(\top_ihp.oisc.regs[45][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1255),
    .D(_01740_),
    .Q_N(_12359_),
    .Q(\top_ihp.oisc.regs[45][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1303),
    .D(_01741_),
    .Q_N(_12358_),
    .Q(\top_ihp.oisc.regs[45][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1272),
    .D(_01742_),
    .Q_N(_12357_),
    .Q(\top_ihp.oisc.regs[45][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1276),
    .D(_01743_),
    .Q_N(_12356_),
    .Q(\top_ihp.oisc.regs[45][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1243),
    .D(_01744_),
    .Q_N(_12355_),
    .Q(\top_ihp.oisc.regs[45][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1236),
    .D(_01745_),
    .Q_N(_12354_),
    .Q(\top_ihp.oisc.regs[45][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_01746_),
    .Q_N(_12353_),
    .Q(\top_ihp.oisc.regs[45][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1180),
    .D(_01747_),
    .Q_N(_12352_),
    .Q(\top_ihp.oisc.regs[45][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1138),
    .D(_01748_),
    .Q_N(_12351_),
    .Q(\top_ihp.oisc.regs[45][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1179),
    .D(_01749_),
    .Q_N(_12350_),
    .Q(\top_ihp.oisc.regs[45][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1190),
    .D(_01750_),
    .Q_N(_12349_),
    .Q(\top_ihp.oisc.regs[45][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1144),
    .D(_01751_),
    .Q_N(_12348_),
    .Q(\top_ihp.oisc.regs[45][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1185),
    .D(_01752_),
    .Q_N(_12347_),
    .Q(\top_ihp.oisc.regs[45][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1178),
    .D(_01753_),
    .Q_N(_12346_),
    .Q(\top_ihp.oisc.regs[45][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1168),
    .D(_01754_),
    .Q_N(_12345_),
    .Q(\top_ihp.oisc.regs[45][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1167),
    .D(_01755_),
    .Q_N(_12344_),
    .Q(\top_ihp.oisc.regs[45][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1188),
    .D(_01756_),
    .Q_N(_12343_),
    .Q(\top_ihp.oisc.regs[45][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1283),
    .D(_01757_),
    .Q_N(_12342_),
    .Q(\top_ihp.oisc.regs[45][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1138),
    .D(_01758_),
    .Q_N(_12341_),
    .Q(\top_ihp.oisc.regs[45][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1267),
    .D(_01759_),
    .Q_N(_12340_),
    .Q(\top_ihp.oisc.regs[45][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1219),
    .D(_01760_),
    .Q_N(_12339_),
    .Q(\top_ihp.oisc.regs[45][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1160),
    .D(_01761_),
    .Q_N(_12338_),
    .Q(\top_ihp.oisc.regs[45][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1149),
    .D(_01762_),
    .Q_N(_12337_),
    .Q(\top_ihp.oisc.regs[45][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[45][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1214),
    .D(_01763_),
    .Q_N(_12336_),
    .Q(\top_ihp.oisc.regs[45][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1279),
    .D(_01764_),
    .Q_N(_12335_),
    .Q(\top_ihp.oisc.regs[46][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1140),
    .D(_01765_),
    .Q_N(_12334_),
    .Q(\top_ihp.oisc.regs[46][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1225),
    .D(_01766_),
    .Q_N(_12333_),
    .Q(\top_ihp.oisc.regs[46][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1275),
    .D(_01767_),
    .Q_N(_12332_),
    .Q(\top_ihp.oisc.regs[46][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1298),
    .D(_01768_),
    .Q_N(_12331_),
    .Q(\top_ihp.oisc.regs[46][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1300),
    .D(_01769_),
    .Q_N(_12330_),
    .Q(\top_ihp.oisc.regs[46][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1309),
    .D(_01770_),
    .Q_N(_12329_),
    .Q(\top_ihp.oisc.regs[46][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1309),
    .D(_01771_),
    .Q_N(_12328_),
    .Q(\top_ihp.oisc.regs[46][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1262),
    .D(_01772_),
    .Q_N(_12327_),
    .Q(\top_ihp.oisc.regs[46][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1307),
    .D(_01773_),
    .Q_N(_12326_),
    .Q(\top_ihp.oisc.regs[46][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1277),
    .D(_01774_),
    .Q_N(_12325_),
    .Q(\top_ihp.oisc.regs[46][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1208),
    .D(_01775_),
    .Q_N(_12324_),
    .Q(\top_ihp.oisc.regs[46][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1256),
    .D(_01776_),
    .Q_N(_12323_),
    .Q(\top_ihp.oisc.regs[46][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1231),
    .D(_01777_),
    .Q_N(_12322_),
    .Q(\top_ihp.oisc.regs[46][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1231),
    .D(_01778_),
    .Q_N(_12321_),
    .Q(\top_ihp.oisc.regs[46][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1174),
    .D(_01779_),
    .Q_N(_12320_),
    .Q(\top_ihp.oisc.regs[46][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1138),
    .D(_01780_),
    .Q_N(_12319_),
    .Q(\top_ihp.oisc.regs[46][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1174),
    .D(_01781_),
    .Q_N(_12318_),
    .Q(\top_ihp.oisc.regs[46][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1195),
    .D(_01782_),
    .Q_N(_12317_),
    .Q(\top_ihp.oisc.regs[46][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1147),
    .D(_01783_),
    .Q_N(_12316_),
    .Q(\top_ihp.oisc.regs[46][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1162),
    .D(_01784_),
    .Q_N(_12315_),
    .Q(\top_ihp.oisc.regs[46][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1186),
    .D(_01785_),
    .Q_N(_12314_),
    .Q(\top_ihp.oisc.regs[46][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1183),
    .D(_01786_),
    .Q_N(_12313_),
    .Q(\top_ihp.oisc.regs[46][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1182),
    .D(_01787_),
    .Q_N(_12312_),
    .Q(\top_ihp.oisc.regs[46][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1250),
    .D(_01788_),
    .Q_N(_12311_),
    .Q(\top_ihp.oisc.regs[46][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1273),
    .D(_01789_),
    .Q_N(_12310_),
    .Q(\top_ihp.oisc.regs[46][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1113),
    .D(_01790_),
    .Q_N(_12309_),
    .Q(\top_ihp.oisc.regs[46][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1213),
    .D(_01791_),
    .Q_N(_12308_),
    .Q(\top_ihp.oisc.regs[46][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1219),
    .D(_01792_),
    .Q_N(_12307_),
    .Q(\top_ihp.oisc.regs[46][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1159),
    .D(_01793_),
    .Q_N(_12306_),
    .Q(\top_ihp.oisc.regs[46][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1159),
    .D(_01794_),
    .Q_N(_12305_),
    .Q(\top_ihp.oisc.regs[46][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[46][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1268),
    .D(_01795_),
    .Q_N(_12304_),
    .Q(\top_ihp.oisc.regs[46][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1279),
    .D(_01796_),
    .Q_N(_12303_),
    .Q(\top_ihp.oisc.regs[47][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1140),
    .D(_01797_),
    .Q_N(_12302_),
    .Q(\top_ihp.oisc.regs[47][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1221),
    .D(_01798_),
    .Q_N(_12301_),
    .Q(\top_ihp.oisc.regs[47][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1279),
    .D(_01799_),
    .Q_N(_12300_),
    .Q(\top_ihp.oisc.regs[47][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1248),
    .D(_01800_),
    .Q_N(_12299_),
    .Q(\top_ihp.oisc.regs[47][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1307),
    .D(_01801_),
    .Q_N(_12298_),
    .Q(\top_ihp.oisc.regs[47][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1298),
    .D(_01802_),
    .Q_N(_12297_),
    .Q(\top_ihp.oisc.regs[47][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1309),
    .D(_01803_),
    .Q_N(_12296_),
    .Q(\top_ihp.oisc.regs[47][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1248),
    .D(_01804_),
    .Q_N(_12295_),
    .Q(\top_ihp.oisc.regs[47][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1309),
    .D(_01805_),
    .Q_N(_12294_),
    .Q(\top_ihp.oisc.regs[47][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1273),
    .D(_01806_),
    .Q_N(_12293_),
    .Q(\top_ihp.oisc.regs[47][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1222),
    .D(_01807_),
    .Q_N(_12292_),
    .Q(\top_ihp.oisc.regs[47][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1256),
    .D(_01808_),
    .Q_N(_12291_),
    .Q(\top_ihp.oisc.regs[47][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_100_clk),
    .RESET_B(net1248),
    .D(_01809_),
    .Q_N(_12290_),
    .Q(\top_ihp.oisc.regs[47][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1190),
    .D(_01810_),
    .Q_N(_12289_),
    .Q(\top_ihp.oisc.regs[47][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1256),
    .D(_01811_),
    .Q_N(_12288_),
    .Q(\top_ihp.oisc.regs[47][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1142),
    .D(_01812_),
    .Q_N(_12287_),
    .Q(\top_ihp.oisc.regs[47][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_73_clk),
    .RESET_B(net1190),
    .D(_01813_),
    .Q_N(_12286_),
    .Q(\top_ihp.oisc.regs[47][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1179),
    .D(_01814_),
    .Q_N(_12285_),
    .Q(\top_ihp.oisc.regs[47][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1148),
    .D(_01815_),
    .Q_N(_12284_),
    .Q(\top_ihp.oisc.regs[47][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1163),
    .D(_01816_),
    .Q_N(_12283_),
    .Q(\top_ihp.oisc.regs[47][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1189),
    .D(_01817_),
    .Q_N(_12282_),
    .Q(\top_ihp.oisc.regs[47][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1169),
    .D(_01818_),
    .Q_N(_12281_),
    .Q(\top_ihp.oisc.regs[47][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1182),
    .D(_01819_),
    .Q_N(_12280_),
    .Q(\top_ihp.oisc.regs[47][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1222),
    .D(_01820_),
    .Q_N(_12279_),
    .Q(\top_ihp.oisc.regs[47][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1270),
    .D(_01821_),
    .Q_N(_12278_),
    .Q(\top_ihp.oisc.regs[47][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1155),
    .D(_01822_),
    .Q_N(_12277_),
    .Q(\top_ihp.oisc.regs[47][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1267),
    .D(_01823_),
    .Q_N(_12276_),
    .Q(\top_ihp.oisc.regs[47][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1213),
    .D(_01824_),
    .Q_N(_12275_),
    .Q(\top_ihp.oisc.regs[47][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1149),
    .D(_01825_),
    .Q_N(_12274_),
    .Q(\top_ihp.oisc.regs[47][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1149),
    .D(_01826_),
    .Q_N(_12273_),
    .Q(\top_ihp.oisc.regs[47][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[47][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1212),
    .D(_01827_),
    .Q_N(_12272_),
    .Q(\top_ihp.oisc.regs[47][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1290),
    .D(_01828_),
    .Q_N(_12271_),
    .Q(\top_ihp.oisc.regs[48][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_01829_),
    .Q_N(_12270_),
    .Q(\top_ihp.oisc.regs[48][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1275),
    .D(_01830_),
    .Q_N(_12269_),
    .Q(\top_ihp.oisc.regs[48][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1224),
    .D(_01831_),
    .Q_N(_12268_),
    .Q(\top_ihp.oisc.regs[48][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1248),
    .D(_01832_),
    .Q_N(_12267_),
    .Q(\top_ihp.oisc.regs[48][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1296),
    .D(_01833_),
    .Q_N(_12266_),
    .Q(\top_ihp.oisc.regs[48][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1298),
    .D(_01834_),
    .Q_N(_12265_),
    .Q(\top_ihp.oisc.regs[48][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1307),
    .D(_01835_),
    .Q_N(_12264_),
    .Q(\top_ihp.oisc.regs[48][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1258),
    .D(_01836_),
    .Q_N(_12263_),
    .Q(\top_ihp.oisc.regs[48][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1260),
    .D(_01837_),
    .Q_N(_12262_),
    .Q(\top_ihp.oisc.regs[48][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1273),
    .D(_01838_),
    .Q_N(_12261_),
    .Q(\top_ihp.oisc.regs[48][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1222),
    .D(_01839_),
    .Q_N(_12260_),
    .Q(\top_ihp.oisc.regs[48][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1255),
    .D(_01840_),
    .Q_N(_12259_),
    .Q(\top_ihp.oisc.regs[48][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1246),
    .D(_01841_),
    .Q_N(_12258_),
    .Q(\top_ihp.oisc.regs[48][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1186),
    .D(_01842_),
    .Q_N(_12257_),
    .Q(\top_ihp.oisc.regs[48][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1178),
    .D(_01843_),
    .Q_N(_12256_),
    .Q(\top_ihp.oisc.regs[48][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1139),
    .D(_01844_),
    .Q_N(_12255_),
    .Q(\top_ihp.oisc.regs[48][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1177),
    .D(_01845_),
    .Q_N(_12254_),
    .Q(\top_ihp.oisc.regs[48][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1177),
    .D(_01846_),
    .Q_N(_12253_),
    .Q(\top_ihp.oisc.regs[48][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1288),
    .D(_01847_),
    .Q_N(_12252_),
    .Q(\top_ihp.oisc.regs[48][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1236),
    .D(_01848_),
    .Q_N(_12251_),
    .Q(\top_ihp.oisc.regs[48][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1178),
    .D(_01849_),
    .Q_N(_12250_),
    .Q(\top_ihp.oisc.regs[48][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1168),
    .D(_01850_),
    .Q_N(_12249_),
    .Q(\top_ihp.oisc.regs[48][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1301),
    .D(_01851_),
    .Q_N(_12248_),
    .Q(\top_ihp.oisc.regs[48][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1298),
    .D(_01852_),
    .Q_N(_12247_),
    .Q(\top_ihp.oisc.regs[48][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1288),
    .D(_01853_),
    .Q_N(_12246_),
    .Q(\top_ihp.oisc.regs[48][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1270),
    .D(_01854_),
    .Q_N(_12245_),
    .Q(\top_ihp.oisc.regs[48][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1217),
    .D(_01855_),
    .Q_N(_12244_),
    .Q(\top_ihp.oisc.regs[48][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1213),
    .D(_01856_),
    .Q_N(_12243_),
    .Q(\top_ihp.oisc.regs[48][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1280),
    .D(_01857_),
    .Q_N(_12242_),
    .Q(\top_ihp.oisc.regs[48][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1163),
    .D(_01858_),
    .Q_N(_12241_),
    .Q(\top_ihp.oisc.regs[48][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[48][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1266),
    .D(_01859_),
    .Q_N(_12240_),
    .Q(\top_ihp.oisc.regs[48][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1284),
    .D(_01860_),
    .Q_N(_12239_),
    .Q(\top_ihp.oisc.regs[49][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1153),
    .D(_01861_),
    .Q_N(_12238_),
    .Q(\top_ihp.oisc.regs[49][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1221),
    .D(_01862_),
    .Q_N(_12237_),
    .Q(\top_ihp.oisc.regs[49][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1275),
    .D(_01863_),
    .Q_N(_12236_),
    .Q(\top_ihp.oisc.regs[49][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1300),
    .D(_01864_),
    .Q_N(_12235_),
    .Q(\top_ihp.oisc.regs[49][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1299),
    .D(_01865_),
    .Q_N(_12234_),
    .Q(\top_ihp.oisc.regs[49][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1277),
    .D(_01866_),
    .Q_N(_12233_),
    .Q(\top_ihp.oisc.regs[49][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1307),
    .D(_01867_),
    .Q_N(_12232_),
    .Q(\top_ihp.oisc.regs[49][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1304),
    .D(_01868_),
    .Q_N(_12231_),
    .Q(\top_ihp.oisc.regs[49][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1261),
    .D(_01869_),
    .Q_N(_12230_),
    .Q(\top_ihp.oisc.regs[49][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1277),
    .D(_01870_),
    .Q_N(_12229_),
    .Q(\top_ihp.oisc.regs[49][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1208),
    .D(_01871_),
    .Q_N(_12228_),
    .Q(\top_ihp.oisc.regs[49][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1244),
    .D(_01872_),
    .Q_N(_12227_),
    .Q(\top_ihp.oisc.regs[49][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1239),
    .D(_01873_),
    .Q_N(_12226_),
    .Q(\top_ihp.oisc.regs[49][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1242),
    .D(_01874_),
    .Q_N(_12225_),
    .Q(\top_ihp.oisc.regs[49][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1239),
    .D(_01875_),
    .Q_N(_12224_),
    .Q(\top_ihp.oisc.regs[49][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1152),
    .D(_01876_),
    .Q_N(_12223_),
    .Q(\top_ihp.oisc.regs[49][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1240),
    .D(_01877_),
    .Q_N(_12222_),
    .Q(\top_ihp.oisc.regs[49][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1189),
    .D(_01878_),
    .Q_N(_12221_),
    .Q(\top_ihp.oisc.regs[49][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1284),
    .D(_01879_),
    .Q_N(_12220_),
    .Q(\top_ihp.oisc.regs[49][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1207),
    .D(_01880_),
    .Q_N(_12219_),
    .Q(\top_ihp.oisc.regs[49][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1183),
    .D(_01881_),
    .Q_N(_12218_),
    .Q(\top_ihp.oisc.regs[49][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1296),
    .D(_01882_),
    .Q_N(_12217_),
    .Q(\top_ihp.oisc.regs[49][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1184),
    .D(_01883_),
    .Q_N(_12216_),
    .Q(\top_ihp.oisc.regs[49][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1230),
    .D(_01884_),
    .Q_N(_12215_),
    .Q(\top_ihp.oisc.regs[49][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1283),
    .D(_01885_),
    .Q_N(_12214_),
    .Q(\top_ihp.oisc.regs[49][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1285),
    .D(_01886_),
    .Q_N(_12213_),
    .Q(\top_ihp.oisc.regs[49][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1286),
    .D(_01887_),
    .Q_N(_12212_),
    .Q(\top_ihp.oisc.regs[49][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1218),
    .D(_01888_),
    .Q_N(_12211_),
    .Q(\top_ihp.oisc.regs[49][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1160),
    .D(_01889_),
    .Q_N(_12210_),
    .Q(\top_ihp.oisc.regs[49][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1211),
    .D(_01890_),
    .Q_N(_12209_),
    .Q(\top_ihp.oisc.regs[49][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[49][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1217),
    .D(_01891_),
    .Q_N(_12208_),
    .Q(\top_ihp.oisc.regs[49][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1326),
    .D(_01892_),
    .Q_N(_12207_),
    .Q(\top_ihp.oisc.regs[4][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1326),
    .D(_01893_),
    .Q_N(_12206_),
    .Q(\top_ihp.oisc.regs[4][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1332),
    .D(_01894_),
    .Q_N(_12205_),
    .Q(\top_ihp.oisc.regs[4][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1332),
    .D(_01895_),
    .Q_N(_12204_),
    .Q(\top_ihp.oisc.regs[4][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1351),
    .D(_01896_),
    .Q_N(_12203_),
    .Q(\top_ihp.oisc.regs[4][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1358),
    .D(_01897_),
    .Q_N(_12202_),
    .Q(\top_ihp.oisc.regs[4][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1358),
    .D(_01898_),
    .Q_N(_12201_),
    .Q(\top_ihp.oisc.regs[4][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1351),
    .D(_01899_),
    .Q_N(_12200_),
    .Q(\top_ihp.oisc.regs[4][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1351),
    .D(_01900_),
    .Q_N(_12199_),
    .Q(\top_ihp.oisc.regs[4][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1358),
    .D(_01901_),
    .Q_N(_12198_),
    .Q(\top_ihp.oisc.regs[4][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1332),
    .D(_01902_),
    .Q_N(_12197_),
    .Q(\top_ihp.oisc.regs[4][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1333),
    .D(_01903_),
    .Q_N(_12196_),
    .Q(\top_ihp.oisc.regs[4][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1358),
    .D(_01904_),
    .Q_N(_12195_),
    .Q(\top_ihp.oisc.regs[4][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1358),
    .D(_01905_),
    .Q_N(_12194_),
    .Q(\top_ihp.oisc.regs[4][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1359),
    .D(_01906_),
    .Q_N(_12193_),
    .Q(\top_ihp.oisc.regs[4][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1359),
    .D(_01907_),
    .Q_N(_12192_),
    .Q(\top_ihp.oisc.regs[4][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1325),
    .D(_01908_),
    .Q_N(_12191_),
    .Q(\top_ihp.oisc.regs[4][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_140_clk),
    .RESET_B(net1359),
    .D(_01909_),
    .Q_N(_12190_),
    .Q(\top_ihp.oisc.regs[4][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_120_clk),
    .RESET_B(net1358),
    .D(_01910_),
    .Q_N(_12189_),
    .Q(\top_ihp.oisc.regs[4][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1332),
    .D(_01911_),
    .Q_N(_12188_),
    .Q(\top_ihp.oisc.regs[4][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_204_clk),
    .RESET_B(net1333),
    .D(_01912_),
    .Q_N(_12187_),
    .Q(\top_ihp.oisc.regs[4][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_117_clk),
    .RESET_B(net1351),
    .D(_01913_),
    .Q_N(_12186_),
    .Q(\top_ihp.oisc.regs[4][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1351),
    .D(_01914_),
    .Q_N(_12185_),
    .Q(\top_ihp.oisc.regs[4][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1352),
    .D(_01915_),
    .Q_N(_12184_),
    .Q(\top_ihp.oisc.regs[4][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1352),
    .D(_01916_),
    .Q_N(_12183_),
    .Q(\top_ihp.oisc.regs[4][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1327),
    .D(_01917_),
    .Q_N(_12182_),
    .Q(\top_ihp.oisc.regs[4][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1328),
    .D(_01918_),
    .Q_N(_12181_),
    .Q(\top_ihp.oisc.regs[4][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1327),
    .D(_01919_),
    .Q_N(_12180_),
    .Q(\top_ihp.oisc.regs[4][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1329),
    .D(_01920_),
    .Q_N(_12179_),
    .Q(\top_ihp.oisc.regs[4][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1352),
    .D(_01921_),
    .Q_N(_12178_),
    .Q(\top_ihp.oisc.regs[4][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_201_clk),
    .RESET_B(net1334),
    .D(_01922_),
    .Q_N(_12177_),
    .Q(\top_ihp.oisc.regs[4][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[4][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1329),
    .D(_01923_),
    .Q_N(_12176_),
    .Q(\top_ihp.oisc.regs[4][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1289),
    .D(_01924_),
    .Q_N(_12175_),
    .Q(\top_ihp.oisc.regs[50][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1145),
    .D(_01925_),
    .Q_N(_12174_),
    .Q(\top_ihp.oisc.regs[50][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1214),
    .D(_01926_),
    .Q_N(_12173_),
    .Q(\top_ihp.oisc.regs[50][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1279),
    .D(_01927_),
    .Q_N(_12172_),
    .Q(\top_ihp.oisc.regs[50][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1312),
    .D(_01928_),
    .Q_N(_12171_),
    .Q(\top_ihp.oisc.regs[50][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1303),
    .D(_01929_),
    .Q_N(_12170_),
    .Q(\top_ihp.oisc.regs[50][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1251),
    .D(_01930_),
    .Q_N(_12169_),
    .Q(\top_ihp.oisc.regs[50][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1316),
    .D(_01931_),
    .Q_N(_12168_),
    .Q(\top_ihp.oisc.regs[50][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1258),
    .D(_01932_),
    .Q_N(_12167_),
    .Q(\top_ihp.oisc.regs[50][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1308),
    .D(_01933_),
    .Q_N(_12166_),
    .Q(\top_ihp.oisc.regs[50][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1313),
    .D(_01934_),
    .Q_N(_12165_),
    .Q(\top_ihp.oisc.regs[50][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1204),
    .D(_01935_),
    .Q_N(_12164_),
    .Q(\top_ihp.oisc.regs[50][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1246),
    .D(_01936_),
    .Q_N(_12163_),
    .Q(\top_ihp.oisc.regs[50][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1316),
    .D(_01937_),
    .Q_N(_12162_),
    .Q(\top_ihp.oisc.regs[50][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_01938_),
    .Q_N(_12161_),
    .Q(\top_ihp.oisc.regs[50][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1318),
    .D(_01939_),
    .Q_N(_12160_),
    .Q(\top_ihp.oisc.regs[50][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1143),
    .D(_01940_),
    .Q_N(_12159_),
    .Q(\top_ihp.oisc.regs[50][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1148),
    .D(_01941_),
    .Q_N(_12158_),
    .Q(\top_ihp.oisc.regs[50][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1192),
    .D(_01942_),
    .Q_N(_12157_),
    .Q(\top_ihp.oisc.regs[50][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1158),
    .D(_01943_),
    .Q_N(_12156_),
    .Q(\top_ihp.oisc.regs[50][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1162),
    .D(_01944_),
    .Q_N(_12155_),
    .Q(\top_ihp.oisc.regs[50][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_95_clk),
    .RESET_B(net1183),
    .D(_01945_),
    .Q_N(_12154_),
    .Q(\top_ihp.oisc.regs[50][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_01946_),
    .Q_N(_12153_),
    .Q(\top_ihp.oisc.regs[50][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1182),
    .D(_01947_),
    .Q_N(_12152_),
    .Q(\top_ihp.oisc.regs[50][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1234),
    .D(_01948_),
    .Q_N(_12151_),
    .Q(\top_ihp.oisc.regs[50][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1271),
    .D(_01949_),
    .Q_N(_12150_),
    .Q(\top_ihp.oisc.regs[50][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1143),
    .D(_01950_),
    .Q_N(_12149_),
    .Q(\top_ihp.oisc.regs[50][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1198),
    .D(_01951_),
    .Q_N(_12148_),
    .Q(\top_ihp.oisc.regs[50][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1201),
    .D(_01952_),
    .Q_N(_12147_),
    .Q(\top_ihp.oisc.regs[50][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1222),
    .D(_01953_),
    .Q_N(_12146_),
    .Q(\top_ihp.oisc.regs[50][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1209),
    .D(_01954_),
    .Q_N(_12145_),
    .Q(\top_ihp.oisc.regs[50][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[50][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1220),
    .D(_01955_),
    .Q_N(_12144_),
    .Q(\top_ihp.oisc.regs[50][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1281),
    .D(_01956_),
    .Q_N(_12143_),
    .Q(\top_ihp.oisc.regs[51][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1153),
    .D(_01957_),
    .Q_N(_12142_),
    .Q(\top_ihp.oisc.regs[51][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1214),
    .D(_01958_),
    .Q_N(_12141_),
    .Q(\top_ihp.oisc.regs[51][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_280_clk),
    .RESET_B(net1279),
    .D(_01959_),
    .Q_N(_12140_),
    .Q(\top_ihp.oisc.regs[51][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1312),
    .D(_01960_),
    .Q_N(_12139_),
    .Q(\top_ihp.oisc.regs[51][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1300),
    .D(_01961_),
    .Q_N(_12138_),
    .Q(\top_ihp.oisc.regs[51][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_199_clk),
    .RESET_B(net1280),
    .D(_01962_),
    .Q_N(_12137_),
    .Q(\top_ihp.oisc.regs[51][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1317),
    .D(_01963_),
    .Q_N(_12136_),
    .Q(\top_ihp.oisc.regs[51][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1259),
    .D(_01964_),
    .Q_N(_12135_),
    .Q(\top_ihp.oisc.regs[51][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1261),
    .D(_01965_),
    .Q_N(_12134_),
    .Q(\top_ihp.oisc.regs[51][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1269),
    .D(_01966_),
    .Q_N(_12133_),
    .Q(\top_ihp.oisc.regs[51][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1208),
    .D(_01967_),
    .Q_N(_12132_),
    .Q(\top_ihp.oisc.regs[51][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1241),
    .D(_01968_),
    .Q_N(_12131_),
    .Q(\top_ihp.oisc.regs[51][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1237),
    .D(_01969_),
    .Q_N(_12130_),
    .Q(\top_ihp.oisc.regs[51][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1191),
    .D(_01970_),
    .Q_N(_12129_),
    .Q(\top_ihp.oisc.regs[51][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1318),
    .D(_01971_),
    .Q_N(_12128_),
    .Q(\top_ihp.oisc.regs[51][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1153),
    .D(_01972_),
    .Q_N(_12127_),
    .Q(\top_ihp.oisc.regs[51][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1239),
    .D(_01973_),
    .Q_N(_12126_),
    .Q(\top_ihp.oisc.regs[51][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1190),
    .D(_01974_),
    .Q_N(_12125_),
    .Q(\top_ihp.oisc.regs[51][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1158),
    .D(_01975_),
    .Q_N(_12124_),
    .Q(\top_ihp.oisc.regs[51][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1162),
    .D(_01976_),
    .Q_N(_12123_),
    .Q(\top_ihp.oisc.regs[51][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1312),
    .D(_01977_),
    .Q_N(_12122_),
    .Q(\top_ihp.oisc.regs[51][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_97_clk),
    .RESET_B(net1183),
    .D(_01978_),
    .Q_N(_12121_),
    .Q(\top_ihp.oisc.regs[51][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1182),
    .D(_01979_),
    .Q_N(_12120_),
    .Q(\top_ihp.oisc.regs[51][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1231),
    .D(_01980_),
    .Q_N(_12119_),
    .Q(\top_ihp.oisc.regs[51][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1271),
    .D(_01981_),
    .Q_N(_12118_),
    .Q(\top_ihp.oisc.regs[51][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1155),
    .D(_01982_),
    .Q_N(_12117_),
    .Q(\top_ihp.oisc.regs[51][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1213),
    .D(_01983_),
    .Q_N(_12116_),
    .Q(\top_ihp.oisc.regs[51][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1212),
    .D(_01984_),
    .Q_N(_12115_),
    .Q(\top_ihp.oisc.regs[51][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1159),
    .D(_01985_),
    .Q_N(_12114_),
    .Q(\top_ihp.oisc.regs[51][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1207),
    .D(_01986_),
    .Q_N(_12113_),
    .Q(\top_ihp.oisc.regs[51][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[51][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1272),
    .D(_01987_),
    .Q_N(_12112_),
    .Q(\top_ihp.oisc.regs[51][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1289),
    .D(_01988_),
    .Q_N(_12111_),
    .Q(\top_ihp.oisc.regs[52][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1154),
    .D(_01989_),
    .Q_N(_12110_),
    .Q(\top_ihp.oisc.regs[52][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1210),
    .D(_01990_),
    .Q_N(_12109_),
    .Q(\top_ihp.oisc.regs[52][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1224),
    .D(_01991_),
    .Q_N(_12108_),
    .Q(\top_ihp.oisc.regs[52][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1248),
    .D(_01992_),
    .Q_N(_12107_),
    .Q(\top_ihp.oisc.regs[52][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1318),
    .D(_01993_),
    .Q_N(_12106_),
    .Q(\top_ihp.oisc.regs[52][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1297),
    .D(_01994_),
    .Q_N(_12105_),
    .Q(\top_ihp.oisc.regs[52][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1318),
    .D(_01995_),
    .Q_N(_12104_),
    .Q(\top_ihp.oisc.regs[52][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1321),
    .D(_01996_),
    .Q_N(_12103_),
    .Q(\top_ihp.oisc.regs[52][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1306),
    .D(_01997_),
    .Q_N(_12102_),
    .Q(\top_ihp.oisc.regs[52][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1280),
    .D(_01998_),
    .Q_N(_12101_),
    .Q(\top_ihp.oisc.regs[52][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1210),
    .D(_01999_),
    .Q_N(_12100_),
    .Q(\top_ihp.oisc.regs[52][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_86_clk),
    .RESET_B(net1255),
    .D(_02000_),
    .Q_N(_12099_),
    .Q(\top_ihp.oisc.regs[52][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1243),
    .D(_02001_),
    .Q_N(_12098_),
    .Q(\top_ihp.oisc.regs[52][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1189),
    .D(_02002_),
    .Q_N(_12097_),
    .Q(\top_ihp.oisc.regs[52][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1195),
    .D(_02003_),
    .Q_N(_12096_),
    .Q(\top_ihp.oisc.regs[52][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1143),
    .D(_02004_),
    .Q_N(_12095_),
    .Q(\top_ihp.oisc.regs[52][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1239),
    .D(_02005_),
    .Q_N(_12094_),
    .Q(\top_ihp.oisc.regs[52][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1195),
    .D(_02006_),
    .Q_N(_12093_),
    .Q(\top_ihp.oisc.regs[52][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1145),
    .D(_02007_),
    .Q_N(_12092_),
    .Q(\top_ihp.oisc.regs[52][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1185),
    .D(_02008_),
    .Q_N(_12091_),
    .Q(\top_ihp.oisc.regs[52][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1192),
    .D(_02009_),
    .Q_N(_12090_),
    .Q(\top_ihp.oisc.regs[52][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1183),
    .D(_02010_),
    .Q_N(_12089_),
    .Q(\top_ihp.oisc.regs[52][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1234),
    .D(_02011_),
    .Q_N(_12088_),
    .Q(\top_ihp.oisc.regs[52][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1229),
    .D(_02012_),
    .Q_N(_12087_),
    .Q(\top_ihp.oisc.regs[52][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_262_clk),
    .RESET_B(net1283),
    .D(_02013_),
    .Q_N(_12086_),
    .Q(\top_ihp.oisc.regs[52][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_313_clk),
    .RESET_B(net1151),
    .D(_02014_),
    .Q_N(_12085_),
    .Q(\top_ihp.oisc.regs[52][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1199),
    .D(_02015_),
    .Q_N(_12084_),
    .Q(\top_ihp.oisc.regs[52][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1204),
    .D(_02016_),
    .Q_N(_12083_),
    .Q(\top_ihp.oisc.regs[52][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1160),
    .D(_02017_),
    .Q_N(_12082_),
    .Q(\top_ihp.oisc.regs[52][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1209),
    .D(_02018_),
    .Q_N(_12081_),
    .Q(\top_ihp.oisc.regs[52][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[52][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_268_clk),
    .RESET_B(net1268),
    .D(_02019_),
    .Q_N(_12080_),
    .Q(\top_ihp.oisc.regs[52][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1284),
    .D(_02020_),
    .Q_N(_12079_),
    .Q(\top_ihp.oisc.regs[53][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_02021_),
    .Q_N(_12078_),
    .Q(\top_ihp.oisc.regs[53][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1214),
    .D(_02022_),
    .Q_N(_12077_),
    .Q(\top_ihp.oisc.regs[53][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1218),
    .D(_02023_),
    .Q_N(_12076_),
    .Q(\top_ihp.oisc.regs[53][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1295),
    .D(_02024_),
    .Q_N(_12075_),
    .Q(\top_ihp.oisc.regs[53][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1303),
    .D(_02025_),
    .Q_N(_12074_),
    .Q(\top_ihp.oisc.regs[53][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_112_clk),
    .RESET_B(net1295),
    .D(_02026_),
    .Q_N(_12073_),
    .Q(\top_ihp.oisc.regs[53][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1303),
    .D(_02027_),
    .Q_N(_12072_),
    .Q(\top_ihp.oisc.regs[53][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1249),
    .D(_02028_),
    .Q_N(_12071_),
    .Q(\top_ihp.oisc.regs[53][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1260),
    .D(_02029_),
    .Q_N(_12070_),
    .Q(\top_ihp.oisc.regs[53][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1268),
    .D(_02030_),
    .Q_N(_12069_),
    .Q(\top_ihp.oisc.regs[53][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1287),
    .D(_02031_),
    .Q_N(_12068_),
    .Q(\top_ihp.oisc.regs[53][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_91_clk),
    .RESET_B(net1242),
    .D(_02032_),
    .Q_N(_12067_),
    .Q(\top_ihp.oisc.regs[53][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1236),
    .D(_02033_),
    .Q_N(_12066_),
    .Q(\top_ihp.oisc.regs[53][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_90_clk),
    .RESET_B(net1239),
    .D(_02034_),
    .Q_N(_12065_),
    .Q(\top_ihp.oisc.regs[53][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_92_clk),
    .RESET_B(net1195),
    .D(_02035_),
    .Q_N(_12064_),
    .Q(\top_ihp.oisc.regs[53][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1143),
    .D(_02036_),
    .Q_N(_12063_),
    .Q(\top_ihp.oisc.regs[53][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1189),
    .D(_02037_),
    .Q_N(_12062_),
    .Q(\top_ihp.oisc.regs[53][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_87_clk),
    .RESET_B(net1260),
    .D(_02038_),
    .Q_N(_12061_),
    .Q(\top_ihp.oisc.regs[53][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1144),
    .D(_02039_),
    .Q_N(_12060_),
    .Q(\top_ihp.oisc.regs[53][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1156),
    .D(_02040_),
    .Q_N(_12059_),
    .Q(\top_ihp.oisc.regs[53][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1183),
    .D(_02041_),
    .Q_N(_12058_),
    .Q(\top_ihp.oisc.regs[53][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1184),
    .D(_02042_),
    .Q_N(_12057_),
    .Q(\top_ihp.oisc.regs[53][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1184),
    .D(_02043_),
    .Q_N(_12056_),
    .Q(\top_ihp.oisc.regs[53][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1229),
    .D(_02044_),
    .Q_N(_12055_),
    .Q(\top_ihp.oisc.regs[53][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1271),
    .D(_02045_),
    .Q_N(_12054_),
    .Q(\top_ihp.oisc.regs[53][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1286),
    .D(_02046_),
    .Q_N(_12053_),
    .Q(\top_ihp.oisc.regs[53][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1286),
    .D(_02047_),
    .Q_N(_12052_),
    .Q(\top_ihp.oisc.regs[53][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1203),
    .D(_02048_),
    .Q_N(_12051_),
    .Q(\top_ihp.oisc.regs[53][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1159),
    .D(_02049_),
    .Q_N(_12050_),
    .Q(\top_ihp.oisc.regs[53][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1206),
    .D(_02050_),
    .Q_N(_12049_),
    .Q(\top_ihp.oisc.regs[53][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[53][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1201),
    .D(_02051_),
    .Q_N(_12048_),
    .Q(\top_ihp.oisc.regs[53][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1279),
    .D(_02052_),
    .Q_N(_12047_),
    .Q(\top_ihp.oisc.regs[54][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1139),
    .D(_02053_),
    .Q_N(_12046_),
    .Q(\top_ihp.oisc.regs[54][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1221),
    .D(_02054_),
    .Q_N(_12045_),
    .Q(\top_ihp.oisc.regs[54][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1219),
    .D(_02055_),
    .Q_N(_12044_),
    .Q(\top_ihp.oisc.regs[54][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1252),
    .D(_02056_),
    .Q_N(_12043_),
    .Q(\top_ihp.oisc.regs[54][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1317),
    .D(_02057_),
    .Q_N(_12042_),
    .Q(\top_ihp.oisc.regs[54][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1261),
    .D(_02058_),
    .Q_N(_12041_),
    .Q(\top_ihp.oisc.regs[54][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1309),
    .D(_02059_),
    .Q_N(_12040_),
    .Q(\top_ihp.oisc.regs[54][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1321),
    .D(_02060_),
    .Q_N(_12039_),
    .Q(\top_ihp.oisc.regs[54][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1310),
    .D(_02061_),
    .Q_N(_12038_),
    .Q(\top_ihp.oisc.regs[54][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_107_clk),
    .RESET_B(net1301),
    .D(_02062_),
    .Q_N(_12037_),
    .Q(\top_ihp.oisc.regs[54][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1278),
    .D(_02063_),
    .Q_N(_12036_),
    .Q(\top_ihp.oisc.regs[54][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1257),
    .D(_02064_),
    .Q_N(_12035_),
    .Q(\top_ihp.oisc.regs[54][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1321),
    .D(_02065_),
    .Q_N(_12034_),
    .Q(\top_ihp.oisc.regs[54][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1179),
    .D(_02066_),
    .Q_N(_12033_),
    .Q(\top_ihp.oisc.regs[54][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1180),
    .D(_02067_),
    .Q_N(_12032_),
    .Q(\top_ihp.oisc.regs[54][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1138),
    .D(_02068_),
    .Q_N(_12031_),
    .Q(\top_ihp.oisc.regs[54][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1163),
    .D(_02069_),
    .Q_N(_12030_),
    .Q(\top_ihp.oisc.regs[54][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1177),
    .D(_02070_),
    .Q_N(_12029_),
    .Q(\top_ihp.oisc.regs[54][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1148),
    .D(_02071_),
    .Q_N(_12028_),
    .Q(\top_ihp.oisc.regs[54][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_269_clk),
    .RESET_B(net1269),
    .D(_02072_),
    .Q_N(_12027_),
    .Q(\top_ihp.oisc.regs[54][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1178),
    .D(_02073_),
    .Q_N(_12026_),
    .Q(\top_ihp.oisc.regs[54][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1169),
    .D(_02074_),
    .Q_N(_12025_),
    .Q(\top_ihp.oisc.regs[54][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1250),
    .D(_02075_),
    .Q_N(_12024_),
    .Q(\top_ihp.oisc.regs[54][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1250),
    .D(_02076_),
    .Q_N(_12023_),
    .Q(\top_ihp.oisc.regs[54][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1266),
    .D(_02077_),
    .Q_N(_12022_),
    .Q(\top_ihp.oisc.regs[54][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1139),
    .D(_02078_),
    .Q_N(_12021_),
    .Q(\top_ihp.oisc.regs[54][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1198),
    .D(_02079_),
    .Q_N(_12020_),
    .Q(\top_ihp.oisc.regs[54][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1217),
    .D(_02080_),
    .Q_N(_12019_),
    .Q(\top_ihp.oisc.regs[54][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net1149),
    .D(_02081_),
    .Q_N(_12018_),
    .Q(\top_ihp.oisc.regs[54][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1209),
    .D(_02082_),
    .Q_N(_12017_),
    .Q(\top_ihp.oisc.regs[54][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[54][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1202),
    .D(_02083_),
    .Q_N(_12016_),
    .Q(\top_ihp.oisc.regs[54][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1281),
    .D(_02084_),
    .Q_N(_12015_),
    .Q(\top_ihp.oisc.regs[55][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_318_clk),
    .RESET_B(net1157),
    .D(_02085_),
    .Q_N(_12014_),
    .Q(\top_ihp.oisc.regs[55][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_281_clk),
    .RESET_B(net1275),
    .D(_02086_),
    .Q_N(_12013_),
    .Q(\top_ihp.oisc.regs[55][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1290),
    .D(_02087_),
    .Q_N(_12012_),
    .Q(\top_ihp.oisc.regs[55][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1249),
    .D(_02088_),
    .Q_N(_12011_),
    .Q(\top_ihp.oisc.regs[55][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1319),
    .D(_02089_),
    .Q_N(_12010_),
    .Q(\top_ihp.oisc.regs[55][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1251),
    .D(_02090_),
    .Q_N(_12009_),
    .Q(\top_ihp.oisc.regs[55][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1319),
    .D(_02091_),
    .Q_N(_12008_),
    .Q(\top_ihp.oisc.regs[55][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1262),
    .D(_02092_),
    .Q_N(_12007_),
    .Q(\top_ihp.oisc.regs[55][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1309),
    .D(_02093_),
    .Q_N(_12006_),
    .Q(\top_ihp.oisc.regs[55][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1281),
    .D(_02094_),
    .Q_N(_12005_),
    .Q(\top_ihp.oisc.regs[55][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1208),
    .D(_02095_),
    .Q_N(_12004_),
    .Q(\top_ihp.oisc.regs[55][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1245),
    .D(_02096_),
    .Q_N(_12003_),
    .Q(\top_ihp.oisc.regs[55][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1245),
    .D(_02097_),
    .Q_N(_12002_),
    .Q(\top_ihp.oisc.regs[55][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1180),
    .D(_02098_),
    .Q_N(_12001_),
    .Q(\top_ihp.oisc.regs[55][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1174),
    .D(_02099_),
    .Q_N(_12000_),
    .Q(\top_ihp.oisc.regs[55][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1113),
    .D(_02100_),
    .Q_N(_11999_),
    .Q(\top_ihp.oisc.regs[55][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1193),
    .D(_02101_),
    .Q_N(_11998_),
    .Q(\top_ihp.oisc.regs[55][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1180),
    .D(_02102_),
    .Q_N(_11997_),
    .Q(\top_ihp.oisc.regs[55][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1145),
    .D(_02103_),
    .Q_N(_11996_),
    .Q(\top_ihp.oisc.regs[55][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1207),
    .D(_02104_),
    .Q_N(_11995_),
    .Q(\top_ihp.oisc.regs[55][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1174),
    .D(_02105_),
    .Q_N(_11994_),
    .Q(\top_ihp.oisc.regs[55][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1171),
    .D(_02106_),
    .Q_N(_11993_),
    .Q(\top_ihp.oisc.regs[55][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1250),
    .D(_02107_),
    .Q_N(_11992_),
    .Q(\top_ihp.oisc.regs[55][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1248),
    .D(_02108_),
    .Q_N(_11991_),
    .Q(\top_ihp.oisc.regs[55][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1266),
    .D(_02109_),
    .Q_N(_11990_),
    .Q(\top_ihp.oisc.regs[55][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1113),
    .D(_02110_),
    .Q_N(_11989_),
    .Q(\top_ihp.oisc.regs[55][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1267),
    .D(_02111_),
    .Q_N(_11988_),
    .Q(\top_ihp.oisc.regs[55][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1201),
    .D(_02112_),
    .Q_N(_11987_),
    .Q(\top_ihp.oisc.regs[55][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1250),
    .D(_02113_),
    .Q_N(_11986_),
    .Q(\top_ihp.oisc.regs[55][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1235),
    .D(_02114_),
    .Q_N(_11985_),
    .Q(\top_ihp.oisc.regs[55][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[55][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1201),
    .D(_02115_),
    .Q_N(_11984_),
    .Q(\top_ihp.oisc.regs[55][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_282_clk),
    .RESET_B(net1281),
    .D(_02116_),
    .Q_N(_11983_),
    .Q(\top_ihp.oisc.regs[56][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1152),
    .D(_02117_),
    .Q_N(_11982_),
    .Q(\top_ihp.oisc.regs[56][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1223),
    .D(_02118_),
    .Q_N(_11981_),
    .Q(\top_ihp.oisc.regs[56][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1227),
    .D(_02119_),
    .Q_N(_11980_),
    .Q(\top_ihp.oisc.regs[56][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1313),
    .D(_02120_),
    .Q_N(_11979_),
    .Q(\top_ihp.oisc.regs[56][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1318),
    .D(_02121_),
    .Q_N(_11978_),
    .Q(\top_ihp.oisc.regs[56][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1317),
    .D(_02122_),
    .Q_N(_11977_),
    .Q(\top_ihp.oisc.regs[56][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1312),
    .D(_02123_),
    .Q_N(_11976_),
    .Q(\top_ihp.oisc.regs[56][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1262),
    .D(_02124_),
    .Q_N(_11975_),
    .Q(\top_ihp.oisc.regs[56][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1317),
    .D(_02125_),
    .Q_N(_11974_),
    .Q(\top_ihp.oisc.regs[56][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1273),
    .D(_02126_),
    .Q_N(_11973_),
    .Q(\top_ihp.oisc.regs[56][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1210),
    .D(_02127_),
    .Q_N(_11972_),
    .Q(\top_ihp.oisc.regs[56][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1256),
    .D(_02128_),
    .Q_N(_11971_),
    .Q(\top_ihp.oisc.regs[56][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1237),
    .D(_02129_),
    .Q_N(_11970_),
    .Q(\top_ihp.oisc.regs[56][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1191),
    .D(_02130_),
    .Q_N(_11969_),
    .Q(\top_ihp.oisc.regs[56][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1194),
    .D(_02131_),
    .Q_N(_11968_),
    .Q(\top_ihp.oisc.regs[56][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1152),
    .D(_02132_),
    .Q_N(_11967_),
    .Q(\top_ihp.oisc.regs[56][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1240),
    .D(_02133_),
    .Q_N(_11966_),
    .Q(\top_ihp.oisc.regs[56][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1179),
    .D(_02134_),
    .Q_N(_11965_),
    .Q(\top_ihp.oisc.regs[56][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1157),
    .D(_02135_),
    .Q_N(_11964_),
    .Q(\top_ihp.oisc.regs[56][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1229),
    .D(_02136_),
    .Q_N(_11963_),
    .Q(\top_ihp.oisc.regs[56][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_76_clk),
    .RESET_B(net1180),
    .D(_02137_),
    .Q_N(_11962_),
    .Q(\top_ihp.oisc.regs[56][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1169),
    .D(_02138_),
    .Q_N(_11961_),
    .Q(\top_ihp.oisc.regs[56][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1235),
    .D(_02139_),
    .Q_N(_11960_),
    .Q(\top_ihp.oisc.regs[56][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1235),
    .D(_02140_),
    .Q_N(_11959_),
    .Q(\top_ihp.oisc.regs[56][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1271),
    .D(_02141_),
    .Q_N(_11958_),
    .Q(\top_ihp.oisc.regs[56][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1270),
    .D(_02142_),
    .Q_N(_11957_),
    .Q(\top_ihp.oisc.regs[56][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1199),
    .D(_02143_),
    .Q_N(_11956_),
    .Q(\top_ihp.oisc.regs[56][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1212),
    .D(_02144_),
    .Q_N(_11955_),
    .Q(\top_ihp.oisc.regs[56][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1162),
    .D(_02145_),
    .Q_N(_11954_),
    .Q(\top_ihp.oisc.regs[56][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1207),
    .D(_02146_),
    .Q_N(_11953_),
    .Q(\top_ihp.oisc.regs[56][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[56][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1220),
    .D(_02147_),
    .Q_N(_11952_),
    .Q(\top_ihp.oisc.regs[56][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1289),
    .D(_02148_),
    .Q_N(_11951_),
    .Q(\top_ihp.oisc.regs[57][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1156),
    .D(_02149_),
    .Q_N(_11950_),
    .Q(\top_ihp.oisc.regs[57][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1215),
    .D(_02150_),
    .Q_N(_11949_),
    .Q(\top_ihp.oisc.regs[57][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1218),
    .D(_02151_),
    .Q_N(_11948_),
    .Q(\top_ihp.oisc.regs[57][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_110_clk),
    .RESET_B(net1314),
    .D(_02152_),
    .Q_N(_11947_),
    .Q(\top_ihp.oisc.regs[57][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_114_clk),
    .RESET_B(net1320),
    .D(_02153_),
    .Q_N(_11946_),
    .Q(\top_ihp.oisc.regs[57][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_02154_),
    .Q_N(_11945_),
    .Q(\top_ihp.oisc.regs[57][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1319),
    .D(_02155_),
    .Q_N(_11944_),
    .Q(\top_ihp.oisc.regs[57][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1262),
    .D(_02156_),
    .Q_N(_11943_),
    .Q(\top_ihp.oisc.regs[57][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1321),
    .D(_02157_),
    .Q_N(_11942_),
    .Q(\top_ihp.oisc.regs[57][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1289),
    .D(_02158_),
    .Q_N(_11941_),
    .Q(\top_ihp.oisc.regs[57][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1203),
    .D(_02159_),
    .Q_N(_11940_),
    .Q(\top_ihp.oisc.regs[57][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1256),
    .D(_02160_),
    .Q_N(_11939_),
    .Q(\top_ihp.oisc.regs[57][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1245),
    .D(_02161_),
    .Q_N(_11938_),
    .Q(\top_ihp.oisc.regs[57][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_80_clk),
    .RESET_B(net1241),
    .D(_02162_),
    .Q_N(_11937_),
    .Q(\top_ihp.oisc.regs[57][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1194),
    .D(_02163_),
    .Q_N(_11936_),
    .Q(\top_ihp.oisc.regs[57][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1154),
    .D(_02164_),
    .Q_N(_11935_),
    .Q(\top_ihp.oisc.regs[57][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_78_clk),
    .RESET_B(net1194),
    .D(_02165_),
    .Q_N(_11934_),
    .Q(\top_ihp.oisc.regs[57][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1314),
    .D(_02166_),
    .Q_N(_11933_),
    .Q(\top_ihp.oisc.regs[57][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1156),
    .D(_02167_),
    .Q_N(_11932_),
    .Q(\top_ihp.oisc.regs[57][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_297_clk),
    .RESET_B(net1157),
    .D(_02168_),
    .Q_N(_11931_),
    .Q(\top_ihp.oisc.regs[57][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_96_clk),
    .RESET_B(net1187),
    .D(_02169_),
    .Q_N(_11930_),
    .Q(\top_ihp.oisc.regs[57][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1186),
    .D(_02170_),
    .Q_N(_11929_),
    .Q(\top_ihp.oisc.regs[57][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1185),
    .D(_02171_),
    .Q_N(_11928_),
    .Q(\top_ihp.oisc.regs[57][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1230),
    .D(_02172_),
    .Q_N(_11927_),
    .Q(\top_ihp.oisc.regs[57][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1270),
    .D(_02173_),
    .Q_N(_11926_),
    .Q(\top_ihp.oisc.regs[57][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_298_clk),
    .RESET_B(net1157),
    .D(_02174_),
    .Q_N(_11925_),
    .Q(\top_ihp.oisc.regs[57][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1199),
    .D(_02175_),
    .Q_N(_11924_),
    .Q(\top_ihp.oisc.regs[57][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_306_clk),
    .RESET_B(net1217),
    .D(_02176_),
    .Q_N(_11923_),
    .Q(\top_ihp.oisc.regs[57][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net1185),
    .D(_02177_),
    .Q_N(_11922_),
    .Q(\top_ihp.oisc.regs[57][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1164),
    .D(_02178_),
    .Q_N(_11921_),
    .Q(\top_ihp.oisc.regs[57][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[57][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1202),
    .D(_02179_),
    .Q_N(_11920_),
    .Q(\top_ihp.oisc.regs[57][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1290),
    .D(_02180_),
    .Q_N(_11919_),
    .Q(\top_ihp.oisc.regs[58][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1140),
    .D(_02181_),
    .Q_N(_11918_),
    .Q(\top_ihp.oisc.regs[58][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1214),
    .D(_02182_),
    .Q_N(_11917_),
    .Q(\top_ihp.oisc.regs[58][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1226),
    .D(_02183_),
    .Q_N(_11916_),
    .Q(\top_ihp.oisc.regs[58][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_102_clk),
    .RESET_B(net1253),
    .D(_02184_),
    .Q_N(_11915_),
    .Q(\top_ihp.oisc.regs[58][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1299),
    .D(_02185_),
    .Q_N(_11914_),
    .Q(\top_ihp.oisc.regs[58][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1309),
    .D(_02186_),
    .Q_N(_11913_),
    .Q(\top_ihp.oisc.regs[58][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1299),
    .D(_02187_),
    .Q_N(_11912_),
    .Q(\top_ihp.oisc.regs[58][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1304),
    .D(_02188_),
    .Q_N(_11911_),
    .Q(\top_ihp.oisc.regs[58][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1304),
    .D(_02189_),
    .Q_N(_11910_),
    .Q(\top_ihp.oisc.regs[58][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1277),
    .D(_02190_),
    .Q_N(_11909_),
    .Q(\top_ihp.oisc.regs[58][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_300_clk),
    .RESET_B(net1203),
    .D(_02191_),
    .Q_N(_11908_),
    .Q(\top_ihp.oisc.regs[58][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1256),
    .D(_02192_),
    .Q_N(_11907_),
    .Q(\top_ihp.oisc.regs[58][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1232),
    .D(_02193_),
    .Q_N(_11906_),
    .Q(\top_ihp.oisc.regs[58][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1173),
    .D(_02194_),
    .Q_N(_11905_),
    .Q(\top_ihp.oisc.regs[58][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1174),
    .D(_02195_),
    .Q_N(_11904_),
    .Q(\top_ihp.oisc.regs[58][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1138),
    .D(_02196_),
    .Q_N(_11903_),
    .Q(\top_ihp.oisc.regs[58][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1172),
    .D(_02197_),
    .Q_N(_11902_),
    .Q(\top_ihp.oisc.regs[58][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_93_clk),
    .RESET_B(net1189),
    .D(_02198_),
    .Q_N(_11901_),
    .Q(\top_ihp.oisc.regs[58][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net1150),
    .D(_02199_),
    .Q_N(_11900_),
    .Q(\top_ihp.oisc.regs[58][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_294_clk),
    .RESET_B(net1162),
    .D(_02200_),
    .Q_N(_11899_),
    .Q(\top_ihp.oisc.regs[58][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1173),
    .D(_02201_),
    .Q_N(_11898_),
    .Q(\top_ihp.oisc.regs[58][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1171),
    .D(_02202_),
    .Q_N(_11897_),
    .Q(\top_ihp.oisc.regs[58][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1166),
    .D(_02203_),
    .Q_N(_11896_),
    .Q(\top_ihp.oisc.regs[58][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1223),
    .D(_02204_),
    .Q_N(_11895_),
    .Q(\top_ihp.oisc.regs[58][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_272_clk),
    .RESET_B(net1288),
    .D(_02205_),
    .Q_N(_11894_),
    .Q(\top_ihp.oisc.regs[58][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_312_clk),
    .RESET_B(net1155),
    .D(_02206_),
    .Q_N(_11893_),
    .Q(\top_ihp.oisc.regs[58][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1267),
    .D(_02207_),
    .Q_N(_11892_),
    .Q(\top_ihp.oisc.regs[58][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1201),
    .D(_02208_),
    .Q_N(_11891_),
    .Q(\top_ihp.oisc.regs[58][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1206),
    .D(_02209_),
    .Q_N(_11890_),
    .Q(\top_ihp.oisc.regs[58][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1235),
    .D(_02210_),
    .Q_N(_11889_),
    .Q(\top_ihp.oisc.regs[58][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[58][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_309_clk),
    .RESET_B(net1202),
    .D(_02211_),
    .Q_N(_11888_),
    .Q(\top_ihp.oisc.regs[58][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1313),
    .D(_02212_),
    .Q_N(_11887_),
    .Q(\top_ihp.oisc.regs[59][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1144),
    .D(_02213_),
    .Q_N(_11886_),
    .Q(\top_ihp.oisc.regs[59][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_291_clk),
    .RESET_B(net1227),
    .D(_02214_),
    .Q_N(_11885_),
    .Q(\top_ihp.oisc.regs[59][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1224),
    .D(_02215_),
    .Q_N(_11884_),
    .Q(\top_ihp.oisc.regs[59][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1295),
    .D(_02216_),
    .Q_N(_11883_),
    .Q(\top_ihp.oisc.regs[59][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1310),
    .D(_02217_),
    .Q_N(_11882_),
    .Q(\top_ihp.oisc.regs[59][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1253),
    .D(_02218_),
    .Q_N(_11881_),
    .Q(\top_ihp.oisc.regs[59][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1304),
    .D(_02219_),
    .Q_N(_11880_),
    .Q(\top_ihp.oisc.regs[59][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1262),
    .D(_02220_),
    .Q_N(_11879_),
    .Q(\top_ihp.oisc.regs[59][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1305),
    .D(_02221_),
    .Q_N(_11878_),
    .Q(\top_ihp.oisc.regs[59][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1272),
    .D(_02222_),
    .Q_N(_11877_),
    .Q(\top_ihp.oisc.regs[59][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1225),
    .D(_02223_),
    .Q_N(_11876_),
    .Q(\top_ihp.oisc.regs[59][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1257),
    .D(_02224_),
    .Q_N(_11875_),
    .Q(\top_ihp.oisc.regs[59][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1252),
    .D(_02225_),
    .Q_N(_11874_),
    .Q(\top_ihp.oisc.regs[59][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1173),
    .D(_02226_),
    .Q_N(_11873_),
    .Q(\top_ihp.oisc.regs[59][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1173),
    .D(_02227_),
    .Q_N(_11872_),
    .Q(\top_ihp.oisc.regs[59][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_314_clk),
    .RESET_B(net1142),
    .D(_02228_),
    .Q_N(_11871_),
    .Q(\top_ihp.oisc.regs[59][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1174),
    .D(_02229_),
    .Q_N(_11870_),
    .Q(\top_ihp.oisc.regs[59][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1174),
    .D(_02230_),
    .Q_N(_11869_),
    .Q(\top_ihp.oisc.regs[59][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1285),
    .D(_02231_),
    .Q_N(_11868_),
    .Q(\top_ihp.oisc.regs[59][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net1188),
    .D(_02232_),
    .Q_N(_11867_),
    .Q(\top_ihp.oisc.regs[59][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1173),
    .D(_02233_),
    .Q_N(_11866_),
    .Q(\top_ihp.oisc.regs[59][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_103_clk),
    .RESET_B(net1237),
    .D(_02234_),
    .Q_N(_11865_),
    .Q(\top_ihp.oisc.regs[59][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1166),
    .D(_02235_),
    .Q_N(_11864_),
    .Q(\top_ihp.oisc.regs[59][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net1230),
    .D(_02236_),
    .Q_N(_11863_),
    .Q(\top_ihp.oisc.regs[59][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_264_clk),
    .RESET_B(net1266),
    .D(_02237_),
    .Q_N(_11862_),
    .Q(\top_ihp.oisc.regs[59][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1198),
    .D(_02238_),
    .Q_N(_11861_),
    .Q(\top_ihp.oisc.regs[59][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_259_clk),
    .RESET_B(net1325),
    .D(_02239_),
    .Q_N(_11860_),
    .Q(\top_ihp.oisc.regs[59][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_303_clk),
    .RESET_B(net1218),
    .D(_02240_),
    .Q_N(_11859_),
    .Q(\top_ihp.oisc.regs[59][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net1188),
    .D(_02241_),
    .Q_N(_11858_),
    .Q(\top_ihp.oisc.regs[59][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1301),
    .D(_02242_),
    .Q_N(_11857_),
    .Q(\top_ihp.oisc.regs[59][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[59][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1218),
    .D(_02243_),
    .Q_N(_11856_),
    .Q(\top_ihp.oisc.regs[59][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1376),
    .D(_02244_),
    .Q_N(_11855_),
    .Q(\top_ihp.oisc.regs[5][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1385),
    .D(_02245_),
    .Q_N(_11854_),
    .Q(\top_ihp.oisc.regs[5][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1389),
    .D(_02246_),
    .Q_N(_11853_),
    .Q(\top_ihp.oisc.regs[5][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1341),
    .D(_02247_),
    .Q_N(_11852_),
    .Q(\top_ihp.oisc.regs[5][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_116_clk),
    .RESET_B(net1316),
    .D(_02248_),
    .Q_N(_11851_),
    .Q(\top_ihp.oisc.regs[5][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1321),
    .D(_02249_),
    .Q_N(_11850_),
    .Q(\top_ihp.oisc.regs[5][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_127_clk),
    .RESET_B(net1321),
    .D(_02250_),
    .Q_N(_11849_),
    .Q(\top_ihp.oisc.regs[5][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1321),
    .D(_02251_),
    .Q_N(_11848_),
    .Q(\top_ihp.oisc.regs[5][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1321),
    .D(_02252_),
    .Q_N(_11847_),
    .Q(\top_ihp.oisc.regs[5][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1322),
    .D(_02253_),
    .Q_N(_11846_),
    .Q(\top_ihp.oisc.regs[5][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1332),
    .D(_02254_),
    .Q_N(_11845_),
    .Q(\top_ihp.oisc.regs[5][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1378),
    .D(_02255_),
    .Q_N(_11844_),
    .Q(\top_ihp.oisc.regs[5][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1355),
    .D(_02256_),
    .Q_N(_11843_),
    .Q(\top_ihp.oisc.regs[5][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1322),
    .D(_02257_),
    .Q_N(_11842_),
    .Q(\top_ihp.oisc.regs[5][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_132_clk),
    .RESET_B(net1322),
    .D(_02258_),
    .Q_N(_11841_),
    .Q(\top_ihp.oisc.regs[5][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_133_clk),
    .RESET_B(net1355),
    .D(_02259_),
    .Q_N(_11840_),
    .Q(\top_ihp.oisc.regs[5][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1340),
    .D(_02260_),
    .Q_N(_11839_),
    .Q(\top_ihp.oisc.regs[5][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1320),
    .D(_02261_),
    .Q_N(_11838_),
    .Q(\top_ihp.oisc.regs[5][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_121_clk),
    .RESET_B(net1322),
    .D(_02262_),
    .Q_N(_11837_),
    .Q(\top_ihp.oisc.regs[5][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_276_clk),
    .RESET_B(net1332),
    .D(_02263_),
    .Q_N(_11836_),
    .Q(\top_ihp.oisc.regs[5][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1389),
    .D(_02264_),
    .Q_N(_11835_),
    .Q(\top_ihp.oisc.regs[5][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_122_clk),
    .RESET_B(net1322),
    .D(_02265_),
    .Q_N(_11834_),
    .Q(\top_ihp.oisc.regs[5][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1348),
    .D(_02266_),
    .Q_N(_11833_),
    .Q(\top_ihp.oisc.regs[5][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_196_clk),
    .RESET_B(net1348),
    .D(_02267_),
    .Q_N(_11832_),
    .Q(\top_ihp.oisc.regs[5][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1315),
    .D(_02268_),
    .Q_N(_11831_),
    .Q(\top_ihp.oisc.regs[5][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_253_clk),
    .RESET_B(net1338),
    .D(_02269_),
    .Q_N(_11830_),
    .Q(\top_ihp.oisc.regs[5][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1391),
    .D(_02270_),
    .Q_N(_11829_),
    .Q(\top_ihp.oisc.regs[5][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1329),
    .D(_02271_),
    .Q_N(_11828_),
    .Q(\top_ihp.oisc.regs[5][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1386),
    .D(_02272_),
    .Q_N(_11827_),
    .Q(\top_ihp.oisc.regs[5][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_197_clk),
    .RESET_B(net1315),
    .D(_02273_),
    .Q_N(_11826_),
    .Q(\top_ihp.oisc.regs[5][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_198_clk),
    .RESET_B(net1315),
    .D(_02274_),
    .Q_N(_11825_),
    .Q(\top_ihp.oisc.regs[5][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[5][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1388),
    .D(_02275_),
    .Q_N(_11824_),
    .Q(\top_ihp.oisc.regs[5][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1272),
    .D(_02276_),
    .Q_N(_11823_),
    .Q(\top_ihp.oisc.regs[60][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_316_clk),
    .RESET_B(net1138),
    .D(_02277_),
    .Q_N(_11822_),
    .Q(\top_ihp.oisc.regs[60][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_289_clk),
    .RESET_B(net1223),
    .D(_02278_),
    .Q_N(_11821_),
    .Q(\top_ihp.oisc.regs[60][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_286_clk),
    .RESET_B(net1226),
    .D(_02279_),
    .Q_N(_11820_),
    .Q(\top_ihp.oisc.regs[60][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1297),
    .D(_02280_),
    .Q_N(_11819_),
    .Q(\top_ihp.oisc.regs[60][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_123_clk),
    .RESET_B(net1308),
    .D(_02281_),
    .Q_N(_11818_),
    .Q(\top_ihp.oisc.regs[60][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_106_clk),
    .RESET_B(net1253),
    .D(_02282_),
    .Q_N(_11817_),
    .Q(\top_ihp.oisc.regs[60][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1310),
    .D(_02283_),
    .Q_N(_11816_),
    .Q(\top_ihp.oisc.regs[60][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_84_clk),
    .RESET_B(net1261),
    .D(_02284_),
    .Q_N(_11815_),
    .Q(\top_ihp.oisc.regs[60][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_128_clk),
    .RESET_B(net1310),
    .D(_02285_),
    .Q_N(_11814_),
    .Q(\top_ihp.oisc.regs[60][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_284_clk),
    .RESET_B(net1280),
    .D(_02286_),
    .Q_N(_11813_),
    .Q(\top_ihp.oisc.regs[60][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1223),
    .D(_02287_),
    .Q_N(_11812_),
    .Q(\top_ihp.oisc.regs[60][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_85_clk),
    .RESET_B(net1257),
    .D(_02288_),
    .Q_N(_11811_),
    .Q(\top_ihp.oisc.regs[60][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1232),
    .D(_02289_),
    .Q_N(_11810_),
    .Q(\top_ihp.oisc.regs[60][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1173),
    .D(_02290_),
    .Q_N(_11809_),
    .Q(\top_ihp.oisc.regs[60][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_74_clk),
    .RESET_B(net1173),
    .D(_02291_),
    .Q_N(_11808_),
    .Q(\top_ihp.oisc.regs[60][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1144),
    .D(_02292_),
    .Q_N(_11807_),
    .Q(\top_ihp.oisc.regs[60][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1175),
    .D(_02293_),
    .Q_N(_11806_),
    .Q(\top_ihp.oisc.regs[60][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1172),
    .D(_02294_),
    .Q_N(_11805_),
    .Q(\top_ihp.oisc.regs[60][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_296_clk),
    .RESET_B(net1150),
    .D(_02295_),
    .Q_N(_11804_),
    .Q(\top_ihp.oisc.regs[60][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1188),
    .D(_02296_),
    .Q_N(_11803_),
    .Q(\top_ihp.oisc.regs[60][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1173),
    .D(_02297_),
    .Q_N(_11802_),
    .Q(\top_ihp.oisc.regs[60][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1171),
    .D(_02298_),
    .Q_N(_11801_),
    .Q(\top_ihp.oisc.regs[60][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net1166),
    .D(_02299_),
    .Q_N(_11800_),
    .Q(\top_ihp.oisc.regs[60][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net1229),
    .D(_02300_),
    .Q_N(_11799_),
    .Q(\top_ihp.oisc.regs[60][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_265_clk),
    .RESET_B(net1269),
    .D(_02301_),
    .Q_N(_11798_),
    .Q(\top_ihp.oisc.regs[60][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1138),
    .D(_02302_),
    .Q_N(_11797_),
    .Q(\top_ihp.oisc.regs[60][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1198),
    .D(_02303_),
    .Q_N(_11796_),
    .Q(\top_ihp.oisc.regs[60][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1212),
    .D(_02304_),
    .Q_N(_11795_),
    .Q(\top_ihp.oisc.regs[60][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1148),
    .D(_02305_),
    .Q_N(_11794_),
    .Q(\top_ihp.oisc.regs[60][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_287_clk),
    .RESET_B(net1225),
    .D(_02306_),
    .Q_N(_11793_),
    .Q(\top_ihp.oisc.regs[60][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[60][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1202),
    .D(_02307_),
    .Q_N(_11792_),
    .Q(\top_ihp.oisc.regs[60][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1290),
    .D(_02308_),
    .Q_N(_11791_),
    .Q(\top_ihp.oisc.regs[61][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_319_clk),
    .RESET_B(net1145),
    .D(_02309_),
    .Q_N(_11790_),
    .Q(\top_ihp.oisc.regs[61][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_278_clk),
    .RESET_B(net1292),
    .D(_02310_),
    .Q_N(_11789_),
    .Q(\top_ihp.oisc.regs[61][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_301_clk),
    .RESET_B(net1218),
    .D(_02311_),
    .Q_N(_11788_),
    .Q(\top_ihp.oisc.regs[61][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_101_clk),
    .RESET_B(net1249),
    .D(_02312_),
    .Q_N(_11787_),
    .Q(\top_ihp.oisc.regs[61][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_113_clk),
    .RESET_B(net1308),
    .D(_02313_),
    .Q_N(_11786_),
    .Q(\top_ihp.oisc.regs[61][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1263),
    .D(_02314_),
    .Q_N(_11785_),
    .Q(\top_ihp.oisc.regs[61][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_129_clk),
    .RESET_B(net1310),
    .D(_02315_),
    .Q_N(_11784_),
    .Q(\top_ihp.oisc.regs[61][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1262),
    .D(_02316_),
    .Q_N(_11783_),
    .Q(\top_ihp.oisc.regs[61][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_131_clk),
    .RESET_B(net1310),
    .D(_02317_),
    .Q_N(_11782_),
    .Q(\top_ihp.oisc.regs[61][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_270_clk),
    .RESET_B(net1284),
    .D(_02318_),
    .Q_N(_11781_),
    .Q(\top_ihp.oisc.regs[61][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1200),
    .D(_02319_),
    .Q_N(_11780_),
    .Q(\top_ihp.oisc.regs[61][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1256),
    .D(_02320_),
    .Q_N(_11779_),
    .Q(\top_ihp.oisc.regs[61][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1311),
    .D(_02321_),
    .Q_N(_11778_),
    .Q(\top_ihp.oisc.regs[61][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1191),
    .D(_02322_),
    .Q_N(_11777_),
    .Q(\top_ihp.oisc.regs[61][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_77_clk),
    .RESET_B(net1194),
    .D(_02323_),
    .Q_N(_11776_),
    .Q(\top_ihp.oisc.regs[61][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_260_clk),
    .RESET_B(net1325),
    .D(_02324_),
    .Q_N(_11775_),
    .Q(\top_ihp.oisc.regs[61][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_71_clk),
    .RESET_B(net1177),
    .D(_02325_),
    .Q_N(_11774_),
    .Q(\top_ihp.oisc.regs[61][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_126_clk),
    .RESET_B(net1308),
    .D(_02326_),
    .Q_N(_11773_),
    .Q(\top_ihp.oisc.regs[61][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1285),
    .D(_02327_),
    .Q_N(_11772_),
    .Q(\top_ihp.oisc.regs[61][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_293_clk),
    .RESET_B(net1207),
    .D(_02328_),
    .Q_N(_11771_),
    .Q(\top_ihp.oisc.regs[61][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_70_clk),
    .RESET_B(net1176),
    .D(_02329_),
    .Q_N(_11770_),
    .Q(\top_ihp.oisc.regs[61][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net1168),
    .D(_02330_),
    .Q_N(_11769_),
    .Q(\top_ihp.oisc.regs[61][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1166),
    .D(_02331_),
    .Q_N(_11768_),
    .Q(\top_ihp.oisc.regs[61][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net1251),
    .D(_02332_),
    .Q_N(_11767_),
    .Q(\top_ihp.oisc.regs[61][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1284),
    .D(_02333_),
    .Q_N(_11766_),
    .Q(\top_ihp.oisc.regs[61][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_263_clk),
    .RESET_B(net1270),
    .D(_02334_),
    .Q_N(_11765_),
    .Q(\top_ihp.oisc.regs[61][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_261_clk),
    .RESET_B(net1286),
    .D(_02335_),
    .Q_N(_11764_),
    .Q(\top_ihp.oisc.regs[61][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_308_clk),
    .RESET_B(net1212),
    .D(_02336_),
    .Q_N(_11763_),
    .Q(\top_ihp.oisc.regs[61][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1158),
    .D(_02337_),
    .Q_N(_11762_),
    .Q(\top_ihp.oisc.regs[61][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1149),
    .D(_02338_),
    .Q_N(_11761_),
    .Q(\top_ihp.oisc.regs[61][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[61][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_307_clk),
    .RESET_B(net1220),
    .D(_02339_),
    .Q_N(_11760_),
    .Q(\top_ihp.oisc.regs[61][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1285),
    .D(_02340_),
    .Q_N(_11759_),
    .Q(\top_ihp.oisc.regs[62][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1141),
    .D(_02341_),
    .Q_N(_11758_),
    .Q(\top_ihp.oisc.regs[62][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1227),
    .D(_02342_),
    .Q_N(_11757_),
    .Q(\top_ihp.oisc.regs[62][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1219),
    .D(_02343_),
    .Q_N(_11756_),
    .Q(\top_ihp.oisc.regs[62][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1249),
    .D(_02344_),
    .Q_N(_11755_),
    .Q(\top_ihp.oisc.regs[62][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_124_clk),
    .RESET_B(net1306),
    .D(_02345_),
    .Q_N(_11754_),
    .Q(\top_ihp.oisc.regs[62][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1310),
    .D(_02346_),
    .Q_N(_11753_),
    .Q(\top_ihp.oisc.regs[62][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_111_clk),
    .RESET_B(net1296),
    .D(_02347_),
    .Q_N(_11752_),
    .Q(\top_ihp.oisc.regs[62][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_83_clk),
    .RESET_B(net1262),
    .D(_02348_),
    .Q_N(_11751_),
    .Q(\top_ihp.oisc.regs[62][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_130_clk),
    .RESET_B(net1305),
    .D(_02349_),
    .Q_N(_11750_),
    .Q(\top_ihp.oisc.regs[62][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_108_clk),
    .RESET_B(net1298),
    .D(_02350_),
    .Q_N(_11749_),
    .Q(\top_ihp.oisc.regs[62][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_299_clk),
    .RESET_B(net1205),
    .D(_02351_),
    .Q_N(_11748_),
    .Q(\top_ihp.oisc.regs[62][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1257),
    .D(_02352_),
    .Q_N(_11747_),
    .Q(\top_ihp.oisc.regs[62][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_82_clk),
    .RESET_B(net1257),
    .D(_02353_),
    .Q_N(_11746_),
    .Q(\top_ihp.oisc.regs[62][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_81_clk),
    .RESET_B(net1241),
    .D(_02354_),
    .Q_N(_11745_),
    .Q(\top_ihp.oisc.regs[62][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_75_clk),
    .RESET_B(net1175),
    .D(_02355_),
    .Q_N(_11744_),
    .Q(\top_ihp.oisc.regs[62][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_315_clk),
    .RESET_B(net1139),
    .D(_02356_),
    .Q_N(_11743_),
    .Q(\top_ihp.oisc.regs[62][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1161),
    .D(_02357_),
    .Q_N(_11742_),
    .Q(\top_ihp.oisc.regs[62][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1176),
    .D(_02358_),
    .Q_N(_11741_),
    .Q(\top_ihp.oisc.regs[62][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net1147),
    .D(_02359_),
    .Q_N(_11740_),
    .Q(\top_ihp.oisc.regs[62][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1162),
    .D(_02360_),
    .Q_N(_11739_),
    .Q(\top_ihp.oisc.regs[62][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_94_clk),
    .RESET_B(net1171),
    .D(_02361_),
    .Q_N(_11738_),
    .Q(\top_ihp.oisc.regs[62][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_37_clk),
    .RESET_B(net1171),
    .D(_02362_),
    .Q_N(_11737_),
    .Q(\top_ihp.oisc.regs[62][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net1166),
    .D(_02363_),
    .Q_N(_11736_),
    .Q(\top_ihp.oisc.regs[62][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_104_clk),
    .RESET_B(net1250),
    .D(_02364_),
    .Q_N(_11735_),
    .Q(\top_ihp.oisc.regs[62][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_267_clk),
    .RESET_B(net1273),
    .D(_02365_),
    .Q_N(_11734_),
    .Q(\top_ihp.oisc.regs[62][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1290),
    .D(_02366_),
    .Q_N(_11733_),
    .Q(\top_ihp.oisc.regs[62][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_311_clk),
    .RESET_B(net1199),
    .D(_02367_),
    .Q_N(_11732_),
    .Q(\top_ihp.oisc.regs[62][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_304_clk),
    .RESET_B(net1205),
    .D(_02368_),
    .Q_N(_11731_),
    .Q(\top_ihp.oisc.regs[62][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1150),
    .D(_02369_),
    .Q_N(_11730_),
    .Q(\top_ihp.oisc.regs[62][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net1150),
    .D(_02370_),
    .Q_N(_11729_),
    .Q(\top_ihp.oisc.regs[62][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[62][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_310_clk),
    .RESET_B(net1202),
    .D(_02371_),
    .Q_N(_11728_),
    .Q(\top_ihp.oisc.regs[62][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1291),
    .D(_02372_),
    .Q_N(_11727_),
    .Q(\top_ihp.oisc.regs[63][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1288),
    .D(_02373_),
    .Q_N(_11726_),
    .Q(\top_ihp.oisc.regs[63][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_292_clk),
    .RESET_B(net1221),
    .D(_02374_),
    .Q_N(_11725_),
    .Q(\top_ihp.oisc.regs[63][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_290_clk),
    .RESET_B(net1224),
    .D(_02375_),
    .Q_N(_11724_),
    .Q(\top_ihp.oisc.regs[63][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_105_clk),
    .RESET_B(net1251),
    .D(_02376_),
    .Q_N(_11723_),
    .Q(\top_ihp.oisc.regs[63][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_109_clk),
    .RESET_B(net1314),
    .D(_02377_),
    .Q_N(_11722_),
    .Q(\top_ihp.oisc.regs[63][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_285_clk),
    .RESET_B(net1276),
    .D(_02378_),
    .Q_N(_11721_),
    .Q(\top_ihp.oisc.regs[63][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_115_clk),
    .RESET_B(net1314),
    .D(_02379_),
    .Q_N(_11720_),
    .Q(\top_ihp.oisc.regs[63][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_88_clk),
    .RESET_B(net1258),
    .D(_02380_),
    .Q_N(_11719_),
    .Q(\top_ihp.oisc.regs[63][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_125_clk),
    .RESET_B(net1306),
    .D(_02381_),
    .Q_N(_11718_),
    .Q(\top_ihp.oisc.regs[63][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_283_clk),
    .RESET_B(net1291),
    .D(_02382_),
    .Q_N(_11717_),
    .Q(\top_ihp.oisc.regs[63][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_288_clk),
    .RESET_B(net1210),
    .D(_02383_),
    .Q_N(_11716_),
    .Q(\top_ihp.oisc.regs[63][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_89_clk),
    .RESET_B(net1243),
    .D(_02384_),
    .Q_N(_11715_),
    .Q(\top_ihp.oisc.regs[63][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_99_clk),
    .RESET_B(net1236),
    .D(_02385_),
    .Q_N(_11714_),
    .Q(\top_ihp.oisc.regs[63][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_98_clk),
    .RESET_B(net1232),
    .D(_02386_),
    .Q_N(_11713_),
    .Q(\top_ihp.oisc.regs[63][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_79_clk),
    .RESET_B(net1194),
    .D(_02387_),
    .Q_N(_11712_),
    .Q(\top_ihp.oisc.regs[63][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_317_clk),
    .RESET_B(net1154),
    .D(_02388_),
    .Q_N(_11711_),
    .Q(\top_ihp.oisc.regs[63][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1193),
    .D(_02389_),
    .Q_N(_11710_),
    .Q(\top_ihp.oisc.regs[63][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1191),
    .D(_02390_),
    .Q_N(_11709_),
    .Q(\top_ihp.oisc.regs[63][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_295_clk),
    .RESET_B(net1161),
    .D(_02391_),
    .Q_N(_11708_),
    .Q(\top_ihp.oisc.regs[63][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net1206),
    .D(_02392_),
    .Q_N(_11707_),
    .Q(\top_ihp.oisc.regs[63][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_72_clk),
    .RESET_B(net1191),
    .D(_02393_),
    .Q_N(_11706_),
    .Q(\top_ihp.oisc.regs[63][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net1184),
    .D(_02394_),
    .Q_N(_11705_),
    .Q(\top_ihp.oisc.regs[63][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net1234),
    .D(_02395_),
    .Q_N(_11704_),
    .Q(\top_ihp.oisc.regs[63][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net1206),
    .D(_02396_),
    .Q_N(_11703_),
    .Q(\top_ihp.oisc.regs[63][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_266_clk),
    .RESET_B(net1285),
    .D(_02397_),
    .Q_N(_11702_),
    .Q(\top_ihp.oisc.regs[63][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_279_clk),
    .RESET_B(net1292),
    .D(_02398_),
    .Q_N(_11701_),
    .Q(\top_ihp.oisc.regs[63][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_271_clk),
    .RESET_B(net1287),
    .D(_02399_),
    .Q_N(_11700_),
    .Q(\top_ihp.oisc.regs[63][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_305_clk),
    .RESET_B(net1213),
    .D(_02400_),
    .Q_N(_11699_),
    .Q(\top_ihp.oisc.regs[63][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net1164),
    .D(_02401_),
    .Q_N(_11698_),
    .Q(\top_ihp.oisc.regs[63][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net1209),
    .D(_02402_),
    .Q_N(_11697_),
    .Q(\top_ihp.oisc.regs[63][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[63][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_302_clk),
    .RESET_B(net1215),
    .D(_02403_),
    .Q_N(_11696_),
    .Q(\top_ihp.oisc.regs[63][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1374),
    .D(_02404_),
    .Q_N(_11695_),
    .Q(\top_ihp.oisc.regs[6][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1383),
    .D(_02405_),
    .Q_N(_11694_),
    .Q(\top_ihp.oisc.regs[6][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1380),
    .D(_02406_),
    .Q_N(_11693_),
    .Q(\top_ihp.oisc.regs[6][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1343),
    .D(_02407_),
    .Q_N(_11692_),
    .Q(\top_ihp.oisc.regs[6][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1406),
    .D(_02408_),
    .Q_N(_11691_),
    .Q(\top_ihp.oisc.regs[6][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_02409_),
    .Q_N(_11690_),
    .Q(\top_ihp.oisc.regs[6][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1407),
    .D(_02410_),
    .Q_N(_11689_),
    .Q(\top_ihp.oisc.regs[6][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_118_clk),
    .RESET_B(net1362),
    .D(_02411_),
    .Q_N(_11688_),
    .Q(\top_ihp.oisc.regs[6][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1362),
    .D(_02412_),
    .Q_N(_11687_),
    .Q(\top_ihp.oisc.regs[6][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_02413_),
    .Q_N(_11686_),
    .Q(\top_ihp.oisc.regs[6][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1345),
    .D(_02414_),
    .Q_N(_11685_),
    .Q(\top_ihp.oisc.regs[6][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1382),
    .D(_02415_),
    .Q_N(_11684_),
    .Q(\top_ihp.oisc.regs[6][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_142_clk),
    .RESET_B(net1401),
    .D(_02416_),
    .Q_N(_11683_),
    .Q(\top_ihp.oisc.regs[6][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1369),
    .D(_02417_),
    .Q_N(_11682_),
    .Q(\top_ihp.oisc.regs[6][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_168_clk),
    .RESET_B(net1407),
    .D(_02418_),
    .Q_N(_11681_),
    .Q(\top_ihp.oisc.regs[6][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1411),
    .D(_02419_),
    .Q_N(_11680_),
    .Q(\top_ihp.oisc.regs[6][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1372),
    .D(_02420_),
    .Q_N(_11679_),
    .Q(\top_ihp.oisc.regs[6][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1369),
    .D(_02421_),
    .Q_N(_11678_),
    .Q(\top_ihp.oisc.regs[6][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1412),
    .D(_02422_),
    .Q_N(_11677_),
    .Q(\top_ihp.oisc.regs[6][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_210_clk),
    .RESET_B(net1381),
    .D(_02423_),
    .Q_N(_11676_),
    .Q(\top_ihp.oisc.regs[6][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1392),
    .D(_02424_),
    .Q_N(_11675_),
    .Q(\top_ihp.oisc.regs[6][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1407),
    .D(_02425_),
    .Q_N(_11674_),
    .Q(\top_ihp.oisc.regs[6][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1397),
    .D(_02426_),
    .Q_N(_11673_),
    .Q(\top_ihp.oisc.regs[6][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1363),
    .D(_02427_),
    .Q_N(_11672_),
    .Q(\top_ihp.oisc.regs[6][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_193_clk),
    .RESET_B(net1361),
    .D(_02428_),
    .Q_N(_11671_),
    .Q(\top_ihp.oisc.regs[6][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1336),
    .D(_02429_),
    .Q_N(_11670_),
    .Q(\top_ihp.oisc.regs[6][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1387),
    .D(_02430_),
    .Q_N(_11669_),
    .Q(\top_ihp.oisc.regs[6][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_257_clk),
    .RESET_B(net1337),
    .D(_02431_),
    .Q_N(_11668_),
    .Q(\top_ihp.oisc.regs[6][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_245_clk),
    .RESET_B(net1383),
    .D(_02432_),
    .Q_N(_11667_),
    .Q(\top_ihp.oisc.regs[6][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_182_clk),
    .RESET_B(net1406),
    .D(_02433_),
    .Q_N(_11666_),
    .Q(\top_ihp.oisc.regs[6][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1392),
    .D(_02434_),
    .Q_N(_11665_),
    .Q(\top_ihp.oisc.regs[6][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[6][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1387),
    .D(_02435_),
    .Q_N(_11664_),
    .Q(\top_ihp.oisc.regs[6][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1376),
    .D(_02436_),
    .Q_N(_11663_),
    .Q(\top_ihp.oisc.regs[7][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1384),
    .D(_02437_),
    .Q_N(_11662_),
    .Q(\top_ihp.oisc.regs[7][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1390),
    .D(_02438_),
    .Q_N(_11661_),
    .Q(\top_ihp.oisc.regs[7][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1333),
    .D(_02439_),
    .Q_N(_11660_),
    .Q(\top_ihp.oisc.regs[7][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_186_clk),
    .RESET_B(net1405),
    .D(_02440_),
    .Q_N(_11659_),
    .Q(\top_ihp.oisc.regs[7][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1407),
    .D(_02441_),
    .Q_N(_11658_),
    .Q(\top_ihp.oisc.regs[7][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1404),
    .D(_02442_),
    .Q_N(_11657_),
    .Q(\top_ihp.oisc.regs[7][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1366),
    .D(_02443_),
    .Q_N(_11656_),
    .Q(\top_ihp.oisc.regs[7][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1370),
    .D(_02444_),
    .Q_N(_11655_),
    .Q(\top_ihp.oisc.regs[7][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1370),
    .D(_02445_),
    .Q_N(_11654_),
    .Q(\top_ihp.oisc.regs[7][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1341),
    .D(_02446_),
    .Q_N(_11653_),
    .Q(\top_ihp.oisc.regs[7][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1378),
    .D(_02447_),
    .Q_N(_11652_),
    .Q(\top_ihp.oisc.regs[7][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1370),
    .D(_02448_),
    .Q_N(_11651_),
    .Q(\top_ihp.oisc.regs[7][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1368),
    .D(_02449_),
    .Q_N(_11650_),
    .Q(\top_ihp.oisc.regs[7][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_144_clk),
    .RESET_B(net1412),
    .D(_02450_),
    .Q_N(_11649_),
    .Q(\top_ihp.oisc.regs[7][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_150_clk),
    .RESET_B(net1412),
    .D(_02451_),
    .Q_N(_11648_),
    .Q(\top_ihp.oisc.regs[7][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1377),
    .D(_02452_),
    .Q_N(_11647_),
    .Q(\top_ihp.oisc.regs[7][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1368),
    .D(_02453_),
    .Q_N(_11646_),
    .Q(\top_ihp.oisc.regs[7][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_138_clk),
    .RESET_B(net1368),
    .D(_02454_),
    .Q_N(_11645_),
    .Q(\top_ihp.oisc.regs[7][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_208_clk),
    .RESET_B(net1379),
    .D(_02455_),
    .Q_N(_11644_),
    .Q(\top_ihp.oisc.regs[7][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1390),
    .D(_02456_),
    .Q_N(_11643_),
    .Q(\top_ihp.oisc.regs[7][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_146_clk),
    .RESET_B(net1402),
    .D(_02457_),
    .Q_N(_11642_),
    .Q(\top_ihp.oisc.regs[7][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_188_clk),
    .RESET_B(net1398),
    .D(_02458_),
    .Q_N(_11641_),
    .Q(\top_ihp.oisc.regs[7][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1363),
    .D(_02459_),
    .Q_N(_11640_),
    .Q(\top_ihp.oisc.regs[7][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1361),
    .D(_02460_),
    .Q_N(_11639_),
    .Q(\top_ihp.oisc.regs[7][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_254_clk),
    .RESET_B(net1328),
    .D(_02461_),
    .Q_N(_11638_),
    .Q(\top_ihp.oisc.regs[7][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1389),
    .D(_02462_),
    .Q_N(_11637_),
    .Q(\top_ihp.oisc.regs[7][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1329),
    .D(_02463_),
    .Q_N(_11636_),
    .Q(\top_ihp.oisc.regs[7][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_229_clk),
    .RESET_B(net1386),
    .D(_02464_),
    .Q_N(_11635_),
    .Q(\top_ihp.oisc.regs[7][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1397),
    .D(_02465_),
    .Q_N(_11634_),
    .Q(\top_ihp.oisc.regs[7][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_184_clk),
    .RESET_B(net1397),
    .D(_02466_),
    .Q_N(_11633_),
    .Q(\top_ihp.oisc.regs[7][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[7][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_252_clk),
    .RESET_B(net1340),
    .D(_02467_),
    .Q_N(_11632_),
    .Q(\top_ihp.oisc.regs[7][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_249_clk),
    .RESET_B(net1374),
    .D(_02468_),
    .Q_N(_11631_),
    .Q(\top_ihp.oisc.regs[8][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_250_clk),
    .RESET_B(net1387),
    .D(_02469_),
    .Q_N(_11630_),
    .Q(\top_ihp.oisc.regs[8][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_207_clk),
    .RESET_B(net1380),
    .D(_02470_),
    .Q_N(_11629_),
    .Q(\top_ihp.oisc.regs[8][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_277_clk),
    .RESET_B(net1333),
    .D(_02471_),
    .Q_N(_11628_),
    .Q(\top_ihp.oisc.regs[8][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_192_clk),
    .RESET_B(net1351),
    .D(_02472_),
    .Q_N(_11627_),
    .Q(\top_ihp.oisc.regs[8][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_148_clk),
    .RESET_B(net1403),
    .D(_02473_),
    .Q_N(_11626_),
    .Q(\top_ihp.oisc.regs[8][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_147_clk),
    .RESET_B(net1402),
    .D(_02474_),
    .Q_N(_11625_),
    .Q(\top_ihp.oisc.regs[8][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_136_clk),
    .RESET_B(net1366),
    .D(_02475_),
    .Q_N(_11624_),
    .Q(\top_ihp.oisc.regs[8][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_134_clk),
    .RESET_B(net1360),
    .D(_02476_),
    .Q_N(_11623_),
    .Q(\top_ihp.oisc.regs[8][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_137_clk),
    .RESET_B(net1369),
    .D(_02477_),
    .Q_N(_11622_),
    .Q(\top_ihp.oisc.regs[8][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_203_clk),
    .RESET_B(net1345),
    .D(_02478_),
    .Q_N(_11621_),
    .Q(\top_ihp.oisc.regs[8][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_202_clk),
    .RESET_B(net1346),
    .D(_02479_),
    .Q_N(_11620_),
    .Q(\top_ihp.oisc.regs[8][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_164_clk),
    .RESET_B(net1413),
    .D(_02480_),
    .Q_N(_11619_),
    .Q(\top_ihp.oisc.regs[8][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_190_clk),
    .RESET_B(net1364),
    .D(_02481_),
    .Q_N(_11618_),
    .Q(\top_ihp.oisc.regs[8][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1413),
    .D(_02482_),
    .Q_N(_11617_),
    .Q(\top_ihp.oisc.regs[8][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1414),
    .D(_02483_),
    .Q_N(_11616_),
    .Q(\top_ihp.oisc.regs[8][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_248_clk),
    .RESET_B(net1372),
    .D(_02484_),
    .Q_N(_11615_),
    .Q(\top_ihp.oisc.regs[8][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1400),
    .D(_02485_),
    .Q_N(_11614_),
    .Q(\top_ihp.oisc.regs[8][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1408),
    .D(_02486_),
    .Q_N(_11613_),
    .Q(\top_ihp.oisc.regs[8][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_211_clk),
    .RESET_B(net1381),
    .D(_02487_),
    .Q_N(_11612_),
    .Q(\top_ihp.oisc.regs[8][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_213_clk),
    .RESET_B(net1392),
    .D(_02488_),
    .Q_N(_11611_),
    .Q(\top_ihp.oisc.regs[8][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1410),
    .D(_02489_),
    .Q_N(_11610_),
    .Q(\top_ihp.oisc.regs[8][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_185_clk),
    .RESET_B(net1395),
    .D(_02490_),
    .Q_N(_11609_),
    .Q(\top_ihp.oisc.regs[8][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1363),
    .D(_02491_),
    .Q_N(_11608_),
    .Q(\top_ihp.oisc.regs[8][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_195_clk),
    .RESET_B(net1352),
    .D(_02492_),
    .Q_N(_11607_),
    .Q(\top_ihp.oisc.regs[8][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1337),
    .D(_02493_),
    .Q_N(_11606_),
    .Q(\top_ihp.oisc.regs[8][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1339),
    .D(_02494_),
    .Q_N(_11605_),
    .Q(\top_ihp.oisc.regs[8][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_255_clk),
    .RESET_B(net1339),
    .D(_02495_),
    .Q_N(_11604_),
    .Q(\top_ihp.oisc.regs[8][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_274_clk),
    .RESET_B(net1329),
    .D(_02496_),
    .Q_N(_11603_),
    .Q(\top_ihp.oisc.regs[8][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1410),
    .D(_02497_),
    .Q_N(_11602_),
    .Q(\top_ihp.oisc.regs[8][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_212_clk),
    .RESET_B(net1392),
    .D(_02498_),
    .Q_N(_11601_),
    .Q(\top_ihp.oisc.regs[8][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[8][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_230_clk),
    .RESET_B(net1388),
    .D(_02499_),
    .Q_N(_11600_),
    .Q(\top_ihp.oisc.regs[8][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][0]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1374),
    .D(_02500_),
    .Q_N(_11599_),
    .Q(\top_ihp.oisc.regs[9][0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][10]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1383),
    .D(_02501_),
    .Q_N(_11598_),
    .Q(\top_ihp.oisc.regs[9][10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][11]$_DFFE_PN0P_  (.CLK(clknet_leaf_227_clk),
    .RESET_B(net1389),
    .D(_02502_),
    .Q_N(_11597_),
    .Q(\top_ihp.oisc.regs[9][11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][12]$_DFFE_PN0P_  (.CLK(clknet_leaf_275_clk),
    .RESET_B(net1343),
    .D(_02503_),
    .Q_N(_11596_),
    .Q(\top_ihp.oisc.regs[9][12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][13]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1408),
    .D(_02504_),
    .Q_N(_11595_),
    .Q(\top_ihp.oisc.regs[9][13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][14]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1411),
    .D(_02505_),
    .Q_N(_11594_),
    .Q(\top_ihp.oisc.regs[9][14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][15]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1411),
    .D(_02506_),
    .Q_N(_11593_),
    .Q(\top_ihp.oisc.regs[9][15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][16]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1359),
    .D(_02507_),
    .Q_N(_11592_),
    .Q(\top_ihp.oisc.regs[9][16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][17]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1367),
    .D(_02508_),
    .Q_N(_11591_),
    .Q(\top_ihp.oisc.regs[9][17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][18]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1369),
    .D(_02509_),
    .Q_N(_11590_),
    .Q(\top_ihp.oisc.regs[9][18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][19]$_DFFE_PN0P_  (.CLK(clknet_leaf_205_clk),
    .RESET_B(net1341),
    .D(_02510_),
    .Q_N(_11589_),
    .Q(\top_ihp.oisc.regs[9][19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][1]$_DFFE_PN0P_  (.CLK(clknet_leaf_206_clk),
    .RESET_B(net1378),
    .D(_02511_),
    .Q_N(_11588_),
    .Q(\top_ihp.oisc.regs[9][1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][20]$_DFFE_PN0P_  (.CLK(clknet_leaf_166_clk),
    .RESET_B(net1400),
    .D(_02512_),
    .Q_N(_11587_),
    .Q(\top_ihp.oisc.regs[9][20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][21]$_DFFE_PN0P_  (.CLK(clknet_leaf_119_clk),
    .RESET_B(net1359),
    .D(_02513_),
    .Q_N(_11586_),
    .Q(\top_ihp.oisc.regs[9][21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][22]$_DFFE_PN0P_  (.CLK(clknet_leaf_167_clk),
    .RESET_B(net1412),
    .D(_02514_),
    .Q_N(_11585_),
    .Q(\top_ihp.oisc.regs[9][22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][23]$_DFFE_PN0P_  (.CLK(clknet_leaf_165_clk),
    .RESET_B(net1412),
    .D(_02515_),
    .Q_N(_11584_),
    .Q(\top_ihp.oisc.regs[9][23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][24]$_DFFE_PN0P_  (.CLK(clknet_leaf_256_clk),
    .RESET_B(net1340),
    .D(_02516_),
    .Q_N(_11583_),
    .Q(\top_ihp.oisc.regs[9][24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][25]$_DFFE_PN0P_  (.CLK(clknet_leaf_141_clk),
    .RESET_B(net1359),
    .D(_02517_),
    .Q_N(_11582_),
    .Q(\top_ihp.oisc.regs[9][25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][26]$_DFFE_PN0P_  (.CLK(clknet_leaf_187_clk),
    .RESET_B(net1408),
    .D(_02518_),
    .Q_N(_11581_),
    .Q(\top_ihp.oisc.regs[9][26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][27]$_DFFE_PN0P_  (.CLK(clknet_leaf_228_clk),
    .RESET_B(net1377),
    .D(_02519_),
    .Q_N(_11580_),
    .Q(\top_ihp.oisc.regs[9][27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][28]$_DFFE_PN0P_  (.CLK(clknet_leaf_209_clk),
    .RESET_B(net1390),
    .D(_02520_),
    .Q_N(_11579_),
    .Q(\top_ihp.oisc.regs[9][28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][29]$_DFFE_PN0P_  (.CLK(clknet_leaf_169_clk),
    .RESET_B(net1408),
    .D(_02521_),
    .Q_N(_11578_),
    .Q(\top_ihp.oisc.regs[9][29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][2]$_DFFE_PN0P_  (.CLK(clknet_leaf_191_clk),
    .RESET_B(net1362),
    .D(_02522_),
    .Q_N(_11577_),
    .Q(\top_ihp.oisc.regs[9][2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][30]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1363),
    .D(_02523_),
    .Q_N(_11576_),
    .Q(\top_ihp.oisc.regs[9][30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][31]$_DFFE_PN0P_  (.CLK(clknet_leaf_194_clk),
    .RESET_B(net1352),
    .D(_02524_),
    .Q_N(_11575_),
    .Q(\top_ihp.oisc.regs[9][31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][3]$_DFFE_PN0P_  (.CLK(clknet_leaf_258_clk),
    .RESET_B(net1329),
    .D(_02525_),
    .Q_N(_11574_),
    .Q(\top_ihp.oisc.regs[9][3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][4]$_DFFE_PN0P_  (.CLK(clknet_leaf_247_clk),
    .RESET_B(net1374),
    .D(_02526_),
    .Q_N(_11573_),
    .Q(\top_ihp.oisc.regs[9][4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][5]$_DFFE_PN0P_  (.CLK(clknet_leaf_273_clk),
    .RESET_B(net1335),
    .D(_02527_),
    .Q_N(_11572_),
    .Q(\top_ihp.oisc.regs[9][5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][6]$_DFFE_PN0P_  (.CLK(clknet_leaf_244_clk),
    .RESET_B(net1383),
    .D(_02528_),
    .Q_N(_11571_),
    .Q(\top_ihp.oisc.regs[9][6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][7]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1406),
    .D(_02529_),
    .Q_N(_11570_),
    .Q(\top_ihp.oisc.regs[9][7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][8]$_DFFE_PN0P_  (.CLK(clknet_leaf_183_clk),
    .RESET_B(net1406),
    .D(_02530_),
    .Q_N(_11569_),
    .Q(\top_ihp.oisc.regs[9][8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.regs[9][9]$_DFFE_PN0P_  (.CLK(clknet_leaf_246_clk),
    .RESET_B(net1383),
    .D(_02531_),
    .Q_N(_11568_),
    .Q(\top_ihp.oisc.regs[9][9] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[0]$_DFFE_PN1P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1114),
    .D(_02532_),
    .Q_N(\top_ihp.oisc.state[0] ),
    .Q(_13699_));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1114),
    .D(_02533_),
    .Q_N(_11567_),
    .Q(\top_ihp.oisc.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1114),
    .D(_02534_),
    .Q_N(_00092_),
    .Q(\top_ihp.oisc.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_320_clk),
    .RESET_B(net1114),
    .D(_02535_),
    .Q_N(_00091_),
    .Q(\top_ihp.oisc.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1113),
    .D(_02536_),
    .Q_N(_00093_),
    .Q(\top_ihp.oisc.state[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[5]$_DFF_PN0_  (.CLK(clknet_leaf_322_clk),
    .RESET_B(net1113),
    .D(_00002_),
    .Q_N(_00078_),
    .Q(\top_ihp.oisc.state[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.state[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_321_clk),
    .RESET_B(net1111),
    .D(_02537_),
    .Q_N(_11566_),
    .Q(\top_ihp.oisc.state[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1119),
    .D(_02538_),
    .Q_N(_00222_),
    .Q(\top_ihp.oisc.wb_dat_o[0] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1078),
    .D(_02539_),
    .Q_N(_11565_),
    .Q(\top_ihp.oisc.wb_dat_o[10] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1085),
    .D(_02540_),
    .Q_N(_11564_),
    .Q(\top_ihp.oisc.wb_dat_o[11] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1133),
    .D(_02541_),
    .Q_N(_11563_),
    .Q(\top_ihp.oisc.wb_dat_o[12] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1089),
    .D(_02542_),
    .Q_N(_11562_),
    .Q(\top_ihp.oisc.wb_dat_o[13] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1134),
    .D(_02543_),
    .Q_N(_11561_),
    .Q(\top_ihp.oisc.wb_dat_o[14] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1085),
    .D(_02544_),
    .Q_N(_11560_),
    .Q(\top_ihp.oisc.wb_dat_o[15] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1134),
    .D(_02545_),
    .Q_N(_11559_),
    .Q(\top_ihp.oisc.wb_dat_o[16] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1078),
    .D(_02546_),
    .Q_N(_11558_),
    .Q(\top_ihp.oisc.wb_dat_o[17] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1130),
    .D(_02547_),
    .Q_N(_11557_),
    .Q(\top_ihp.oisc.wb_dat_o[18] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1130),
    .D(_02548_),
    .Q_N(_11556_),
    .Q(\top_ihp.oisc.wb_dat_o[19] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1131),
    .D(_02549_),
    .Q_N(_00223_),
    .Q(\top_ihp.oisc.wb_dat_o[1] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1133),
    .D(_02550_),
    .Q_N(_11555_),
    .Q(\top_ihp.oisc.wb_dat_o[20] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1130),
    .D(_02551_),
    .Q_N(_11554_),
    .Q(\top_ihp.oisc.wb_dat_o[21] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1132),
    .D(_02552_),
    .Q_N(_11553_),
    .Q(\top_ihp.oisc.wb_dat_o[22] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1134),
    .D(_02553_),
    .Q_N(_11552_),
    .Q(\top_ihp.oisc.wb_dat_o[23] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1133),
    .D(_02554_),
    .Q_N(_11551_),
    .Q(\top_ihp.oisc.wb_dat_o[24] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1133),
    .D(_02555_),
    .Q_N(_11550_),
    .Q(\top_ihp.oisc.wb_dat_o[25] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1123),
    .D(_02556_),
    .Q_N(_11549_),
    .Q(\top_ihp.oisc.wb_dat_o[26] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1130),
    .D(_02557_),
    .Q_N(_11548_),
    .Q(\top_ihp.oisc.wb_dat_o[27] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1134),
    .D(_02558_),
    .Q_N(_11547_),
    .Q(\top_ihp.oisc.wb_dat_o[28] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1132),
    .D(_02559_),
    .Q_N(_11546_),
    .Q(\top_ihp.oisc.wb_dat_o[29] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1123),
    .D(_02560_),
    .Q_N(_00224_),
    .Q(\top_ihp.oisc.wb_dat_o[2] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1129),
    .D(_02561_),
    .Q_N(_11545_),
    .Q(\top_ihp.oisc.wb_dat_o[30] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1123),
    .D(_02562_),
    .Q_N(_11544_),
    .Q(\top_ihp.oisc.wb_dat_o[31] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1131),
    .D(_02563_),
    .Q_N(_00225_),
    .Q(\top_ihp.oisc.wb_dat_o[3] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1131),
    .D(_02564_),
    .Q_N(_00226_),
    .Q(\top_ihp.oisc.wb_dat_o[4] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1127),
    .D(_02565_),
    .Q_N(_00227_),
    .Q(\top_ihp.oisc.wb_dat_o[5] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1135),
    .D(_02566_),
    .Q_N(_00228_),
    .Q(\top_ihp.oisc.wb_dat_o[6] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_53_clk),
    .RESET_B(net1123),
    .D(_02567_),
    .Q_N(_00229_),
    .Q(\top_ihp.oisc.wb_dat_o[7] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_38_clk),
    .RESET_B(net1121),
    .D(_02568_),
    .Q_N(_11543_),
    .Q(\top_ihp.oisc.wb_dat_o[8] ));
 sg13g2_dfrbp_1 \top_ihp.oisc.wb_dat_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1134),
    .D(_02569_),
    .Q_N(_13627_),
    .Q(\top_ihp.oisc.wb_dat_o[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1129),
    .D(_00003_),
    .Q_N(_11542_),
    .Q(\top_ihp.wb_ack_coproc ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1089),
    .D(_02570_),
    .Q_N(_11541_),
    .Q(\top_ihp.wb_coproc.dat_o[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1079),
    .D(_02571_),
    .Q_N(_11540_),
    .Q(\top_ihp.wb_coproc.dat_o[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1087),
    .D(_02572_),
    .Q_N(_11539_),
    .Q(\top_ihp.wb_coproc.dat_o[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1078),
    .D(_02573_),
    .Q_N(_11538_),
    .Q(\top_ihp.wb_coproc.dat_o[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1095),
    .D(_02574_),
    .Q_N(_11537_),
    .Q(\top_ihp.wb_coproc.dat_o[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1087),
    .D(_02575_),
    .Q_N(_11536_),
    .Q(\top_ihp.wb_coproc.dat_o[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1079),
    .D(_02576_),
    .Q_N(_11535_),
    .Q(\top_ihp.wb_coproc.dat_o[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_46_clk),
    .RESET_B(net1085),
    .D(_02577_),
    .Q_N(_11534_),
    .Q(\top_ihp.wb_coproc.dat_o[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1087),
    .D(_02578_),
    .Q_N(_11533_),
    .Q(\top_ihp.wb_coproc.dat_o[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_50_clk),
    .RESET_B(net1089),
    .D(_02579_),
    .Q_N(_11532_),
    .Q(\top_ihp.wb_coproc.dat_o[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1095),
    .D(_02580_),
    .Q_N(_11531_),
    .Q(\top_ihp.wb_coproc.dat_o[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1095),
    .D(_02581_),
    .Q_N(_11530_),
    .Q(\top_ihp.wb_coproc.dat_o[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1095),
    .D(_02582_),
    .Q_N(_11529_),
    .Q(\top_ihp.wb_coproc.dat_o[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1096),
    .D(_02583_),
    .Q_N(_11528_),
    .Q(\top_ihp.wb_coproc.dat_o[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1095),
    .D(_02584_),
    .Q_N(_11527_),
    .Q(\top_ihp.wb_coproc.dat_o[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1097),
    .D(_02585_),
    .Q_N(_11526_),
    .Q(\top_ihp.wb_coproc.dat_o[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1097),
    .D(_02586_),
    .Q_N(_11525_),
    .Q(\top_ihp.wb_coproc.dat_o[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_69_clk),
    .RESET_B(net1130),
    .D(_02587_),
    .Q_N(_11524_),
    .Q(\top_ihp.wb_coproc.dat_o[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1130),
    .D(_02588_),
    .Q_N(_11523_),
    .Q(\top_ihp.wb_coproc.dat_o[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1130),
    .D(_02589_),
    .Q_N(_11522_),
    .Q(\top_ihp.wb_coproc.dat_o[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1092),
    .D(_02590_),
    .Q_N(_11521_),
    .Q(\top_ihp.wb_coproc.dat_o[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1097),
    .D(_02591_),
    .Q_N(_11520_),
    .Q(\top_ihp.wb_coproc.dat_o[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1087),
    .D(_02592_),
    .Q_N(_11519_),
    .Q(\top_ihp.wb_coproc.dat_o[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1092),
    .D(_02593_),
    .Q_N(_11518_),
    .Q(\top_ihp.wb_coproc.dat_o[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1098),
    .D(_02594_),
    .Q_N(_11517_),
    .Q(\top_ihp.wb_coproc.dat_o[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1089),
    .D(_02595_),
    .Q_N(_11516_),
    .Q(\top_ihp.wb_coproc.dat_o[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1089),
    .D(_02596_),
    .Q_N(_11515_),
    .Q(\top_ihp.wb_coproc.dat_o[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1095),
    .D(_02597_),
    .Q_N(_11514_),
    .Q(\top_ihp.wb_coproc.dat_o[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1095),
    .D(_02598_),
    .Q_N(_11513_),
    .Q(\top_ihp.wb_coproc.dat_o[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1095),
    .D(_02599_),
    .Q_N(_11512_),
    .Q(\top_ihp.wb_coproc.dat_o[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1096),
    .D(_02600_),
    .Q_N(_11511_),
    .Q(\top_ihp.wb_coproc.dat_o[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.dat_o[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_52_clk),
    .RESET_B(net1127),
    .D(_02601_),
    .Q_N(_11510_),
    .Q(\top_ihp.wb_coproc.dat_o[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1075),
    .D(_02602_),
    .Q_N(_11509_),
    .Q(\top_ihp.wb_coproc.opa[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1075),
    .D(_02603_),
    .Q_N(_00191_),
    .Q(\top_ihp.wb_coproc.opa[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1075),
    .D(_02604_),
    .Q_N(_00192_),
    .Q(\top_ihp.wb_coproc.opa[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1075),
    .D(_02605_),
    .Q_N(_00193_),
    .Q(\top_ihp.wb_coproc.opa[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1080),
    .D(_02606_),
    .Q_N(_00194_),
    .Q(\top_ihp.wb_coproc.opa[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1077),
    .D(_02607_),
    .Q_N(_00195_),
    .Q(\top_ihp.wb_coproc.opa[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1076),
    .D(_02608_),
    .Q_N(_00196_),
    .Q(\top_ihp.wb_coproc.opa[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1078),
    .D(_02609_),
    .Q_N(_00197_),
    .Q(\top_ihp.wb_coproc.opa[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1076),
    .D(_02610_),
    .Q_N(_00198_),
    .Q(\top_ihp.wb_coproc.opa[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1078),
    .D(_02611_),
    .Q_N(_00199_),
    .Q(\top_ihp.wb_coproc.opa[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1094),
    .D(_02612_),
    .Q_N(_00200_),
    .Q(\top_ihp.wb_coproc.opa[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1077),
    .D(_02613_),
    .Q_N(_00211_),
    .Q(\top_ihp.wb_coproc.opa[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1082),
    .D(_02614_),
    .Q_N(_00201_),
    .Q(\top_ihp.wb_coproc.opa[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1082),
    .D(_02615_),
    .Q_N(_00202_),
    .Q(\top_ihp.wb_coproc.opa[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1082),
    .D(_02616_),
    .Q_N(_00203_),
    .Q(\top_ihp.wb_coproc.opa[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1082),
    .D(_02617_),
    .Q_N(_00204_),
    .Q(\top_ihp.wb_coproc.opa[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1082),
    .D(_02618_),
    .Q_N(_00205_),
    .Q(\top_ihp.wb_coproc.opa[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1093),
    .D(_02619_),
    .Q_N(_00206_),
    .Q(\top_ihp.wb_coproc.opa[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1092),
    .D(_02620_),
    .Q_N(_00207_),
    .Q(\top_ihp.wb_coproc.opa[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1093),
    .D(_02621_),
    .Q_N(_00208_),
    .Q(\top_ihp.wb_coproc.opa[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1080),
    .D(_02622_),
    .Q_N(_00209_),
    .Q(\top_ihp.wb_coproc.opa[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1080),
    .D(_02623_),
    .Q_N(_00210_),
    .Q(\top_ihp.wb_coproc.opa[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1077),
    .D(_02624_),
    .Q_N(_00183_),
    .Q(\top_ihp.wb_coproc.opa[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1080),
    .D(_02625_),
    .Q_N(_11508_),
    .Q(\top_ihp.wb_coproc.opa[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1082),
    .D(_02626_),
    .Q_N(_11507_),
    .Q(\top_ihp.wb_coproc.opa[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1077),
    .D(_02627_),
    .Q_N(_00184_),
    .Q(\top_ihp.wb_coproc.opa[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1079),
    .D(_02628_),
    .Q_N(_00185_),
    .Q(\top_ihp.wb_coproc.opa[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1080),
    .D(_02629_),
    .Q_N(_00186_),
    .Q(\top_ihp.wb_coproc.opa[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1080),
    .D(_02630_),
    .Q_N(_00187_),
    .Q(\top_ihp.wb_coproc.opa[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_56_clk),
    .RESET_B(net1082),
    .D(_02631_),
    .Q_N(_00188_),
    .Q(\top_ihp.wb_coproc.opa[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_49_clk),
    .RESET_B(net1087),
    .D(_02632_),
    .Q_N(_00189_),
    .Q(\top_ihp.wb_coproc.opa[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opa[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1087),
    .D(_02633_),
    .Q_N(_00190_),
    .Q(\top_ihp.wb_coproc.opa[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1080),
    .D(_02634_),
    .Q_N(_11506_),
    .Q(\top_ihp.wb_coproc.opb[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1076),
    .D(_02635_),
    .Q_N(_11505_),
    .Q(\top_ihp.wb_coproc.opb[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1075),
    .D(_02636_),
    .Q_N(_11504_),
    .Q(\top_ihp.wb_coproc.opb[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1076),
    .D(_02637_),
    .Q_N(_11503_),
    .Q(\top_ihp.wb_coproc.opb[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1094),
    .D(_02638_),
    .Q_N(_11502_),
    .Q(\top_ihp.wb_coproc.opb[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1077),
    .D(_02639_),
    .Q_N(_11501_),
    .Q(\top_ihp.wb_coproc.opb[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_45_clk),
    .RESET_B(net1076),
    .D(_02640_),
    .Q_N(_11500_),
    .Q(\top_ihp.wb_coproc.opb[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1078),
    .D(_02641_),
    .Q_N(_11499_),
    .Q(\top_ihp.wb_coproc.opb[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1069),
    .D(_02642_),
    .Q_N(_11498_),
    .Q(\top_ihp.wb_coproc.opb[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1078),
    .D(_02643_),
    .Q_N(_11497_),
    .Q(\top_ihp.wb_coproc.opb[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1091),
    .D(_02644_),
    .Q_N(_11496_),
    .Q(\top_ihp.wb_coproc.opb[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1081),
    .D(_02645_),
    .Q_N(_11495_),
    .Q(\top_ihp.wb_coproc.opb[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_59_clk),
    .RESET_B(net1083),
    .D(_02646_),
    .Q_N(_11494_),
    .Q(\top_ihp.wb_coproc.opb[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1092),
    .D(_02647_),
    .Q_N(_11493_),
    .Q(\top_ihp.wb_coproc.opb[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1092),
    .D(_02648_),
    .Q_N(_11492_),
    .Q(\top_ihp.wb_coproc.opb[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1083),
    .D(_02649_),
    .Q_N(_11491_),
    .Q(\top_ihp.wb_coproc.opb[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1092),
    .D(_02650_),
    .Q_N(_11490_),
    .Q(\top_ihp.wb_coproc.opb[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1097),
    .D(_02651_),
    .Q_N(_11489_),
    .Q(\top_ihp.wb_coproc.opb[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1094),
    .D(_02652_),
    .Q_N(_11488_),
    .Q(\top_ihp.wb_coproc.opb[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1093),
    .D(_02653_),
    .Q_N(_11487_),
    .Q(\top_ihp.wb_coproc.opb[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1081),
    .D(_02654_),
    .Q_N(_11486_),
    .Q(\top_ihp.wb_coproc.opb[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1081),
    .D(_02655_),
    .Q_N(_11485_),
    .Q(\top_ihp.wb_coproc.opb[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1080),
    .D(_02656_),
    .Q_N(_00182_),
    .Q(\top_ihp.wb_coproc.opb[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1081),
    .D(_02657_),
    .Q_N(_11484_),
    .Q(\top_ihp.wb_coproc.opb[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_58_clk),
    .RESET_B(net1092),
    .D(_02658_),
    .Q_N(_11483_),
    .Q(\top_ihp.wb_coproc.opb[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1082),
    .D(_02659_),
    .Q_N(_00181_),
    .Q(\top_ihp.wb_coproc.opb[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1079),
    .D(_02660_),
    .Q_N(_00180_),
    .Q(\top_ihp.wb_coproc.opb[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_55_clk),
    .RESET_B(net1094),
    .D(_02661_),
    .Q_N(_11482_),
    .Q(\top_ihp.wb_coproc.opb[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_47_clk),
    .RESET_B(net1079),
    .D(_02662_),
    .Q_N(_11481_),
    .Q(\top_ihp.wb_coproc.opb[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_57_clk),
    .RESET_B(net1094),
    .D(_02663_),
    .Q_N(_11480_),
    .Q(\top_ihp.wb_coproc.opb[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1094),
    .D(_02664_),
    .Q_N(_11479_),
    .Q(\top_ihp.wb_coproc.opb[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_coproc.opb[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_48_clk),
    .RESET_B(net1091),
    .D(_02665_),
    .Q_N(_11478_),
    .Q(\top_ihp.wb_coproc.opb[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1984),
    .D(_02666_),
    .Q_N(_00264_),
    .Q(\top_ihp.wb_emem.bit_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1985),
    .D(_02667_),
    .Q_N(_11477_),
    .Q(\top_ihp.wb_emem.bit_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1986),
    .D(_02668_),
    .Q_N(_11476_),
    .Q(\top_ihp.wb_emem.bit_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1987),
    .D(_02669_),
    .Q_N(_11475_),
    .Q(\top_ihp.wb_emem.bit_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1988),
    .D(_02670_),
    .Q_N(_11474_),
    .Q(\top_ihp.wb_emem.bit_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1989),
    .D(_02671_),
    .Q_N(_11473_),
    .Q(\top_ihp.wb_emem.bit_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1990),
    .D(_02672_),
    .Q_N(_11472_),
    .Q(\top_ihp.wb_emem.bit_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1991),
    .D(_02673_),
    .Q_N(_11471_),
    .Q(\top_ihp.wb_emem.bit_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[0]$_DFFE_NN0P_  (.CLK(net2122),
    .RESET_B(net1119),
    .D(_02674_),
    .Q_N(_00160_),
    .Q(\top_ihp.wb_dati_ram[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[10]$_DFFE_NN0P_  (.CLK(net2121),
    .RESET_B(net1088),
    .D(_02675_),
    .Q_N(_00127_),
    .Q(\top_ihp.wb_dati_ram[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[11]$_DFFE_NN0P_  (.CLK(net2120),
    .RESET_B(net1123),
    .D(_02676_),
    .Q_N(_00130_),
    .Q(\top_ihp.wb_dati_ram[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[12]$_DFFE_NN0P_  (.CLK(net2119),
    .RESET_B(net1125),
    .D(_02677_),
    .Q_N(_00148_),
    .Q(\top_ihp.wb_dati_ram[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[13]$_DFFE_NN0P_  (.CLK(net2118),
    .RESET_B(net1125),
    .D(_02678_),
    .Q_N(_00151_),
    .Q(\top_ihp.wb_dati_ram[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[14]$_DFFE_NN0P_  (.CLK(net2117),
    .RESET_B(net1121),
    .D(_02679_),
    .Q_N(_00154_),
    .Q(\top_ihp.wb_dati_ram[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[15]$_DFFE_NN0P_  (.CLK(net2116),
    .RESET_B(net1121),
    .D(_02680_),
    .Q_N(_00157_),
    .Q(\top_ihp.wb_dati_ram[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[16]$_DFFE_NN0P_  (.CLK(net2115),
    .RESET_B(net1121),
    .D(_02681_),
    .Q_N(_00136_),
    .Q(\top_ihp.wb_dati_ram[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[17]$_DFFE_NN0P_  (.CLK(net2114),
    .RESET_B(net1121),
    .D(_02682_),
    .Q_N(_00139_),
    .Q(\top_ihp.wb_dati_ram[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[18]$_DFFE_NN0P_  (.CLK(net2113),
    .RESET_B(net1121),
    .D(_02683_),
    .Q_N(_00142_),
    .Q(\top_ihp.wb_dati_ram[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[19]$_DFFE_NN0P_  (.CLK(net2112),
    .RESET_B(net1121),
    .D(_02684_),
    .Q_N(_00145_),
    .Q(\top_ihp.wb_dati_ram[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[1]$_DFFE_NN0P_  (.CLK(net2111),
    .RESET_B(net1121),
    .D(_02685_),
    .Q_N(_00163_),
    .Q(\top_ihp.wb_dati_ram[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[20]$_DFFE_NN0P_  (.CLK(net2110),
    .RESET_B(net1129),
    .D(_02686_),
    .Q_N(_00082_),
    .Q(\top_ihp.wb_dati_ram[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[21]$_DFFE_NN0P_  (.CLK(net2109),
    .RESET_B(net1127),
    .D(_02687_),
    .Q_N(_00088_),
    .Q(\top_ihp.wb_dati_ram[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[22]$_DFFE_NN0P_  (.CLK(net2108),
    .RESET_B(net1129),
    .D(_02688_),
    .Q_N(_00085_),
    .Q(\top_ihp.wb_dati_ram[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[23]$_DFFE_NN0P_  (.CLK(net2107),
    .RESET_B(net1088),
    .D(_02689_),
    .Q_N(_00118_),
    .Q(\top_ihp.wb_dati_ram[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[24]$_DFFE_NN0P_  (.CLK(net2106),
    .RESET_B(net1118),
    .D(_02690_),
    .Q_N(_11470_),
    .Q(\top_ihp.wb_dati_ram[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[25]$_DFFE_NN0P_  (.CLK(net2105),
    .RESET_B(net1119),
    .D(_02691_),
    .Q_N(_00231_),
    .Q(\top_ihp.wb_dati_ram[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[26]$_DFFE_NN0P_  (.CLK(net2104),
    .RESET_B(net1119),
    .D(_02692_),
    .Q_N(_00100_),
    .Q(\top_ihp.wb_dati_ram[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[27]$_DFFE_NN0P_  (.CLK(net2103),
    .RESET_B(net1119),
    .D(_02693_),
    .Q_N(_00106_),
    .Q(\top_ihp.wb_dati_ram[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[28]$_DFFE_NN0P_  (.CLK(net2102),
    .RESET_B(net1119),
    .D(_02694_),
    .Q_N(_00103_),
    .Q(\top_ihp.wb_dati_ram[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[29]$_DFFE_NN0P_  (.CLK(net2101),
    .RESET_B(net1119),
    .D(_02695_),
    .Q_N(_00109_),
    .Q(\top_ihp.wb_dati_ram[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[2]$_DFFE_NN0P_  (.CLK(net2100),
    .RESET_B(net1119),
    .D(_02696_),
    .Q_N(_00166_),
    .Q(\top_ihp.wb_dati_ram[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[30]$_DFFE_NN0P_  (.CLK(net2099),
    .RESET_B(net1089),
    .D(_02697_),
    .Q_N(_00112_),
    .Q(\top_ihp.wb_dati_ram[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[31]$_DFFE_NN0P_  (.CLK(net2098),
    .RESET_B(net1090),
    .D(_02698_),
    .Q_N(_00133_),
    .Q(\top_ihp.wb_dati_ram[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[32]$_DFFE_NN0P_  (.CLK(net2097),
    .RESET_B(net1088),
    .D(_02699_),
    .Q_N(_11469_),
    .Q(\top_ihp.wb_emem.cmd[32] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[33]$_DFFE_NN0P_  (.CLK(net2096),
    .RESET_B(net1088),
    .D(_02700_),
    .Q_N(_11468_),
    .Q(\top_ihp.wb_emem.cmd[33] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[34]$_DFFE_NN0P_  (.CLK(net2095),
    .RESET_B(net1090),
    .D(_02701_),
    .Q_N(_11467_),
    .Q(\top_ihp.wb_emem.cmd[34] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[35]$_DFFE_NN0P_  (.CLK(net2094),
    .RESET_B(net1085),
    .D(_02702_),
    .Q_N(_11466_),
    .Q(\top_ihp.wb_emem.cmd[35] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[36]$_DFFE_NN0P_  (.CLK(net2093),
    .RESET_B(net1085),
    .D(_02703_),
    .Q_N(_11465_),
    .Q(\top_ihp.wb_emem.cmd[36] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[37]$_DFFE_NN0P_  (.CLK(net2092),
    .RESET_B(net1085),
    .D(_02704_),
    .Q_N(_11464_),
    .Q(\top_ihp.wb_emem.cmd[37] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[38]$_DFFE_NN0P_  (.CLK(net2091),
    .RESET_B(net1071),
    .D(_02705_),
    .Q_N(_11463_),
    .Q(\top_ihp.wb_emem.cmd[38] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[39]$_DFFE_NN0P_  (.CLK(net2090),
    .RESET_B(net1071),
    .D(_02706_),
    .Q_N(_11462_),
    .Q(\top_ihp.wb_emem.cmd[39] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[3]$_DFFE_NN0P_  (.CLK(net2089),
    .RESET_B(net1089),
    .D(_02707_),
    .Q_N(_00169_),
    .Q(\top_ihp.wb_dati_ram[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[40]$_DFFE_NN0P_  (.CLK(net2088),
    .RESET_B(net1071),
    .D(_02708_),
    .Q_N(_11461_),
    .Q(\top_ihp.wb_emem.cmd[40] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[41]$_DFFE_NN0P_  (.CLK(net2087),
    .RESET_B(net1071),
    .D(_02709_),
    .Q_N(_11460_),
    .Q(\top_ihp.wb_emem.cmd[41] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[42]$_DFFE_NN0P_  (.CLK(net2086),
    .RESET_B(net1071),
    .D(_02710_),
    .Q_N(_11459_),
    .Q(\top_ihp.wb_emem.cmd[42] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[43]$_DFFE_NN0P_  (.CLK(net2085),
    .RESET_B(net1072),
    .D(_02711_),
    .Q_N(_11458_),
    .Q(\top_ihp.wb_emem.cmd[43] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[44]$_DFFE_NN0P_  (.CLK(net2084),
    .RESET_B(net1072),
    .D(_02712_),
    .Q_N(_11457_),
    .Q(\top_ihp.wb_emem.cmd[44] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[45]$_DFFE_NN0P_  (.CLK(net2083),
    .RESET_B(net1072),
    .D(_02713_),
    .Q_N(_11456_),
    .Q(\top_ihp.wb_emem.cmd[45] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[46]$_DFFE_NN0P_  (.CLK(net2082),
    .RESET_B(net1071),
    .D(_02714_),
    .Q_N(_11455_),
    .Q(\top_ihp.wb_emem.cmd[46] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[47]$_DFFE_NN0P_  (.CLK(net2081),
    .RESET_B(net1086),
    .D(_02715_),
    .Q_N(_11454_),
    .Q(\top_ihp.wb_emem.cmd[47] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[48]$_DFFE_NN1P_  (.CLK(net2080),
    .RESET_B(net1088),
    .D(_02716_),
    .Q_N(\top_ihp.wb_emem.cmd[48] ),
    .Q(_00340_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[49]$_DFFE_NN0P_  (.CLK(net2079),
    .RESET_B(net1088),
    .D(_02717_),
    .Q_N(_11453_),
    .Q(\top_ihp.wb_emem.cmd[49] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[4]$_DFFE_NN0P_  (.CLK(net2078),
    .RESET_B(net1096),
    .D(_02718_),
    .Q_N(_00172_),
    .Q(\top_ihp.wb_dati_ram[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[50]$_DFFE_NN0P_  (.CLK(net2077),
    .RESET_B(net1088),
    .D(_02719_),
    .Q_N(_11452_),
    .Q(\top_ihp.wb_emem.cmd[50] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[51]$_DFFE_NN1P_  (.CLK(net2076),
    .RESET_B(net1088),
    .D(_02720_),
    .Q_N(\top_ihp.wb_emem.cmd[51] ),
    .Q(_00341_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[52]$_DFFE_NN1P_  (.CLK(net2075),
    .RESET_B(net1086),
    .D(_02721_),
    .Q_N(\top_ihp.wb_emem.cmd[52] ),
    .Q(_00342_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[53]$_DFFE_NN0P_  (.CLK(net2074),
    .RESET_B(net1086),
    .D(_02722_),
    .Q_N(_11451_),
    .Q(\top_ihp.wb_emem.cmd[53] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[54]$_DFFE_NN0P_  (.CLK(net2073),
    .RESET_B(net1086),
    .D(_02723_),
    .Q_N(_11450_),
    .Q(\top_ihp.wb_emem.cmd[54] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[55]$_DFFE_NN1P_  (.CLK(net2072),
    .RESET_B(net1086),
    .D(_02724_),
    .Q_N(\top_ihp.wb_emem.cmd[55] ),
    .Q(_00343_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[56]$_DFFE_NN0P_  (.CLK(net2071),
    .RESET_B(net1085),
    .D(_02725_),
    .Q_N(_11449_),
    .Q(\top_ihp.wb_emem.cmd[56] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[57]$_DFFE_NN1P_  (.CLK(net2070),
    .RESET_B(net1078),
    .D(_02726_),
    .Q_N(\top_ihp.wb_emem.cmd[57] ),
    .Q(_00344_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[58]$_DFFE_NN1P_  (.CLK(net2069),
    .RESET_B(net1069),
    .D(_02727_),
    .Q_N(\top_ihp.wb_emem.cmd[58] ),
    .Q(_00345_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[59]$_DFFE_NN0P_  (.CLK(net2068),
    .RESET_B(net1071),
    .D(_02728_),
    .Q_N(_11448_),
    .Q(\top_ihp.wb_emem.cmd[59] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[5]$_DFFE_NN0P_  (.CLK(net2067),
    .RESET_B(net1096),
    .D(_02729_),
    .Q_N(_00175_),
    .Q(\top_ihp.wb_dati_ram[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[60]$_DFFE_NN0P_  (.CLK(net2066),
    .RESET_B(net1069),
    .D(_02730_),
    .Q_N(_11447_),
    .Q(\top_ihp.wb_emem.cmd[60] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[61]$_DFFE_NN1P_  (.CLK(net2065),
    .RESET_B(net1070),
    .D(_02731_),
    .Q_N(\top_ihp.wb_emem.cmd[61] ),
    .Q(_00346_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[62]$_DFFE_NN1P_  (.CLK(net2064),
    .RESET_B(net1070),
    .D(_02732_),
    .Q_N(\top_ihp.wb_emem.cmd[62] ),
    .Q(_00347_));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[63]$_DFFE_NN0P_  (.CLK(net2063),
    .RESET_B(net1085),
    .D(_02733_),
    .Q_N(_11446_),
    .Q(\top_ihp.wb_emem.cmd[63] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[6]$_DFFE_NN0P_  (.CLK(net2062),
    .RESET_B(net1089),
    .D(_02734_),
    .Q_N(_00115_),
    .Q(\top_ihp.wb_dati_ram[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[7]$_DFFE_NN0P_  (.CLK(net2061),
    .RESET_B(net1090),
    .D(_02735_),
    .Q_N(_00178_),
    .Q(\top_ihp.wb_dati_ram[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[8]$_DFFE_NN0P_  (.CLK(net2060),
    .RESET_B(net1072),
    .D(_02736_),
    .Q_N(_00121_),
    .Q(\top_ihp.wb_dati_ram[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.cmd[9]$_DFFE_NN0P_  (.CLK(net2059),
    .RESET_B(net1073),
    .D(_02737_),
    .Q_N(_00124_),
    .Q(\top_ihp.wb_dati_ram[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_bit$_DFFE_PP_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1992),
    .D(_02738_),
    .Q_N(_11445_),
    .Q(\top_ihp.wb_emem.last_bit ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.last_wait$_DFFE_PP_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net1993),
    .D(_02739_),
    .Q_N(_11444_),
    .Q(\top_ihp.wb_emem.last_wait ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P_  (.CLK(net2058),
    .RESET_B(net1994),
    .D(_02740_),
    .Q_N(_11443_),
    .Q(\top_ihp.wb_emem.nbits[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P_  (.CLK(net2057),
    .RESET_B(net1995),
    .D(_02741_),
    .Q_N(_11442_),
    .Q(\top_ihp.wb_emem.nbits[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P_  (.CLK(net2056),
    .RESET_B(net1996),
    .D(_02742_),
    .Q_N(_11441_),
    .Q(\top_ihp.wb_emem.nbits[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P_  (.CLK(net2055),
    .RESET_B(net1997),
    .D(_02743_),
    .Q_N(_11440_),
    .Q(\top_ihp.wb_emem.nbits[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[0]$_DFFE_NN0P_  (.CLK(net2054),
    .RESET_B(net1073),
    .D(_02744_),
    .Q_N(_11439_),
    .Q(\top_ihp.wb_emem.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[1]$_DFFE_NN0P_  (.CLK(net2053),
    .RESET_B(net1072),
    .D(_02745_),
    .Q_N(_11438_),
    .Q(\top_ihp.wb_emem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[2]$_DFFE_NN0P_  (.CLK(net2052),
    .RESET_B(net1073),
    .D(_02746_),
    .Q_N(_11437_),
    .Q(\top_ihp.wb_emem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.state[3]$_DFFE_NN0P_  (.CLK(net2051),
    .RESET_B(net1071),
    .D(_02747_),
    .Q_N(\top_ihp.ram_cs_o ),
    .Q(\top_ihp.wb_emem.state[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1998),
    .D(_02748_),
    .Q_N(_00265_),
    .Q(\top_ihp.wb_emem.wait_counter[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_221_clk),
    .RESET_B(net1999),
    .D(_02749_),
    .Q_N(_11436_),
    .Q(\top_ihp.wb_emem.wait_counter[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2000),
    .D(_02750_),
    .Q_N(_11435_),
    .Q(\top_ihp.wb_emem.wait_counter[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2001),
    .D(_02751_),
    .Q_N(_11434_),
    .Q(\top_ihp.wb_emem.wait_counter[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_222_clk),
    .RESET_B(net2002),
    .D(_02752_),
    .Q_N(_11433_),
    .Q(\top_ihp.wb_emem.wait_counter[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2003),
    .D(_02753_),
    .Q_N(_11432_),
    .Q(\top_ihp.wb_emem.wait_counter[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2004),
    .D(_02754_),
    .Q_N(_11431_),
    .Q(\top_ihp.wb_emem.wait_counter[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P_  (.CLK(clknet_leaf_223_clk),
    .RESET_B(net2005),
    .D(_02755_),
    .Q_N(_13628_),
    .Q(\top_ihp.wb_emem.wait_counter[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1118),
    .D(_00004_),
    .Q_N(_00094_),
    .Q(\top_ihp.wb_ack_gpio ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.dat_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_40_clk),
    .RESET_B(net1118),
    .D(_02756_),
    .Q_N(_11430_),
    .Q(\top_ihp.wb_dati_gpio[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1098),
    .D(_02757_),
    .Q_N(_11429_),
    .Q(\top_ihp.gpio_o_1 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[1]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1097),
    .D(_02758_),
    .Q_N(\top_ihp.gpio_o_2 ),
    .Q(_00348_));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1098),
    .D(_02759_),
    .Q_N(_11428_),
    .Q(\top_ihp.gpio_o_3 ));
 sg13g2_dfrbp_1 \top_ihp.wb_gpio.data_o[3]$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1098),
    .D(_02760_),
    .Q_N(\top_ihp.gpio_o_4 ),
    .Q(_00349_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[0]$_DFFE_NN0P_  (.CLK(net2050),
    .RESET_B(net1106),
    .D(_02761_),
    .Q_N(_11427_),
    .Q(\top_ihp.wb_imem.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[1]$_DFFE_NN0P_  (.CLK(net2049),
    .RESET_B(net1107),
    .D(_02762_),
    .Q_N(_11426_),
    .Q(\top_ihp.wb_imem.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[2]$_DFFE_NN0P_  (.CLK(net2048),
    .RESET_B(net1106),
    .D(_02763_),
    .Q_N(_11425_),
    .Q(\top_ihp.wb_imem.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[3]$_DFFE_NN0P_  (.CLK(net2047),
    .RESET_B(net1101),
    .D(_02764_),
    .Q_N(_11424_),
    .Q(\top_ihp.wb_imem.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[4]$_DFFE_NN0P_  (.CLK(net2046),
    .RESET_B(net1102),
    .D(_02765_),
    .Q_N(_11423_),
    .Q(\top_ihp.wb_imem.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.bits_left[5]$_DFFE_NN0P_  (.CLK(net2045),
    .RESET_B(net1101),
    .D(_02766_),
    .Q_N(_11422_),
    .Q(\top_ihp.wb_imem.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[0]$_DFFE_NN0P_  (.CLK(net2044),
    .RESET_B(net1118),
    .D(_02767_),
    .Q_N(_00159_),
    .Q(\top_ihp.wb_dati_rom[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[10]$_DFFE_NN0P_  (.CLK(net2043),
    .RESET_B(net1107),
    .D(_02768_),
    .Q_N(_00126_),
    .Q(\top_ihp.wb_dati_rom[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[11]$_DFFE_NN0P_  (.CLK(net2042),
    .RESET_B(net1107),
    .D(_02769_),
    .Q_N(_00129_),
    .Q(\top_ihp.wb_dati_rom[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[12]$_DFFE_NN0P_  (.CLK(net2041),
    .RESET_B(net1107),
    .D(_02770_),
    .Q_N(_00147_),
    .Q(\top_ihp.wb_dati_rom[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[13]$_DFFE_NN0P_  (.CLK(net2040),
    .RESET_B(net1108),
    .D(_02771_),
    .Q_N(_00150_),
    .Q(\top_ihp.wb_dati_rom[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[14]$_DFFE_NN0P_  (.CLK(net2039),
    .RESET_B(net1108),
    .D(_02772_),
    .Q_N(_00153_),
    .Q(\top_ihp.wb_dati_rom[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[15]$_DFFE_NN0P_  (.CLK(net2038),
    .RESET_B(net1108),
    .D(_02773_),
    .Q_N(_00156_),
    .Q(\top_ihp.wb_dati_rom[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[16]$_DFFE_NN0P_  (.CLK(net2037),
    .RESET_B(net1120),
    .D(_02774_),
    .Q_N(_00135_),
    .Q(\top_ihp.wb_dati_rom[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[17]$_DFFE_NN0P_  (.CLK(net2036),
    .RESET_B(net1108),
    .D(_02775_),
    .Q_N(_00138_),
    .Q(\top_ihp.wb_dati_rom[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[18]$_DFFE_NN0P_  (.CLK(net2035),
    .RESET_B(net1129),
    .D(_02776_),
    .Q_N(_00141_),
    .Q(\top_ihp.wb_dati_rom[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[19]$_DFFE_NN0P_  (.CLK(net2034),
    .RESET_B(net1129),
    .D(_02777_),
    .Q_N(_00144_),
    .Q(\top_ihp.wb_dati_rom[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[1]$_DFFE_NN0P_  (.CLK(net2033),
    .RESET_B(net1120),
    .D(_02778_),
    .Q_N(_00162_),
    .Q(\top_ihp.wb_dati_rom[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[20]$_DFFE_NN0P_  (.CLK(net2032),
    .RESET_B(net1129),
    .D(_02779_),
    .Q_N(_00081_),
    .Q(\top_ihp.wb_dati_rom[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[21]$_DFFE_NN0P_  (.CLK(net2031),
    .RESET_B(net1136),
    .D(_02780_),
    .Q_N(_00087_),
    .Q(\top_ihp.wb_dati_rom[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[22]$_DFFE_NN0P_  (.CLK(net2030),
    .RESET_B(net1129),
    .D(_02781_),
    .Q_N(_00084_),
    .Q(\top_ihp.wb_dati_rom[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[23]$_DFFE_NN0P_  (.CLK(net2029),
    .RESET_B(net1120),
    .D(_02782_),
    .Q_N(_00117_),
    .Q(\top_ihp.wb_dati_rom[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[24]$_DFFE_NN0P_  (.CLK(net2028),
    .RESET_B(net1118),
    .D(_02783_),
    .Q_N(_11421_),
    .Q(\top_ihp.wb_dati_rom[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[25]$_DFFE_NN0P_  (.CLK(net2027),
    .RESET_B(net1118),
    .D(_02784_),
    .Q_N(_00230_),
    .Q(\top_ihp.wb_dati_rom[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[26]$_DFFE_NN0P_  (.CLK(net2026),
    .RESET_B(net1106),
    .D(_02785_),
    .Q_N(_00099_),
    .Q(\top_ihp.wb_dati_rom[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[27]$_DFFE_NN0P_  (.CLK(net2025),
    .RESET_B(net1106),
    .D(_02786_),
    .Q_N(_00105_),
    .Q(\top_ihp.wb_dati_rom[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[28]$_DFFE_NN0P_  (.CLK(net2024),
    .RESET_B(net1106),
    .D(_02787_),
    .Q_N(_00102_),
    .Q(\top_ihp.wb_dati_rom[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[29]$_DFFE_NN0P_  (.CLK(net2023),
    .RESET_B(net1107),
    .D(_02788_),
    .Q_N(_00108_),
    .Q(\top_ihp.wb_dati_rom[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[2]$_DFFE_NN0P_  (.CLK(net2022),
    .RESET_B(net1120),
    .D(_02789_),
    .Q_N(_00165_),
    .Q(\top_ihp.wb_dati_rom[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[30]$_DFFE_NN0P_  (.CLK(net2021),
    .RESET_B(net1106),
    .D(_02790_),
    .Q_N(_00111_),
    .Q(\top_ihp.wb_dati_rom[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[31]$_DFFE_NN0P_  (.CLK(net2020),
    .RESET_B(net1106),
    .D(_02791_),
    .Q_N(_00132_),
    .Q(\top_ihp.wb_dati_rom[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[3]$_DFFE_NN0P_  (.CLK(net2019),
    .RESET_B(net1120),
    .D(_02792_),
    .Q_N(_00168_),
    .Q(\top_ihp.wb_dati_rom[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[4]$_DFFE_NN0P_  (.CLK(net2018),
    .RESET_B(net1120),
    .D(_02793_),
    .Q_N(_00171_),
    .Q(\top_ihp.wb_dati_rom[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[5]$_DFFE_NN0P_  (.CLK(net2017),
    .RESET_B(net1120),
    .D(_02794_),
    .Q_N(_00174_),
    .Q(\top_ihp.wb_dati_rom[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[6]$_DFFE_NN0P_  (.CLK(net2016),
    .RESET_B(net1120),
    .D(_02795_),
    .Q_N(_00114_),
    .Q(\top_ihp.wb_dati_rom[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[7]$_DFFE_NN0P_  (.CLK(net2015),
    .RESET_B(net1109),
    .D(_02796_),
    .Q_N(_00177_),
    .Q(\top_ihp.wb_dati_rom[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[8]$_DFFE_NN0P_  (.CLK(net2014),
    .RESET_B(net1107),
    .D(_02797_),
    .Q_N(_00120_),
    .Q(\top_ihp.wb_dati_rom[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.cmd[9]$_DFFE_NN0P_  (.CLK(net2013),
    .RESET_B(net1107),
    .D(_02798_),
    .Q_N(_00123_),
    .Q(\top_ihp.wb_dati_rom[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.spi_cs_o$_DFFE_NN1P_  (.CLK(net2012),
    .RESET_B(net1097),
    .D(_02799_),
    .Q_N(\top_ihp.rom_cs_o ),
    .Q(_00350_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[0]$_DFF_NN1_  (.CLK(net2011),
    .RESET_B(net1118),
    .D(_00355_),
    .Q_N(\top_ihp.wb_imem.state[0] ),
    .Q(_13700_));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[1]$_DFF_NN0_  (.CLK(net2010),
    .RESET_B(net1108),
    .D(_00000_),
    .Q_N(_00095_),
    .Q(\top_ihp.wb_imem.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_imem.state[2]$_DFF_NN0_  (.CLK(net2009),
    .RESET_B(net1118),
    .D(_00001_),
    .Q_N(_13629_),
    .Q(\top_ihp.wb_imem.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.ack_o$_DFF_PN0_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1131),
    .D(_13703_),
    .Q_N(_11420_),
    .Q(\top_ihp.wb_ack_spi ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1133),
    .D(_02800_),
    .Q_N(_11419_),
    .Q(\top_ihp.wb_spi.bits_left[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1133),
    .D(_02801_),
    .Q_N(_11418_),
    .Q(\top_ihp.wb_spi.bits_left[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1133),
    .D(_02802_),
    .Q_N(_11417_),
    .Q(\top_ihp.wb_spi.bits_left[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1131),
    .D(_02803_),
    .Q_N(_11416_),
    .Q(\top_ihp.wb_spi.bits_left[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_66_clk),
    .RESET_B(net1132),
    .D(_02804_),
    .Q_N(_11415_),
    .Q(\top_ihp.wb_spi.bits_left[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.bits_left[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1131),
    .D(_02805_),
    .Q_N(_11414_),
    .Q(\top_ihp.wb_spi.bits_left[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1124),
    .D(_02806_),
    .Q_N(_11413_),
    .Q(\top_ihp.wb_dati_spi[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[10]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1126),
    .D(_02807_),
    .Q_N(_00143_),
    .Q(\top_ihp.wb_dati_spi[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[11]$_DFFE_PN0P_  (.CLK(clknet_leaf_65_clk),
    .RESET_B(net1126),
    .D(_02808_),
    .Q_N(_00146_),
    .Q(\top_ihp.wb_dati_spi[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[12]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1131),
    .D(_02809_),
    .Q_N(_00083_),
    .Q(\top_ihp.wb_dati_spi[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[13]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1126),
    .D(_02810_),
    .Q_N(_00089_),
    .Q(\top_ihp.wb_dati_spi[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[14]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1126),
    .D(_02811_),
    .Q_N(_00086_),
    .Q(\top_ihp.wb_dati_spi[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[15]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1126),
    .D(_02812_),
    .Q_N(_00119_),
    .Q(\top_ihp.wb_dati_spi[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[16]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1098),
    .D(_02813_),
    .Q_N(_00122_),
    .Q(\top_ihp.wb_dati_spi[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[17]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1098),
    .D(_02814_),
    .Q_N(_00125_),
    .Q(\top_ihp.wb_dati_spi[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[18]$_DFFE_PN0P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1098),
    .D(_02815_),
    .Q_N(_00128_),
    .Q(\top_ihp.wb_dati_spi[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[19]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1124),
    .D(_02816_),
    .Q_N(_00131_),
    .Q(\top_ihp.wb_dati_spi[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1124),
    .D(_02817_),
    .Q_N(_00232_),
    .Q(\top_ihp.wb_dati_spi[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[20]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1124),
    .D(_02818_),
    .Q_N(_00149_),
    .Q(\top_ihp.wb_dati_spi[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[21]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1124),
    .D(_02819_),
    .Q_N(_00152_),
    .Q(\top_ihp.wb_dati_spi[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[22]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1126),
    .D(_02820_),
    .Q_N(_00155_),
    .Q(\top_ihp.wb_dati_spi[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[23]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1126),
    .D(_02821_),
    .Q_N(_00158_),
    .Q(\top_ihp.wb_dati_spi[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[24]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1128),
    .D(_02822_),
    .Q_N(_00161_),
    .Q(\top_ihp.wb_dati_spi[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[25]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1127),
    .D(_02823_),
    .Q_N(_00164_),
    .Q(\top_ihp.wb_dati_spi[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[26]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1131),
    .D(_02824_),
    .Q_N(_00167_),
    .Q(\top_ihp.wb_dati_spi[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[27]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1130),
    .D(_02825_),
    .Q_N(_00170_),
    .Q(\top_ihp.wb_dati_spi[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[28]$_DFFE_PN0P_  (.CLK(clknet_leaf_68_clk),
    .RESET_B(net1127),
    .D(_02826_),
    .Q_N(_00173_),
    .Q(\top_ihp.wb_dati_spi[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[29]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1127),
    .D(_02827_),
    .Q_N(_00176_),
    .Q(\top_ihp.wb_dati_spi[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_64_clk),
    .RESET_B(net1124),
    .D(_02828_),
    .Q_N(_00101_),
    .Q(\top_ihp.wb_dati_spi[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[30]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1127),
    .D(_02829_),
    .Q_N(_00116_),
    .Q(\top_ihp.wb_dati_spi[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[31]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1096),
    .D(_02830_),
    .Q_N(_00179_),
    .Q(\top_ihp.wb_dati_spi[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1124),
    .D(_02831_),
    .Q_N(_00107_),
    .Q(\top_ihp.wb_dati_spi[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1124),
    .D(_02832_),
    .Q_N(_00104_),
    .Q(\top_ihp.wb_dati_spi[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1123),
    .D(_02833_),
    .Q_N(_00110_),
    .Q(\top_ihp.wb_dati_spi[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_54_clk),
    .RESET_B(net1123),
    .D(_02834_),
    .Q_N(_00113_),
    .Q(\top_ihp.wb_dati_spi[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1123),
    .D(_02835_),
    .Q_N(_00134_),
    .Q(\top_ihp.wb_dati_spi[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[8]$_DFFE_PN0P_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1125),
    .D(_02836_),
    .Q_N(_00137_),
    .Q(\top_ihp.wb_dati_spi[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.cmd[9]$_DFFE_PN0P_  (.CLK(clknet_leaf_63_clk),
    .RESET_B(net1126),
    .D(_02837_),
    .Q_N(_00140_),
    .Q(\top_ihp.wb_dati_spi[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[0]$_DFF_NN0_  (.CLK(net2008),
    .RESET_B(net1097),
    .D(_11386_),
    .Q_N(_11386_),
    .Q(\top_ihp.wb_spi.spi_clk_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_clk_cnt[1]$_DFF_NN0_  (.CLK(net2007),
    .RESET_B(net1097),
    .D(_00266_),
    .Q_N(_11412_),
    .Q(\top_ihp.spi_clk_o ));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_1$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1092),
    .D(_02838_),
    .Q_N(\top_ihp.spi_cs_o_1 ),
    .Q(_00351_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_2$_DFFE_PN1P_  (.CLK(clknet_leaf_62_clk),
    .RESET_B(net1093),
    .D(_02839_),
    .Q_N(\top_ihp.spi_cs_o_2 ),
    .Q(_00352_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.spi_cs_o_3$_DFFE_PN1P_  (.CLK(clknet_leaf_61_clk),
    .RESET_B(net1093),
    .D(_02840_),
    .Q_N(\top_ihp.spi_cs_o_3 ),
    .Q(_00353_));
 sg13g2_dfrbp_1 \top_ihp.wb_spi.state$_DFF_PN0_  (.CLK(clknet_leaf_67_clk),
    .RESET_B(net1132),
    .D(_13704_),
    .Q_N(_00096_),
    .Q(\top_ihp.wb_spi.state ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net2006),
    .D(_02841_),
    .Q_N(_00080_),
    .Q(\top_ihp.wb_ack_uart ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1069),
    .D(_02842_),
    .Q_N(_11411_),
    .Q(\top_ihp.wb_uart.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.state[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1069),
    .D(_02843_),
    .Q_N(_11410_),
    .Q(\top_ihp.wb_uart.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1070),
    .D(_02844_),
    .Q_N(_00220_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1070),
    .D(_02845_),
    .Q_N(_11409_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1070),
    .D(_02846_),
    .Q_N(_11408_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1070),
    .D(_02847_),
    .Q_N(_13630_),
    .Q(\top_ihp.wb_uart.uart_rx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1420),
    .D(_00005_),
    .Q_N(_13631_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1419),
    .D(_00006_),
    .Q_N(_13632_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1415),
    .D(_00007_),
    .Q_N(_13633_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_172_clk),
    .RESET_B(net1415),
    .D(_00008_),
    .Q_N(_13634_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1415),
    .D(_00009_),
    .Q_N(_13635_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1416),
    .D(_00010_),
    .Q_N(_13636_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_159_clk),
    .RESET_B(net1415),
    .D(_00011_),
    .Q_N(_13637_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1416),
    .D(_00012_),
    .Q_N(_13638_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1416),
    .D(_00013_),
    .Q_N(_13639_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1417),
    .D(_00014_),
    .Q_N(_13640_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1417),
    .D(_00015_),
    .Q_N(_13641_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1420),
    .D(_00016_),
    .Q_N(_13642_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1417),
    .D(_00017_),
    .Q_N(_13643_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1417),
    .D(_00018_),
    .Q_N(_13644_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1416),
    .D(_00019_),
    .Q_N(_13645_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1416),
    .D(_00020_),
    .Q_N(_13646_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_155_clk),
    .RESET_B(net1416),
    .D(_00021_),
    .Q_N(_13647_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1416),
    .D(_00022_),
    .Q_N(_13648_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_156_clk),
    .RESET_B(net1416),
    .D(_00023_),
    .Q_N(_13649_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1415),
    .D(_00024_),
    .Q_N(_13650_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1415),
    .D(_00025_),
    .Q_N(_13651_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_160_clk),
    .RESET_B(net1418),
    .D(_00026_),
    .Q_N(_13652_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1420),
    .D(_00027_),
    .Q_N(_13653_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1415),
    .D(_00028_),
    .Q_N(_13654_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_161_clk),
    .RESET_B(net1415),
    .D(_00029_),
    .Q_N(_13655_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_217_clk),
    .RESET_B(net1420),
    .D(_00030_),
    .Q_N(_13656_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1419),
    .D(_00031_),
    .Q_N(_13657_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_179_clk),
    .RESET_B(net1419),
    .D(_00032_),
    .Q_N(_00097_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1419),
    .D(_00033_),
    .Q_N(_13658_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_178_clk),
    .RESET_B(net1419),
    .D(_00034_),
    .Q_N(_13659_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_177_clk),
    .RESET_B(net1419),
    .D(_00035_),
    .Q_N(_13660_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_173_clk),
    .RESET_B(net1419),
    .D(_00036_),
    .Q_N(_11407_),
    .Q(\top_ihp.wb_uart.uart_rx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1072),
    .D(_02848_),
    .Q_N(_11406_),
    .Q(\top_ihp.wb_dati_uart[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1072),
    .D(_02849_),
    .Q_N(_11405_),
    .Q(\top_ihp.wb_dati_uart[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1074),
    .D(_02850_),
    .Q_N(_11404_),
    .Q(\top_ihp.wb_dati_uart[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net1072),
    .D(_02851_),
    .Q_N(_11403_),
    .Q(\top_ihp.wb_dati_uart[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net1074),
    .D(_02852_),
    .Q_N(_11402_),
    .Q(\top_ihp.wb_dati_uart[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1101),
    .D(_02853_),
    .Q_N(_11401_),
    .Q(\top_ihp.wb_dati_uart[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net1101),
    .D(_02854_),
    .Q_N(_11400_),
    .Q(\top_ihp.wb_dati_uart[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net1106),
    .D(_02855_),
    .Q_N(_11399_),
    .Q(\top_ihp.wb_dati_uart[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.rx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1066),
    .D(_02856_),
    .Q_N(_13661_),
    .Q(\top_ihp.wb_uart.rx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1069),
    .D(\top_ihp.wb_uart.uart_rx.next_state[0] ),
    .Q_N(_13662_),
    .Q(\top_ihp.wb_uart.uart_rx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1069),
    .D(\top_ihp.wb_uart.uart_rx.next_state[1] ),
    .Q_N(_13663_),
    .Q(\top_ihp.wb_uart.uart_rx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_rx.state[2]$_DFF_PN0_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net1070),
    .D(\top_ihp.wb_uart.uart_rx.next_state[2] ),
    .Q_N(_00098_),
    .Q(\top_ihp.wb_uart.uart_rx.state[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1066),
    .D(_02857_),
    .Q_N(_11398_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1066),
    .D(_02858_),
    .Q_N(_11397_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1066),
    .D(_02859_),
    .Q_N(_00221_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.bit_cnt[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1066),
    .D(_02860_),
    .Q_N(_13664_),
    .Q(\top_ihp.wb_uart.uart_tx.bit_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[0]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1063),
    .D(_00037_),
    .Q_N(_13665_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[10]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00038_),
    .Q_N(_13666_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[10] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[11]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00039_),
    .Q_N(_13667_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[11] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[12]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00040_),
    .Q_N(_13668_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[12] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[13]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1062),
    .D(_00041_),
    .Q_N(_13669_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[13] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[14]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1062),
    .D(_00042_),
    .Q_N(_13670_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[14] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[15]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1062),
    .D(_00043_),
    .Q_N(_13671_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[15] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[16]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1062),
    .D(_00044_),
    .Q_N(_13672_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[16] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[17]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1063),
    .D(_00045_),
    .Q_N(_13673_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[17] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[18]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1063),
    .D(_00046_),
    .Q_N(_13674_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[18] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[19]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1063),
    .D(_00047_),
    .Q_N(_13675_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[19] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[1]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1063),
    .D(_00048_),
    .Q_N(_13676_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[20]$_DFF_PN0_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net1064),
    .D(_00049_),
    .Q_N(_13677_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[20] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[21]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1065),
    .D(_00050_),
    .Q_N(_13678_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[21] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[22]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1065),
    .D(_00051_),
    .Q_N(_13679_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[22] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[23]$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00052_),
    .Q_N(_13680_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[23] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[24]$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00053_),
    .Q_N(_13681_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[24] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[25]$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00054_),
    .Q_N(_13682_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[25] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[26]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1065),
    .D(_00055_),
    .Q_N(_13683_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[26] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[27]$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00056_),
    .Q_N(_13684_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[27] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[28]$_DFF_PN0_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net1065),
    .D(_00057_),
    .Q_N(_13685_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[28] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[29]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1068),
    .D(_00058_),
    .Q_N(_13686_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[29] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[2]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1063),
    .D(_00059_),
    .Q_N(_13687_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[30]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1068),
    .D(_00060_),
    .Q_N(_13688_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[30] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[31]$_DFF_PN0_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net1068),
    .D(_00061_),
    .Q_N(_13689_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[31] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[3]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1061),
    .D(_00062_),
    .Q_N(_13690_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[4]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1063),
    .D(_00063_),
    .Q_N(_13691_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[5]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1063),
    .D(_00064_),
    .Q_N(_13692_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[6]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00065_),
    .Q_N(_13693_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[7]$_DFF_PN0_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net1061),
    .D(_00066_),
    .Q_N(_13694_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[8]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00067_),
    .Q_N(_13695_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[8] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.cycle_cnt[9]$_DFF_PN0_  (.CLK(clknet_leaf_326_clk),
    .RESET_B(net1061),
    .D(_00068_),
    .Q_N(_13696_),
    .Q(\top_ihp.wb_uart.uart_tx.cycle_cnt[9] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[0]$_DFF_PN0_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1066),
    .D(\top_ihp.wb_uart.uart_tx.next_state[0] ),
    .Q_N(_13697_),
    .Q(\top_ihp.wb_uart.uart_tx.state[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.state[1]$_DFF_PN0_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1067),
    .D(\top_ihp.wb_uart.uart_tx.next_state[1] ),
    .Q_N(_11396_),
    .Q(\top_ihp.wb_uart.uart_tx.state[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[0]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1075),
    .D(_02861_),
    .Q_N(_11395_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[0] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[1]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1066),
    .D(_02862_),
    .Q_N(_11394_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[1] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[2]$_DFFE_PN0P_  (.CLK(clknet_leaf_43_clk),
    .RESET_B(net1075),
    .D(_02863_),
    .Q_N(_11393_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[2] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[3]$_DFFE_PN0P_  (.CLK(clknet_leaf_44_clk),
    .RESET_B(net1075),
    .D(_02864_),
    .Q_N(_11392_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[3] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[4]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1069),
    .D(_02865_),
    .Q_N(_11391_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[4] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[5]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1067),
    .D(_02866_),
    .Q_N(_11390_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[5] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[6]$_DFFE_PN0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net1066),
    .D(_02867_),
    .Q_N(_11389_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[6] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_latch[7]$_DFFE_PN0P_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net1067),
    .D(_02868_),
    .Q_N(_11388_),
    .Q(\top_ihp.wb_uart.uart_tx.tx_data_latch[7] ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_data_ready$_DFFE_PN0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net1067),
    .D(_02869_),
    .Q_N(_11387_),
    .Q(\top_ihp.wb_uart.tx_ready ));
 sg13g2_dfrbp_1 \top_ihp.wb_uart.uart_tx.tx_reg$_DFF_PN1_  (.CLK(clknet_leaf_60_clk),
    .RESET_B(net1081),
    .D(_00356_),
    .Q_N(\top_ihp.tx ),
    .Q(_13701_));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[1]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[2]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[3]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[5]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uio_out[0]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uio_out[1]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uio_out[2]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uio_out[3]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uio_out[4]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uio_out[5]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uio_out[6]));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uio_out[7]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[0]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[1]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[2]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[3]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[4]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[5]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[6]));
 sg13g2_buf_1 output25 (.A(net25),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout26 (.A(_02978_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_02937_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_11149_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_10974_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_10460_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_10450_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_06559_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_05946_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_05623_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_03312_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_03262_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_03019_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_02976_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_02924_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_11303_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_11225_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_11222_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_11220_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_11219_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_11192_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_11155_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_11147_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_11102_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_10991_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_10917_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_10888_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_10855_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_10813_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_10688_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_10649_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_10600_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_10568_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_10509_),
    .X(net58));
 sg13g2_buf_4 fanout59 (.X(net59),
    .A(_10429_));
 sg13g2_buf_2 fanout60 (.A(_10274_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_10090_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_10051_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_10010_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_09889_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_06403_),
    .X(net65));
 sg13g2_buf_4 fanout66 (.X(net66),
    .A(_06383_));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_06334_));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_06294_));
 sg13g2_buf_4 fanout69 (.X(net69),
    .A(_06235_));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_06233_));
 sg13g2_buf_4 fanout71 (.X(net71),
    .A(_05980_));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_05786_));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_05749_));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_05739_));
 sg13g2_buf_2 fanout75 (.A(_05668_),
    .X(net75));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_05659_));
 sg13g2_buf_2 fanout77 (.A(_05652_),
    .X(net77));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_05637_));
 sg13g2_buf_2 fanout79 (.A(_03310_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_03275_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_03266_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_03264_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_03258_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_03254_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_03250_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_03244_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_03074_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_02946_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_02939_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_02932_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_02929_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_02927_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_02921_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_02917_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_02915_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_02913_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_11296_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_11293_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_11291_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_11290_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_11284_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_11262_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_11256_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_11221_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_11203_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_11151_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_11122_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_11115_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_11109_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_11107_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_11104_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_11098_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_11094_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_11091_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_11089_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_10941_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_10940_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_10932_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_10845_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_10834_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_10804_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_10779_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_10776_));
 sg13g2_buf_2 fanout124 (.A(_10773_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_10745_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_10742_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_10740_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_10739_),
    .X(net128));
 sg13g2_buf_4 fanout129 (.X(net129),
    .A(_10738_));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(_10704_));
 sg13g2_buf_2 fanout131 (.A(_10687_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_10648_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_10626_),
    .X(net133));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(_10599_));
 sg13g2_buf_2 fanout135 (.A(_10567_),
    .X(net135));
 sg13g2_buf_2 fanout136 (.A(_10500_),
    .X(net136));
 sg13g2_buf_2 fanout137 (.A(_10362_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_10343_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_10319_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_10206_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_10089_),
    .X(net141));
 sg13g2_buf_4 fanout142 (.X(net142),
    .A(_10009_));
 sg13g2_buf_2 fanout143 (.A(_09888_),
    .X(net143));
 sg13g2_buf_2 fanout144 (.A(_08912_),
    .X(net144));
 sg13g2_buf_2 fanout145 (.A(_08884_),
    .X(net145));
 sg13g2_buf_2 fanout146 (.A(_08863_),
    .X(net146));
 sg13g2_buf_2 fanout147 (.A(_08780_),
    .X(net147));
 sg13g2_buf_2 fanout148 (.A(_08753_),
    .X(net148));
 sg13g2_buf_2 fanout149 (.A(_08732_),
    .X(net149));
 sg13g2_buf_2 fanout150 (.A(_06506_),
    .X(net150));
 sg13g2_buf_2 fanout151 (.A(_06354_),
    .X(net151));
 sg13g2_buf_4 fanout152 (.X(net152),
    .A(_06308_));
 sg13g2_buf_4 fanout153 (.X(net153),
    .A(_06148_));
 sg13g2_buf_4 fanout154 (.X(net154),
    .A(_06117_));
 sg13g2_buf_4 fanout155 (.X(net155),
    .A(_06035_));
 sg13g2_buf_4 fanout156 (.X(net156),
    .A(_05978_));
 sg13g2_buf_2 fanout157 (.A(_05970_),
    .X(net157));
 sg13g2_buf_4 fanout158 (.X(net158),
    .A(_05948_));
 sg13g2_buf_2 fanout159 (.A(_05945_),
    .X(net159));
 sg13g2_buf_2 fanout160 (.A(_05922_),
    .X(net160));
 sg13g2_buf_4 fanout161 (.X(net161),
    .A(_05909_));
 sg13g2_buf_4 fanout162 (.X(net162),
    .A(_05831_));
 sg13g2_buf_2 fanout163 (.A(_05829_),
    .X(net163));
 sg13g2_buf_4 fanout164 (.X(net164),
    .A(_05818_));
 sg13g2_buf_2 fanout165 (.A(_05795_),
    .X(net165));
 sg13g2_buf_2 fanout166 (.A(_05789_),
    .X(net166));
 sg13g2_buf_2 fanout167 (.A(_05784_),
    .X(net167));
 sg13g2_buf_2 fanout168 (.A(_05778_),
    .X(net168));
 sg13g2_buf_4 fanout169 (.X(net169),
    .A(_05771_));
 sg13g2_buf_4 fanout170 (.X(net170),
    .A(_05768_));
 sg13g2_buf_2 fanout171 (.A(_05767_),
    .X(net171));
 sg13g2_buf_2 fanout172 (.A(_05761_),
    .X(net172));
 sg13g2_buf_4 fanout173 (.X(net173),
    .A(_05748_));
 sg13g2_buf_2 fanout174 (.A(_05747_),
    .X(net174));
 sg13g2_buf_2 fanout175 (.A(_05732_),
    .X(net175));
 sg13g2_buf_4 fanout176 (.X(net176),
    .A(_05717_));
 sg13g2_buf_2 fanout177 (.A(_05712_),
    .X(net177));
 sg13g2_buf_4 fanout178 (.X(net178),
    .A(_05669_));
 sg13g2_buf_4 fanout179 (.X(net179),
    .A(_05666_));
 sg13g2_buf_4 fanout180 (.X(net180),
    .A(_05661_));
 sg13g2_buf_4 fanout181 (.X(net181),
    .A(_05658_));
 sg13g2_buf_2 fanout182 (.A(_05651_),
    .X(net182));
 sg13g2_buf_4 fanout183 (.X(net183),
    .A(_05649_));
 sg13g2_buf_4 fanout184 (.X(net184),
    .A(_05642_));
 sg13g2_buf_4 fanout185 (.X(net185),
    .A(_05636_));
 sg13g2_buf_4 fanout186 (.X(net186),
    .A(_05634_));
 sg13g2_buf_4 fanout187 (.X(net187),
    .A(_05632_));
 sg13g2_buf_4 fanout188 (.X(net188),
    .A(_05630_));
 sg13g2_buf_4 fanout189 (.X(net189),
    .A(_05628_));
 sg13g2_buf_4 fanout190 (.X(net190),
    .A(_05626_));
 sg13g2_buf_2 fanout191 (.A(_05486_),
    .X(net191));
 sg13g2_buf_4 fanout192 (.X(net192),
    .A(_05472_));
 sg13g2_buf_4 fanout193 (.X(net193),
    .A(_05466_));
 sg13g2_buf_2 fanout194 (.A(_05338_),
    .X(net194));
 sg13g2_buf_2 fanout195 (.A(_05328_),
    .X(net195));
 sg13g2_buf_4 fanout196 (.X(net196),
    .A(_04310_));
 sg13g2_buf_4 fanout197 (.X(net197),
    .A(_04309_));
 sg13g2_buf_4 fanout198 (.X(net198),
    .A(_04308_));
 sg13g2_buf_4 fanout199 (.X(net199),
    .A(_04305_));
 sg13g2_buf_4 fanout200 (.X(net200),
    .A(_04304_));
 sg13g2_buf_4 fanout201 (.X(net201),
    .A(_04303_));
 sg13g2_buf_4 fanout202 (.X(net202),
    .A(_04178_));
 sg13g2_buf_4 fanout203 (.X(net203),
    .A(_04087_));
 sg13g2_buf_4 fanout204 (.X(net204),
    .A(_03920_));
 sg13g2_buf_2 fanout205 (.A(_03283_),
    .X(net205));
 sg13g2_buf_2 fanout206 (.A(_03271_),
    .X(net206));
 sg13g2_buf_2 fanout207 (.A(_03268_),
    .X(net207));
 sg13g2_buf_2 fanout208 (.A(_03256_),
    .X(net208));
 sg13g2_buf_2 fanout209 (.A(_03127_),
    .X(net209));
 sg13g2_buf_2 fanout210 (.A(_02944_),
    .X(net210));
 sg13g2_buf_2 fanout211 (.A(_02935_),
    .X(net211));
 sg13g2_buf_2 fanout212 (.A(_02919_),
    .X(net212));
 sg13g2_buf_2 fanout213 (.A(_11380_),
    .X(net213));
 sg13g2_buf_2 fanout214 (.A(_11368_),
    .X(net214));
 sg13g2_buf_2 fanout215 (.A(_11364_),
    .X(net215));
 sg13g2_buf_4 fanout216 (.X(net216),
    .A(_11361_));
 sg13g2_buf_2 fanout217 (.A(_11342_),
    .X(net217));
 sg13g2_buf_2 fanout218 (.A(_11340_),
    .X(net218));
 sg13g2_buf_2 fanout219 (.A(_11330_),
    .X(net219));
 sg13g2_buf_4 fanout220 (.X(net220),
    .A(_11329_));
 sg13g2_buf_2 fanout221 (.A(_11314_),
    .X(net221));
 sg13g2_buf_2 fanout222 (.A(_11311_),
    .X(net222));
 sg13g2_buf_2 fanout223 (.A(_11301_),
    .X(net223));
 sg13g2_buf_2 fanout224 (.A(_11300_),
    .X(net224));
 sg13g2_buf_4 fanout225 (.X(net225),
    .A(_11299_));
 sg13g2_buf_2 fanout226 (.A(_11292_),
    .X(net226));
 sg13g2_buf_2 fanout227 (.A(_11275_),
    .X(net227));
 sg13g2_buf_2 fanout228 (.A(_11272_),
    .X(net228));
 sg13g2_buf_2 fanout229 (.A(_11268_),
    .X(net229));
 sg13g2_buf_2 fanout230 (.A(_11267_),
    .X(net230));
 sg13g2_buf_4 fanout231 (.X(net231),
    .A(_11261_));
 sg13g2_buf_2 fanout232 (.A(_11211_),
    .X(net232));
 sg13g2_buf_2 fanout233 (.A(_11165_),
    .X(net233));
 sg13g2_buf_2 fanout234 (.A(_11120_),
    .X(net234));
 sg13g2_buf_2 fanout235 (.A(_11112_),
    .X(net235));
 sg13g2_buf_2 fanout236 (.A(_11096_),
    .X(net236));
 sg13g2_buf_2 fanout237 (.A(_11066_),
    .X(net237));
 sg13g2_buf_2 fanout238 (.A(_11065_),
    .X(net238));
 sg13g2_buf_2 fanout239 (.A(_11054_),
    .X(net239));
 sg13g2_buf_2 fanout240 (.A(_11053_),
    .X(net240));
 sg13g2_buf_4 fanout241 (.X(net241),
    .A(_11050_));
 sg13g2_buf_2 fanout242 (.A(_11033_),
    .X(net242));
 sg13g2_buf_2 fanout243 (.A(_11031_),
    .X(net243));
 sg13g2_buf_2 fanout244 (.A(_11022_),
    .X(net244));
 sg13g2_buf_2 fanout245 (.A(_11021_),
    .X(net245));
 sg13g2_buf_4 fanout246 (.X(net246),
    .A(_11020_));
 sg13g2_buf_2 fanout247 (.A(_11005_),
    .X(net247));
 sg13g2_buf_2 fanout248 (.A(_11002_),
    .X(net248));
 sg13g2_buf_2 fanout249 (.A(_10993_),
    .X(net249));
 sg13g2_buf_2 fanout250 (.A(_10992_),
    .X(net250));
 sg13g2_buf_4 fanout251 (.X(net251),
    .A(_10990_));
 sg13g2_buf_2 fanout252 (.A(_10965_),
    .X(net252));
 sg13g2_buf_2 fanout253 (.A(_10953_),
    .X(net253));
 sg13g2_buf_2 fanout254 (.A(_10931_),
    .X(net254));
 sg13g2_buf_4 fanout255 (.X(net255),
    .A(_10819_));
 sg13g2_buf_2 fanout256 (.A(_10812_),
    .X(net256));
 sg13g2_buf_4 fanout257 (.X(net257),
    .A(_10808_));
 sg13g2_buf_2 fanout258 (.A(_10807_),
    .X(net258));
 sg13g2_buf_2 fanout259 (.A(_10801_),
    .X(net259));
 sg13g2_buf_2 fanout260 (.A(_10797_),
    .X(net260));
 sg13g2_buf_2 fanout261 (.A(_10796_),
    .X(net261));
 sg13g2_buf_2 fanout262 (.A(_10772_),
    .X(net262));
 sg13g2_buf_2 fanout263 (.A(_10765_),
    .X(net263));
 sg13g2_buf_2 fanout264 (.A(_10741_),
    .X(net264));
 sg13g2_buf_2 fanout265 (.A(_10737_),
    .X(net265));
 sg13g2_buf_2 fanout266 (.A(_10674_),
    .X(net266));
 sg13g2_buf_2 fanout267 (.A(_10625_),
    .X(net267));
 sg13g2_buf_2 fanout268 (.A(_10533_),
    .X(net268));
 sg13g2_buf_4 fanout269 (.X(net269),
    .A(_10467_));
 sg13g2_buf_2 fanout270 (.A(_10416_),
    .X(net270));
 sg13g2_buf_2 fanout271 (.A(_10393_),
    .X(net271));
 sg13g2_buf_2 fanout272 (.A(_10380_),
    .X(net272));
 sg13g2_buf_2 fanout273 (.A(_10361_),
    .X(net273));
 sg13g2_buf_4 fanout274 (.X(net274),
    .A(_10318_));
 sg13g2_buf_2 fanout275 (.A(_10246_),
    .X(net275));
 sg13g2_buf_2 fanout276 (.A(_10205_),
    .X(net276));
 sg13g2_buf_2 fanout277 (.A(_10159_),
    .X(net277));
 sg13g2_buf_2 fanout278 (.A(_10122_),
    .X(net278));
 sg13g2_buf_2 fanout279 (.A(_06287_),
    .X(net279));
 sg13g2_buf_2 fanout280 (.A(_06276_),
    .X(net280));
 sg13g2_buf_2 fanout281 (.A(_06256_),
    .X(net281));
 sg13g2_buf_4 fanout282 (.X(net282),
    .A(_06158_));
 sg13g2_buf_4 fanout283 (.X(net283),
    .A(_06138_));
 sg13g2_buf_4 fanout284 (.X(net284),
    .A(_06113_));
 sg13g2_buf_2 fanout285 (.A(_06108_),
    .X(net285));
 sg13g2_buf_4 fanout286 (.X(net286),
    .A(_06066_));
 sg13g2_buf_2 fanout287 (.A(_05975_),
    .X(net287));
 sg13g2_buf_4 fanout288 (.X(net288),
    .A(_05968_));
 sg13g2_buf_4 fanout289 (.X(net289),
    .A(_05926_));
 sg13g2_buf_2 fanout290 (.A(_05901_),
    .X(net290));
 sg13g2_buf_2 fanout291 (.A(_05892_),
    .X(net291));
 sg13g2_buf_2 fanout292 (.A(_05876_),
    .X(net292));
 sg13g2_buf_4 fanout293 (.X(net293),
    .A(_05861_));
 sg13g2_buf_2 fanout294 (.A(_05859_),
    .X(net294));
 sg13g2_buf_2 fanout295 (.A(_05828_),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_05821_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_05809_),
    .X(net297));
 sg13g2_buf_2 fanout298 (.A(_05796_),
    .X(net298));
 sg13g2_buf_2 fanout299 (.A(_05788_),
    .X(net299));
 sg13g2_buf_4 fanout300 (.X(net300),
    .A(_05782_));
 sg13g2_buf_4 fanout301 (.X(net301),
    .A(_05779_));
 sg13g2_buf_2 fanout302 (.A(_05774_),
    .X(net302));
 sg13g2_buf_4 fanout303 (.X(net303),
    .A(_05772_));
 sg13g2_buf_2 fanout304 (.A(_05762_),
    .X(net304));
 sg13g2_buf_4 fanout305 (.X(net305),
    .A(_05759_));
 sg13g2_buf_2 fanout306 (.A(_05758_),
    .X(net306));
 sg13g2_buf_2 fanout307 (.A(_05752_),
    .X(net307));
 sg13g2_buf_4 fanout308 (.X(net308),
    .A(_05751_));
 sg13g2_buf_4 fanout309 (.X(net309),
    .A(_05745_));
 sg13g2_buf_2 fanout310 (.A(_05744_),
    .X(net310));
 sg13g2_buf_4 fanout311 (.X(net311),
    .A(_05742_));
 sg13g2_buf_4 fanout312 (.X(net312),
    .A(_05730_));
 sg13g2_buf_2 fanout313 (.A(_05727_),
    .X(net313));
 sg13g2_buf_2 fanout314 (.A(_05723_),
    .X(net314));
 sg13g2_buf_4 fanout315 (.X(net315),
    .A(_05720_));
 sg13g2_buf_4 fanout316 (.X(net316),
    .A(_05715_));
 sg13g2_buf_2 fanout317 (.A(_05705_),
    .X(net317));
 sg13g2_buf_2 fanout318 (.A(_05688_),
    .X(net318));
 sg13g2_buf_4 fanout319 (.X(net319),
    .A(_05686_));
 sg13g2_buf_2 fanout320 (.A(_05681_),
    .X(net320));
 sg13g2_buf_4 fanout321 (.X(net321),
    .A(_05665_));
 sg13g2_buf_4 fanout322 (.X(net322),
    .A(_05663_));
 sg13g2_buf_4 fanout323 (.X(net323),
    .A(_05655_));
 sg13g2_buf_2 fanout324 (.A(_05648_),
    .X(net324));
 sg13g2_buf_4 fanout325 (.X(net325),
    .A(_05645_));
 sg13g2_buf_4 fanout326 (.X(net326),
    .A(_05641_));
 sg13g2_buf_2 fanout327 (.A(_05640_),
    .X(net327));
 sg13g2_buf_2 fanout328 (.A(_05633_),
    .X(net328));
 sg13g2_buf_2 fanout329 (.A(_05627_),
    .X(net329));
 sg13g2_buf_2 fanout330 (.A(_05616_),
    .X(net330));
 sg13g2_buf_2 fanout331 (.A(_05612_),
    .X(net331));
 sg13g2_buf_4 fanout332 (.X(net332),
    .A(_05501_));
 sg13g2_buf_2 fanout333 (.A(_05494_),
    .X(net333));
 sg13g2_buf_2 fanout334 (.A(_05485_),
    .X(net334));
 sg13g2_buf_2 fanout335 (.A(_05422_),
    .X(net335));
 sg13g2_buf_2 fanout336 (.A(_05403_),
    .X(net336));
 sg13g2_buf_2 fanout337 (.A(_05382_),
    .X(net337));
 sg13g2_buf_2 fanout338 (.A(_05327_),
    .X(net338));
 sg13g2_buf_2 fanout339 (.A(_05311_),
    .X(net339));
 sg13g2_buf_2 fanout340 (.A(_05130_),
    .X(net340));
 sg13g2_buf_2 fanout341 (.A(_03604_),
    .X(net341));
 sg13g2_buf_2 fanout342 (.A(_03592_),
    .X(net342));
 sg13g2_buf_2 fanout343 (.A(_03281_),
    .X(net343));
 sg13g2_buf_2 fanout344 (.A(_03163_),
    .X(net344));
 sg13g2_buf_2 fanout345 (.A(_03159_),
    .X(net345));
 sg13g2_buf_2 fanout346 (.A(_03158_),
    .X(net346));
 sg13g2_buf_4 fanout347 (.X(net347),
    .A(_03153_));
 sg13g2_buf_2 fanout348 (.A(_03125_),
    .X(net348));
 sg13g2_buf_2 fanout349 (.A(_03122_),
    .X(net349));
 sg13g2_buf_2 fanout350 (.A(_03060_),
    .X(net350));
 sg13g2_buf_2 fanout351 (.A(_03056_),
    .X(net351));
 sg13g2_buf_2 fanout352 (.A(_03055_),
    .X(net352));
 sg13g2_buf_2 fanout353 (.A(_03033_),
    .X(net353));
 sg13g2_buf_2 fanout354 (.A(_03030_),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(_03021_),
    .X(net355));
 sg13g2_buf_2 fanout356 (.A(_03020_),
    .X(net356));
 sg13g2_buf_4 fanout357 (.X(net357),
    .A(_03018_));
 sg13g2_buf_2 fanout358 (.A(_03000_),
    .X(net358));
 sg13g2_buf_2 fanout359 (.A(_02997_),
    .X(net359));
 sg13g2_buf_2 fanout360 (.A(_02988_),
    .X(net360));
 sg13g2_buf_2 fanout361 (.A(_02987_),
    .X(net361));
 sg13g2_buf_4 fanout362 (.X(net362),
    .A(_02986_));
 sg13g2_buf_2 fanout363 (.A(_02967_),
    .X(net363));
 sg13g2_buf_2 fanout364 (.A(_02965_),
    .X(net364));
 sg13g2_buf_2 fanout365 (.A(_02954_),
    .X(net365));
 sg13g2_buf_2 fanout366 (.A(_02953_),
    .X(net366));
 sg13g2_buf_4 fanout367 (.X(net367),
    .A(_02950_));
 sg13g2_buf_2 fanout368 (.A(_02930_),
    .X(net368));
 sg13g2_buf_2 fanout369 (.A(_02925_),
    .X(net369));
 sg13g2_buf_2 fanout370 (.A(_02910_),
    .X(net370));
 sg13g2_buf_2 fanout371 (.A(_02909_),
    .X(net371));
 sg13g2_buf_4 fanout372 (.X(net372),
    .A(_02908_));
 sg13g2_buf_2 fanout373 (.A(_02887_),
    .X(net373));
 sg13g2_buf_2 fanout374 (.A(_02884_),
    .X(net374));
 sg13g2_buf_2 fanout375 (.A(_02883_),
    .X(net375));
 sg13g2_buf_4 fanout376 (.X(net376),
    .A(_02878_));
 sg13g2_buf_2 fanout377 (.A(_11365_),
    .X(net377));
 sg13g2_buf_2 fanout378 (.A(_11363_),
    .X(net378));
 sg13g2_buf_2 fanout379 (.A(_11331_),
    .X(net379));
 sg13g2_buf_2 fanout380 (.A(_11328_),
    .X(net380));
 sg13g2_buf_2 fanout381 (.A(_11298_),
    .X(net381));
 sg13g2_buf_2 fanout382 (.A(_11281_),
    .X(net382));
 sg13g2_buf_2 fanout383 (.A(_11260_),
    .X(net383));
 sg13g2_buf_2 fanout384 (.A(_11237_),
    .X(net384));
 sg13g2_buf_2 fanout385 (.A(_11234_),
    .X(net385));
 sg13g2_buf_2 fanout386 (.A(_11233_),
    .X(net386));
 sg13g2_buf_2 fanout387 (.A(_11228_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(_11019_),
    .X(net388));
 sg13g2_buf_2 fanout389 (.A(_10989_),
    .X(net389));
 sg13g2_buf_2 fanout390 (.A(_10961_),
    .X(net390));
 sg13g2_buf_2 fanout391 (.A(_10954_),
    .X(net391));
 sg13g2_buf_2 fanout392 (.A(_10952_),
    .X(net392));
 sg13g2_buf_2 fanout393 (.A(_10925_),
    .X(net393));
 sg13g2_buf_2 fanout394 (.A(_10922_),
    .X(net394));
 sg13g2_buf_2 fanout395 (.A(_10921_),
    .X(net395));
 sg13g2_buf_4 fanout396 (.X(net396),
    .A(_10818_));
 sg13g2_buf_2 fanout397 (.A(_10810_),
    .X(net397));
 sg13g2_buf_2 fanout398 (.A(_10800_),
    .X(net398));
 sg13g2_buf_2 fanout399 (.A(_10798_),
    .X(net399));
 sg13g2_buf_2 fanout400 (.A(_10726_),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(_10662_),
    .X(net401));
 sg13g2_buf_4 fanout402 (.X(net402),
    .A(_10441_));
 sg13g2_buf_2 fanout403 (.A(_10415_),
    .X(net403));
 sg13g2_buf_2 fanout404 (.A(_10277_),
    .X(net404));
 sg13g2_buf_2 fanout405 (.A(_10275_),
    .X(net405));
 sg13g2_buf_2 fanout406 (.A(_10224_),
    .X(net406));
 sg13g2_buf_2 fanout407 (.A(_10171_),
    .X(net407));
 sg13g2_buf_2 fanout408 (.A(_10011_),
    .X(net408));
 sg13g2_buf_2 fanout409 (.A(_09944_),
    .X(net409));
 sg13g2_buf_2 fanout410 (.A(_06240_),
    .X(net410));
 sg13g2_buf_2 fanout411 (.A(_06070_),
    .X(net411));
 sg13g2_buf_4 fanout412 (.X(net412),
    .A(_06053_));
 sg13g2_buf_2 fanout413 (.A(_05998_),
    .X(net413));
 sg13g2_buf_2 fanout414 (.A(_05956_),
    .X(net414));
 sg13g2_buf_4 fanout415 (.X(net415),
    .A(_05931_));
 sg13g2_buf_2 fanout416 (.A(_05914_),
    .X(net416));
 sg13g2_buf_4 fanout417 (.X(net417),
    .A(_05890_));
 sg13g2_buf_4 fanout418 (.X(net418),
    .A(_05887_));
 sg13g2_buf_2 fanout419 (.A(_05878_),
    .X(net419));
 sg13g2_buf_2 fanout420 (.A(_05847_),
    .X(net420));
 sg13g2_buf_4 fanout421 (.X(net421),
    .A(_05799_));
 sg13g2_buf_4 fanout422 (.X(net422),
    .A(_05776_));
 sg13g2_buf_4 fanout423 (.X(net423),
    .A(_05734_));
 sg13g2_buf_2 fanout424 (.A(_05729_),
    .X(net424));
 sg13g2_buf_4 fanout425 (.X(net425),
    .A(_05725_));
 sg13g2_buf_2 fanout426 (.A(_05714_),
    .X(net426));
 sg13g2_buf_2 fanout427 (.A(_05709_),
    .X(net427));
 sg13g2_buf_2 fanout428 (.A(_05685_),
    .X(net428));
 sg13g2_buf_2 fanout429 (.A(_05683_),
    .X(net429));
 sg13g2_buf_4 fanout430 (.X(net430),
    .A(_05662_));
 sg13g2_buf_4 fanout431 (.X(net431),
    .A(_05654_));
 sg13g2_buf_2 fanout432 (.A(_05646_),
    .X(net432));
 sg13g2_buf_4 fanout433 (.X(net433),
    .A(_05644_));
 sg13g2_buf_2 fanout434 (.A(_05578_),
    .X(net434));
 sg13g2_buf_4 fanout435 (.X(net435),
    .A(_05520_));
 sg13g2_buf_4 fanout436 (.X(net436),
    .A(_05507_));
 sg13g2_buf_2 fanout437 (.A(_05504_),
    .X(net437));
 sg13g2_buf_2 fanout438 (.A(_05496_),
    .X(net438));
 sg13g2_buf_2 fanout439 (.A(_05489_),
    .X(net439));
 sg13g2_buf_4 fanout440 (.X(net440),
    .A(_05479_));
 sg13g2_buf_2 fanout441 (.A(_05460_),
    .X(net441));
 sg13g2_buf_2 fanout442 (.A(_05456_),
    .X(net442));
 sg13g2_buf_2 fanout443 (.A(_05454_),
    .X(net443));
 sg13g2_buf_4 fanout444 (.X(net444),
    .A(_05451_));
 sg13g2_buf_2 fanout445 (.A(_05437_),
    .X(net445));
 sg13g2_buf_4 fanout446 (.X(net446),
    .A(_05430_));
 sg13g2_buf_2 fanout447 (.A(_05415_),
    .X(net447));
 sg13g2_buf_2 fanout448 (.A(_05397_),
    .X(net448));
 sg13g2_buf_2 fanout449 (.A(_05390_),
    .X(net449));
 sg13g2_buf_4 fanout450 (.X(net450),
    .A(_05388_));
 sg13g2_buf_2 fanout451 (.A(_05384_),
    .X(net451));
 sg13g2_buf_4 fanout452 (.X(net452),
    .A(_05310_));
 sg13g2_buf_2 fanout453 (.A(_04982_),
    .X(net453));
 sg13g2_buf_2 fanout454 (.A(_04970_),
    .X(net454));
 sg13g2_buf_2 fanout455 (.A(_04930_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_04918_),
    .X(net456));
 sg13g2_buf_2 fanout457 (.A(_04877_),
    .X(net457));
 sg13g2_buf_2 fanout458 (.A(_04874_),
    .X(net458));
 sg13g2_buf_2 fanout459 (.A(_04869_),
    .X(net459));
 sg13g2_buf_2 fanout460 (.A(_04782_),
    .X(net460));
 sg13g2_buf_2 fanout461 (.A(_04734_),
    .X(net461));
 sg13g2_buf_2 fanout462 (.A(_03694_),
    .X(net462));
 sg13g2_buf_2 fanout463 (.A(_03691_),
    .X(net463));
 sg13g2_buf_2 fanout464 (.A(_03690_),
    .X(net464));
 sg13g2_buf_4 fanout465 (.X(net465),
    .A(_03685_));
 sg13g2_buf_2 fanout466 (.A(_03666_),
    .X(net466));
 sg13g2_buf_2 fanout467 (.A(_03664_),
    .X(net467));
 sg13g2_buf_2 fanout468 (.A(_03654_),
    .X(net468));
 sg13g2_buf_4 fanout469 (.X(net469),
    .A(_03653_));
 sg13g2_buf_2 fanout470 (.A(_03632_),
    .X(net470));
 sg13g2_buf_2 fanout471 (.A(_03629_),
    .X(net471));
 sg13g2_buf_2 fanout472 (.A(_03628_),
    .X(net472));
 sg13g2_buf_4 fanout473 (.X(net473),
    .A(_03623_));
 sg13g2_buf_2 fanout474 (.A(_03600_),
    .X(net474));
 sg13g2_buf_2 fanout475 (.A(_03593_),
    .X(net475));
 sg13g2_buf_2 fanout476 (.A(_03591_),
    .X(net476));
 sg13g2_buf_2 fanout477 (.A(_03575_),
    .X(net477));
 sg13g2_buf_2 fanout478 (.A(_03572_),
    .X(net478));
 sg13g2_buf_2 fanout479 (.A(_03563_),
    .X(net479));
 sg13g2_buf_2 fanout480 (.A(_03562_),
    .X(net480));
 sg13g2_buf_4 fanout481 (.X(net481),
    .A(_03561_));
 sg13g2_buf_2 fanout482 (.A(_03536_),
    .X(net482));
 sg13g2_buf_2 fanout483 (.A(_03533_),
    .X(net483));
 sg13g2_buf_2 fanout484 (.A(_03507_),
    .X(net484));
 sg13g2_buf_2 fanout485 (.A(_03504_),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_03503_),
    .X(net486));
 sg13g2_buf_4 fanout487 (.X(net487),
    .A(_03498_));
 sg13g2_buf_2 fanout488 (.A(_03483_),
    .X(net488));
 sg13g2_buf_2 fanout489 (.A(_03480_),
    .X(net489));
 sg13g2_buf_2 fanout490 (.A(_03471_),
    .X(net490));
 sg13g2_buf_2 fanout491 (.A(_03470_),
    .X(net491));
 sg13g2_buf_4 fanout492 (.X(net492),
    .A(_03469_));
 sg13g2_buf_2 fanout493 (.A(_03448_),
    .X(net493));
 sg13g2_buf_2 fanout494 (.A(_03445_),
    .X(net494));
 sg13g2_buf_2 fanout495 (.A(_03444_),
    .X(net495));
 sg13g2_buf_2 fanout496 (.A(_03425_),
    .X(net496));
 sg13g2_buf_2 fanout497 (.A(_03422_),
    .X(net497));
 sg13g2_buf_2 fanout498 (.A(_03413_),
    .X(net498));
 sg13g2_buf_2 fanout499 (.A(_03412_),
    .X(net499));
 sg13g2_buf_4 fanout500 (.X(net500),
    .A(_03411_));
 sg13g2_buf_2 fanout501 (.A(_03394_),
    .X(net501));
 sg13g2_buf_2 fanout502 (.A(_03392_),
    .X(net502));
 sg13g2_buf_2 fanout503 (.A(_03382_),
    .X(net503));
 sg13g2_buf_2 fanout504 (.A(_03381_),
    .X(net504));
 sg13g2_buf_2 fanout505 (.A(_03357_),
    .X(net505));
 sg13g2_buf_2 fanout506 (.A(_03354_),
    .X(net506));
 sg13g2_buf_2 fanout507 (.A(_03353_),
    .X(net507));
 sg13g2_buf_2 fanout508 (.A(_03348_),
    .X(net508));
 sg13g2_buf_2 fanout509 (.A(_03333_),
    .X(net509));
 sg13g2_buf_2 fanout510 (.A(_03330_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_03321_),
    .X(net511));
 sg13g2_buf_2 fanout512 (.A(_03320_),
    .X(net512));
 sg13g2_buf_4 fanout513 (.X(net513),
    .A(_03319_));
 sg13g2_buf_2 fanout514 (.A(_03303_),
    .X(net514));
 sg13g2_buf_2 fanout515 (.A(_03302_),
    .X(net515));
 sg13g2_buf_2 fanout516 (.A(_03291_),
    .X(net516));
 sg13g2_buf_2 fanout517 (.A(_03290_),
    .X(net517));
 sg13g2_buf_4 fanout518 (.X(net518),
    .A(_03287_));
 sg13g2_buf_2 fanout519 (.A(_03251_),
    .X(net519));
 sg13g2_buf_2 fanout520 (.A(_03247_),
    .X(net520));
 sg13g2_buf_2 fanout521 (.A(_03220_),
    .X(net521));
 sg13g2_buf_2 fanout522 (.A(_03217_),
    .X(net522));
 sg13g2_buf_2 fanout523 (.A(_03216_),
    .X(net523));
 sg13g2_buf_2 fanout524 (.A(_03211_),
    .X(net524));
 sg13g2_buf_2 fanout525 (.A(_03196_),
    .X(net525));
 sg13g2_buf_2 fanout526 (.A(_03193_),
    .X(net526));
 sg13g2_buf_2 fanout527 (.A(_03184_),
    .X(net527));
 sg13g2_buf_2 fanout528 (.A(_03183_),
    .X(net528));
 sg13g2_buf_4 fanout529 (.X(net529),
    .A(_03182_));
 sg13g2_buf_2 fanout530 (.A(_03152_),
    .X(net530));
 sg13g2_buf_2 fanout531 (.A(_03123_),
    .X(net531));
 sg13g2_buf_2 fanout532 (.A(_03121_),
    .X(net532));
 sg13g2_buf_2 fanout533 (.A(_03115_),
    .X(net533));
 sg13g2_buf_2 fanout534 (.A(_03095_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_03093_),
    .X(net535));
 sg13g2_buf_2 fanout536 (.A(_03083_),
    .X(net536));
 sg13g2_buf_4 fanout537 (.X(net537),
    .A(_03082_));
 sg13g2_buf_2 fanout538 (.A(_03050_),
    .X(net538));
 sg13g2_buf_2 fanout539 (.A(_03017_),
    .X(net539));
 sg13g2_buf_2 fanout540 (.A(_02882_),
    .X(net540));
 sg13g2_buf_2 fanout541 (.A(_02877_),
    .X(net541));
 sg13g2_buf_2 fanout542 (.A(_11232_),
    .X(net542));
 sg13g2_buf_2 fanout543 (.A(_11227_),
    .X(net543));
 sg13g2_buf_2 fanout544 (.A(_11207_),
    .X(net544));
 sg13g2_buf_2 fanout545 (.A(_11204_),
    .X(net545));
 sg13g2_buf_2 fanout546 (.A(_11194_),
    .X(net546));
 sg13g2_buf_2 fanout547 (.A(_11193_),
    .X(net547));
 sg13g2_buf_4 fanout548 (.X(net548),
    .A(_11191_));
 sg13g2_buf_2 fanout549 (.A(_11172_),
    .X(net549));
 sg13g2_buf_2 fanout550 (.A(_11170_),
    .X(net550));
 sg13g2_buf_2 fanout551 (.A(_11159_),
    .X(net551));
 sg13g2_buf_4 fanout552 (.X(net552),
    .A(_11158_));
 sg13g2_buf_2 fanout553 (.A(_11140_),
    .X(net553));
 sg13g2_buf_2 fanout554 (.A(_11137_),
    .X(net554));
 sg13g2_buf_2 fanout555 (.A(_11128_),
    .X(net555));
 sg13g2_buf_2 fanout556 (.A(_11127_),
    .X(net556));
 sg13g2_buf_4 fanout557 (.X(net557),
    .A(_11126_));
 sg13g2_buf_2 fanout558 (.A(_11105_),
    .X(net558));
 sg13g2_buf_2 fanout559 (.A(_11100_),
    .X(net559));
 sg13g2_buf_2 fanout560 (.A(_11086_),
    .X(net560));
 sg13g2_buf_2 fanout561 (.A(_11085_),
    .X(net561));
 sg13g2_buf_4 fanout562 (.X(net562),
    .A(_11084_));
 sg13g2_buf_2 fanout563 (.A(_10920_),
    .X(net563));
 sg13g2_buf_4 fanout564 (.X(net564),
    .A(_10916_));
 sg13g2_buf_2 fanout565 (.A(_10899_),
    .X(net565));
 sg13g2_buf_2 fanout566 (.A(_10896_),
    .X(net566));
 sg13g2_buf_2 fanout567 (.A(_10886_),
    .X(net567));
 sg13g2_buf_2 fanout568 (.A(_10885_),
    .X(net568));
 sg13g2_buf_4 fanout569 (.X(net569),
    .A(_10884_));
 sg13g2_buf_2 fanout570 (.A(_10866_),
    .X(net570));
 sg13g2_buf_2 fanout571 (.A(_10864_),
    .X(net571));
 sg13g2_buf_2 fanout572 (.A(_10853_),
    .X(net572));
 sg13g2_buf_2 fanout573 (.A(_10852_),
    .X(net573));
 sg13g2_buf_4 fanout574 (.X(net574),
    .A(_10836_));
 sg13g2_buf_2 fanout575 (.A(_10829_),
    .X(net575));
 sg13g2_buf_2 fanout576 (.A(_10828_),
    .X(net576));
 sg13g2_buf_4 fanout577 (.X(net577),
    .A(_10827_));
 sg13g2_buf_4 fanout578 (.X(net578),
    .A(_10805_));
 sg13g2_buf_4 fanout579 (.X(net579),
    .A(_10794_));
 sg13g2_buf_2 fanout580 (.A(_10791_),
    .X(net580));
 sg13g2_buf_2 fanout581 (.A(_10790_),
    .X(net581));
 sg13g2_buf_2 fanout582 (.A(_10767_),
    .X(net582));
 sg13g2_buf_2 fanout583 (.A(_10763_),
    .X(net583));
 sg13g2_buf_4 fanout584 (.X(net584),
    .A(_10755_));
 sg13g2_buf_2 fanout585 (.A(_10752_),
    .X(net585));
 sg13g2_buf_2 fanout586 (.A(_10727_),
    .X(net586));
 sg13g2_buf_2 fanout587 (.A(_10719_),
    .X(net587));
 sg13g2_buf_2 fanout588 (.A(_10714_),
    .X(net588));
 sg13g2_buf_2 fanout589 (.A(_10702_),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(_10701_),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(_10052_),
    .X(net591));
 sg13g2_buf_2 fanout592 (.A(_09943_),
    .X(net592));
 sg13g2_buf_2 fanout593 (.A(_08859_),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(_06433_),
    .X(net594));
 sg13g2_buf_4 fanout595 (.X(net595),
    .A(_06162_));
 sg13g2_buf_2 fanout596 (.A(_06143_),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_06134_),
    .X(net597));
 sg13g2_buf_2 fanout598 (.A(_05938_),
    .X(net598));
 sg13g2_buf_4 fanout599 (.X(net599),
    .A(_05889_));
 sg13g2_buf_2 fanout600 (.A(_05851_),
    .X(net600));
 sg13g2_buf_2 fanout601 (.A(_05845_),
    .X(net601));
 sg13g2_buf_2 fanout602 (.A(_05832_),
    .X(net602));
 sg13g2_buf_4 fanout603 (.X(net603),
    .A(_05820_));
 sg13g2_buf_2 fanout604 (.A(_05806_),
    .X(net604));
 sg13g2_buf_4 fanout605 (.X(net605),
    .A(_05710_));
 sg13g2_buf_4 fanout606 (.X(net606),
    .A(_05696_));
 sg13g2_buf_2 fanout607 (.A(_05676_),
    .X(net607));
 sg13g2_buf_2 fanout608 (.A(_05674_),
    .X(net608));
 sg13g2_buf_4 fanout609 (.X(net609),
    .A(_05590_));
 sg13g2_buf_2 fanout610 (.A(_05565_),
    .X(net610));
 sg13g2_buf_2 fanout611 (.A(_05503_),
    .X(net611));
 sg13g2_buf_2 fanout612 (.A(_05469_),
    .X(net612));
 sg13g2_buf_2 fanout613 (.A(_05404_),
    .X(net613));
 sg13g2_buf_4 fanout614 (.X(net614),
    .A(_05360_));
 sg13g2_buf_2 fanout615 (.A(_05342_),
    .X(net615));
 sg13g2_buf_2 fanout616 (.A(_04809_),
    .X(net616));
 sg13g2_buf_2 fanout617 (.A(_04769_),
    .X(net617));
 sg13g2_buf_2 fanout618 (.A(_04733_),
    .X(net618));
 sg13g2_buf_2 fanout619 (.A(_04731_),
    .X(net619));
 sg13g2_buf_2 fanout620 (.A(_04106_),
    .X(net620));
 sg13g2_buf_2 fanout621 (.A(_04083_),
    .X(net621));
 sg13g2_buf_2 fanout622 (.A(_04021_),
    .X(net622));
 sg13g2_buf_2 fanout623 (.A(_04018_),
    .X(net623));
 sg13g2_buf_2 fanout624 (.A(_03914_),
    .X(net624));
 sg13g2_buf_2 fanout625 (.A(_03908_),
    .X(net625));
 sg13g2_buf_2 fanout626 (.A(_03689_),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(_03684_),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(_03655_),
    .X(net628));
 sg13g2_buf_2 fanout629 (.A(_03652_),
    .X(net629));
 sg13g2_buf_2 fanout630 (.A(_03627_),
    .X(net630));
 sg13g2_buf_2 fanout631 (.A(_03622_),
    .X(net631));
 sg13g2_buf_2 fanout632 (.A(_03534_),
    .X(net632));
 sg13g2_buf_2 fanout633 (.A(_03532_),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(_03528_),
    .X(net634));
 sg13g2_buf_2 fanout635 (.A(_03502_),
    .X(net635));
 sg13g2_buf_2 fanout636 (.A(_03497_),
    .X(net636));
 sg13g2_buf_2 fanout637 (.A(_03468_),
    .X(net637));
 sg13g2_buf_2 fanout638 (.A(_03443_),
    .X(net638));
 sg13g2_buf_4 fanout639 (.X(net639),
    .A(_03439_));
 sg13g2_buf_4 fanout640 (.X(net640),
    .A(_03377_));
 sg13g2_buf_2 fanout641 (.A(_03352_),
    .X(net641));
 sg13g2_buf_2 fanout642 (.A(_03347_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(_03318_),
    .X(net643));
 sg13g2_buf_2 fanout644 (.A(_03248_),
    .X(net644));
 sg13g2_buf_2 fanout645 (.A(_03246_),
    .X(net645));
 sg13g2_buf_2 fanout646 (.A(_03241_),
    .X(net646));
 sg13g2_buf_2 fanout647 (.A(_03215_),
    .X(net647));
 sg13g2_buf_2 fanout648 (.A(_03210_),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(_03181_),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(_03114_),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(_03084_),
    .X(net651));
 sg13g2_buf_2 fanout652 (.A(_03081_),
    .X(net652));
 sg13g2_buf_2 fanout653 (.A(_03049_),
    .X(net653));
 sg13g2_buf_2 fanout654 (.A(_11190_),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_11160_),
    .X(net655));
 sg13g2_buf_2 fanout656 (.A(_11157_),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(_11083_),
    .X(net657));
 sg13g2_buf_2 fanout658 (.A(_10883_),
    .X(net658));
 sg13g2_buf_2 fanout659 (.A(_10826_),
    .X(net659));
 sg13g2_buf_2 fanout660 (.A(_10789_),
    .X(net660));
 sg13g2_buf_2 fanout661 (.A(_10753_),
    .X(net661));
 sg13g2_buf_2 fanout662 (.A(_10751_),
    .X(net662));
 sg13g2_buf_1 fanout663 (.A(_10169_),
    .X(net663));
 sg13g2_buf_2 fanout664 (.A(_07946_),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_07743_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(_07724_),
    .X(net666));
 sg13g2_buf_2 fanout667 (.A(_07637_),
    .X(net667));
 sg13g2_buf_4 fanout668 (.X(net668),
    .A(_06260_));
 sg13g2_buf_4 fanout669 (.X(net669),
    .A(_06119_));
 sg13g2_buf_2 fanout670 (.A(_06021_),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(_06003_),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(_05934_),
    .X(net672));
 sg13g2_buf_4 fanout673 (.X(net673),
    .A(_05802_));
 sg13g2_buf_2 fanout674 (.A(_05678_),
    .X(net674));
 sg13g2_buf_4 fanout675 (.X(net675),
    .A(_05572_));
 sg13g2_buf_2 fanout676 (.A(_05566_),
    .X(net676));
 sg13g2_buf_4 fanout677 (.X(net677),
    .A(_05564_));
 sg13g2_buf_2 fanout678 (.A(_05529_),
    .X(net678));
 sg13g2_buf_4 fanout679 (.X(net679),
    .A(_05508_));
 sg13g2_buf_2 fanout680 (.A(_05386_),
    .X(net680));
 sg13g2_buf_4 fanout681 (.X(net681),
    .A(_05363_));
 sg13g2_buf_4 fanout682 (.X(net682),
    .A(_05359_));
 sg13g2_buf_2 fanout683 (.A(_05344_),
    .X(net683));
 sg13g2_buf_4 fanout684 (.X(net684),
    .A(_05341_));
 sg13g2_buf_2 fanout685 (.A(_05282_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(_04725_),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(_03824_),
    .X(net687));
 sg13g2_buf_2 fanout688 (.A(_03527_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(_03438_),
    .X(net689));
 sg13g2_buf_2 fanout690 (.A(_03240_),
    .X(net690));
 sg13g2_buf_4 fanout691 (.X(net691),
    .A(_10849_));
 sg13g2_buf_2 fanout692 (.A(_09915_),
    .X(net692));
 sg13g2_buf_2 fanout693 (.A(_06390_),
    .X(net693));
 sg13g2_buf_2 fanout694 (.A(_06163_),
    .X(net694));
 sg13g2_buf_2 fanout695 (.A(_06160_),
    .X(net695));
 sg13g2_buf_2 fanout696 (.A(_06009_),
    .X(net696));
 sg13g2_buf_2 fanout697 (.A(_05932_),
    .X(net697));
 sg13g2_buf_2 fanout698 (.A(_05871_),
    .X(net698));
 sg13g2_buf_2 fanout699 (.A(_05810_),
    .X(net699));
 sg13g2_buf_2 fanout700 (.A(_05599_),
    .X(net700));
 sg13g2_buf_4 fanout701 (.X(net701),
    .A(_05530_));
 sg13g2_buf_2 fanout702 (.A(_05417_),
    .X(net702));
 sg13g2_buf_2 fanout703 (.A(_05400_),
    .X(net703));
 sg13g2_buf_4 fanout704 (.X(net704),
    .A(_05362_));
 sg13g2_buf_2 fanout705 (.A(_05358_),
    .X(net705));
 sg13g2_buf_4 fanout706 (.X(net706),
    .A(_05343_));
 sg13g2_buf_2 fanout707 (.A(_05331_),
    .X(net707));
 sg13g2_buf_2 fanout708 (.A(_05292_),
    .X(net708));
 sg13g2_buf_4 fanout709 (.X(net709),
    .A(_05272_));
 sg13g2_buf_2 fanout710 (.A(_05148_),
    .X(net710));
 sg13g2_buf_2 fanout711 (.A(_04105_),
    .X(net711));
 sg13g2_buf_2 fanout712 (.A(_04104_),
    .X(net712));
 sg13g2_buf_2 fanout713 (.A(_04017_),
    .X(net713));
 sg13g2_buf_2 fanout714 (.A(_04015_),
    .X(net714));
 sg13g2_buf_2 fanout715 (.A(_03902_),
    .X(net715));
 sg13g2_buf_2 fanout716 (.A(_03899_),
    .X(net716));
 sg13g2_buf_2 fanout717 (.A(_03823_),
    .X(net717));
 sg13g2_buf_4 fanout718 (.X(net718),
    .A(_03733_));
 sg13g2_buf_2 fanout719 (.A(_03717_),
    .X(net719));
 sg13g2_buf_2 fanout720 (.A(_06312_),
    .X(net720));
 sg13g2_buf_2 fanout721 (.A(_06056_),
    .X(net721));
 sg13g2_buf_2 fanout722 (.A(_05575_),
    .X(net722));
 sg13g2_buf_2 fanout723 (.A(_05426_),
    .X(net723));
 sg13g2_buf_2 fanout724 (.A(_05353_),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(_05142_),
    .X(net725));
 sg13g2_buf_2 fanout726 (.A(_05119_),
    .X(net726));
 sg13g2_buf_2 fanout727 (.A(_05118_),
    .X(net727));
 sg13g2_buf_2 fanout728 (.A(_03716_),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(_03079_),
    .X(net729));
 sg13g2_buf_2 fanout730 (.A(_10586_),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(_10100_),
    .X(net731));
 sg13g2_buf_2 fanout732 (.A(_09720_),
    .X(net732));
 sg13g2_buf_2 fanout733 (.A(_07636_),
    .X(net733));
 sg13g2_buf_4 fanout734 (.X(net734),
    .A(_05509_));
 sg13g2_buf_2 fanout735 (.A(_05154_),
    .X(net735));
 sg13g2_buf_2 fanout736 (.A(_05147_),
    .X(net736));
 sg13g2_buf_4 fanout737 (.X(net737),
    .A(_05132_));
 sg13g2_buf_2 fanout738 (.A(_05109_),
    .X(net738));
 sg13g2_buf_2 fanout739 (.A(_03715_),
    .X(net739));
 sg13g2_buf_2 fanout740 (.A(_10696_),
    .X(net740));
 sg13g2_buf_2 fanout741 (.A(_07635_),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(_05433_),
    .X(net742));
 sg13g2_buf_2 fanout743 (.A(_05365_),
    .X(net743));
 sg13g2_buf_2 fanout744 (.A(_05183_),
    .X(net744));
 sg13g2_buf_2 fanout745 (.A(_05146_),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(_04897_),
    .X(net746));
 sg13g2_buf_2 fanout747 (.A(_03737_),
    .X(net747));
 sg13g2_buf_4 fanout748 (.X(net748),
    .A(_03714_));
 sg13g2_buf_2 fanout749 (.A(_10477_),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(_08982_),
    .X(net750));
 sg13g2_buf_2 fanout751 (.A(_08981_),
    .X(net751));
 sg13g2_buf_4 fanout752 (.X(net752),
    .A(_07720_));
 sg13g2_buf_2 fanout753 (.A(_07716_),
    .X(net753));
 sg13g2_buf_2 fanout754 (.A(_07684_),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(_07678_),
    .X(net755));
 sg13g2_buf_2 fanout756 (.A(_07625_),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(_07590_),
    .X(net757));
 sg13g2_buf_2 fanout758 (.A(_07572_),
    .X(net758));
 sg13g2_buf_2 fanout759 (.A(_04937_),
    .X(net759));
 sg13g2_buf_2 fanout760 (.A(_04896_),
    .X(net760));
 sg13g2_buf_2 fanout761 (.A(_04643_),
    .X(net761));
 sg13g2_buf_2 fanout762 (.A(_04472_),
    .X(net762));
 sg13g2_buf_2 fanout763 (.A(_08980_),
    .X(net763));
 sg13g2_buf_2 fanout764 (.A(_07772_),
    .X(net764));
 sg13g2_buf_2 fanout765 (.A(_07719_),
    .X(net765));
 sg13g2_buf_2 fanout766 (.A(_07718_),
    .X(net766));
 sg13g2_buf_2 fanout767 (.A(_07682_),
    .X(net767));
 sg13g2_buf_2 fanout768 (.A(_07680_),
    .X(net768));
 sg13g2_buf_2 fanout769 (.A(_07657_),
    .X(net769));
 sg13g2_buf_2 fanout770 (.A(_07649_),
    .X(net770));
 sg13g2_buf_2 fanout771 (.A(_07646_),
    .X(net771));
 sg13g2_buf_2 fanout772 (.A(_07640_),
    .X(net772));
 sg13g2_buf_2 fanout773 (.A(_07624_),
    .X(net773));
 sg13g2_buf_2 fanout774 (.A(_07594_),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(_07589_),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(_07571_),
    .X(net776));
 sg13g2_buf_2 fanout777 (.A(_04882_),
    .X(net777));
 sg13g2_buf_2 fanout778 (.A(_04642_),
    .X(net778));
 sg13g2_buf_2 fanout779 (.A(_04485_),
    .X(net779));
 sg13g2_buf_2 fanout780 (.A(_04476_),
    .X(net780));
 sg13g2_buf_2 fanout781 (.A(_04469_),
    .X(net781));
 sg13g2_buf_2 fanout782 (.A(_04457_),
    .X(net782));
 sg13g2_buf_2 fanout783 (.A(_04423_),
    .X(net783));
 sg13g2_buf_2 fanout784 (.A(_04416_),
    .X(net784));
 sg13g2_buf_2 fanout785 (.A(_04410_),
    .X(net785));
 sg13g2_buf_2 fanout786 (.A(_04387_),
    .X(net786));
 sg13g2_buf_2 fanout787 (.A(_04381_),
    .X(net787));
 sg13g2_buf_2 fanout788 (.A(_04375_),
    .X(net788));
 sg13g2_buf_2 fanout789 (.A(_04357_),
    .X(net789));
 sg13g2_buf_2 fanout790 (.A(_09822_),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(_09817_),
    .X(net791));
 sg13g2_buf_2 fanout792 (.A(_09668_),
    .X(net792));
 sg13g2_buf_2 fanout793 (.A(_09003_),
    .X(net793));
 sg13g2_buf_2 fanout794 (.A(\top_ihp.oisc.reg_rb[2] ),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(_08581_),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(_08548_),
    .X(net796));
 sg13g2_buf_2 fanout797 (.A(_08441_),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(_08424_),
    .X(net798));
 sg13g2_buf_2 fanout799 (.A(_07795_),
    .X(net799));
 sg13g2_buf_4 fanout800 (.X(net800),
    .A(_07767_));
 sg13g2_buf_2 fanout801 (.A(_07728_),
    .X(net801));
 sg13g2_buf_4 fanout802 (.X(net802),
    .A(_07704_));
 sg13g2_buf_4 fanout803 (.X(net803),
    .A(_07700_));
 sg13g2_buf_2 fanout804 (.A(_07681_),
    .X(net804));
 sg13g2_buf_2 fanout805 (.A(_07673_),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(_07671_),
    .X(net806));
 sg13g2_buf_4 fanout807 (.X(net807),
    .A(_07639_));
 sg13g2_buf_4 fanout808 (.X(net808),
    .A(_07583_));
 sg13g2_buf_2 fanout809 (.A(_07577_),
    .X(net809));
 sg13g2_buf_4 fanout810 (.X(net810),
    .A(_07570_));
 sg13g2_buf_2 fanout811 (.A(_04467_),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(_04434_),
    .X(net812));
 sg13g2_buf_2 fanout813 (.A(_04432_),
    .X(net813));
 sg13g2_buf_2 fanout814 (.A(_04427_),
    .X(net814));
 sg13g2_buf_2 fanout815 (.A(_04420_),
    .X(net815));
 sg13g2_buf_2 fanout816 (.A(_04394_),
    .X(net816));
 sg13g2_buf_2 fanout817 (.A(_04392_),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(_04366_),
    .X(net818));
 sg13g2_buf_2 fanout819 (.A(_04364_),
    .X(net819));
 sg13g2_buf_2 fanout820 (.A(_04360_),
    .X(net820));
 sg13g2_buf_2 fanout821 (.A(_10536_),
    .X(net821));
 sg13g2_buf_2 fanout822 (.A(_10331_),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(_09853_),
    .X(net823));
 sg13g2_buf_2 fanout824 (.A(_09833_),
    .X(net824));
 sg13g2_buf_2 fanout825 (.A(_09830_),
    .X(net825));
 sg13g2_buf_2 fanout826 (.A(_09821_),
    .X(net826));
 sg13g2_buf_2 fanout827 (.A(_09816_),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(_09139_),
    .X(net828));
 sg13g2_buf_2 fanout829 (.A(_09011_),
    .X(net829));
 sg13g2_buf_2 fanout830 (.A(_08999_),
    .X(net830));
 sg13g2_buf_2 fanout831 (.A(_08440_),
    .X(net831));
 sg13g2_buf_2 fanout832 (.A(_08418_),
    .X(net832));
 sg13g2_buf_2 fanout833 (.A(_07769_),
    .X(net833));
 sg13g2_buf_2 fanout834 (.A(_07733_),
    .X(net834));
 sg13g2_buf_4 fanout835 (.X(net835),
    .A(_07713_));
 sg13g2_buf_2 fanout836 (.A(_07628_),
    .X(net836));
 sg13g2_buf_2 fanout837 (.A(_07602_),
    .X(net837));
 sg13g2_buf_2 fanout838 (.A(_07599_),
    .X(net838));
 sg13g2_buf_2 fanout839 (.A(_07568_),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(_05373_),
    .X(net840));
 sg13g2_buf_4 fanout841 (.X(net841),
    .A(_05303_));
 sg13g2_buf_2 fanout842 (.A(_04675_),
    .X(net842));
 sg13g2_buf_2 fanout843 (.A(_04363_),
    .X(net843));
 sg13g2_buf_2 fanout844 (.A(_04359_),
    .X(net844));
 sg13g2_buf_2 fanout845 (.A(_09815_),
    .X(net845));
 sg13g2_buf_2 fanout846 (.A(_08958_),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(_07761_),
    .X(net847));
 sg13g2_buf_2 fanout848 (.A(_07754_),
    .X(net848));
 sg13g2_buf_2 fanout849 (.A(_07726_),
    .X(net849));
 sg13g2_buf_2 fanout850 (.A(_07692_),
    .X(net850));
 sg13g2_buf_2 fanout851 (.A(_07674_),
    .X(net851));
 sg13g2_buf_2 fanout852 (.A(_07627_),
    .X(net852));
 sg13g2_buf_2 fanout853 (.A(_07582_),
    .X(net853));
 sg13g2_buf_2 fanout854 (.A(_04772_),
    .X(net854));
 sg13g2_buf_2 fanout855 (.A(_04771_),
    .X(net855));
 sg13g2_buf_2 fanout856 (.A(_04758_),
    .X(net856));
 sg13g2_buf_2 fanout857 (.A(_04754_),
    .X(net857));
 sg13g2_buf_2 fanout858 (.A(_10152_),
    .X(net858));
 sg13g2_buf_2 fanout859 (.A(_09829_),
    .X(net859));
 sg13g2_buf_2 fanout860 (.A(_09122_),
    .X(net860));
 sg13g2_buf_2 fanout861 (.A(_08945_),
    .X(net861));
 sg13g2_buf_2 fanout862 (.A(_08595_),
    .X(net862));
 sg13g2_buf_2 fanout863 (.A(_07712_),
    .X(net863));
 sg13g2_buf_2 fanout864 (.A(_07691_),
    .X(net864));
 sg13g2_buf_2 fanout865 (.A(_07581_),
    .X(net865));
 sg13g2_buf_2 fanout866 (.A(_04723_),
    .X(net866));
 sg13g2_buf_4 fanout867 (.X(net867),
    .A(_03779_));
 sg13g2_buf_2 fanout868 (.A(_03761_),
    .X(net868));
 sg13g2_buf_2 fanout869 (.A(_03759_),
    .X(net869));
 sg13g2_buf_4 fanout870 (.X(net870),
    .A(_03756_));
 sg13g2_buf_2 fanout871 (.A(_03727_),
    .X(net871));
 sg13g2_buf_2 fanout872 (.A(_10229_),
    .X(net872));
 sg13g2_buf_2 fanout873 (.A(_10110_),
    .X(net873));
 sg13g2_buf_2 fanout874 (.A(_10054_),
    .X(net874));
 sg13g2_buf_2 fanout875 (.A(_10042_),
    .X(net875));
 sg13g2_buf_2 fanout876 (.A(_09884_),
    .X(net876));
 sg13g2_buf_2 fanout877 (.A(_09873_),
    .X(net877));
 sg13g2_buf_2 fanout878 (.A(_09828_),
    .X(net878));
 sg13g2_buf_2 fanout879 (.A(_09818_),
    .X(net879));
 sg13g2_buf_2 fanout880 (.A(_09786_),
    .X(net880));
 sg13g2_buf_2 fanout881 (.A(_09341_),
    .X(net881));
 sg13g2_buf_2 fanout882 (.A(_09313_),
    .X(net882));
 sg13g2_buf_2 fanout883 (.A(_09259_),
    .X(net883));
 sg13g2_buf_2 fanout884 (.A(_09223_),
    .X(net884));
 sg13g2_buf_2 fanout885 (.A(_09153_),
    .X(net885));
 sg13g2_buf_2 fanout886 (.A(_09064_),
    .X(net886));
 sg13g2_buf_2 fanout887 (.A(_09059_),
    .X(net887));
 sg13g2_buf_2 fanout888 (.A(_09054_),
    .X(net888));
 sg13g2_buf_2 fanout889 (.A(_09025_),
    .X(net889));
 sg13g2_buf_2 fanout890 (.A(_09006_),
    .X(net890));
 sg13g2_buf_2 fanout891 (.A(_08965_),
    .X(net891));
 sg13g2_buf_2 fanout892 (.A(_08211_),
    .X(net892));
 sg13g2_buf_2 fanout893 (.A(_07695_),
    .X(net893));
 sg13g2_buf_2 fanout894 (.A(_04487_),
    .X(net894));
 sg13g2_buf_2 fanout895 (.A(_04483_),
    .X(net895));
 sg13g2_buf_2 fanout896 (.A(_04318_),
    .X(net896));
 sg13g2_buf_2 fanout897 (.A(_03929_),
    .X(net897));
 sg13g2_buf_2 fanout898 (.A(_03851_),
    .X(net898));
 sg13g2_buf_2 fanout899 (.A(_03840_),
    .X(net899));
 sg13g2_buf_2 fanout900 (.A(_03755_),
    .X(net900));
 sg13g2_buf_2 fanout901 (.A(_10155_),
    .X(net901));
 sg13g2_buf_2 fanout902 (.A(_10003_),
    .X(net902));
 sg13g2_buf_2 fanout903 (.A(_09877_),
    .X(net903));
 sg13g2_buf_2 fanout904 (.A(_09827_),
    .X(net904));
 sg13g2_buf_2 fanout905 (.A(_09825_),
    .X(net905));
 sg13g2_buf_2 fanout906 (.A(_09814_),
    .X(net906));
 sg13g2_buf_2 fanout907 (.A(_09785_),
    .X(net907));
 sg13g2_buf_2 fanout908 (.A(_09267_),
    .X(net908));
 sg13g2_buf_2 fanout909 (.A(_09256_),
    .X(net909));
 sg13g2_buf_2 fanout910 (.A(_09251_),
    .X(net910));
 sg13g2_buf_2 fanout911 (.A(_09248_),
    .X(net911));
 sg13g2_buf_2 fanout912 (.A(_09231_),
    .X(net912));
 sg13g2_buf_2 fanout913 (.A(_09226_),
    .X(net913));
 sg13g2_buf_2 fanout914 (.A(_09212_),
    .X(net914));
 sg13g2_buf_2 fanout915 (.A(_09205_),
    .X(net915));
 sg13g2_buf_2 fanout916 (.A(_09198_),
    .X(net916));
 sg13g2_buf_2 fanout917 (.A(_09155_),
    .X(net917));
 sg13g2_buf_2 fanout918 (.A(_09143_),
    .X(net918));
 sg13g2_buf_2 fanout919 (.A(_09128_),
    .X(net919));
 sg13g2_buf_2 fanout920 (.A(_09119_),
    .X(net920));
 sg13g2_buf_2 fanout921 (.A(_09117_),
    .X(net921));
 sg13g2_buf_2 fanout922 (.A(_09108_),
    .X(net922));
 sg13g2_buf_2 fanout923 (.A(_09107_),
    .X(net923));
 sg13g2_buf_2 fanout924 (.A(_09095_),
    .X(net924));
 sg13g2_buf_2 fanout925 (.A(_09080_),
    .X(net925));
 sg13g2_buf_2 fanout926 (.A(_09077_),
    .X(net926));
 sg13g2_buf_2 fanout927 (.A(_09063_),
    .X(net927));
 sg13g2_buf_2 fanout928 (.A(_09053_),
    .X(net928));
 sg13g2_buf_2 fanout929 (.A(_09051_),
    .X(net929));
 sg13g2_buf_2 fanout930 (.A(_09044_),
    .X(net930));
 sg13g2_buf_2 fanout931 (.A(_09030_),
    .X(net931));
 sg13g2_buf_2 fanout932 (.A(_09024_),
    .X(net932));
 sg13g2_buf_2 fanout933 (.A(_09018_),
    .X(net933));
 sg13g2_buf_2 fanout934 (.A(_08420_),
    .X(net934));
 sg13g2_buf_4 fanout935 (.X(net935),
    .A(_07643_));
 sg13g2_buf_2 fanout936 (.A(_04960_),
    .X(net936));
 sg13g2_buf_2 fanout937 (.A(_04863_),
    .X(net937));
 sg13g2_buf_2 fanout938 (.A(_04482_),
    .X(net938));
 sg13g2_buf_2 fanout939 (.A(_03982_),
    .X(net939));
 sg13g2_buf_2 fanout940 (.A(_03889_),
    .X(net940));
 sg13g2_buf_2 fanout941 (.A(_03855_),
    .X(net941));
 sg13g2_buf_2 fanout942 (.A(_03848_),
    .X(net942));
 sg13g2_buf_2 fanout943 (.A(_03839_),
    .X(net943));
 sg13g2_buf_2 fanout944 (.A(_03835_),
    .X(net944));
 sg13g2_buf_2 fanout945 (.A(_03833_),
    .X(net945));
 sg13g2_buf_2 fanout946 (.A(_03830_),
    .X(net946));
 sg13g2_buf_2 fanout947 (.A(_03827_),
    .X(net947));
 sg13g2_buf_2 fanout948 (.A(_03728_),
    .X(net948));
 sg13g2_buf_2 fanout949 (.A(_10116_),
    .X(net949));
 sg13g2_buf_2 fanout950 (.A(_10092_),
    .X(net950));
 sg13g2_buf_2 fanout951 (.A(_09982_),
    .X(net951));
 sg13g2_buf_2 fanout952 (.A(_09871_),
    .X(net952));
 sg13g2_buf_2 fanout953 (.A(_09850_),
    .X(net953));
 sg13g2_buf_2 fanout954 (.A(_09848_),
    .X(net954));
 sg13g2_buf_2 fanout955 (.A(_09846_),
    .X(net955));
 sg13g2_buf_2 fanout956 (.A(_09824_),
    .X(net956));
 sg13g2_buf_2 fanout957 (.A(_09813_),
    .X(net957));
 sg13g2_buf_2 fanout958 (.A(_09789_),
    .X(net958));
 sg13g2_buf_2 fanout959 (.A(_09779_),
    .X(net959));
 sg13g2_buf_2 fanout960 (.A(_09671_),
    .X(net960));
 sg13g2_buf_2 fanout961 (.A(_09296_),
    .X(net961));
 sg13g2_buf_2 fanout962 (.A(_09175_),
    .X(net962));
 sg13g2_buf_2 fanout963 (.A(_09142_),
    .X(net963));
 sg13g2_buf_2 fanout964 (.A(_09127_),
    .X(net964));
 sg13g2_buf_2 fanout965 (.A(_09116_),
    .X(net965));
 sg13g2_buf_2 fanout966 (.A(_09113_),
    .X(net966));
 sg13g2_buf_2 fanout967 (.A(_09096_),
    .X(net967));
 sg13g2_buf_2 fanout968 (.A(_09092_),
    .X(net968));
 sg13g2_buf_2 fanout969 (.A(_09083_),
    .X(net969));
 sg13g2_buf_2 fanout970 (.A(_09078_),
    .X(net970));
 sg13g2_buf_2 fanout971 (.A(_09068_),
    .X(net971));
 sg13g2_buf_2 fanout972 (.A(_09062_),
    .X(net972));
 sg13g2_buf_2 fanout973 (.A(_09056_),
    .X(net973));
 sg13g2_buf_2 fanout974 (.A(_09048_),
    .X(net974));
 sg13g2_buf_2 fanout975 (.A(_09041_),
    .X(net975));
 sg13g2_buf_2 fanout976 (.A(_09039_),
    .X(net976));
 sg13g2_buf_2 fanout977 (.A(_09036_),
    .X(net977));
 sg13g2_buf_2 fanout978 (.A(_09033_),
    .X(net978));
 sg13g2_buf_2 fanout979 (.A(_09023_),
    .X(net979));
 sg13g2_buf_2 fanout980 (.A(_09017_),
    .X(net980));
 sg13g2_buf_2 fanout981 (.A(_09014_),
    .X(net981));
 sg13g2_buf_2 fanout982 (.A(_09000_),
    .X(net982));
 sg13g2_buf_2 fanout983 (.A(_08436_),
    .X(net983));
 sg13g2_buf_2 fanout984 (.A(_08419_),
    .X(net984));
 sg13g2_buf_4 fanout985 (.X(net985),
    .A(_07642_));
 sg13g2_buf_2 fanout986 (.A(_04920_),
    .X(net986));
 sg13g2_buf_2 fanout987 (.A(_04906_),
    .X(net987));
 sg13g2_buf_2 fanout988 (.A(_04902_),
    .X(net988));
 sg13g2_buf_2 fanout989 (.A(_04901_),
    .X(net989));
 sg13g2_buf_2 fanout990 (.A(_04026_),
    .X(net990));
 sg13g2_buf_2 fanout991 (.A(_03879_),
    .X(net991));
 sg13g2_buf_2 fanout992 (.A(_03869_),
    .X(net992));
 sg13g2_buf_2 fanout993 (.A(_03860_),
    .X(net993));
 sg13g2_buf_2 fanout994 (.A(_03850_),
    .X(net994));
 sg13g2_buf_2 fanout995 (.A(_03847_),
    .X(net995));
 sg13g2_buf_2 fanout996 (.A(_03842_),
    .X(net996));
 sg13g2_buf_2 fanout997 (.A(_03832_),
    .X(net997));
 sg13g2_buf_2 fanout998 (.A(_03829_),
    .X(net998));
 sg13g2_buf_2 fanout999 (.A(_09999_),
    .X(net999));
 sg13g2_buf_2 fanout1000 (.A(_09924_),
    .X(net1000));
 sg13g2_buf_2 fanout1001 (.A(_09860_),
    .X(net1001));
 sg13g2_buf_2 fanout1002 (.A(_09823_),
    .X(net1002));
 sg13g2_buf_2 fanout1003 (.A(_09811_),
    .X(net1003));
 sg13g2_buf_2 fanout1004 (.A(_09804_),
    .X(net1004));
 sg13g2_buf_2 fanout1005 (.A(_09793_),
    .X(net1005));
 sg13g2_buf_2 fanout1006 (.A(_09791_),
    .X(net1006));
 sg13g2_buf_2 fanout1007 (.A(_09788_),
    .X(net1007));
 sg13g2_buf_2 fanout1008 (.A(_09670_),
    .X(net1008));
 sg13g2_buf_2 fanout1009 (.A(_09126_),
    .X(net1009));
 sg13g2_buf_2 fanout1010 (.A(_09106_),
    .X(net1010));
 sg13g2_buf_2 fanout1011 (.A(_09067_),
    .X(net1011));
 sg13g2_buf_2 fanout1012 (.A(_09065_),
    .X(net1012));
 sg13g2_buf_2 fanout1013 (.A(_09046_),
    .X(net1013));
 sg13g2_buf_2 fanout1014 (.A(_09038_),
    .X(net1014));
 sg13g2_buf_2 fanout1015 (.A(_09035_),
    .X(net1015));
 sg13g2_buf_2 fanout1016 (.A(_09027_),
    .X(net1016));
 sg13g2_buf_2 fanout1017 (.A(_09022_),
    .X(net1017));
 sg13g2_buf_2 fanout1018 (.A(_09020_),
    .X(net1018));
 sg13g2_buf_2 fanout1019 (.A(_09013_),
    .X(net1019));
 sg13g2_buf_2 fanout1020 (.A(_08985_),
    .X(net1020));
 sg13g2_buf_2 fanout1021 (.A(_08964_),
    .X(net1021));
 sg13g2_buf_2 fanout1022 (.A(_08952_),
    .X(net1022));
 sg13g2_buf_2 fanout1023 (.A(_08949_),
    .X(net1023));
 sg13g2_buf_2 fanout1024 (.A(_08942_),
    .X(net1024));
 sg13g2_buf_2 fanout1025 (.A(_08658_),
    .X(net1025));
 sg13g2_buf_2 fanout1026 (.A(_08546_),
    .X(net1026));
 sg13g2_buf_2 fanout1027 (.A(_08435_),
    .X(net1027));
 sg13g2_buf_2 fanout1028 (.A(_08413_),
    .X(net1028));
 sg13g2_buf_2 fanout1029 (.A(_08366_),
    .X(net1029));
 sg13g2_buf_2 fanout1030 (.A(_08260_),
    .X(net1030));
 sg13g2_buf_2 fanout1031 (.A(_08217_),
    .X(net1031));
 sg13g2_buf_2 fanout1032 (.A(_08200_),
    .X(net1032));
 sg13g2_buf_2 fanout1033 (.A(_03825_),
    .X(net1033));
 sg13g2_buf_2 fanout1034 (.A(_03753_),
    .X(net1034));
 sg13g2_buf_2 fanout1035 (.A(_09810_),
    .X(net1035));
 sg13g2_buf_2 fanout1036 (.A(_09790_),
    .X(net1036));
 sg13g2_buf_2 fanout1037 (.A(_09782_),
    .X(net1037));
 sg13g2_buf_2 fanout1038 (.A(_09028_),
    .X(net1038));
 sg13g2_buf_2 fanout1039 (.A(_09019_),
    .X(net1039));
 sg13g2_buf_2 fanout1040 (.A(_09015_),
    .X(net1040));
 sg13g2_buf_4 fanout1041 (.X(net1041),
    .A(_08993_));
 sg13g2_buf_2 fanout1042 (.A(_08710_),
    .X(net1042));
 sg13g2_buf_2 fanout1043 (.A(_08709_),
    .X(net1043));
 sg13g2_buf_2 fanout1044 (.A(_08708_),
    .X(net1044));
 sg13g2_buf_4 fanout1045 (.X(net1045),
    .A(_08557_));
 sg13g2_buf_2 fanout1046 (.A(_08450_),
    .X(net1046));
 sg13g2_buf_2 fanout1047 (.A(_08394_),
    .X(net1047));
 sg13g2_buf_2 fanout1048 (.A(_08380_),
    .X(net1048));
 sg13g2_buf_2 fanout1049 (.A(_08338_),
    .X(net1049));
 sg13g2_buf_2 fanout1050 (.A(_08329_),
    .X(net1050));
 sg13g2_buf_2 fanout1051 (.A(_08285_),
    .X(net1051));
 sg13g2_buf_4 fanout1052 (.X(net1052),
    .A(_08274_));
 sg13g2_buf_4 fanout1053 (.X(net1053),
    .A(_08262_));
 sg13g2_buf_2 fanout1054 (.A(_08261_),
    .X(net1054));
 sg13g2_buf_2 fanout1055 (.A(_08256_),
    .X(net1055));
 sg13g2_buf_2 fanout1056 (.A(_08228_),
    .X(net1056));
 sg13g2_buf_2 fanout1057 (.A(_08227_),
    .X(net1057));
 sg13g2_buf_2 fanout1058 (.A(_08223_),
    .X(net1058));
 sg13g2_buf_2 fanout1059 (.A(_08221_),
    .X(net1059));
 sg13g2_buf_2 fanout1060 (.A(_08669_),
    .X(net1060));
 sg13g2_buf_4 fanout1061 (.X(net1061),
    .A(net1064));
 sg13g2_buf_2 fanout1062 (.A(net1064),
    .X(net1062));
 sg13g2_buf_4 fanout1063 (.X(net1063),
    .A(net1064));
 sg13g2_buf_1 fanout1064 (.A(net1074),
    .X(net1064));
 sg13g2_buf_4 fanout1065 (.X(net1065),
    .A(net1068));
 sg13g2_buf_4 fanout1066 (.X(net1066),
    .A(net1068));
 sg13g2_buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sg13g2_buf_2 fanout1068 (.A(net1074),
    .X(net1068));
 sg13g2_buf_4 fanout1069 (.X(net1069),
    .A(net1070));
 sg13g2_buf_4 fanout1070 (.X(net1070),
    .A(net1074));
 sg13g2_buf_4 fanout1071 (.X(net1071),
    .A(net1073));
 sg13g2_buf_4 fanout1072 (.X(net1072),
    .A(net1073));
 sg13g2_buf_2 fanout1073 (.A(net1074),
    .X(net1073));
 sg13g2_buf_2 fanout1074 (.A(net1137),
    .X(net1074));
 sg13g2_buf_4 fanout1075 (.X(net1075),
    .A(net1076));
 sg13g2_buf_2 fanout1076 (.A(net1077),
    .X(net1076));
 sg13g2_buf_2 fanout1077 (.A(net1084),
    .X(net1077));
 sg13g2_buf_4 fanout1078 (.X(net1078),
    .A(net1084));
 sg13g2_buf_2 fanout1079 (.A(net1084),
    .X(net1079));
 sg13g2_buf_4 fanout1080 (.X(net1080),
    .A(net1083));
 sg13g2_buf_2 fanout1081 (.A(net1083),
    .X(net1081));
 sg13g2_buf_4 fanout1082 (.X(net1082),
    .A(net1083));
 sg13g2_buf_2 fanout1083 (.A(net1084),
    .X(net1083));
 sg13g2_buf_1 fanout1084 (.A(net1100),
    .X(net1084));
 sg13g2_buf_4 fanout1085 (.X(net1085),
    .A(net1087));
 sg13g2_buf_2 fanout1086 (.A(net1087),
    .X(net1086));
 sg13g2_buf_4 fanout1087 (.X(net1087),
    .A(net1091));
 sg13g2_buf_4 fanout1088 (.X(net1088),
    .A(net1090));
 sg13g2_buf_4 fanout1089 (.X(net1089),
    .A(net1090));
 sg13g2_buf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sg13g2_buf_1 fanout1091 (.A(net1100),
    .X(net1091));
 sg13g2_buf_4 fanout1092 (.X(net1092),
    .A(net1094));
 sg13g2_buf_2 fanout1093 (.A(net1094),
    .X(net1093));
 sg13g2_buf_4 fanout1094 (.X(net1094),
    .A(net1100));
 sg13g2_buf_4 fanout1095 (.X(net1095),
    .A(net1099));
 sg13g2_buf_2 fanout1096 (.A(net1099),
    .X(net1096));
 sg13g2_buf_4 fanout1097 (.X(net1097),
    .A(net1099));
 sg13g2_buf_4 fanout1098 (.X(net1098),
    .A(net1099));
 sg13g2_buf_1 fanout1099 (.A(net1100),
    .X(net1099));
 sg13g2_buf_1 fanout1100 (.A(net1137),
    .X(net1100));
 sg13g2_buf_4 fanout1101 (.X(net1101),
    .A(net1103));
 sg13g2_buf_2 fanout1102 (.A(net1103),
    .X(net1102));
 sg13g2_buf_1 fanout1103 (.A(net1109),
    .X(net1103));
 sg13g2_buf_4 fanout1104 (.X(net1104),
    .A(net1109));
 sg13g2_buf_2 fanout1105 (.A(net1109),
    .X(net1105));
 sg13g2_buf_4 fanout1106 (.X(net1106),
    .A(net1107));
 sg13g2_buf_4 fanout1107 (.X(net1107),
    .A(net1108));
 sg13g2_buf_4 fanout1108 (.X(net1108),
    .A(net1109));
 sg13g2_buf_2 fanout1109 (.A(net1137),
    .X(net1109));
 sg13g2_buf_4 fanout1110 (.X(net1110),
    .A(net1111));
 sg13g2_buf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sg13g2_buf_4 fanout1112 (.X(net1112),
    .A(net1117));
 sg13g2_buf_4 fanout1113 (.X(net1113),
    .A(net1114));
 sg13g2_buf_2 fanout1114 (.A(net1117),
    .X(net1114));
 sg13g2_buf_4 fanout1115 (.X(net1115),
    .A(net1117));
 sg13g2_buf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sg13g2_buf_1 fanout1117 (.A(net1137),
    .X(net1117));
 sg13g2_buf_4 fanout1118 (.X(net1118),
    .A(net1122));
 sg13g2_buf_4 fanout1119 (.X(net1119),
    .A(net1122));
 sg13g2_buf_4 fanout1120 (.X(net1120),
    .A(net1122));
 sg13g2_buf_4 fanout1121 (.X(net1121),
    .A(net1122));
 sg13g2_buf_1 fanout1122 (.A(net1128),
    .X(net1122));
 sg13g2_buf_4 fanout1123 (.X(net1123),
    .A(net1125));
 sg13g2_buf_4 fanout1124 (.X(net1124),
    .A(net1125));
 sg13g2_buf_2 fanout1125 (.A(net1128),
    .X(net1125));
 sg13g2_buf_4 fanout1126 (.X(net1126),
    .A(net1127));
 sg13g2_buf_4 fanout1127 (.X(net1127),
    .A(net1128));
 sg13g2_buf_1 fanout1128 (.A(net1136),
    .X(net1128));
 sg13g2_buf_4 fanout1129 (.X(net1129),
    .A(net1136));
 sg13g2_buf_4 fanout1130 (.X(net1130),
    .A(net1132));
 sg13g2_buf_4 fanout1131 (.X(net1131),
    .A(net1132));
 sg13g2_buf_2 fanout1132 (.A(net1135),
    .X(net1132));
 sg13g2_buf_4 fanout1133 (.X(net1133),
    .A(net1135));
 sg13g2_buf_2 fanout1134 (.A(net1135),
    .X(net1134));
 sg13g2_buf_1 fanout1135 (.A(net1136),
    .X(net1135));
 sg13g2_buf_1 fanout1136 (.A(net1137),
    .X(net1136));
 sg13g2_buf_1 fanout1137 (.A(net1),
    .X(net1137));
 sg13g2_buf_4 fanout1138 (.X(net1138),
    .A(net1141));
 sg13g2_buf_2 fanout1139 (.A(net1141),
    .X(net1139));
 sg13g2_buf_4 fanout1140 (.X(net1140),
    .A(net1141));
 sg13g2_buf_1 fanout1141 (.A(net1165),
    .X(net1141));
 sg13g2_buf_4 fanout1142 (.X(net1142),
    .A(net1146));
 sg13g2_buf_2 fanout1143 (.A(net1146),
    .X(net1143));
 sg13g2_buf_4 fanout1144 (.X(net1144),
    .A(net1146));
 sg13g2_buf_2 fanout1145 (.A(net1146),
    .X(net1145));
 sg13g2_buf_1 fanout1146 (.A(net1165),
    .X(net1146));
 sg13g2_buf_4 fanout1147 (.X(net1147),
    .A(net1149));
 sg13g2_buf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sg13g2_buf_4 fanout1149 (.X(net1149),
    .A(net1150));
 sg13g2_buf_2 fanout1150 (.A(net1165),
    .X(net1150));
 sg13g2_buf_4 fanout1151 (.X(net1151),
    .A(net1153));
 sg13g2_buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sg13g2_buf_4 fanout1153 (.X(net1153),
    .A(net1157));
 sg13g2_buf_4 fanout1154 (.X(net1154),
    .A(net1156));
 sg13g2_buf_2 fanout1155 (.A(net1156),
    .X(net1155));
 sg13g2_buf_4 fanout1156 (.X(net1156),
    .A(net1157));
 sg13g2_buf_2 fanout1157 (.A(net1165),
    .X(net1157));
 sg13g2_buf_4 fanout1158 (.X(net1158),
    .A(net1161));
 sg13g2_buf_4 fanout1159 (.X(net1159),
    .A(net1161));
 sg13g2_buf_2 fanout1160 (.A(net1161),
    .X(net1160));
 sg13g2_buf_2 fanout1161 (.A(net1164),
    .X(net1161));
 sg13g2_buf_4 fanout1162 (.X(net1162),
    .A(net1163));
 sg13g2_buf_4 fanout1163 (.X(net1163),
    .A(net1164));
 sg13g2_buf_1 fanout1164 (.A(net1165),
    .X(net1164));
 sg13g2_buf_1 fanout1165 (.A(net1265),
    .X(net1165));
 sg13g2_buf_4 fanout1166 (.X(net1166),
    .A(net1170));
 sg13g2_buf_2 fanout1167 (.A(net1170),
    .X(net1167));
 sg13g2_buf_4 fanout1168 (.X(net1168),
    .A(net1170));
 sg13g2_buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sg13g2_buf_1 fanout1170 (.A(net1197),
    .X(net1170));
 sg13g2_buf_4 fanout1171 (.X(net1171),
    .A(net1197));
 sg13g2_buf_4 fanout1172 (.X(net1172),
    .A(net1176));
 sg13g2_buf_4 fanout1173 (.X(net1173),
    .A(net1175));
 sg13g2_buf_4 fanout1174 (.X(net1174),
    .A(net1175));
 sg13g2_buf_1 fanout1175 (.A(net1176),
    .X(net1175));
 sg13g2_buf_1 fanout1176 (.A(net1181),
    .X(net1176));
 sg13g2_buf_4 fanout1177 (.X(net1177),
    .A(net1181));
 sg13g2_buf_2 fanout1178 (.A(net1181),
    .X(net1178));
 sg13g2_buf_4 fanout1179 (.X(net1179),
    .A(net1180));
 sg13g2_buf_4 fanout1180 (.X(net1180),
    .A(net1181));
 sg13g2_buf_1 fanout1181 (.A(net1197),
    .X(net1181));
 sg13g2_buf_4 fanout1182 (.X(net1182),
    .A(net1184));
 sg13g2_buf_4 fanout1183 (.X(net1183),
    .A(net1184));
 sg13g2_buf_2 fanout1184 (.A(net1197),
    .X(net1184));
 sg13g2_buf_4 fanout1185 (.X(net1185),
    .A(net1188));
 sg13g2_buf_4 fanout1186 (.X(net1186),
    .A(net1187));
 sg13g2_buf_4 fanout1187 (.X(net1187),
    .A(net1188));
 sg13g2_buf_2 fanout1188 (.A(net1197),
    .X(net1188));
 sg13g2_buf_4 fanout1189 (.X(net1189),
    .A(net1192));
 sg13g2_buf_4 fanout1190 (.X(net1190),
    .A(net1192));
 sg13g2_buf_4 fanout1191 (.X(net1191),
    .A(net1192));
 sg13g2_buf_2 fanout1192 (.A(net1196),
    .X(net1192));
 sg13g2_buf_4 fanout1193 (.X(net1193),
    .A(net1196));
 sg13g2_buf_2 fanout1194 (.A(net1196),
    .X(net1194));
 sg13g2_buf_4 fanout1195 (.X(net1195),
    .A(net1196));
 sg13g2_buf_1 fanout1196 (.A(net1197),
    .X(net1196));
 sg13g2_buf_1 fanout1197 (.A(net1265),
    .X(net1197));
 sg13g2_buf_4 fanout1198 (.X(net1198),
    .A(net1200));
 sg13g2_buf_2 fanout1199 (.A(net1200),
    .X(net1199));
 sg13g2_buf_4 fanout1200 (.X(net1200),
    .A(net1205));
 sg13g2_buf_4 fanout1201 (.X(net1201),
    .A(net1204));
 sg13g2_buf_2 fanout1202 (.A(net1204),
    .X(net1202));
 sg13g2_buf_4 fanout1203 (.X(net1203),
    .A(net1204));
 sg13g2_buf_2 fanout1204 (.A(net1205),
    .X(net1204));
 sg13g2_buf_1 fanout1205 (.A(net1211),
    .X(net1205));
 sg13g2_buf_4 fanout1206 (.X(net1206),
    .A(net1207));
 sg13g2_buf_4 fanout1207 (.X(net1207),
    .A(net1211));
 sg13g2_buf_4 fanout1208 (.X(net1208),
    .A(net1210));
 sg13g2_buf_4 fanout1209 (.X(net1209),
    .A(net1210));
 sg13g2_buf_2 fanout1210 (.A(net1211),
    .X(net1210));
 sg13g2_buf_1 fanout1211 (.A(net1265),
    .X(net1211));
 sg13g2_buf_4 fanout1212 (.X(net1212),
    .A(net1216));
 sg13g2_buf_4 fanout1213 (.X(net1213),
    .A(net1216));
 sg13g2_buf_4 fanout1214 (.X(net1214),
    .A(net1216));
 sg13g2_buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sg13g2_buf_1 fanout1216 (.A(net1228),
    .X(net1216));
 sg13g2_buf_4 fanout1217 (.X(net1217),
    .A(net1220));
 sg13g2_buf_4 fanout1218 (.X(net1218),
    .A(net1220));
 sg13g2_buf_2 fanout1219 (.A(net1220),
    .X(net1219));
 sg13g2_buf_2 fanout1220 (.A(net1228),
    .X(net1220));
 sg13g2_buf_4 fanout1221 (.X(net1221),
    .A(net1223));
 sg13g2_buf_4 fanout1222 (.X(net1222),
    .A(net1223));
 sg13g2_buf_4 fanout1223 (.X(net1223),
    .A(net1228));
 sg13g2_buf_4 fanout1224 (.X(net1224),
    .A(net1227));
 sg13g2_buf_4 fanout1225 (.X(net1225),
    .A(net1227));
 sg13g2_buf_2 fanout1226 (.A(net1227),
    .X(net1226));
 sg13g2_buf_2 fanout1227 (.A(net1228),
    .X(net1227));
 sg13g2_buf_1 fanout1228 (.A(net1265),
    .X(net1228));
 sg13g2_buf_4 fanout1229 (.X(net1229),
    .A(net1233));
 sg13g2_buf_2 fanout1230 (.A(net1233),
    .X(net1230));
 sg13g2_buf_4 fanout1231 (.X(net1231),
    .A(net1233));
 sg13g2_buf_2 fanout1232 (.A(net1233),
    .X(net1232));
 sg13g2_buf_1 fanout1233 (.A(net1247),
    .X(net1233));
 sg13g2_buf_4 fanout1234 (.X(net1234),
    .A(net1238));
 sg13g2_buf_2 fanout1235 (.A(net1238),
    .X(net1235));
 sg13g2_buf_4 fanout1236 (.X(net1236),
    .A(net1238));
 sg13g2_buf_2 fanout1237 (.A(net1238),
    .X(net1237));
 sg13g2_buf_1 fanout1238 (.A(net1247),
    .X(net1238));
 sg13g2_buf_4 fanout1239 (.X(net1239),
    .A(net1242));
 sg13g2_buf_4 fanout1240 (.X(net1240),
    .A(net1241));
 sg13g2_buf_4 fanout1241 (.X(net1241),
    .A(net1242));
 sg13g2_buf_2 fanout1242 (.A(net1247),
    .X(net1242));
 sg13g2_buf_4 fanout1243 (.X(net1243),
    .A(net1246));
 sg13g2_buf_4 fanout1244 (.X(net1244),
    .A(net1246));
 sg13g2_buf_4 fanout1245 (.X(net1245),
    .A(net1246));
 sg13g2_buf_2 fanout1246 (.A(net1247),
    .X(net1246));
 sg13g2_buf_1 fanout1247 (.A(net1264),
    .X(net1247));
 sg13g2_buf_4 fanout1248 (.X(net1248),
    .A(net1254));
 sg13g2_buf_2 fanout1249 (.A(net1254),
    .X(net1249));
 sg13g2_buf_4 fanout1250 (.X(net1250),
    .A(net1254));
 sg13g2_buf_4 fanout1251 (.X(net1251),
    .A(net1253));
 sg13g2_buf_4 fanout1252 (.X(net1252),
    .A(net1253));
 sg13g2_buf_4 fanout1253 (.X(net1253),
    .A(net1254));
 sg13g2_buf_1 fanout1254 (.A(net1264),
    .X(net1254));
 sg13g2_buf_4 fanout1255 (.X(net1255),
    .A(net1258));
 sg13g2_buf_4 fanout1256 (.X(net1256),
    .A(net1257));
 sg13g2_buf_4 fanout1257 (.X(net1257),
    .A(net1258));
 sg13g2_buf_2 fanout1258 (.A(net1264),
    .X(net1258));
 sg13g2_buf_4 fanout1259 (.X(net1259),
    .A(net1263));
 sg13g2_buf_2 fanout1260 (.A(net1263),
    .X(net1260));
 sg13g2_buf_4 fanout1261 (.X(net1261),
    .A(net1263));
 sg13g2_buf_4 fanout1262 (.X(net1262),
    .A(net1263));
 sg13g2_buf_2 fanout1263 (.A(net1264),
    .X(net1263));
 sg13g2_buf_1 fanout1264 (.A(net1265),
    .X(net1264));
 sg13g2_buf_1 fanout1265 (.A(net1),
    .X(net1265));
 sg13g2_buf_4 fanout1266 (.X(net1266),
    .A(net1269));
 sg13g2_buf_4 fanout1267 (.X(net1267),
    .A(net1269));
 sg13g2_buf_4 fanout1268 (.X(net1268),
    .A(net1269));
 sg13g2_buf_2 fanout1269 (.A(net1282),
    .X(net1269));
 sg13g2_buf_4 fanout1270 (.X(net1270),
    .A(net1274));
 sg13g2_buf_2 fanout1271 (.A(net1274),
    .X(net1271));
 sg13g2_buf_4 fanout1272 (.X(net1272),
    .A(net1274));
 sg13g2_buf_2 fanout1273 (.A(net1274),
    .X(net1273));
 sg13g2_buf_1 fanout1274 (.A(net1282),
    .X(net1274));
 sg13g2_buf_4 fanout1275 (.X(net1275),
    .A(net1278));
 sg13g2_buf_4 fanout1276 (.X(net1276),
    .A(net1278));
 sg13g2_buf_2 fanout1277 (.A(net1278),
    .X(net1277));
 sg13g2_buf_2 fanout1278 (.A(net1282),
    .X(net1278));
 sg13g2_buf_4 fanout1279 (.X(net1279),
    .A(net1281));
 sg13g2_buf_4 fanout1280 (.X(net1280),
    .A(net1281));
 sg13g2_buf_2 fanout1281 (.A(net1282),
    .X(net1281));
 sg13g2_buf_1 fanout1282 (.A(net1294),
    .X(net1282));
 sg13g2_buf_4 fanout1283 (.X(net1283),
    .A(net1285));
 sg13g2_buf_4 fanout1284 (.X(net1284),
    .A(net1285));
 sg13g2_buf_4 fanout1285 (.X(net1285),
    .A(net1294));
 sg13g2_buf_4 fanout1286 (.X(net1286),
    .A(net1288));
 sg13g2_buf_4 fanout1287 (.X(net1287),
    .A(net1288));
 sg13g2_buf_4 fanout1288 (.X(net1288),
    .A(net1294));
 sg13g2_buf_4 fanout1289 (.X(net1289),
    .A(net1291));
 sg13g2_buf_2 fanout1290 (.A(net1291),
    .X(net1290));
 sg13g2_buf_2 fanout1291 (.A(net1293),
    .X(net1291));
 sg13g2_buf_4 fanout1292 (.X(net1292),
    .A(net1293));
 sg13g2_buf_2 fanout1293 (.A(net1294),
    .X(net1293));
 sg13g2_buf_1 fanout1294 (.A(net1421),
    .X(net1294));
 sg13g2_buf_4 fanout1295 (.X(net1295),
    .A(net1302));
 sg13g2_buf_2 fanout1296 (.A(net1302),
    .X(net1296));
 sg13g2_buf_4 fanout1297 (.X(net1297),
    .A(net1302));
 sg13g2_buf_4 fanout1298 (.X(net1298),
    .A(net1301));
 sg13g2_buf_4 fanout1299 (.X(net1299),
    .A(net1301));
 sg13g2_buf_2 fanout1300 (.A(net1301),
    .X(net1300));
 sg13g2_buf_2 fanout1301 (.A(net1302),
    .X(net1301));
 sg13g2_buf_1 fanout1302 (.A(net1324),
    .X(net1302));
 sg13g2_buf_4 fanout1303 (.X(net1303),
    .A(net1306));
 sg13g2_buf_4 fanout1304 (.X(net1304),
    .A(net1305));
 sg13g2_buf_4 fanout1305 (.X(net1305),
    .A(net1306));
 sg13g2_buf_2 fanout1306 (.A(net1324),
    .X(net1306));
 sg13g2_buf_4 fanout1307 (.X(net1307),
    .A(net1311));
 sg13g2_buf_2 fanout1308 (.A(net1311),
    .X(net1308));
 sg13g2_buf_4 fanout1309 (.X(net1309),
    .A(net1310));
 sg13g2_buf_4 fanout1310 (.X(net1310),
    .A(net1311));
 sg13g2_buf_1 fanout1311 (.A(net1324),
    .X(net1311));
 sg13g2_buf_4 fanout1312 (.X(net1312),
    .A(net1316));
 sg13g2_buf_4 fanout1313 (.X(net1313),
    .A(net1316));
 sg13g2_buf_4 fanout1314 (.X(net1314),
    .A(net1315));
 sg13g2_buf_4 fanout1315 (.X(net1315),
    .A(net1316));
 sg13g2_buf_4 fanout1316 (.X(net1316),
    .A(net1323));
 sg13g2_buf_4 fanout1317 (.X(net1317),
    .A(net1319));
 sg13g2_buf_4 fanout1318 (.X(net1318),
    .A(net1323));
 sg13g2_buf_2 fanout1319 (.A(net1323),
    .X(net1319));
 sg13g2_buf_4 fanout1320 (.X(net1320),
    .A(net1322));
 sg13g2_buf_4 fanout1321 (.X(net1321),
    .A(net1322));
 sg13g2_buf_4 fanout1322 (.X(net1322),
    .A(net1323));
 sg13g2_buf_1 fanout1323 (.A(net1324),
    .X(net1323));
 sg13g2_buf_1 fanout1324 (.A(net1421),
    .X(net1324));
 sg13g2_buf_4 fanout1325 (.X(net1325),
    .A(net1327));
 sg13g2_buf_4 fanout1326 (.X(net1326),
    .A(net1327));
 sg13g2_buf_2 fanout1327 (.A(net1335),
    .X(net1327));
 sg13g2_buf_4 fanout1328 (.X(net1328),
    .A(net1329));
 sg13g2_buf_4 fanout1329 (.X(net1329),
    .A(net1335));
 sg13g2_buf_4 fanout1330 (.X(net1330),
    .A(net1334));
 sg13g2_buf_4 fanout1331 (.X(net1331),
    .A(net1334));
 sg13g2_buf_4 fanout1332 (.X(net1332),
    .A(net1333));
 sg13g2_buf_4 fanout1333 (.X(net1333),
    .A(net1334));
 sg13g2_buf_1 fanout1334 (.A(net1335),
    .X(net1334));
 sg13g2_buf_1 fanout1335 (.A(net1371),
    .X(net1335));
 sg13g2_buf_4 fanout1336 (.X(net1336),
    .A(net1338));
 sg13g2_buf_2 fanout1337 (.A(net1338),
    .X(net1337));
 sg13g2_buf_2 fanout1338 (.A(net1347),
    .X(net1338));
 sg13g2_buf_4 fanout1339 (.X(net1339),
    .A(net1340));
 sg13g2_buf_4 fanout1340 (.X(net1340),
    .A(net1347));
 sg13g2_buf_4 fanout1341 (.X(net1341),
    .A(net1343));
 sg13g2_buf_4 fanout1342 (.X(net1342),
    .A(net1343));
 sg13g2_buf_2 fanout1343 (.A(net1347),
    .X(net1343));
 sg13g2_buf_4 fanout1344 (.X(net1344),
    .A(net1346));
 sg13g2_buf_4 fanout1345 (.X(net1345),
    .A(net1346));
 sg13g2_buf_2 fanout1346 (.A(net1347),
    .X(net1346));
 sg13g2_buf_1 fanout1347 (.A(net1371),
    .X(net1347));
 sg13g2_buf_4 fanout1348 (.X(net1348),
    .A(net1349));
 sg13g2_buf_4 fanout1349 (.X(net1349),
    .A(net1353));
 sg13g2_buf_2 fanout1350 (.A(net1353),
    .X(net1350));
 sg13g2_buf_4 fanout1351 (.X(net1351),
    .A(net1353));
 sg13g2_buf_4 fanout1352 (.X(net1352),
    .A(net1353));
 sg13g2_buf_2 fanout1353 (.A(net1360),
    .X(net1353));
 sg13g2_buf_4 fanout1354 (.X(net1354),
    .A(net1357));
 sg13g2_buf_4 fanout1355 (.X(net1355),
    .A(net1357));
 sg13g2_buf_2 fanout1356 (.A(net1357),
    .X(net1356));
 sg13g2_buf_2 fanout1357 (.A(net1360),
    .X(net1357));
 sg13g2_buf_4 fanout1358 (.X(net1358),
    .A(net1359));
 sg13g2_buf_4 fanout1359 (.X(net1359),
    .A(net1360));
 sg13g2_buf_1 fanout1360 (.A(net1371),
    .X(net1360));
 sg13g2_buf_4 fanout1361 (.X(net1361),
    .A(net1365));
 sg13g2_buf_2 fanout1362 (.A(net1365),
    .X(net1362));
 sg13g2_buf_4 fanout1363 (.X(net1363),
    .A(net1365));
 sg13g2_buf_4 fanout1364 (.X(net1364),
    .A(net1365));
 sg13g2_buf_1 fanout1365 (.A(net1371),
    .X(net1365));
 sg13g2_buf_4 fanout1366 (.X(net1366),
    .A(net1367));
 sg13g2_buf_4 fanout1367 (.X(net1367),
    .A(net1370));
 sg13g2_buf_4 fanout1368 (.X(net1368),
    .A(net1369));
 sg13g2_buf_4 fanout1369 (.X(net1369),
    .A(net1370));
 sg13g2_buf_2 fanout1370 (.A(net1371),
    .X(net1370));
 sg13g2_buf_1 fanout1371 (.A(net1421),
    .X(net1371));
 sg13g2_buf_4 fanout1372 (.X(net1372),
    .A(net1373));
 sg13g2_buf_4 fanout1373 (.X(net1373),
    .A(net1377));
 sg13g2_buf_4 fanout1374 (.X(net1374),
    .A(net1376));
 sg13g2_buf_2 fanout1375 (.A(net1376),
    .X(net1375));
 sg13g2_buf_4 fanout1376 (.X(net1376),
    .A(net1377));
 sg13g2_buf_2 fanout1377 (.A(net1393),
    .X(net1377));
 sg13g2_buf_4 fanout1378 (.X(net1378),
    .A(net1379));
 sg13g2_buf_4 fanout1379 (.X(net1379),
    .A(net1382));
 sg13g2_buf_4 fanout1380 (.X(net1380),
    .A(net1382));
 sg13g2_buf_2 fanout1381 (.A(net1382),
    .X(net1381));
 sg13g2_buf_2 fanout1382 (.A(net1393),
    .X(net1382));
 sg13g2_buf_4 fanout1383 (.X(net1383),
    .A(net1384));
 sg13g2_buf_4 fanout1384 (.X(net1384),
    .A(net1386));
 sg13g2_buf_4 fanout1385 (.X(net1385),
    .A(net1386));
 sg13g2_buf_2 fanout1386 (.A(net1388),
    .X(net1386));
 sg13g2_buf_4 fanout1387 (.X(net1387),
    .A(net1388));
 sg13g2_buf_2 fanout1388 (.A(net1393),
    .X(net1388));
 sg13g2_buf_4 fanout1389 (.X(net1389),
    .A(net1390));
 sg13g2_buf_4 fanout1390 (.X(net1390),
    .A(net1392));
 sg13g2_buf_4 fanout1391 (.X(net1391),
    .A(net1392));
 sg13g2_buf_2 fanout1392 (.A(net1393),
    .X(net1392));
 sg13g2_buf_1 fanout1393 (.A(net1421),
    .X(net1393));
 sg13g2_buf_4 fanout1394 (.X(net1394),
    .A(net1395));
 sg13g2_buf_4 fanout1395 (.X(net1395),
    .A(net1398));
 sg13g2_buf_4 fanout1396 (.X(net1396),
    .A(net1397));
 sg13g2_buf_4 fanout1397 (.X(net1397),
    .A(net1398));
 sg13g2_buf_2 fanout1398 (.A(net1414),
    .X(net1398));
 sg13g2_buf_4 fanout1399 (.X(net1399),
    .A(net1404));
 sg13g2_buf_4 fanout1400 (.X(net1400),
    .A(net1404));
 sg13g2_buf_4 fanout1401 (.X(net1401),
    .A(net1403));
 sg13g2_buf_4 fanout1402 (.X(net1402),
    .A(net1403));
 sg13g2_buf_2 fanout1403 (.A(net1404),
    .X(net1403));
 sg13g2_buf_2 fanout1404 (.A(net1414),
    .X(net1404));
 sg13g2_buf_4 fanout1405 (.X(net1405),
    .A(net1409));
 sg13g2_buf_2 fanout1406 (.A(net1409),
    .X(net1406));
 sg13g2_buf_4 fanout1407 (.X(net1407),
    .A(net1409));
 sg13g2_buf_2 fanout1408 (.A(net1409),
    .X(net1408));
 sg13g2_buf_1 fanout1409 (.A(net1410),
    .X(net1409));
 sg13g2_buf_2 fanout1410 (.A(net1414),
    .X(net1410));
 sg13g2_buf_4 fanout1411 (.X(net1411),
    .A(net1412));
 sg13g2_buf_4 fanout1412 (.X(net1412),
    .A(net1413));
 sg13g2_buf_4 fanout1413 (.X(net1413),
    .A(net1414));
 sg13g2_buf_2 fanout1414 (.A(net1421),
    .X(net1414));
 sg13g2_buf_4 fanout1415 (.X(net1415),
    .A(net1418));
 sg13g2_buf_4 fanout1416 (.X(net1416),
    .A(net1418));
 sg13g2_buf_2 fanout1417 (.A(net1418),
    .X(net1417));
 sg13g2_buf_1 fanout1418 (.A(net1419),
    .X(net1418));
 sg13g2_buf_4 fanout1419 (.X(net1419),
    .A(net1420));
 sg13g2_buf_2 fanout1420 (.A(net1421),
    .X(net1420));
 sg13g2_buf_2 fanout1421 (.A(net1),
    .X(net1421));
 sg13g2_tiehi _24827__1422 (.L_HI(net1422));
 sg13g2_tiehi _24828__1423 (.L_HI(net1423));
 sg13g2_tiehi _24829__1424 (.L_HI(net1424));
 sg13g2_tiehi _24830__1425 (.L_HI(net1425));
 sg13g2_tiehi _24831__1426 (.L_HI(net1426));
 sg13g2_tiehi _24832__1427 (.L_HI(net1427));
 sg13g2_tiehi _24833__1428 (.L_HI(net1428));
 sg13g2_tiehi _24834__1429 (.L_HI(net1429));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[0]$_DFF_P__1430  (.L_HI(net1430));
 sg13g2_tiehi \top_ihp.oisc.mem_addr_lowbits[1]$_DFF_P__1431  (.L_HI(net1431));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[0]$_DFFE_PP__1432  (.L_HI(net1432));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[1]$_DFFE_PP__1433  (.L_HI(net1433));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[2]$_DFFE_PP__1434  (.L_HI(net1434));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[3]$_DFFE_PP__1435  (.L_HI(net1435));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[4]$_DFFE_PP__1436  (.L_HI(net1436));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[5]$_DFFE_PP__1437  (.L_HI(net1437));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[6]$_DFFE_PP__1438  (.L_HI(net1438));
 sg13g2_tiehi \top_ihp.oisc.micro_pc[7]$_DFFE_PP__1439  (.L_HI(net1439));
 sg13g2_tiehi \top_ihp.oisc.regs[16][0]$_DFFE_PP__1440  (.L_HI(net1440));
 sg13g2_tiehi \top_ihp.oisc.regs[16][10]$_DFFE_PP__1441  (.L_HI(net1441));
 sg13g2_tiehi \top_ihp.oisc.regs[16][11]$_DFFE_PP__1442  (.L_HI(net1442));
 sg13g2_tiehi \top_ihp.oisc.regs[16][12]$_DFFE_PP__1443  (.L_HI(net1443));
 sg13g2_tiehi \top_ihp.oisc.regs[16][13]$_DFFE_PP__1444  (.L_HI(net1444));
 sg13g2_tiehi \top_ihp.oisc.regs[16][14]$_DFFE_PP__1445  (.L_HI(net1445));
 sg13g2_tiehi \top_ihp.oisc.regs[16][15]$_DFFE_PP__1446  (.L_HI(net1446));
 sg13g2_tiehi \top_ihp.oisc.regs[16][16]$_DFFE_PP__1447  (.L_HI(net1447));
 sg13g2_tiehi \top_ihp.oisc.regs[16][17]$_DFFE_PP__1448  (.L_HI(net1448));
 sg13g2_tiehi \top_ihp.oisc.regs[16][18]$_DFFE_PP__1449  (.L_HI(net1449));
 sg13g2_tiehi \top_ihp.oisc.regs[16][19]$_DFFE_PP__1450  (.L_HI(net1450));
 sg13g2_tiehi \top_ihp.oisc.regs[16][1]$_DFFE_PP__1451  (.L_HI(net1451));
 sg13g2_tiehi \top_ihp.oisc.regs[16][20]$_DFFE_PP__1452  (.L_HI(net1452));
 sg13g2_tiehi \top_ihp.oisc.regs[16][21]$_DFFE_PP__1453  (.L_HI(net1453));
 sg13g2_tiehi \top_ihp.oisc.regs[16][22]$_DFFE_PP__1454  (.L_HI(net1454));
 sg13g2_tiehi \top_ihp.oisc.regs[16][23]$_DFFE_PP__1455  (.L_HI(net1455));
 sg13g2_tiehi \top_ihp.oisc.regs[16][24]$_DFFE_PP__1456  (.L_HI(net1456));
 sg13g2_tiehi \top_ihp.oisc.regs[16][25]$_DFFE_PP__1457  (.L_HI(net1457));
 sg13g2_tiehi \top_ihp.oisc.regs[16][26]$_DFFE_PP__1458  (.L_HI(net1458));
 sg13g2_tiehi \top_ihp.oisc.regs[16][27]$_DFFE_PP__1459  (.L_HI(net1459));
 sg13g2_tiehi \top_ihp.oisc.regs[16][28]$_DFFE_PP__1460  (.L_HI(net1460));
 sg13g2_tiehi \top_ihp.oisc.regs[16][29]$_DFFE_PP__1461  (.L_HI(net1461));
 sg13g2_tiehi \top_ihp.oisc.regs[16][2]$_DFFE_PP__1462  (.L_HI(net1462));
 sg13g2_tiehi \top_ihp.oisc.regs[16][30]$_DFFE_PP__1463  (.L_HI(net1463));
 sg13g2_tiehi \top_ihp.oisc.regs[16][31]$_DFFE_PP__1464  (.L_HI(net1464));
 sg13g2_tiehi \top_ihp.oisc.regs[16][3]$_DFFE_PP__1465  (.L_HI(net1465));
 sg13g2_tiehi \top_ihp.oisc.regs[16][4]$_DFFE_PP__1466  (.L_HI(net1466));
 sg13g2_tiehi \top_ihp.oisc.regs[16][5]$_DFFE_PP__1467  (.L_HI(net1467));
 sg13g2_tiehi \top_ihp.oisc.regs[16][6]$_DFFE_PP__1468  (.L_HI(net1468));
 sg13g2_tiehi \top_ihp.oisc.regs[16][7]$_DFFE_PP__1469  (.L_HI(net1469));
 sg13g2_tiehi \top_ihp.oisc.regs[16][8]$_DFFE_PP__1470  (.L_HI(net1470));
 sg13g2_tiehi \top_ihp.oisc.regs[16][9]$_DFFE_PP__1471  (.L_HI(net1471));
 sg13g2_tiehi \top_ihp.oisc.regs[17][0]$_DFFE_PP__1472  (.L_HI(net1472));
 sg13g2_tiehi \top_ihp.oisc.regs[17][10]$_DFFE_PP__1473  (.L_HI(net1473));
 sg13g2_tiehi \top_ihp.oisc.regs[17][11]$_DFFE_PP__1474  (.L_HI(net1474));
 sg13g2_tiehi \top_ihp.oisc.regs[17][12]$_DFFE_PP__1475  (.L_HI(net1475));
 sg13g2_tiehi \top_ihp.oisc.regs[17][13]$_DFFE_PP__1476  (.L_HI(net1476));
 sg13g2_tiehi \top_ihp.oisc.regs[17][14]$_DFFE_PP__1477  (.L_HI(net1477));
 sg13g2_tiehi \top_ihp.oisc.regs[17][15]$_DFFE_PP__1478  (.L_HI(net1478));
 sg13g2_tiehi \top_ihp.oisc.regs[17][16]$_DFFE_PP__1479  (.L_HI(net1479));
 sg13g2_tiehi \top_ihp.oisc.regs[17][17]$_DFFE_PP__1480  (.L_HI(net1480));
 sg13g2_tiehi \top_ihp.oisc.regs[17][18]$_DFFE_PP__1481  (.L_HI(net1481));
 sg13g2_tiehi \top_ihp.oisc.regs[17][19]$_DFFE_PP__1482  (.L_HI(net1482));
 sg13g2_tiehi \top_ihp.oisc.regs[17][1]$_DFFE_PP__1483  (.L_HI(net1483));
 sg13g2_tiehi \top_ihp.oisc.regs[17][20]$_DFFE_PP__1484  (.L_HI(net1484));
 sg13g2_tiehi \top_ihp.oisc.regs[17][21]$_DFFE_PP__1485  (.L_HI(net1485));
 sg13g2_tiehi \top_ihp.oisc.regs[17][22]$_DFFE_PP__1486  (.L_HI(net1486));
 sg13g2_tiehi \top_ihp.oisc.regs[17][23]$_DFFE_PP__1487  (.L_HI(net1487));
 sg13g2_tiehi \top_ihp.oisc.regs[17][24]$_DFFE_PP__1488  (.L_HI(net1488));
 sg13g2_tiehi \top_ihp.oisc.regs[17][25]$_DFFE_PP__1489  (.L_HI(net1489));
 sg13g2_tiehi \top_ihp.oisc.regs[17][26]$_DFFE_PP__1490  (.L_HI(net1490));
 sg13g2_tiehi \top_ihp.oisc.regs[17][27]$_DFFE_PP__1491  (.L_HI(net1491));
 sg13g2_tiehi \top_ihp.oisc.regs[17][28]$_DFFE_PP__1492  (.L_HI(net1492));
 sg13g2_tiehi \top_ihp.oisc.regs[17][29]$_DFFE_PP__1493  (.L_HI(net1493));
 sg13g2_tiehi \top_ihp.oisc.regs[17][2]$_DFFE_PP__1494  (.L_HI(net1494));
 sg13g2_tiehi \top_ihp.oisc.regs[17][30]$_DFFE_PP__1495  (.L_HI(net1495));
 sg13g2_tiehi \top_ihp.oisc.regs[17][31]$_DFFE_PP__1496  (.L_HI(net1496));
 sg13g2_tiehi \top_ihp.oisc.regs[17][3]$_DFFE_PP__1497  (.L_HI(net1497));
 sg13g2_tiehi \top_ihp.oisc.regs[17][4]$_DFFE_PP__1498  (.L_HI(net1498));
 sg13g2_tiehi \top_ihp.oisc.regs[17][5]$_DFFE_PP__1499  (.L_HI(net1499));
 sg13g2_tiehi \top_ihp.oisc.regs[17][6]$_DFFE_PP__1500  (.L_HI(net1500));
 sg13g2_tiehi \top_ihp.oisc.regs[17][7]$_DFFE_PP__1501  (.L_HI(net1501));
 sg13g2_tiehi \top_ihp.oisc.regs[17][8]$_DFFE_PP__1502  (.L_HI(net1502));
 sg13g2_tiehi \top_ihp.oisc.regs[17][9]$_DFFE_PP__1503  (.L_HI(net1503));
 sg13g2_tiehi \top_ihp.oisc.regs[18][0]$_DFFE_PP__1504  (.L_HI(net1504));
 sg13g2_tiehi \top_ihp.oisc.regs[18][10]$_DFFE_PP__1505  (.L_HI(net1505));
 sg13g2_tiehi \top_ihp.oisc.regs[18][11]$_DFFE_PP__1506  (.L_HI(net1506));
 sg13g2_tiehi \top_ihp.oisc.regs[18][12]$_DFFE_PP__1507  (.L_HI(net1507));
 sg13g2_tiehi \top_ihp.oisc.regs[18][13]$_DFFE_PP__1508  (.L_HI(net1508));
 sg13g2_tiehi \top_ihp.oisc.regs[18][14]$_DFFE_PP__1509  (.L_HI(net1509));
 sg13g2_tiehi \top_ihp.oisc.regs[18][15]$_DFFE_PP__1510  (.L_HI(net1510));
 sg13g2_tiehi \top_ihp.oisc.regs[18][16]$_DFFE_PP__1511  (.L_HI(net1511));
 sg13g2_tiehi \top_ihp.oisc.regs[18][17]$_DFFE_PP__1512  (.L_HI(net1512));
 sg13g2_tiehi \top_ihp.oisc.regs[18][18]$_DFFE_PP__1513  (.L_HI(net1513));
 sg13g2_tiehi \top_ihp.oisc.regs[18][19]$_DFFE_PP__1514  (.L_HI(net1514));
 sg13g2_tiehi \top_ihp.oisc.regs[18][1]$_DFFE_PP__1515  (.L_HI(net1515));
 sg13g2_tiehi \top_ihp.oisc.regs[18][20]$_DFFE_PP__1516  (.L_HI(net1516));
 sg13g2_tiehi \top_ihp.oisc.regs[18][21]$_DFFE_PP__1517  (.L_HI(net1517));
 sg13g2_tiehi \top_ihp.oisc.regs[18][22]$_DFFE_PP__1518  (.L_HI(net1518));
 sg13g2_tiehi \top_ihp.oisc.regs[18][23]$_DFFE_PP__1519  (.L_HI(net1519));
 sg13g2_tiehi \top_ihp.oisc.regs[18][24]$_DFFE_PP__1520  (.L_HI(net1520));
 sg13g2_tiehi \top_ihp.oisc.regs[18][25]$_DFFE_PP__1521  (.L_HI(net1521));
 sg13g2_tiehi \top_ihp.oisc.regs[18][26]$_DFFE_PP__1522  (.L_HI(net1522));
 sg13g2_tiehi \top_ihp.oisc.regs[18][27]$_DFFE_PP__1523  (.L_HI(net1523));
 sg13g2_tiehi \top_ihp.oisc.regs[18][28]$_DFFE_PP__1524  (.L_HI(net1524));
 sg13g2_tiehi \top_ihp.oisc.regs[18][29]$_DFFE_PP__1525  (.L_HI(net1525));
 sg13g2_tiehi \top_ihp.oisc.regs[18][2]$_DFFE_PP__1526  (.L_HI(net1526));
 sg13g2_tiehi \top_ihp.oisc.regs[18][30]$_DFFE_PP__1527  (.L_HI(net1527));
 sg13g2_tiehi \top_ihp.oisc.regs[18][31]$_DFFE_PP__1528  (.L_HI(net1528));
 sg13g2_tiehi \top_ihp.oisc.regs[18][3]$_DFFE_PP__1529  (.L_HI(net1529));
 sg13g2_tiehi \top_ihp.oisc.regs[18][4]$_DFFE_PP__1530  (.L_HI(net1530));
 sg13g2_tiehi \top_ihp.oisc.regs[18][5]$_DFFE_PP__1531  (.L_HI(net1531));
 sg13g2_tiehi \top_ihp.oisc.regs[18][6]$_DFFE_PP__1532  (.L_HI(net1532));
 sg13g2_tiehi \top_ihp.oisc.regs[18][7]$_DFFE_PP__1533  (.L_HI(net1533));
 sg13g2_tiehi \top_ihp.oisc.regs[18][8]$_DFFE_PP__1534  (.L_HI(net1534));
 sg13g2_tiehi \top_ihp.oisc.regs[18][9]$_DFFE_PP__1535  (.L_HI(net1535));
 sg13g2_tiehi \top_ihp.oisc.regs[19][0]$_DFFE_PP__1536  (.L_HI(net1536));
 sg13g2_tiehi \top_ihp.oisc.regs[19][10]$_DFFE_PP__1537  (.L_HI(net1537));
 sg13g2_tiehi \top_ihp.oisc.regs[19][11]$_DFFE_PP__1538  (.L_HI(net1538));
 sg13g2_tiehi \top_ihp.oisc.regs[19][12]$_DFFE_PP__1539  (.L_HI(net1539));
 sg13g2_tiehi \top_ihp.oisc.regs[19][13]$_DFFE_PP__1540  (.L_HI(net1540));
 sg13g2_tiehi \top_ihp.oisc.regs[19][14]$_DFFE_PP__1541  (.L_HI(net1541));
 sg13g2_tiehi \top_ihp.oisc.regs[19][15]$_DFFE_PP__1542  (.L_HI(net1542));
 sg13g2_tiehi \top_ihp.oisc.regs[19][16]$_DFFE_PP__1543  (.L_HI(net1543));
 sg13g2_tiehi \top_ihp.oisc.regs[19][17]$_DFFE_PP__1544  (.L_HI(net1544));
 sg13g2_tiehi \top_ihp.oisc.regs[19][18]$_DFFE_PP__1545  (.L_HI(net1545));
 sg13g2_tiehi \top_ihp.oisc.regs[19][19]$_DFFE_PP__1546  (.L_HI(net1546));
 sg13g2_tiehi \top_ihp.oisc.regs[19][1]$_DFFE_PP__1547  (.L_HI(net1547));
 sg13g2_tiehi \top_ihp.oisc.regs[19][20]$_DFFE_PP__1548  (.L_HI(net1548));
 sg13g2_tiehi \top_ihp.oisc.regs[19][21]$_DFFE_PP__1549  (.L_HI(net1549));
 sg13g2_tiehi \top_ihp.oisc.regs[19][22]$_DFFE_PP__1550  (.L_HI(net1550));
 sg13g2_tiehi \top_ihp.oisc.regs[19][23]$_DFFE_PP__1551  (.L_HI(net1551));
 sg13g2_tiehi \top_ihp.oisc.regs[19][24]$_DFFE_PP__1552  (.L_HI(net1552));
 sg13g2_tiehi \top_ihp.oisc.regs[19][25]$_DFFE_PP__1553  (.L_HI(net1553));
 sg13g2_tiehi \top_ihp.oisc.regs[19][26]$_DFFE_PP__1554  (.L_HI(net1554));
 sg13g2_tiehi \top_ihp.oisc.regs[19][27]$_DFFE_PP__1555  (.L_HI(net1555));
 sg13g2_tiehi \top_ihp.oisc.regs[19][28]$_DFFE_PP__1556  (.L_HI(net1556));
 sg13g2_tiehi \top_ihp.oisc.regs[19][29]$_DFFE_PP__1557  (.L_HI(net1557));
 sg13g2_tiehi \top_ihp.oisc.regs[19][2]$_DFFE_PP__1558  (.L_HI(net1558));
 sg13g2_tiehi \top_ihp.oisc.regs[19][30]$_DFFE_PP__1559  (.L_HI(net1559));
 sg13g2_tiehi \top_ihp.oisc.regs[19][31]$_DFFE_PP__1560  (.L_HI(net1560));
 sg13g2_tiehi \top_ihp.oisc.regs[19][3]$_DFFE_PP__1561  (.L_HI(net1561));
 sg13g2_tiehi \top_ihp.oisc.regs[19][4]$_DFFE_PP__1562  (.L_HI(net1562));
 sg13g2_tiehi \top_ihp.oisc.regs[19][5]$_DFFE_PP__1563  (.L_HI(net1563));
 sg13g2_tiehi \top_ihp.oisc.regs[19][6]$_DFFE_PP__1564  (.L_HI(net1564));
 sg13g2_tiehi \top_ihp.oisc.regs[19][7]$_DFFE_PP__1565  (.L_HI(net1565));
 sg13g2_tiehi \top_ihp.oisc.regs[19][8]$_DFFE_PP__1566  (.L_HI(net1566));
 sg13g2_tiehi \top_ihp.oisc.regs[19][9]$_DFFE_PP__1567  (.L_HI(net1567));
 sg13g2_tiehi \top_ihp.oisc.regs[20][0]$_DFFE_PP__1568  (.L_HI(net1568));
 sg13g2_tiehi \top_ihp.oisc.regs[20][10]$_DFFE_PP__1569  (.L_HI(net1569));
 sg13g2_tiehi \top_ihp.oisc.regs[20][11]$_DFFE_PP__1570  (.L_HI(net1570));
 sg13g2_tiehi \top_ihp.oisc.regs[20][12]$_DFFE_PP__1571  (.L_HI(net1571));
 sg13g2_tiehi \top_ihp.oisc.regs[20][13]$_DFFE_PP__1572  (.L_HI(net1572));
 sg13g2_tiehi \top_ihp.oisc.regs[20][14]$_DFFE_PP__1573  (.L_HI(net1573));
 sg13g2_tiehi \top_ihp.oisc.regs[20][15]$_DFFE_PP__1574  (.L_HI(net1574));
 sg13g2_tiehi \top_ihp.oisc.regs[20][16]$_DFFE_PP__1575  (.L_HI(net1575));
 sg13g2_tiehi \top_ihp.oisc.regs[20][17]$_DFFE_PP__1576  (.L_HI(net1576));
 sg13g2_tiehi \top_ihp.oisc.regs[20][18]$_DFFE_PP__1577  (.L_HI(net1577));
 sg13g2_tiehi \top_ihp.oisc.regs[20][19]$_DFFE_PP__1578  (.L_HI(net1578));
 sg13g2_tiehi \top_ihp.oisc.regs[20][1]$_DFFE_PP__1579  (.L_HI(net1579));
 sg13g2_tiehi \top_ihp.oisc.regs[20][20]$_DFFE_PP__1580  (.L_HI(net1580));
 sg13g2_tiehi \top_ihp.oisc.regs[20][21]$_DFFE_PP__1581  (.L_HI(net1581));
 sg13g2_tiehi \top_ihp.oisc.regs[20][22]$_DFFE_PP__1582  (.L_HI(net1582));
 sg13g2_tiehi \top_ihp.oisc.regs[20][23]$_DFFE_PP__1583  (.L_HI(net1583));
 sg13g2_tiehi \top_ihp.oisc.regs[20][24]$_DFFE_PP__1584  (.L_HI(net1584));
 sg13g2_tiehi \top_ihp.oisc.regs[20][25]$_DFFE_PP__1585  (.L_HI(net1585));
 sg13g2_tiehi \top_ihp.oisc.regs[20][26]$_DFFE_PP__1586  (.L_HI(net1586));
 sg13g2_tiehi \top_ihp.oisc.regs[20][27]$_DFFE_PP__1587  (.L_HI(net1587));
 sg13g2_tiehi \top_ihp.oisc.regs[20][28]$_DFFE_PP__1588  (.L_HI(net1588));
 sg13g2_tiehi \top_ihp.oisc.regs[20][29]$_DFFE_PP__1589  (.L_HI(net1589));
 sg13g2_tiehi \top_ihp.oisc.regs[20][2]$_DFFE_PP__1590  (.L_HI(net1590));
 sg13g2_tiehi \top_ihp.oisc.regs[20][30]$_DFFE_PP__1591  (.L_HI(net1591));
 sg13g2_tiehi \top_ihp.oisc.regs[20][31]$_DFFE_PP__1592  (.L_HI(net1592));
 sg13g2_tiehi \top_ihp.oisc.regs[20][3]$_DFFE_PP__1593  (.L_HI(net1593));
 sg13g2_tiehi \top_ihp.oisc.regs[20][4]$_DFFE_PP__1594  (.L_HI(net1594));
 sg13g2_tiehi \top_ihp.oisc.regs[20][5]$_DFFE_PP__1595  (.L_HI(net1595));
 sg13g2_tiehi \top_ihp.oisc.regs[20][6]$_DFFE_PP__1596  (.L_HI(net1596));
 sg13g2_tiehi \top_ihp.oisc.regs[20][7]$_DFFE_PP__1597  (.L_HI(net1597));
 sg13g2_tiehi \top_ihp.oisc.regs[20][8]$_DFFE_PP__1598  (.L_HI(net1598));
 sg13g2_tiehi \top_ihp.oisc.regs[20][9]$_DFFE_PP__1599  (.L_HI(net1599));
 sg13g2_tiehi \top_ihp.oisc.regs[21][0]$_DFFE_PP__1600  (.L_HI(net1600));
 sg13g2_tiehi \top_ihp.oisc.regs[21][10]$_DFFE_PP__1601  (.L_HI(net1601));
 sg13g2_tiehi \top_ihp.oisc.regs[21][11]$_DFFE_PP__1602  (.L_HI(net1602));
 sg13g2_tiehi \top_ihp.oisc.regs[21][12]$_DFFE_PP__1603  (.L_HI(net1603));
 sg13g2_tiehi \top_ihp.oisc.regs[21][13]$_DFFE_PP__1604  (.L_HI(net1604));
 sg13g2_tiehi \top_ihp.oisc.regs[21][14]$_DFFE_PP__1605  (.L_HI(net1605));
 sg13g2_tiehi \top_ihp.oisc.regs[21][15]$_DFFE_PP__1606  (.L_HI(net1606));
 sg13g2_tiehi \top_ihp.oisc.regs[21][16]$_DFFE_PP__1607  (.L_HI(net1607));
 sg13g2_tiehi \top_ihp.oisc.regs[21][17]$_DFFE_PP__1608  (.L_HI(net1608));
 sg13g2_tiehi \top_ihp.oisc.regs[21][18]$_DFFE_PP__1609  (.L_HI(net1609));
 sg13g2_tiehi \top_ihp.oisc.regs[21][19]$_DFFE_PP__1610  (.L_HI(net1610));
 sg13g2_tiehi \top_ihp.oisc.regs[21][1]$_DFFE_PP__1611  (.L_HI(net1611));
 sg13g2_tiehi \top_ihp.oisc.regs[21][20]$_DFFE_PP__1612  (.L_HI(net1612));
 sg13g2_tiehi \top_ihp.oisc.regs[21][21]$_DFFE_PP__1613  (.L_HI(net1613));
 sg13g2_tiehi \top_ihp.oisc.regs[21][22]$_DFFE_PP__1614  (.L_HI(net1614));
 sg13g2_tiehi \top_ihp.oisc.regs[21][23]$_DFFE_PP__1615  (.L_HI(net1615));
 sg13g2_tiehi \top_ihp.oisc.regs[21][24]$_DFFE_PP__1616  (.L_HI(net1616));
 sg13g2_tiehi \top_ihp.oisc.regs[21][25]$_DFFE_PP__1617  (.L_HI(net1617));
 sg13g2_tiehi \top_ihp.oisc.regs[21][26]$_DFFE_PP__1618  (.L_HI(net1618));
 sg13g2_tiehi \top_ihp.oisc.regs[21][27]$_DFFE_PP__1619  (.L_HI(net1619));
 sg13g2_tiehi \top_ihp.oisc.regs[21][28]$_DFFE_PP__1620  (.L_HI(net1620));
 sg13g2_tiehi \top_ihp.oisc.regs[21][29]$_DFFE_PP__1621  (.L_HI(net1621));
 sg13g2_tiehi \top_ihp.oisc.regs[21][2]$_DFFE_PP__1622  (.L_HI(net1622));
 sg13g2_tiehi \top_ihp.oisc.regs[21][30]$_DFFE_PP__1623  (.L_HI(net1623));
 sg13g2_tiehi \top_ihp.oisc.regs[21][31]$_DFFE_PP__1624  (.L_HI(net1624));
 sg13g2_tiehi \top_ihp.oisc.regs[21][3]$_DFFE_PP__1625  (.L_HI(net1625));
 sg13g2_tiehi \top_ihp.oisc.regs[21][4]$_DFFE_PP__1626  (.L_HI(net1626));
 sg13g2_tiehi \top_ihp.oisc.regs[21][5]$_DFFE_PP__1627  (.L_HI(net1627));
 sg13g2_tiehi \top_ihp.oisc.regs[21][6]$_DFFE_PP__1628  (.L_HI(net1628));
 sg13g2_tiehi \top_ihp.oisc.regs[21][7]$_DFFE_PP__1629  (.L_HI(net1629));
 sg13g2_tiehi \top_ihp.oisc.regs[21][8]$_DFFE_PP__1630  (.L_HI(net1630));
 sg13g2_tiehi \top_ihp.oisc.regs[21][9]$_DFFE_PP__1631  (.L_HI(net1631));
 sg13g2_tiehi \top_ihp.oisc.regs[22][0]$_DFFE_PP__1632  (.L_HI(net1632));
 sg13g2_tiehi \top_ihp.oisc.regs[22][10]$_DFFE_PP__1633  (.L_HI(net1633));
 sg13g2_tiehi \top_ihp.oisc.regs[22][11]$_DFFE_PP__1634  (.L_HI(net1634));
 sg13g2_tiehi \top_ihp.oisc.regs[22][12]$_DFFE_PP__1635  (.L_HI(net1635));
 sg13g2_tiehi \top_ihp.oisc.regs[22][13]$_DFFE_PP__1636  (.L_HI(net1636));
 sg13g2_tiehi \top_ihp.oisc.regs[22][14]$_DFFE_PP__1637  (.L_HI(net1637));
 sg13g2_tiehi \top_ihp.oisc.regs[22][15]$_DFFE_PP__1638  (.L_HI(net1638));
 sg13g2_tiehi \top_ihp.oisc.regs[22][16]$_DFFE_PP__1639  (.L_HI(net1639));
 sg13g2_tiehi \top_ihp.oisc.regs[22][17]$_DFFE_PP__1640  (.L_HI(net1640));
 sg13g2_tiehi \top_ihp.oisc.regs[22][18]$_DFFE_PP__1641  (.L_HI(net1641));
 sg13g2_tiehi \top_ihp.oisc.regs[22][19]$_DFFE_PP__1642  (.L_HI(net1642));
 sg13g2_tiehi \top_ihp.oisc.regs[22][1]$_DFFE_PP__1643  (.L_HI(net1643));
 sg13g2_tiehi \top_ihp.oisc.regs[22][20]$_DFFE_PP__1644  (.L_HI(net1644));
 sg13g2_tiehi \top_ihp.oisc.regs[22][21]$_DFFE_PP__1645  (.L_HI(net1645));
 sg13g2_tiehi \top_ihp.oisc.regs[22][22]$_DFFE_PP__1646  (.L_HI(net1646));
 sg13g2_tiehi \top_ihp.oisc.regs[22][23]$_DFFE_PP__1647  (.L_HI(net1647));
 sg13g2_tiehi \top_ihp.oisc.regs[22][24]$_DFFE_PP__1648  (.L_HI(net1648));
 sg13g2_tiehi \top_ihp.oisc.regs[22][25]$_DFFE_PP__1649  (.L_HI(net1649));
 sg13g2_tiehi \top_ihp.oisc.regs[22][26]$_DFFE_PP__1650  (.L_HI(net1650));
 sg13g2_tiehi \top_ihp.oisc.regs[22][27]$_DFFE_PP__1651  (.L_HI(net1651));
 sg13g2_tiehi \top_ihp.oisc.regs[22][28]$_DFFE_PP__1652  (.L_HI(net1652));
 sg13g2_tiehi \top_ihp.oisc.regs[22][29]$_DFFE_PP__1653  (.L_HI(net1653));
 sg13g2_tiehi \top_ihp.oisc.regs[22][2]$_DFFE_PP__1654  (.L_HI(net1654));
 sg13g2_tiehi \top_ihp.oisc.regs[22][30]$_DFFE_PP__1655  (.L_HI(net1655));
 sg13g2_tiehi \top_ihp.oisc.regs[22][31]$_DFFE_PP__1656  (.L_HI(net1656));
 sg13g2_tiehi \top_ihp.oisc.regs[22][3]$_DFFE_PP__1657  (.L_HI(net1657));
 sg13g2_tiehi \top_ihp.oisc.regs[22][4]$_DFFE_PP__1658  (.L_HI(net1658));
 sg13g2_tiehi \top_ihp.oisc.regs[22][5]$_DFFE_PP__1659  (.L_HI(net1659));
 sg13g2_tiehi \top_ihp.oisc.regs[22][6]$_DFFE_PP__1660  (.L_HI(net1660));
 sg13g2_tiehi \top_ihp.oisc.regs[22][7]$_DFFE_PP__1661  (.L_HI(net1661));
 sg13g2_tiehi \top_ihp.oisc.regs[22][8]$_DFFE_PP__1662  (.L_HI(net1662));
 sg13g2_tiehi \top_ihp.oisc.regs[22][9]$_DFFE_PP__1663  (.L_HI(net1663));
 sg13g2_tiehi \top_ihp.oisc.regs[23][0]$_DFFE_PP__1664  (.L_HI(net1664));
 sg13g2_tiehi \top_ihp.oisc.regs[23][10]$_DFFE_PP__1665  (.L_HI(net1665));
 sg13g2_tiehi \top_ihp.oisc.regs[23][11]$_DFFE_PP__1666  (.L_HI(net1666));
 sg13g2_tiehi \top_ihp.oisc.regs[23][12]$_DFFE_PP__1667  (.L_HI(net1667));
 sg13g2_tiehi \top_ihp.oisc.regs[23][13]$_DFFE_PP__1668  (.L_HI(net1668));
 sg13g2_tiehi \top_ihp.oisc.regs[23][14]$_DFFE_PP__1669  (.L_HI(net1669));
 sg13g2_tiehi \top_ihp.oisc.regs[23][15]$_DFFE_PP__1670  (.L_HI(net1670));
 sg13g2_tiehi \top_ihp.oisc.regs[23][16]$_DFFE_PP__1671  (.L_HI(net1671));
 sg13g2_tiehi \top_ihp.oisc.regs[23][17]$_DFFE_PP__1672  (.L_HI(net1672));
 sg13g2_tiehi \top_ihp.oisc.regs[23][18]$_DFFE_PP__1673  (.L_HI(net1673));
 sg13g2_tiehi \top_ihp.oisc.regs[23][19]$_DFFE_PP__1674  (.L_HI(net1674));
 sg13g2_tiehi \top_ihp.oisc.regs[23][1]$_DFFE_PP__1675  (.L_HI(net1675));
 sg13g2_tiehi \top_ihp.oisc.regs[23][20]$_DFFE_PP__1676  (.L_HI(net1676));
 sg13g2_tiehi \top_ihp.oisc.regs[23][21]$_DFFE_PP__1677  (.L_HI(net1677));
 sg13g2_tiehi \top_ihp.oisc.regs[23][22]$_DFFE_PP__1678  (.L_HI(net1678));
 sg13g2_tiehi \top_ihp.oisc.regs[23][23]$_DFFE_PP__1679  (.L_HI(net1679));
 sg13g2_tiehi \top_ihp.oisc.regs[23][24]$_DFFE_PP__1680  (.L_HI(net1680));
 sg13g2_tiehi \top_ihp.oisc.regs[23][25]$_DFFE_PP__1681  (.L_HI(net1681));
 sg13g2_tiehi \top_ihp.oisc.regs[23][26]$_DFFE_PP__1682  (.L_HI(net1682));
 sg13g2_tiehi \top_ihp.oisc.regs[23][27]$_DFFE_PP__1683  (.L_HI(net1683));
 sg13g2_tiehi \top_ihp.oisc.regs[23][28]$_DFFE_PP__1684  (.L_HI(net1684));
 sg13g2_tiehi \top_ihp.oisc.regs[23][29]$_DFFE_PP__1685  (.L_HI(net1685));
 sg13g2_tiehi \top_ihp.oisc.regs[23][2]$_DFFE_PP__1686  (.L_HI(net1686));
 sg13g2_tiehi \top_ihp.oisc.regs[23][30]$_DFFE_PP__1687  (.L_HI(net1687));
 sg13g2_tiehi \top_ihp.oisc.regs[23][31]$_DFFE_PP__1688  (.L_HI(net1688));
 sg13g2_tiehi \top_ihp.oisc.regs[23][3]$_DFFE_PP__1689  (.L_HI(net1689));
 sg13g2_tiehi \top_ihp.oisc.regs[23][4]$_DFFE_PP__1690  (.L_HI(net1690));
 sg13g2_tiehi \top_ihp.oisc.regs[23][5]$_DFFE_PP__1691  (.L_HI(net1691));
 sg13g2_tiehi \top_ihp.oisc.regs[23][6]$_DFFE_PP__1692  (.L_HI(net1692));
 sg13g2_tiehi \top_ihp.oisc.regs[23][7]$_DFFE_PP__1693  (.L_HI(net1693));
 sg13g2_tiehi \top_ihp.oisc.regs[23][8]$_DFFE_PP__1694  (.L_HI(net1694));
 sg13g2_tiehi \top_ihp.oisc.regs[23][9]$_DFFE_PP__1695  (.L_HI(net1695));
 sg13g2_tiehi \top_ihp.oisc.regs[24][0]$_DFFE_PP__1696  (.L_HI(net1696));
 sg13g2_tiehi \top_ihp.oisc.regs[24][10]$_DFFE_PP__1697  (.L_HI(net1697));
 sg13g2_tiehi \top_ihp.oisc.regs[24][11]$_DFFE_PP__1698  (.L_HI(net1698));
 sg13g2_tiehi \top_ihp.oisc.regs[24][12]$_DFFE_PP__1699  (.L_HI(net1699));
 sg13g2_tiehi \top_ihp.oisc.regs[24][13]$_DFFE_PP__1700  (.L_HI(net1700));
 sg13g2_tiehi \top_ihp.oisc.regs[24][14]$_DFFE_PP__1701  (.L_HI(net1701));
 sg13g2_tiehi \top_ihp.oisc.regs[24][15]$_DFFE_PP__1702  (.L_HI(net1702));
 sg13g2_tiehi \top_ihp.oisc.regs[24][16]$_DFFE_PP__1703  (.L_HI(net1703));
 sg13g2_tiehi \top_ihp.oisc.regs[24][17]$_DFFE_PP__1704  (.L_HI(net1704));
 sg13g2_tiehi \top_ihp.oisc.regs[24][18]$_DFFE_PP__1705  (.L_HI(net1705));
 sg13g2_tiehi \top_ihp.oisc.regs[24][19]$_DFFE_PP__1706  (.L_HI(net1706));
 sg13g2_tiehi \top_ihp.oisc.regs[24][1]$_DFFE_PP__1707  (.L_HI(net1707));
 sg13g2_tiehi \top_ihp.oisc.regs[24][20]$_DFFE_PP__1708  (.L_HI(net1708));
 sg13g2_tiehi \top_ihp.oisc.regs[24][21]$_DFFE_PP__1709  (.L_HI(net1709));
 sg13g2_tiehi \top_ihp.oisc.regs[24][22]$_DFFE_PP__1710  (.L_HI(net1710));
 sg13g2_tiehi \top_ihp.oisc.regs[24][23]$_DFFE_PP__1711  (.L_HI(net1711));
 sg13g2_tiehi \top_ihp.oisc.regs[24][24]$_DFFE_PP__1712  (.L_HI(net1712));
 sg13g2_tiehi \top_ihp.oisc.regs[24][25]$_DFFE_PP__1713  (.L_HI(net1713));
 sg13g2_tiehi \top_ihp.oisc.regs[24][26]$_DFFE_PP__1714  (.L_HI(net1714));
 sg13g2_tiehi \top_ihp.oisc.regs[24][27]$_DFFE_PP__1715  (.L_HI(net1715));
 sg13g2_tiehi \top_ihp.oisc.regs[24][28]$_DFFE_PP__1716  (.L_HI(net1716));
 sg13g2_tiehi \top_ihp.oisc.regs[24][29]$_DFFE_PP__1717  (.L_HI(net1717));
 sg13g2_tiehi \top_ihp.oisc.regs[24][2]$_DFFE_PP__1718  (.L_HI(net1718));
 sg13g2_tiehi \top_ihp.oisc.regs[24][30]$_DFFE_PP__1719  (.L_HI(net1719));
 sg13g2_tiehi \top_ihp.oisc.regs[24][31]$_DFFE_PP__1720  (.L_HI(net1720));
 sg13g2_tiehi \top_ihp.oisc.regs[24][3]$_DFFE_PP__1721  (.L_HI(net1721));
 sg13g2_tiehi \top_ihp.oisc.regs[24][4]$_DFFE_PP__1722  (.L_HI(net1722));
 sg13g2_tiehi \top_ihp.oisc.regs[24][5]$_DFFE_PP__1723  (.L_HI(net1723));
 sg13g2_tiehi \top_ihp.oisc.regs[24][6]$_DFFE_PP__1724  (.L_HI(net1724));
 sg13g2_tiehi \top_ihp.oisc.regs[24][7]$_DFFE_PP__1725  (.L_HI(net1725));
 sg13g2_tiehi \top_ihp.oisc.regs[24][8]$_DFFE_PP__1726  (.L_HI(net1726));
 sg13g2_tiehi \top_ihp.oisc.regs[24][9]$_DFFE_PP__1727  (.L_HI(net1727));
 sg13g2_tiehi \top_ihp.oisc.regs[25][0]$_DFFE_PP__1728  (.L_HI(net1728));
 sg13g2_tiehi \top_ihp.oisc.regs[25][10]$_DFFE_PP__1729  (.L_HI(net1729));
 sg13g2_tiehi \top_ihp.oisc.regs[25][11]$_DFFE_PP__1730  (.L_HI(net1730));
 sg13g2_tiehi \top_ihp.oisc.regs[25][12]$_DFFE_PP__1731  (.L_HI(net1731));
 sg13g2_tiehi \top_ihp.oisc.regs[25][13]$_DFFE_PP__1732  (.L_HI(net1732));
 sg13g2_tiehi \top_ihp.oisc.regs[25][14]$_DFFE_PP__1733  (.L_HI(net1733));
 sg13g2_tiehi \top_ihp.oisc.regs[25][15]$_DFFE_PP__1734  (.L_HI(net1734));
 sg13g2_tiehi \top_ihp.oisc.regs[25][16]$_DFFE_PP__1735  (.L_HI(net1735));
 sg13g2_tiehi \top_ihp.oisc.regs[25][17]$_DFFE_PP__1736  (.L_HI(net1736));
 sg13g2_tiehi \top_ihp.oisc.regs[25][18]$_DFFE_PP__1737  (.L_HI(net1737));
 sg13g2_tiehi \top_ihp.oisc.regs[25][19]$_DFFE_PP__1738  (.L_HI(net1738));
 sg13g2_tiehi \top_ihp.oisc.regs[25][1]$_DFFE_PP__1739  (.L_HI(net1739));
 sg13g2_tiehi \top_ihp.oisc.regs[25][20]$_DFFE_PP__1740  (.L_HI(net1740));
 sg13g2_tiehi \top_ihp.oisc.regs[25][21]$_DFFE_PP__1741  (.L_HI(net1741));
 sg13g2_tiehi \top_ihp.oisc.regs[25][22]$_DFFE_PP__1742  (.L_HI(net1742));
 sg13g2_tiehi \top_ihp.oisc.regs[25][23]$_DFFE_PP__1743  (.L_HI(net1743));
 sg13g2_tiehi \top_ihp.oisc.regs[25][24]$_DFFE_PP__1744  (.L_HI(net1744));
 sg13g2_tiehi \top_ihp.oisc.regs[25][25]$_DFFE_PP__1745  (.L_HI(net1745));
 sg13g2_tiehi \top_ihp.oisc.regs[25][26]$_DFFE_PP__1746  (.L_HI(net1746));
 sg13g2_tiehi \top_ihp.oisc.regs[25][27]$_DFFE_PP__1747  (.L_HI(net1747));
 sg13g2_tiehi \top_ihp.oisc.regs[25][28]$_DFFE_PP__1748  (.L_HI(net1748));
 sg13g2_tiehi \top_ihp.oisc.regs[25][29]$_DFFE_PP__1749  (.L_HI(net1749));
 sg13g2_tiehi \top_ihp.oisc.regs[25][2]$_DFFE_PP__1750  (.L_HI(net1750));
 sg13g2_tiehi \top_ihp.oisc.regs[25][30]$_DFFE_PP__1751  (.L_HI(net1751));
 sg13g2_tiehi \top_ihp.oisc.regs[25][31]$_DFFE_PP__1752  (.L_HI(net1752));
 sg13g2_tiehi \top_ihp.oisc.regs[25][3]$_DFFE_PP__1753  (.L_HI(net1753));
 sg13g2_tiehi \top_ihp.oisc.regs[25][4]$_DFFE_PP__1754  (.L_HI(net1754));
 sg13g2_tiehi \top_ihp.oisc.regs[25][5]$_DFFE_PP__1755  (.L_HI(net1755));
 sg13g2_tiehi \top_ihp.oisc.regs[25][6]$_DFFE_PP__1756  (.L_HI(net1756));
 sg13g2_tiehi \top_ihp.oisc.regs[25][7]$_DFFE_PP__1757  (.L_HI(net1757));
 sg13g2_tiehi \top_ihp.oisc.regs[25][8]$_DFFE_PP__1758  (.L_HI(net1758));
 sg13g2_tiehi \top_ihp.oisc.regs[25][9]$_DFFE_PP__1759  (.L_HI(net1759));
 sg13g2_tiehi \top_ihp.oisc.regs[26][0]$_DFFE_PP__1760  (.L_HI(net1760));
 sg13g2_tiehi \top_ihp.oisc.regs[26][10]$_DFFE_PP__1761  (.L_HI(net1761));
 sg13g2_tiehi \top_ihp.oisc.regs[26][11]$_DFFE_PP__1762  (.L_HI(net1762));
 sg13g2_tiehi \top_ihp.oisc.regs[26][12]$_DFFE_PP__1763  (.L_HI(net1763));
 sg13g2_tiehi \top_ihp.oisc.regs[26][13]$_DFFE_PP__1764  (.L_HI(net1764));
 sg13g2_tiehi \top_ihp.oisc.regs[26][14]$_DFFE_PP__1765  (.L_HI(net1765));
 sg13g2_tiehi \top_ihp.oisc.regs[26][15]$_DFFE_PP__1766  (.L_HI(net1766));
 sg13g2_tiehi \top_ihp.oisc.regs[26][16]$_DFFE_PP__1767  (.L_HI(net1767));
 sg13g2_tiehi \top_ihp.oisc.regs[26][17]$_DFFE_PP__1768  (.L_HI(net1768));
 sg13g2_tiehi \top_ihp.oisc.regs[26][18]$_DFFE_PP__1769  (.L_HI(net1769));
 sg13g2_tiehi \top_ihp.oisc.regs[26][19]$_DFFE_PP__1770  (.L_HI(net1770));
 sg13g2_tiehi \top_ihp.oisc.regs[26][1]$_DFFE_PP__1771  (.L_HI(net1771));
 sg13g2_tiehi \top_ihp.oisc.regs[26][20]$_DFFE_PP__1772  (.L_HI(net1772));
 sg13g2_tiehi \top_ihp.oisc.regs[26][21]$_DFFE_PP__1773  (.L_HI(net1773));
 sg13g2_tiehi \top_ihp.oisc.regs[26][22]$_DFFE_PP__1774  (.L_HI(net1774));
 sg13g2_tiehi \top_ihp.oisc.regs[26][23]$_DFFE_PP__1775  (.L_HI(net1775));
 sg13g2_tiehi \top_ihp.oisc.regs[26][24]$_DFFE_PP__1776  (.L_HI(net1776));
 sg13g2_tiehi \top_ihp.oisc.regs[26][25]$_DFFE_PP__1777  (.L_HI(net1777));
 sg13g2_tiehi \top_ihp.oisc.regs[26][26]$_DFFE_PP__1778  (.L_HI(net1778));
 sg13g2_tiehi \top_ihp.oisc.regs[26][27]$_DFFE_PP__1779  (.L_HI(net1779));
 sg13g2_tiehi \top_ihp.oisc.regs[26][28]$_DFFE_PP__1780  (.L_HI(net1780));
 sg13g2_tiehi \top_ihp.oisc.regs[26][29]$_DFFE_PP__1781  (.L_HI(net1781));
 sg13g2_tiehi \top_ihp.oisc.regs[26][2]$_DFFE_PP__1782  (.L_HI(net1782));
 sg13g2_tiehi \top_ihp.oisc.regs[26][30]$_DFFE_PP__1783  (.L_HI(net1783));
 sg13g2_tiehi \top_ihp.oisc.regs[26][31]$_DFFE_PP__1784  (.L_HI(net1784));
 sg13g2_tiehi \top_ihp.oisc.regs[26][3]$_DFFE_PP__1785  (.L_HI(net1785));
 sg13g2_tiehi \top_ihp.oisc.regs[26][4]$_DFFE_PP__1786  (.L_HI(net1786));
 sg13g2_tiehi \top_ihp.oisc.regs[26][5]$_DFFE_PP__1787  (.L_HI(net1787));
 sg13g2_tiehi \top_ihp.oisc.regs[26][6]$_DFFE_PP__1788  (.L_HI(net1788));
 sg13g2_tiehi \top_ihp.oisc.regs[26][7]$_DFFE_PP__1789  (.L_HI(net1789));
 sg13g2_tiehi \top_ihp.oisc.regs[26][8]$_DFFE_PP__1790  (.L_HI(net1790));
 sg13g2_tiehi \top_ihp.oisc.regs[26][9]$_DFFE_PP__1791  (.L_HI(net1791));
 sg13g2_tiehi \top_ihp.oisc.regs[27][0]$_DFFE_PP__1792  (.L_HI(net1792));
 sg13g2_tiehi \top_ihp.oisc.regs[27][10]$_DFFE_PP__1793  (.L_HI(net1793));
 sg13g2_tiehi \top_ihp.oisc.regs[27][11]$_DFFE_PP__1794  (.L_HI(net1794));
 sg13g2_tiehi \top_ihp.oisc.regs[27][12]$_DFFE_PP__1795  (.L_HI(net1795));
 sg13g2_tiehi \top_ihp.oisc.regs[27][13]$_DFFE_PP__1796  (.L_HI(net1796));
 sg13g2_tiehi \top_ihp.oisc.regs[27][14]$_DFFE_PP__1797  (.L_HI(net1797));
 sg13g2_tiehi \top_ihp.oisc.regs[27][15]$_DFFE_PP__1798  (.L_HI(net1798));
 sg13g2_tiehi \top_ihp.oisc.regs[27][16]$_DFFE_PP__1799  (.L_HI(net1799));
 sg13g2_tiehi \top_ihp.oisc.regs[27][17]$_DFFE_PP__1800  (.L_HI(net1800));
 sg13g2_tiehi \top_ihp.oisc.regs[27][18]$_DFFE_PP__1801  (.L_HI(net1801));
 sg13g2_tiehi \top_ihp.oisc.regs[27][19]$_DFFE_PP__1802  (.L_HI(net1802));
 sg13g2_tiehi \top_ihp.oisc.regs[27][1]$_DFFE_PP__1803  (.L_HI(net1803));
 sg13g2_tiehi \top_ihp.oisc.regs[27][20]$_DFFE_PP__1804  (.L_HI(net1804));
 sg13g2_tiehi \top_ihp.oisc.regs[27][21]$_DFFE_PP__1805  (.L_HI(net1805));
 sg13g2_tiehi \top_ihp.oisc.regs[27][22]$_DFFE_PP__1806  (.L_HI(net1806));
 sg13g2_tiehi \top_ihp.oisc.regs[27][23]$_DFFE_PP__1807  (.L_HI(net1807));
 sg13g2_tiehi \top_ihp.oisc.regs[27][24]$_DFFE_PP__1808  (.L_HI(net1808));
 sg13g2_tiehi \top_ihp.oisc.regs[27][25]$_DFFE_PP__1809  (.L_HI(net1809));
 sg13g2_tiehi \top_ihp.oisc.regs[27][26]$_DFFE_PP__1810  (.L_HI(net1810));
 sg13g2_tiehi \top_ihp.oisc.regs[27][27]$_DFFE_PP__1811  (.L_HI(net1811));
 sg13g2_tiehi \top_ihp.oisc.regs[27][28]$_DFFE_PP__1812  (.L_HI(net1812));
 sg13g2_tiehi \top_ihp.oisc.regs[27][29]$_DFFE_PP__1813  (.L_HI(net1813));
 sg13g2_tiehi \top_ihp.oisc.regs[27][2]$_DFFE_PP__1814  (.L_HI(net1814));
 sg13g2_tiehi \top_ihp.oisc.regs[27][30]$_DFFE_PP__1815  (.L_HI(net1815));
 sg13g2_tiehi \top_ihp.oisc.regs[27][31]$_DFFE_PP__1816  (.L_HI(net1816));
 sg13g2_tiehi \top_ihp.oisc.regs[27][3]$_DFFE_PP__1817  (.L_HI(net1817));
 sg13g2_tiehi \top_ihp.oisc.regs[27][4]$_DFFE_PP__1818  (.L_HI(net1818));
 sg13g2_tiehi \top_ihp.oisc.regs[27][5]$_DFFE_PP__1819  (.L_HI(net1819));
 sg13g2_tiehi \top_ihp.oisc.regs[27][6]$_DFFE_PP__1820  (.L_HI(net1820));
 sg13g2_tiehi \top_ihp.oisc.regs[27][7]$_DFFE_PP__1821  (.L_HI(net1821));
 sg13g2_tiehi \top_ihp.oisc.regs[27][8]$_DFFE_PP__1822  (.L_HI(net1822));
 sg13g2_tiehi \top_ihp.oisc.regs[27][9]$_DFFE_PP__1823  (.L_HI(net1823));
 sg13g2_tiehi \top_ihp.oisc.regs[28][0]$_DFFE_PP__1824  (.L_HI(net1824));
 sg13g2_tiehi \top_ihp.oisc.regs[28][10]$_DFFE_PP__1825  (.L_HI(net1825));
 sg13g2_tiehi \top_ihp.oisc.regs[28][11]$_DFFE_PP__1826  (.L_HI(net1826));
 sg13g2_tiehi \top_ihp.oisc.regs[28][12]$_DFFE_PP__1827  (.L_HI(net1827));
 sg13g2_tiehi \top_ihp.oisc.regs[28][13]$_DFFE_PP__1828  (.L_HI(net1828));
 sg13g2_tiehi \top_ihp.oisc.regs[28][14]$_DFFE_PP__1829  (.L_HI(net1829));
 sg13g2_tiehi \top_ihp.oisc.regs[28][15]$_DFFE_PP__1830  (.L_HI(net1830));
 sg13g2_tiehi \top_ihp.oisc.regs[28][16]$_DFFE_PP__1831  (.L_HI(net1831));
 sg13g2_tiehi \top_ihp.oisc.regs[28][17]$_DFFE_PP__1832  (.L_HI(net1832));
 sg13g2_tiehi \top_ihp.oisc.regs[28][18]$_DFFE_PP__1833  (.L_HI(net1833));
 sg13g2_tiehi \top_ihp.oisc.regs[28][19]$_DFFE_PP__1834  (.L_HI(net1834));
 sg13g2_tiehi \top_ihp.oisc.regs[28][1]$_DFFE_PP__1835  (.L_HI(net1835));
 sg13g2_tiehi \top_ihp.oisc.regs[28][20]$_DFFE_PP__1836  (.L_HI(net1836));
 sg13g2_tiehi \top_ihp.oisc.regs[28][21]$_DFFE_PP__1837  (.L_HI(net1837));
 sg13g2_tiehi \top_ihp.oisc.regs[28][22]$_DFFE_PP__1838  (.L_HI(net1838));
 sg13g2_tiehi \top_ihp.oisc.regs[28][23]$_DFFE_PP__1839  (.L_HI(net1839));
 sg13g2_tiehi \top_ihp.oisc.regs[28][24]$_DFFE_PP__1840  (.L_HI(net1840));
 sg13g2_tiehi \top_ihp.oisc.regs[28][25]$_DFFE_PP__1841  (.L_HI(net1841));
 sg13g2_tiehi \top_ihp.oisc.regs[28][26]$_DFFE_PP__1842  (.L_HI(net1842));
 sg13g2_tiehi \top_ihp.oisc.regs[28][27]$_DFFE_PP__1843  (.L_HI(net1843));
 sg13g2_tiehi \top_ihp.oisc.regs[28][28]$_DFFE_PP__1844  (.L_HI(net1844));
 sg13g2_tiehi \top_ihp.oisc.regs[28][29]$_DFFE_PP__1845  (.L_HI(net1845));
 sg13g2_tiehi \top_ihp.oisc.regs[28][2]$_DFFE_PP__1846  (.L_HI(net1846));
 sg13g2_tiehi \top_ihp.oisc.regs[28][30]$_DFFE_PP__1847  (.L_HI(net1847));
 sg13g2_tiehi \top_ihp.oisc.regs[28][31]$_DFFE_PP__1848  (.L_HI(net1848));
 sg13g2_tiehi \top_ihp.oisc.regs[28][3]$_DFFE_PP__1849  (.L_HI(net1849));
 sg13g2_tiehi \top_ihp.oisc.regs[28][4]$_DFFE_PP__1850  (.L_HI(net1850));
 sg13g2_tiehi \top_ihp.oisc.regs[28][5]$_DFFE_PP__1851  (.L_HI(net1851));
 sg13g2_tiehi \top_ihp.oisc.regs[28][6]$_DFFE_PP__1852  (.L_HI(net1852));
 sg13g2_tiehi \top_ihp.oisc.regs[28][7]$_DFFE_PP__1853  (.L_HI(net1853));
 sg13g2_tiehi \top_ihp.oisc.regs[28][8]$_DFFE_PP__1854  (.L_HI(net1854));
 sg13g2_tiehi \top_ihp.oisc.regs[28][9]$_DFFE_PP__1855  (.L_HI(net1855));
 sg13g2_tiehi \top_ihp.oisc.regs[29][0]$_DFFE_PP__1856  (.L_HI(net1856));
 sg13g2_tiehi \top_ihp.oisc.regs[29][10]$_DFFE_PP__1857  (.L_HI(net1857));
 sg13g2_tiehi \top_ihp.oisc.regs[29][11]$_DFFE_PP__1858  (.L_HI(net1858));
 sg13g2_tiehi \top_ihp.oisc.regs[29][12]$_DFFE_PP__1859  (.L_HI(net1859));
 sg13g2_tiehi \top_ihp.oisc.regs[29][13]$_DFFE_PP__1860  (.L_HI(net1860));
 sg13g2_tiehi \top_ihp.oisc.regs[29][14]$_DFFE_PP__1861  (.L_HI(net1861));
 sg13g2_tiehi \top_ihp.oisc.regs[29][15]$_DFFE_PP__1862  (.L_HI(net1862));
 sg13g2_tiehi \top_ihp.oisc.regs[29][16]$_DFFE_PP__1863  (.L_HI(net1863));
 sg13g2_tiehi \top_ihp.oisc.regs[29][17]$_DFFE_PP__1864  (.L_HI(net1864));
 sg13g2_tiehi \top_ihp.oisc.regs[29][18]$_DFFE_PP__1865  (.L_HI(net1865));
 sg13g2_tiehi \top_ihp.oisc.regs[29][19]$_DFFE_PP__1866  (.L_HI(net1866));
 sg13g2_tiehi \top_ihp.oisc.regs[29][1]$_DFFE_PP__1867  (.L_HI(net1867));
 sg13g2_tiehi \top_ihp.oisc.regs[29][20]$_DFFE_PP__1868  (.L_HI(net1868));
 sg13g2_tiehi \top_ihp.oisc.regs[29][21]$_DFFE_PP__1869  (.L_HI(net1869));
 sg13g2_tiehi \top_ihp.oisc.regs[29][22]$_DFFE_PP__1870  (.L_HI(net1870));
 sg13g2_tiehi \top_ihp.oisc.regs[29][23]$_DFFE_PP__1871  (.L_HI(net1871));
 sg13g2_tiehi \top_ihp.oisc.regs[29][24]$_DFFE_PP__1872  (.L_HI(net1872));
 sg13g2_tiehi \top_ihp.oisc.regs[29][25]$_DFFE_PP__1873  (.L_HI(net1873));
 sg13g2_tiehi \top_ihp.oisc.regs[29][26]$_DFFE_PP__1874  (.L_HI(net1874));
 sg13g2_tiehi \top_ihp.oisc.regs[29][27]$_DFFE_PP__1875  (.L_HI(net1875));
 sg13g2_tiehi \top_ihp.oisc.regs[29][28]$_DFFE_PP__1876  (.L_HI(net1876));
 sg13g2_tiehi \top_ihp.oisc.regs[29][29]$_DFFE_PP__1877  (.L_HI(net1877));
 sg13g2_tiehi \top_ihp.oisc.regs[29][2]$_DFFE_PP__1878  (.L_HI(net1878));
 sg13g2_tiehi \top_ihp.oisc.regs[29][30]$_DFFE_PP__1879  (.L_HI(net1879));
 sg13g2_tiehi \top_ihp.oisc.regs[29][31]$_DFFE_PP__1880  (.L_HI(net1880));
 sg13g2_tiehi \top_ihp.oisc.regs[29][3]$_DFFE_PP__1881  (.L_HI(net1881));
 sg13g2_tiehi \top_ihp.oisc.regs[29][4]$_DFFE_PP__1882  (.L_HI(net1882));
 sg13g2_tiehi \top_ihp.oisc.regs[29][5]$_DFFE_PP__1883  (.L_HI(net1883));
 sg13g2_tiehi \top_ihp.oisc.regs[29][6]$_DFFE_PP__1884  (.L_HI(net1884));
 sg13g2_tiehi \top_ihp.oisc.regs[29][7]$_DFFE_PP__1885  (.L_HI(net1885));
 sg13g2_tiehi \top_ihp.oisc.regs[29][8]$_DFFE_PP__1886  (.L_HI(net1886));
 sg13g2_tiehi \top_ihp.oisc.regs[29][9]$_DFFE_PP__1887  (.L_HI(net1887));
 sg13g2_tiehi \top_ihp.oisc.regs[30][0]$_DFFE_PP__1888  (.L_HI(net1888));
 sg13g2_tiehi \top_ihp.oisc.regs[30][10]$_DFFE_PP__1889  (.L_HI(net1889));
 sg13g2_tiehi \top_ihp.oisc.regs[30][11]$_DFFE_PP__1890  (.L_HI(net1890));
 sg13g2_tiehi \top_ihp.oisc.regs[30][12]$_DFFE_PP__1891  (.L_HI(net1891));
 sg13g2_tiehi \top_ihp.oisc.regs[30][13]$_DFFE_PP__1892  (.L_HI(net1892));
 sg13g2_tiehi \top_ihp.oisc.regs[30][14]$_DFFE_PP__1893  (.L_HI(net1893));
 sg13g2_tiehi \top_ihp.oisc.regs[30][15]$_DFFE_PP__1894  (.L_HI(net1894));
 sg13g2_tiehi \top_ihp.oisc.regs[30][16]$_DFFE_PP__1895  (.L_HI(net1895));
 sg13g2_tiehi \top_ihp.oisc.regs[30][17]$_DFFE_PP__1896  (.L_HI(net1896));
 sg13g2_tiehi \top_ihp.oisc.regs[30][18]$_DFFE_PP__1897  (.L_HI(net1897));
 sg13g2_tiehi \top_ihp.oisc.regs[30][19]$_DFFE_PP__1898  (.L_HI(net1898));
 sg13g2_tiehi \top_ihp.oisc.regs[30][1]$_DFFE_PP__1899  (.L_HI(net1899));
 sg13g2_tiehi \top_ihp.oisc.regs[30][20]$_DFFE_PP__1900  (.L_HI(net1900));
 sg13g2_tiehi \top_ihp.oisc.regs[30][21]$_DFFE_PP__1901  (.L_HI(net1901));
 sg13g2_tiehi \top_ihp.oisc.regs[30][22]$_DFFE_PP__1902  (.L_HI(net1902));
 sg13g2_tiehi \top_ihp.oisc.regs[30][23]$_DFFE_PP__1903  (.L_HI(net1903));
 sg13g2_tiehi \top_ihp.oisc.regs[30][24]$_DFFE_PP__1904  (.L_HI(net1904));
 sg13g2_tiehi \top_ihp.oisc.regs[30][25]$_DFFE_PP__1905  (.L_HI(net1905));
 sg13g2_tiehi \top_ihp.oisc.regs[30][26]$_DFFE_PP__1906  (.L_HI(net1906));
 sg13g2_tiehi \top_ihp.oisc.regs[30][27]$_DFFE_PP__1907  (.L_HI(net1907));
 sg13g2_tiehi \top_ihp.oisc.regs[30][28]$_DFFE_PP__1908  (.L_HI(net1908));
 sg13g2_tiehi \top_ihp.oisc.regs[30][29]$_DFFE_PP__1909  (.L_HI(net1909));
 sg13g2_tiehi \top_ihp.oisc.regs[30][2]$_DFFE_PP__1910  (.L_HI(net1910));
 sg13g2_tiehi \top_ihp.oisc.regs[30][30]$_DFFE_PP__1911  (.L_HI(net1911));
 sg13g2_tiehi \top_ihp.oisc.regs[30][31]$_DFFE_PP__1912  (.L_HI(net1912));
 sg13g2_tiehi \top_ihp.oisc.regs[30][3]$_DFFE_PP__1913  (.L_HI(net1913));
 sg13g2_tiehi \top_ihp.oisc.regs[30][4]$_DFFE_PP__1914  (.L_HI(net1914));
 sg13g2_tiehi \top_ihp.oisc.regs[30][5]$_DFFE_PP__1915  (.L_HI(net1915));
 sg13g2_tiehi \top_ihp.oisc.regs[30][6]$_DFFE_PP__1916  (.L_HI(net1916));
 sg13g2_tiehi \top_ihp.oisc.regs[30][7]$_DFFE_PP__1917  (.L_HI(net1917));
 sg13g2_tiehi \top_ihp.oisc.regs[30][8]$_DFFE_PP__1918  (.L_HI(net1918));
 sg13g2_tiehi \top_ihp.oisc.regs[30][9]$_DFFE_PP__1919  (.L_HI(net1919));
 sg13g2_tiehi \top_ihp.oisc.regs[31][0]$_DFFE_PP__1920  (.L_HI(net1920));
 sg13g2_tiehi \top_ihp.oisc.regs[31][10]$_DFFE_PP__1921  (.L_HI(net1921));
 sg13g2_tiehi \top_ihp.oisc.regs[31][11]$_DFFE_PP__1922  (.L_HI(net1922));
 sg13g2_tiehi \top_ihp.oisc.regs[31][12]$_DFFE_PP__1923  (.L_HI(net1923));
 sg13g2_tiehi \top_ihp.oisc.regs[31][13]$_DFFE_PP__1924  (.L_HI(net1924));
 sg13g2_tiehi \top_ihp.oisc.regs[31][14]$_DFFE_PP__1925  (.L_HI(net1925));
 sg13g2_tiehi \top_ihp.oisc.regs[31][15]$_DFFE_PP__1926  (.L_HI(net1926));
 sg13g2_tiehi \top_ihp.oisc.regs[31][16]$_DFFE_PP__1927  (.L_HI(net1927));
 sg13g2_tiehi \top_ihp.oisc.regs[31][17]$_DFFE_PP__1928  (.L_HI(net1928));
 sg13g2_tiehi \top_ihp.oisc.regs[31][18]$_DFFE_PP__1929  (.L_HI(net1929));
 sg13g2_tiehi \top_ihp.oisc.regs[31][19]$_DFFE_PP__1930  (.L_HI(net1930));
 sg13g2_tiehi \top_ihp.oisc.regs[31][1]$_DFFE_PP__1931  (.L_HI(net1931));
 sg13g2_tiehi \top_ihp.oisc.regs[31][20]$_DFFE_PP__1932  (.L_HI(net1932));
 sg13g2_tiehi \top_ihp.oisc.regs[31][21]$_DFFE_PP__1933  (.L_HI(net1933));
 sg13g2_tiehi \top_ihp.oisc.regs[31][22]$_DFFE_PP__1934  (.L_HI(net1934));
 sg13g2_tiehi \top_ihp.oisc.regs[31][23]$_DFFE_PP__1935  (.L_HI(net1935));
 sg13g2_tiehi \top_ihp.oisc.regs[31][24]$_DFFE_PP__1936  (.L_HI(net1936));
 sg13g2_tiehi \top_ihp.oisc.regs[31][25]$_DFFE_PP__1937  (.L_HI(net1937));
 sg13g2_tiehi \top_ihp.oisc.regs[31][26]$_DFFE_PP__1938  (.L_HI(net1938));
 sg13g2_tiehi \top_ihp.oisc.regs[31][27]$_DFFE_PP__1939  (.L_HI(net1939));
 sg13g2_tiehi \top_ihp.oisc.regs[31][28]$_DFFE_PP__1940  (.L_HI(net1940));
 sg13g2_tiehi \top_ihp.oisc.regs[31][29]$_DFFE_PP__1941  (.L_HI(net1941));
 sg13g2_tiehi \top_ihp.oisc.regs[31][2]$_DFFE_PP__1942  (.L_HI(net1942));
 sg13g2_tiehi \top_ihp.oisc.regs[31][30]$_DFFE_PP__1943  (.L_HI(net1943));
 sg13g2_tiehi \top_ihp.oisc.regs[31][31]$_DFFE_PP__1944  (.L_HI(net1944));
 sg13g2_tiehi \top_ihp.oisc.regs[31][3]$_DFFE_PP__1945  (.L_HI(net1945));
 sg13g2_tiehi \top_ihp.oisc.regs[31][4]$_DFFE_PP__1946  (.L_HI(net1946));
 sg13g2_tiehi \top_ihp.oisc.regs[31][5]$_DFFE_PP__1947  (.L_HI(net1947));
 sg13g2_tiehi \top_ihp.oisc.regs[31][6]$_DFFE_PP__1948  (.L_HI(net1948));
 sg13g2_tiehi \top_ihp.oisc.regs[31][7]$_DFFE_PP__1949  (.L_HI(net1949));
 sg13g2_tiehi \top_ihp.oisc.regs[31][8]$_DFFE_PP__1950  (.L_HI(net1950));
 sg13g2_tiehi \top_ihp.oisc.regs[31][9]$_DFFE_PP__1951  (.L_HI(net1951));
 sg13g2_tiehi \top_ihp.oisc.regs[32][0]$_DFFE_PP__1952  (.L_HI(net1952));
 sg13g2_tiehi \top_ihp.oisc.regs[32][10]$_DFFE_PP__1953  (.L_HI(net1953));
 sg13g2_tiehi \top_ihp.oisc.regs[32][11]$_DFFE_PP__1954  (.L_HI(net1954));
 sg13g2_tiehi \top_ihp.oisc.regs[32][12]$_DFFE_PP__1955  (.L_HI(net1955));
 sg13g2_tiehi \top_ihp.oisc.regs[32][13]$_DFFE_PP__1956  (.L_HI(net1956));
 sg13g2_tiehi \top_ihp.oisc.regs[32][14]$_DFFE_PP__1957  (.L_HI(net1957));
 sg13g2_tiehi \top_ihp.oisc.regs[32][15]$_DFFE_PP__1958  (.L_HI(net1958));
 sg13g2_tiehi \top_ihp.oisc.regs[32][16]$_DFFE_PP__1959  (.L_HI(net1959));
 sg13g2_tiehi \top_ihp.oisc.regs[32][17]$_DFFE_PP__1960  (.L_HI(net1960));
 sg13g2_tiehi \top_ihp.oisc.regs[32][18]$_DFFE_PP__1961  (.L_HI(net1961));
 sg13g2_tiehi \top_ihp.oisc.regs[32][19]$_DFFE_PP__1962  (.L_HI(net1962));
 sg13g2_tiehi \top_ihp.oisc.regs[32][1]$_DFFE_PP__1963  (.L_HI(net1963));
 sg13g2_tiehi \top_ihp.oisc.regs[32][20]$_DFFE_PP__1964  (.L_HI(net1964));
 sg13g2_tiehi \top_ihp.oisc.regs[32][21]$_DFFE_PP__1965  (.L_HI(net1965));
 sg13g2_tiehi \top_ihp.oisc.regs[32][22]$_DFFE_PP__1966  (.L_HI(net1966));
 sg13g2_tiehi \top_ihp.oisc.regs[32][23]$_DFFE_PP__1967  (.L_HI(net1967));
 sg13g2_tiehi \top_ihp.oisc.regs[32][24]$_DFFE_PP__1968  (.L_HI(net1968));
 sg13g2_tiehi \top_ihp.oisc.regs[32][25]$_DFFE_PP__1969  (.L_HI(net1969));
 sg13g2_tiehi \top_ihp.oisc.regs[32][26]$_DFFE_PP__1970  (.L_HI(net1970));
 sg13g2_tiehi \top_ihp.oisc.regs[32][27]$_DFFE_PP__1971  (.L_HI(net1971));
 sg13g2_tiehi \top_ihp.oisc.regs[32][28]$_DFFE_PP__1972  (.L_HI(net1972));
 sg13g2_tiehi \top_ihp.oisc.regs[32][29]$_DFFE_PP__1973  (.L_HI(net1973));
 sg13g2_tiehi \top_ihp.oisc.regs[32][2]$_DFFE_PP__1974  (.L_HI(net1974));
 sg13g2_tiehi \top_ihp.oisc.regs[32][30]$_DFFE_PP__1975  (.L_HI(net1975));
 sg13g2_tiehi \top_ihp.oisc.regs[32][31]$_DFFE_PP__1976  (.L_HI(net1976));
 sg13g2_tiehi \top_ihp.oisc.regs[32][3]$_DFFE_PP__1977  (.L_HI(net1977));
 sg13g2_tiehi \top_ihp.oisc.regs[32][4]$_DFFE_PP__1978  (.L_HI(net1978));
 sg13g2_tiehi \top_ihp.oisc.regs[32][5]$_DFFE_PP__1979  (.L_HI(net1979));
 sg13g2_tiehi \top_ihp.oisc.regs[32][6]$_DFFE_PP__1980  (.L_HI(net1980));
 sg13g2_tiehi \top_ihp.oisc.regs[32][7]$_DFFE_PP__1981  (.L_HI(net1981));
 sg13g2_tiehi \top_ihp.oisc.regs[32][8]$_DFFE_PP__1982  (.L_HI(net1982));
 sg13g2_tiehi \top_ihp.oisc.regs[32][9]$_DFFE_PP__1983  (.L_HI(net1983));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[0]$_SDFFCE_PN0P__1984  (.L_HI(net1984));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[1]$_SDFFCE_PN0P__1985  (.L_HI(net1985));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[2]$_SDFFCE_PN0P__1986  (.L_HI(net1986));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[3]$_SDFFCE_PN0P__1987  (.L_HI(net1987));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[4]$_SDFFCE_PN0P__1988  (.L_HI(net1988));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[5]$_SDFFCE_PN0P__1989  (.L_HI(net1989));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[6]$_SDFFCE_PN0P__1990  (.L_HI(net1990));
 sg13g2_tiehi \top_ihp.wb_emem.bit_counter[7]$_SDFFCE_PN0P__1991  (.L_HI(net1991));
 sg13g2_tiehi \top_ihp.wb_emem.last_bit$_DFFE_PP__1992  (.L_HI(net1992));
 sg13g2_tiehi \top_ihp.wb_emem.last_wait$_DFFE_PP__1993  (.L_HI(net1993));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[3]$_SDFFCE_NP1P__1994  (.L_HI(net1994));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[4]$_SDFFCE_NP0P__1995  (.L_HI(net1995));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[5]$_SDFFCE_NP0P__1996  (.L_HI(net1996));
 sg13g2_tiehi \top_ihp.wb_emem.nbits[6]$_SDFFCE_NP0P__1997  (.L_HI(net1997));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[0]$_SDFFCE_PN0P__1998  (.L_HI(net1998));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[1]$_SDFFCE_PN0P__1999  (.L_HI(net1999));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[2]$_SDFFCE_PN0P__2000  (.L_HI(net2000));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[3]$_SDFFCE_PN0P__2001  (.L_HI(net2001));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[4]$_SDFFCE_PN0P__2002  (.L_HI(net2002));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[5]$_SDFFCE_PN0P__2003  (.L_HI(net2003));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[6]$_SDFFCE_PN0P__2004  (.L_HI(net2004));
 sg13g2_tiehi \top_ihp.wb_emem.wait_counter[7]$_SDFFCE_PN0P__2005  (.L_HI(net2005));
 sg13g2_tiehi \top_ihp.wb_uart.ack_o$_SDFFCE_PP0P__2006  (.L_HI(net2006));
 sg13g2_inv_1 net1791_2 (.Y(net2008),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 net1791_3 (.Y(net2009),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net1791_4 (.Y(net2010),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net1791_5 (.Y(net2011),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net1791_6 (.Y(net2012),
    .A(clknet_leaf_62_clk));
 sg13g2_inv_1 net1791_7 (.Y(net2013),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net1791_8 (.Y(net2014),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net1791_9 (.Y(net2015),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net1791_10 (.Y(net2016),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net1791_11 (.Y(net2017),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net1791_12 (.Y(net2018),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net1791_13 (.Y(net2019),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net1791_14 (.Y(net2020),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net1791_15 (.Y(net2021),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 net1791_16 (.Y(net2022),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net1791_17 (.Y(net2023),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 net1791_18 (.Y(net2024),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 net1791_19 (.Y(net2025),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 net1791_20 (.Y(net2026),
    .A(clknet_leaf_17_clk));
 sg13g2_inv_1 net1791_21 (.Y(net2027),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net2027_22 (.Y(net2028),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net2027_23 (.Y(net2029),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_24 (.Y(net2030),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_25 (.Y(net2031),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 net2027_26 (.Y(net2032),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_27 (.Y(net2033),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net2027_28 (.Y(net2034),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_29 (.Y(net2035),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_30 (.Y(net2036),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_31 (.Y(net2037),
    .A(clknet_leaf_39_clk));
 sg13g2_inv_1 net2027_32 (.Y(net2038),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net2027_33 (.Y(net2039),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net2027_34 (.Y(net2040),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net2027_35 (.Y(net2041),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net2027_36 (.Y(net2042),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net2027_37 (.Y(net2043),
    .A(clknet_leaf_16_clk));
 sg13g2_inv_1 net2027_38 (.Y(net2044),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net2027_39 (.Y(net2045),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 net2027_40 (.Y(net2046),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 net2027_41 (.Y(net2047),
    .A(clknet_leaf_3_clk));
 sg13g2_inv_1 net2027_42 (.Y(net2048),
    .A(clknet_leaf_5_clk));
 sg13g2_inv_1 net2027_43 (.Y(net2049),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net2027_44 (.Y(net2050),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 net2027_45 (.Y(net2051),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net2027_46 (.Y(net2052),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 net2027_47 (.Y(net2053),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 net2027_48 (.Y(net2054),
    .A(clknet_leaf_10_clk));
 sg13g2_inv_1 net2027_49 (.Y(net2055),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 net2027_50 (.Y(net2056),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 net2027_51 (.Y(net2057),
    .A(clknet_leaf_7_clk));
 sg13g2_inv_1 net2027_52 (.Y(net2058),
    .A(clknet_leaf_6_clk));
 sg13g2_inv_1 net2027_53 (.Y(net2059),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_54 (.Y(net2060),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_55 (.Y(net2061),
    .A(clknet_leaf_47_clk));
 sg13g2_inv_1 net2027_56 (.Y(net2062),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 net2027_57 (.Y(net2063),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net2027_58 (.Y(net2064),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net2027_59 (.Y(net2065),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net2027_60 (.Y(net2066),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net2027_61 (.Y(net2067),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_62 (.Y(net2068),
    .A(clknet_leaf_11_clk));
 sg13g2_inv_1 net2027_63 (.Y(net2069),
    .A(clknet_leaf_13_clk));
 sg13g2_inv_1 net2027_64 (.Y(net2070),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net2027_65 (.Y(net2071),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_66 (.Y(net2072),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_67 (.Y(net2073),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 net2027_68 (.Y(net2074),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 net2027_69 (.Y(net2075),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 net2027_70 (.Y(net2076),
    .A(clknet_leaf_46_clk));
 sg13g2_inv_1 net2027_71 (.Y(net2077),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_72 (.Y(net2078),
    .A(clknet_leaf_56_clk));
 sg13g2_inv_1 net2027_73 (.Y(net2079),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_74 (.Y(net2080),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_75 (.Y(net2081),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_76 (.Y(net2082),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_77 (.Y(net2083),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_78 (.Y(net2084),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_79 (.Y(net2085),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_80 (.Y(net2086),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net2027_81 (.Y(net2087),
    .A(clknet_leaf_15_clk));
 sg13g2_inv_1 net2027_82 (.Y(net2088),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_83 (.Y(net2089),
    .A(clknet_leaf_49_clk));
 sg13g2_inv_1 net2027_84 (.Y(net2090),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_85 (.Y(net2091),
    .A(clknet_leaf_14_clk));
 sg13g2_inv_1 net2027_86 (.Y(net2092),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_87 (.Y(net2093),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_88 (.Y(net2094),
    .A(clknet_leaf_43_clk));
 sg13g2_inv_1 net2027_89 (.Y(net2095),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_90 (.Y(net2096),
    .A(clknet_leaf_42_clk));
 sg13g2_inv_1 net2027_91 (.Y(net2097),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_92 (.Y(net2098),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_93 (.Y(net2099),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_94 (.Y(net2100),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_95 (.Y(net2101),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_96 (.Y(net2102),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_97 (.Y(net2103),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_98 (.Y(net2104),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_99 (.Y(net2105),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_100 (.Y(net2106),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net2027_101 (.Y(net2107),
    .A(clknet_leaf_40_clk));
 sg13g2_inv_1 net2027_102 (.Y(net2108),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 net2027_103 (.Y(net2109),
    .A(clknet_leaf_52_clk));
 sg13g2_inv_1 net2027_104 (.Y(net2110),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_105 (.Y(net2111),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_106 (.Y(net2112),
    .A(clknet_leaf_37_clk));
 sg13g2_inv_1 net2027_107 (.Y(net2113),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net2027_108 (.Y(net2114),
    .A(clknet_leaf_50_clk));
 sg13g2_inv_1 net2027_109 (.Y(net2115),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_110 (.Y(net2116),
    .A(clknet_leaf_38_clk));
 sg13g2_inv_1 net2027_111 (.Y(net2117),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_112 (.Y(net2118),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net2027_113 (.Y(net2119),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net2027_114 (.Y(net2120),
    .A(clknet_leaf_53_clk));
 sg13g2_inv_1 net2027_115 (.Y(net2121),
    .A(clknet_leaf_41_clk));
 sg13g2_inv_1 net2027_116 (.Y(net2122),
    .A(clknet_leaf_51_clk));
 sg13g2_inv_1 net2027_117 (.Y(net2123),
    .A(clknet_leaf_61_clk));
 sg13g2_inv_1 net2027_118 (.Y(net2124),
    .A(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_6_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_6_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_6_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_6_7__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_37_clk));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_38_clk));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_39_clk));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_40_clk));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_41_clk));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_42_clk));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_6_5__leaf_clk),
    .X(clknet_leaf_43_clk));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_44_clk));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_45_clk));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_46_clk));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_47_clk));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_48_clk));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_6_16__leaf_clk),
    .X(clknet_leaf_49_clk));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_50_clk));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_52_clk));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_6_18__leaf_clk),
    .X(clknet_leaf_53_clk));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_54_clk));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_55_clk));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_6_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_58_clk));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_59_clk));
 sg13g2_buf_8 clkbuf_leaf_60_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_60_clk));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_61_clk));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_6_21__leaf_clk),
    .X(clknet_leaf_62_clk));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_63_clk));
 sg13g2_buf_8 clkbuf_leaf_64_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_64_clk));
 sg13g2_buf_8 clkbuf_leaf_65_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_65_clk));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_66_clk));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_67_clk));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_6_20__leaf_clk),
    .X(clknet_leaf_68_clk));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_69_clk));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_70_clk));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_71_clk));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_72_clk));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_73_clk));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_74_clk));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_75_clk));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_6_23__leaf_clk),
    .X(clknet_leaf_76_clk));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_77_clk));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_78_clk));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_79_clk));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_80_clk));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_6_29__leaf_clk),
    .X(clknet_leaf_81_clk));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_82_clk));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_83_clk));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_84_clk));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_85_clk));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_86_clk));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_87_clk));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_88_clk));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_89_clk));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_90_clk));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_91_clk));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_6_28__leaf_clk),
    .X(clknet_leaf_92_clk));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_6_22__leaf_clk),
    .X(clknet_leaf_93_clk));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_94_clk));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_6_19__leaf_clk),
    .X(clknet_leaf_95_clk));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_96_clk));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_97_clk));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_98_clk));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_6_25__leaf_clk),
    .X(clknet_leaf_99_clk));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_100_clk));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_101_clk));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_102_clk));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_103_clk));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_6_24__leaf_clk),
    .X(clknet_leaf_104_clk));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_105_clk));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_106_clk));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_107_clk));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_108_clk));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_109_clk));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_110_clk));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_6_26__leaf_clk),
    .X(clknet_leaf_111_clk));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_112_clk));
 sg13g2_buf_8 clkbuf_leaf_113_clk (.A(clknet_6_27__leaf_clk),
    .X(clknet_leaf_113_clk));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_114_clk));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_115_clk));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_116_clk));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_117_clk));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_118_clk));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_119_clk));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_120_clk));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_121_clk));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_122_clk));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_6_49__leaf_clk),
    .X(clknet_leaf_123_clk));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_124_clk));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_6_30__leaf_clk),
    .X(clknet_leaf_125_clk));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_126_clk));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_127_clk));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_128_clk));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_129_clk));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_6_31__leaf_clk),
    .X(clknet_leaf_130_clk));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_131_clk));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_132_clk));
 sg13g2_buf_8 clkbuf_leaf_133_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_133_clk));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_134_clk));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_6_53__leaf_clk),
    .X(clknet_leaf_135_clk));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_136_clk));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_137_clk));
 sg13g2_buf_8 clkbuf_leaf_138_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_138_clk));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_139_clk));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_6_52__leaf_clk),
    .X(clknet_leaf_140_clk));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_141_clk));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_142_clk));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_143_clk));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_144_clk));
 sg13g2_buf_8 clkbuf_leaf_145_clk (.A(clknet_6_54__leaf_clk),
    .X(clknet_leaf_145_clk));
 sg13g2_buf_8 clkbuf_leaf_146_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_146_clk));
 sg13g2_buf_8 clkbuf_leaf_147_clk (.A(clknet_6_55__leaf_clk),
    .X(clknet_leaf_147_clk));
 sg13g2_buf_8 clkbuf_leaf_148_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_148_clk));
 sg13g2_buf_8 clkbuf_leaf_149_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_149_clk));
 sg13g2_buf_8 clkbuf_leaf_150_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_150_clk));
 sg13g2_buf_8 clkbuf_leaf_151_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_151_clk));
 sg13g2_buf_8 clkbuf_leaf_152_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_152_clk));
 sg13g2_buf_8 clkbuf_leaf_153_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_153_clk));
 sg13g2_buf_8 clkbuf_leaf_154_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_154_clk));
 sg13g2_buf_8 clkbuf_leaf_155_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_155_clk));
 sg13g2_buf_8 clkbuf_leaf_156_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_156_clk));
 sg13g2_buf_8 clkbuf_leaf_157_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_157_clk));
 sg13g2_buf_8 clkbuf_leaf_158_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_158_clk));
 sg13g2_buf_8 clkbuf_leaf_159_clk (.A(clknet_6_63__leaf_clk),
    .X(clknet_leaf_159_clk));
 sg13g2_buf_8 clkbuf_leaf_160_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_160_clk));
 sg13g2_buf_8 clkbuf_leaf_161_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_161_clk));
 sg13g2_buf_8 clkbuf_leaf_162_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_162_clk));
 sg13g2_buf_8 clkbuf_leaf_163_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_163_clk));
 sg13g2_buf_8 clkbuf_leaf_164_clk (.A(clknet_6_60__leaf_clk),
    .X(clknet_leaf_164_clk));
 sg13g2_buf_8 clkbuf_leaf_165_clk (.A(clknet_6_61__leaf_clk),
    .X(clknet_leaf_165_clk));
 sg13g2_buf_8 clkbuf_leaf_166_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_166_clk));
 sg13g2_buf_8 clkbuf_leaf_167_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_167_clk));
 sg13g2_buf_8 clkbuf_leaf_168_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_168_clk));
 sg13g2_buf_8 clkbuf_leaf_169_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_169_clk));
 sg13g2_buf_8 clkbuf_leaf_170_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_170_clk));
 sg13g2_buf_8 clkbuf_leaf_171_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_171_clk));
 sg13g2_buf_8 clkbuf_leaf_172_clk (.A(clknet_6_62__leaf_clk),
    .X(clknet_leaf_172_clk));
 sg13g2_buf_8 clkbuf_leaf_173_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_173_clk));
 sg13g2_buf_8 clkbuf_leaf_174_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_174_clk));
 sg13g2_buf_8 clkbuf_leaf_175_clk (.A(clknet_6_59__leaf_clk),
    .X(clknet_leaf_175_clk));
 sg13g2_buf_8 clkbuf_leaf_176_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_176_clk));
 sg13g2_buf_8 clkbuf_leaf_177_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_177_clk));
 sg13g2_buf_8 clkbuf_leaf_178_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_178_clk));
 sg13g2_buf_8 clkbuf_leaf_179_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_179_clk));
 sg13g2_buf_8 clkbuf_leaf_180_clk (.A(clknet_6_58__leaf_clk),
    .X(clknet_leaf_180_clk));
 sg13g2_buf_8 clkbuf_leaf_181_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_181_clk));
 sg13g2_buf_8 clkbuf_leaf_182_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_182_clk));
 sg13g2_buf_8 clkbuf_leaf_183_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_183_clk));
 sg13g2_buf_8 clkbuf_leaf_184_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_184_clk));
 sg13g2_buf_8 clkbuf_leaf_185_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_185_clk));
 sg13g2_buf_8 clkbuf_leaf_186_clk (.A(clknet_6_56__leaf_clk),
    .X(clknet_leaf_186_clk));
 sg13g2_buf_8 clkbuf_leaf_187_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_187_clk));
 sg13g2_buf_8 clkbuf_leaf_188_clk (.A(clknet_6_57__leaf_clk),
    .X(clknet_leaf_188_clk));
 sg13g2_buf_8 clkbuf_leaf_189_clk (.A(clknet_6_51__leaf_clk),
    .X(clknet_leaf_189_clk));
 sg13g2_buf_8 clkbuf_leaf_190_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_190_clk));
 sg13g2_buf_8 clkbuf_leaf_191_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_191_clk));
 sg13g2_buf_8 clkbuf_leaf_192_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_192_clk));
 sg13g2_buf_8 clkbuf_leaf_193_clk (.A(clknet_6_50__leaf_clk),
    .X(clknet_leaf_193_clk));
 sg13g2_buf_8 clkbuf_leaf_194_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_194_clk));
 sg13g2_buf_8 clkbuf_leaf_195_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_195_clk));
 sg13g2_buf_8 clkbuf_leaf_196_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_196_clk));
 sg13g2_buf_8 clkbuf_leaf_197_clk (.A(clknet_6_48__leaf_clk),
    .X(clknet_leaf_197_clk));
 sg13g2_buf_8 clkbuf_leaf_198_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_198_clk));
 sg13g2_buf_8 clkbuf_leaf_199_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_199_clk));
 sg13g2_buf_8 clkbuf_leaf_200_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_200_clk));
 sg13g2_buf_8 clkbuf_leaf_201_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_201_clk));
 sg13g2_buf_8 clkbuf_leaf_202_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_202_clk));
 sg13g2_buf_8 clkbuf_leaf_203_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_203_clk));
 sg13g2_buf_8 clkbuf_leaf_204_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_204_clk));
 sg13g2_buf_8 clkbuf_leaf_205_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_205_clk));
 sg13g2_buf_8 clkbuf_leaf_206_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_206_clk));
 sg13g2_buf_8 clkbuf_leaf_207_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_207_clk));
 sg13g2_buf_8 clkbuf_leaf_208_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_208_clk));
 sg13g2_buf_8 clkbuf_leaf_209_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_209_clk));
 sg13g2_buf_8 clkbuf_leaf_210_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_210_clk));
 sg13g2_buf_8 clkbuf_leaf_211_clk (.A(clknet_6_39__leaf_clk),
    .X(clknet_leaf_211_clk));
 sg13g2_buf_8 clkbuf_leaf_212_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_212_clk));
 sg13g2_buf_8 clkbuf_leaf_213_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_213_clk));
 sg13g2_buf_8 clkbuf_leaf_214_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_214_clk));
 sg13g2_buf_8 clkbuf_leaf_215_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_215_clk));
 sg13g2_buf_8 clkbuf_leaf_216_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_216_clk));
 sg13g2_buf_8 clkbuf_leaf_217_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_217_clk));
 sg13g2_buf_8 clkbuf_leaf_218_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_218_clk));
 sg13g2_buf_8 clkbuf_leaf_219_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_219_clk));
 sg13g2_buf_8 clkbuf_leaf_220_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_220_clk));
 sg13g2_buf_8 clkbuf_leaf_221_clk (.A(clknet_6_47__leaf_clk),
    .X(clknet_leaf_221_clk));
 sg13g2_buf_8 clkbuf_leaf_222_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_222_clk));
 sg13g2_buf_8 clkbuf_leaf_223_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_223_clk));
 sg13g2_buf_8 clkbuf_leaf_224_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_224_clk));
 sg13g2_buf_8 clkbuf_leaf_225_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_225_clk));
 sg13g2_buf_8 clkbuf_leaf_226_clk (.A(clknet_6_45__leaf_clk),
    .X(clknet_leaf_226_clk));
 sg13g2_buf_8 clkbuf_leaf_227_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_227_clk));
 sg13g2_buf_8 clkbuf_leaf_228_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_228_clk));
 sg13g2_buf_8 clkbuf_leaf_229_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_229_clk));
 sg13g2_buf_8 clkbuf_leaf_230_clk (.A(clknet_6_44__leaf_clk),
    .X(clknet_leaf_230_clk));
 sg13g2_buf_8 clkbuf_leaf_231_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_231_clk));
 sg13g2_buf_8 clkbuf_leaf_232_clk (.A(clknet_6_46__leaf_clk),
    .X(clknet_leaf_232_clk));
 sg13g2_buf_8 clkbuf_leaf_233_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_233_clk));
 sg13g2_buf_8 clkbuf_leaf_234_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_234_clk));
 sg13g2_buf_8 clkbuf_leaf_235_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_235_clk));
 sg13g2_buf_8 clkbuf_leaf_236_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_236_clk));
 sg13g2_buf_8 clkbuf_leaf_237_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_237_clk));
 sg13g2_buf_8 clkbuf_leaf_238_clk (.A(clknet_6_43__leaf_clk),
    .X(clknet_leaf_238_clk));
 sg13g2_buf_8 clkbuf_leaf_239_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_239_clk));
 sg13g2_buf_8 clkbuf_leaf_240_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_240_clk));
 sg13g2_buf_8 clkbuf_leaf_241_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_241_clk));
 sg13g2_buf_8 clkbuf_leaf_242_clk (.A(clknet_6_42__leaf_clk),
    .X(clknet_leaf_242_clk));
 sg13g2_buf_8 clkbuf_leaf_243_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_243_clk));
 sg13g2_buf_8 clkbuf_leaf_244_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_244_clk));
 sg13g2_buf_8 clkbuf_leaf_245_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_245_clk));
 sg13g2_buf_8 clkbuf_leaf_246_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_246_clk));
 sg13g2_buf_8 clkbuf_leaf_247_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_247_clk));
 sg13g2_buf_8 clkbuf_leaf_248_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_248_clk));
 sg13g2_buf_8 clkbuf_leaf_249_clk (.A(clknet_6_40__leaf_clk),
    .X(clknet_leaf_249_clk));
 sg13g2_buf_8 clkbuf_leaf_250_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_250_clk));
 sg13g2_buf_8 clkbuf_leaf_251_clk (.A(clknet_6_41__leaf_clk),
    .X(clknet_leaf_251_clk));
 sg13g2_buf_8 clkbuf_leaf_252_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_252_clk));
 sg13g2_buf_8 clkbuf_leaf_253_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_253_clk));
 sg13g2_buf_8 clkbuf_leaf_254_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_254_clk));
 sg13g2_buf_8 clkbuf_leaf_255_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_255_clk));
 sg13g2_buf_8 clkbuf_leaf_256_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_256_clk));
 sg13g2_buf_8 clkbuf_leaf_257_clk (.A(clknet_6_35__leaf_clk),
    .X(clknet_leaf_257_clk));
 sg13g2_buf_8 clkbuf_leaf_258_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_258_clk));
 sg13g2_buf_8 clkbuf_leaf_259_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_259_clk));
 sg13g2_buf_8 clkbuf_leaf_260_clk (.A(clknet_6_34__leaf_clk),
    .X(clknet_leaf_260_clk));
 sg13g2_buf_8 clkbuf_leaf_261_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_261_clk));
 sg13g2_buf_8 clkbuf_leaf_262_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_262_clk));
 sg13g2_buf_8 clkbuf_leaf_263_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_263_clk));
 sg13g2_buf_8 clkbuf_leaf_264_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_264_clk));
 sg13g2_buf_8 clkbuf_leaf_265_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_265_clk));
 sg13g2_buf_8 clkbuf_leaf_266_clk (.A(clknet_6_32__leaf_clk),
    .X(clknet_leaf_266_clk));
 sg13g2_buf_8 clkbuf_leaf_267_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_267_clk));
 sg13g2_buf_8 clkbuf_leaf_268_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_268_clk));
 sg13g2_buf_8 clkbuf_leaf_269_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_269_clk));
 sg13g2_buf_8 clkbuf_leaf_270_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_270_clk));
 sg13g2_buf_8 clkbuf_leaf_271_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_271_clk));
 sg13g2_buf_8 clkbuf_leaf_272_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_272_clk));
 sg13g2_buf_8 clkbuf_leaf_273_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_273_clk));
 sg13g2_buf_8 clkbuf_leaf_274_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_274_clk));
 sg13g2_buf_8 clkbuf_leaf_275_clk (.A(clknet_6_38__leaf_clk),
    .X(clknet_leaf_275_clk));
 sg13g2_buf_8 clkbuf_leaf_276_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_276_clk));
 sg13g2_buf_8 clkbuf_leaf_277_clk (.A(clknet_6_36__leaf_clk),
    .X(clknet_leaf_277_clk));
 sg13g2_buf_8 clkbuf_leaf_278_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_278_clk));
 sg13g2_buf_8 clkbuf_leaf_279_clk (.A(clknet_6_33__leaf_clk),
    .X(clknet_leaf_279_clk));
 sg13g2_buf_8 clkbuf_leaf_280_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_280_clk));
 sg13g2_buf_8 clkbuf_leaf_281_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_281_clk));
 sg13g2_buf_8 clkbuf_leaf_282_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_282_clk));
 sg13g2_buf_8 clkbuf_leaf_283_clk (.A(clknet_6_37__leaf_clk),
    .X(clknet_leaf_283_clk));
 sg13g2_buf_8 clkbuf_leaf_284_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_284_clk));
 sg13g2_buf_8 clkbuf_leaf_285_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_285_clk));
 sg13g2_buf_8 clkbuf_leaf_286_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_286_clk));
 sg13g2_buf_8 clkbuf_leaf_287_clk (.A(clknet_6_15__leaf_clk),
    .X(clknet_leaf_287_clk));
 sg13g2_buf_8 clkbuf_leaf_288_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_288_clk));
 sg13g2_buf_8 clkbuf_leaf_289_clk (.A(clknet_6_13__leaf_clk),
    .X(clknet_leaf_289_clk));
 sg13g2_buf_8 clkbuf_leaf_290_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_290_clk));
 sg13g2_buf_8 clkbuf_leaf_291_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_291_clk));
 sg13g2_buf_8 clkbuf_leaf_292_clk (.A(clknet_6_14__leaf_clk),
    .X(clknet_leaf_292_clk));
 sg13g2_buf_8 clkbuf_leaf_293_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_293_clk));
 sg13g2_buf_8 clkbuf_leaf_294_clk (.A(clknet_6_12__leaf_clk),
    .X(clknet_leaf_294_clk));
 sg13g2_buf_8 clkbuf_leaf_295_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_295_clk));
 sg13g2_buf_8 clkbuf_leaf_296_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_296_clk));
 sg13g2_buf_8 clkbuf_leaf_297_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_297_clk));
 sg13g2_buf_8 clkbuf_leaf_298_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_298_clk));
 sg13g2_buf_8 clkbuf_leaf_299_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_299_clk));
 sg13g2_buf_8 clkbuf_leaf_300_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_300_clk));
 sg13g2_buf_8 clkbuf_leaf_301_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_301_clk));
 sg13g2_buf_8 clkbuf_leaf_302_clk (.A(clknet_6_11__leaf_clk),
    .X(clknet_leaf_302_clk));
 sg13g2_buf_8 clkbuf_leaf_303_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_303_clk));
 sg13g2_buf_8 clkbuf_leaf_304_clk (.A(clknet_6_9__leaf_clk),
    .X(clknet_leaf_304_clk));
 sg13g2_buf_8 clkbuf_leaf_305_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_305_clk));
 sg13g2_buf_8 clkbuf_leaf_306_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_306_clk));
 sg13g2_buf_8 clkbuf_leaf_307_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_307_clk));
 sg13g2_buf_8 clkbuf_leaf_308_clk (.A(clknet_6_10__leaf_clk),
    .X(clknet_leaf_308_clk));
 sg13g2_buf_8 clkbuf_leaf_309_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_309_clk));
 sg13g2_buf_8 clkbuf_leaf_310_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_310_clk));
 sg13g2_buf_8 clkbuf_leaf_311_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_311_clk));
 sg13g2_buf_8 clkbuf_leaf_312_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_312_clk));
 sg13g2_buf_8 clkbuf_leaf_313_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_313_clk));
 sg13g2_buf_8 clkbuf_leaf_314_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_314_clk));
 sg13g2_buf_8 clkbuf_leaf_315_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_315_clk));
 sg13g2_buf_8 clkbuf_leaf_316_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_316_clk));
 sg13g2_buf_8 clkbuf_leaf_317_clk (.A(clknet_6_8__leaf_clk),
    .X(clknet_leaf_317_clk));
 sg13g2_buf_8 clkbuf_leaf_318_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_318_clk));
 sg13g2_buf_8 clkbuf_leaf_319_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_319_clk));
 sg13g2_buf_8 clkbuf_leaf_320_clk (.A(clknet_6_3__leaf_clk),
    .X(clknet_leaf_320_clk));
 sg13g2_buf_8 clkbuf_leaf_321_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_321_clk));
 sg13g2_buf_8 clkbuf_leaf_322_clk (.A(clknet_6_2__leaf_clk),
    .X(clknet_leaf_322_clk));
 sg13g2_buf_8 clkbuf_leaf_323_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_323_clk));
 sg13g2_buf_8 clkbuf_leaf_324_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_324_clk));
 sg13g2_buf_8 clkbuf_leaf_325_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_325_clk));
 sg13g2_buf_8 clkbuf_leaf_326_clk (.A(clknet_6_0__leaf_clk),
    .X(clknet_leaf_326_clk));
 sg13g2_buf_4 clkbuf_0_clk (.X(clknet_0_clk),
    .A(clk));
 sg13g2_buf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sg13g2_buf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sg13g2_buf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sg13g2_buf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sg13g2_buf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sg13g2_buf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sg13g2_buf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sg13g2_buf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_0__f_clk (.X(clknet_6_0__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_1__f_clk (.X(clknet_6_1__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_2__f_clk (.X(clknet_6_2__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_3__f_clk (.X(clknet_6_3__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_4__f_clk (.X(clknet_6_4__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_5__f_clk (.X(clknet_6_5__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_6__f_clk (.X(clknet_6_6__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_7__f_clk (.X(clknet_6_7__leaf_clk),
    .A(clknet_3_0_0_clk));
 sg13g2_buf_4 clkbuf_6_8__f_clk (.X(clknet_6_8__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_9__f_clk (.X(clknet_6_9__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_10__f_clk (.X(clknet_6_10__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_11__f_clk (.X(clknet_6_11__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_12__f_clk (.X(clknet_6_12__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_13__f_clk (.X(clknet_6_13__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_14__f_clk (.X(clknet_6_14__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_15__f_clk (.X(clknet_6_15__leaf_clk),
    .A(clknet_3_1_0_clk));
 sg13g2_buf_4 clkbuf_6_16__f_clk (.X(clknet_6_16__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_17__f_clk (.X(clknet_6_17__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_18__f_clk (.X(clknet_6_18__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_19__f_clk (.X(clknet_6_19__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_20__f_clk (.X(clknet_6_20__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_21__f_clk (.X(clknet_6_21__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_22__f_clk (.X(clknet_6_22__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_23__f_clk (.X(clknet_6_23__leaf_clk),
    .A(clknet_3_2_0_clk));
 sg13g2_buf_4 clkbuf_6_24__f_clk (.X(clknet_6_24__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_25__f_clk (.X(clknet_6_25__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_26__f_clk (.X(clknet_6_26__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_27__f_clk (.X(clknet_6_27__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_28__f_clk (.X(clknet_6_28__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_29__f_clk (.X(clknet_6_29__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_30__f_clk (.X(clknet_6_30__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_31__f_clk (.X(clknet_6_31__leaf_clk),
    .A(clknet_3_3_0_clk));
 sg13g2_buf_4 clkbuf_6_32__f_clk (.X(clknet_6_32__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_33__f_clk (.X(clknet_6_33__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_34__f_clk (.X(clknet_6_34__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_35__f_clk (.X(clknet_6_35__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_36__f_clk (.X(clknet_6_36__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_37__f_clk (.X(clknet_6_37__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_38__f_clk (.X(clknet_6_38__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_39__f_clk (.X(clknet_6_39__leaf_clk),
    .A(clknet_3_4_0_clk));
 sg13g2_buf_4 clkbuf_6_40__f_clk (.X(clknet_6_40__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_41__f_clk (.X(clknet_6_41__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_42__f_clk (.X(clknet_6_42__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_43__f_clk (.X(clknet_6_43__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_44__f_clk (.X(clknet_6_44__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_45__f_clk (.X(clknet_6_45__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_46__f_clk (.X(clknet_6_46__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_47__f_clk (.X(clknet_6_47__leaf_clk),
    .A(clknet_3_5_0_clk));
 sg13g2_buf_4 clkbuf_6_48__f_clk (.X(clknet_6_48__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_49__f_clk (.X(clknet_6_49__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_50__f_clk (.X(clknet_6_50__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_51__f_clk (.X(clknet_6_51__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_52__f_clk (.X(clknet_6_52__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_53__f_clk (.X(clknet_6_53__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_54__f_clk (.X(clknet_6_54__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_55__f_clk (.X(clknet_6_55__leaf_clk),
    .A(clknet_3_6_0_clk));
 sg13g2_buf_4 clkbuf_6_56__f_clk (.X(clknet_6_56__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_57__f_clk (.X(clknet_6_57__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_58__f_clk (.X(clknet_6_58__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_59__f_clk (.X(clknet_6_59__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_60__f_clk (.X(clknet_6_60__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_61__f_clk (.X(clknet_6_61__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_62__f_clk (.X(clknet_6_62__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_4 clkbuf_6_63__f_clk (.X(clknet_6_63__leaf_clk),
    .A(clknet_3_7_0_clk));
 sg13g2_buf_8 clkload0 (.A(clknet_6_1__leaf_clk));
 sg13g2_buf_8 clkload1 (.A(clknet_6_2__leaf_clk));
 sg13g2_buf_8 clkload2 (.A(clknet_6_3__leaf_clk));
 sg13g2_buf_8 clkload3 (.A(clknet_6_4__leaf_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_6_5__leaf_clk));
 sg13g2_buf_8 clkload5 (.A(clknet_6_6__leaf_clk));
 sg13g2_buf_8 clkload6 (.A(clknet_6_7__leaf_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_6_9__leaf_clk));
 sg13g2_buf_8 clkload8 (.A(clknet_6_10__leaf_clk));
 sg13g2_buf_8 clkload9 (.A(clknet_6_11__leaf_clk));
 sg13g2_buf_8 clkload10 (.A(clknet_6_12__leaf_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_6_13__leaf_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_6_14__leaf_clk));
 sg13g2_buf_8 clkload13 (.A(clknet_6_15__leaf_clk));
 sg13g2_buf_8 clkload14 (.A(clknet_6_17__leaf_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_6_18__leaf_clk));
 sg13g2_buf_8 clkload16 (.A(clknet_6_19__leaf_clk));
 sg13g2_buf_8 clkload17 (.A(clknet_6_20__leaf_clk));
 sg13g2_buf_8 clkload18 (.A(clknet_6_21__leaf_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_6_22__leaf_clk));
 sg13g2_buf_8 clkload20 (.A(clknet_6_23__leaf_clk));
 sg13g2_buf_8 clkload21 (.A(clknet_6_25__leaf_clk));
 sg13g2_buf_8 clkload22 (.A(clknet_6_26__leaf_clk));
 sg13g2_buf_8 clkload23 (.A(clknet_6_27__leaf_clk));
 sg13g2_buf_8 clkload24 (.A(clknet_6_28__leaf_clk));
 sg13g2_buf_8 clkload25 (.A(clknet_6_29__leaf_clk));
 sg13g2_buf_8 clkload26 (.A(clknet_6_30__leaf_clk));
 sg13g2_buf_8 clkload27 (.A(clknet_6_31__leaf_clk));
 sg13g2_buf_8 clkload28 (.A(clknet_6_33__leaf_clk));
 sg13g2_buf_8 clkload29 (.A(clknet_6_34__leaf_clk));
 sg13g2_buf_8 clkload30 (.A(clknet_6_35__leaf_clk));
 sg13g2_buf_8 clkload31 (.A(clknet_6_36__leaf_clk));
 sg13g2_buf_8 clkload32 (.A(clknet_6_37__leaf_clk));
 sg13g2_buf_8 clkload33 (.A(clknet_6_38__leaf_clk));
 sg13g2_buf_8 clkload34 (.A(clknet_6_39__leaf_clk));
 sg13g2_buf_8 clkload35 (.A(clknet_6_41__leaf_clk));
 sg13g2_buf_8 clkload36 (.A(clknet_6_42__leaf_clk));
 sg13g2_buf_8 clkload37 (.A(clknet_6_43__leaf_clk));
 sg13g2_buf_8 clkload38 (.A(clknet_6_44__leaf_clk));
 sg13g2_buf_8 clkload39 (.A(clknet_6_45__leaf_clk));
 sg13g2_buf_8 clkload40 (.A(clknet_6_46__leaf_clk));
 sg13g2_buf_8 clkload41 (.A(clknet_6_47__leaf_clk));
 sg13g2_buf_8 clkload42 (.A(clknet_6_49__leaf_clk));
 sg13g2_buf_8 clkload43 (.A(clknet_6_50__leaf_clk));
 sg13g2_buf_8 clkload44 (.A(clknet_6_51__leaf_clk));
 sg13g2_buf_8 clkload45 (.A(clknet_6_52__leaf_clk));
 sg13g2_buf_8 clkload46 (.A(clknet_6_53__leaf_clk));
 sg13g2_buf_8 clkload47 (.A(clknet_6_54__leaf_clk));
 sg13g2_buf_8 clkload48 (.A(clknet_6_55__leaf_clk));
 sg13g2_inv_4 clkload49 (.A(clknet_leaf_325_clk));
 sg13g2_inv_2 clkload50 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload51 (.A(clknet_leaf_57_clk));
 sg13g2_inv_2 clkload52 (.A(clknet_leaf_37_clk));
 sg13g2_inv_4 clkload53 (.A(clknet_leaf_199_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_00356_));
 sg13g2_antennanp ANTENNA_2 (.A(_00410_));
 sg13g2_antennanp ANTENNA_3 (.A(_00422_));
 sg13g2_antennanp ANTENNA_4 (.A(_00425_));
 sg13g2_antennanp ANTENNA_5 (.A(_00432_));
 sg13g2_antennanp ANTENNA_6 (.A(_00443_));
 sg13g2_antennanp ANTENNA_7 (.A(_00443_));
 sg13g2_antennanp ANTENNA_8 (.A(_02799_));
 sg13g2_antennanp ANTENNA_9 (.A(_02799_));
 sg13g2_antennanp ANTENNA_10 (.A(_02924_));
 sg13g2_antennanp ANTENNA_11 (.A(_02924_));
 sg13g2_antennanp ANTENNA_12 (.A(_02924_));
 sg13g2_antennanp ANTENNA_13 (.A(_02924_));
 sg13g2_antennanp ANTENNA_14 (.A(_02935_));
 sg13g2_antennanp ANTENNA_15 (.A(_02935_));
 sg13g2_antennanp ANTENNA_16 (.A(_02935_));
 sg13g2_antennanp ANTENNA_17 (.A(_02946_));
 sg13g2_antennanp ANTENNA_18 (.A(_02946_));
 sg13g2_antennanp ANTENNA_19 (.A(_02946_));
 sg13g2_antennanp ANTENNA_20 (.A(_02946_));
 sg13g2_antennanp ANTENNA_21 (.A(_03019_));
 sg13g2_antennanp ANTENNA_22 (.A(_03019_));
 sg13g2_antennanp ANTENNA_23 (.A(_03019_));
 sg13g2_antennanp ANTENNA_24 (.A(_03019_));
 sg13g2_antennanp ANTENNA_25 (.A(_03055_));
 sg13g2_antennanp ANTENNA_26 (.A(_03055_));
 sg13g2_antennanp ANTENNA_27 (.A(_03055_));
 sg13g2_antennanp ANTENNA_28 (.A(_03060_));
 sg13g2_antennanp ANTENNA_29 (.A(_03060_));
 sg13g2_antennanp ANTENNA_30 (.A(_03060_));
 sg13g2_antennanp ANTENNA_31 (.A(_03079_));
 sg13g2_antennanp ANTENNA_32 (.A(_03079_));
 sg13g2_antennanp ANTENNA_33 (.A(_03079_));
 sg13g2_antennanp ANTENNA_34 (.A(_03079_));
 sg13g2_antennanp ANTENNA_35 (.A(_03184_));
 sg13g2_antennanp ANTENNA_36 (.A(_03184_));
 sg13g2_antennanp ANTENNA_37 (.A(_03184_));
 sg13g2_antennanp ANTENNA_38 (.A(_03184_));
 sg13g2_antennanp ANTENNA_39 (.A(_03184_));
 sg13g2_antennanp ANTENNA_40 (.A(_03268_));
 sg13g2_antennanp ANTENNA_41 (.A(_03268_));
 sg13g2_antennanp ANTENNA_42 (.A(_03268_));
 sg13g2_antennanp ANTENNA_43 (.A(_03684_));
 sg13g2_antennanp ANTENNA_44 (.A(_03684_));
 sg13g2_antennanp ANTENNA_45 (.A(_03714_));
 sg13g2_antennanp ANTENNA_46 (.A(_03714_));
 sg13g2_antennanp ANTENNA_47 (.A(_03714_));
 sg13g2_antennanp ANTENNA_48 (.A(_03760_));
 sg13g2_antennanp ANTENNA_49 (.A(_03760_));
 sg13g2_antennanp ANTENNA_50 (.A(_03760_));
 sg13g2_antennanp ANTENNA_51 (.A(_03760_));
 sg13g2_antennanp ANTENNA_52 (.A(_03760_));
 sg13g2_antennanp ANTENNA_53 (.A(_03760_));
 sg13g2_antennanp ANTENNA_54 (.A(_03776_));
 sg13g2_antennanp ANTENNA_55 (.A(_03776_));
 sg13g2_antennanp ANTENNA_56 (.A(_03776_));
 sg13g2_antennanp ANTENNA_57 (.A(_03776_));
 sg13g2_antennanp ANTENNA_58 (.A(_03776_));
 sg13g2_antennanp ANTENNA_59 (.A(_03776_));
 sg13g2_antennanp ANTENNA_60 (.A(_04617_));
 sg13g2_antennanp ANTENNA_61 (.A(_04617_));
 sg13g2_antennanp ANTENNA_62 (.A(_04617_));
 sg13g2_antennanp ANTENNA_63 (.A(_04617_));
 sg13g2_antennanp ANTENNA_64 (.A(_04617_));
 sg13g2_antennanp ANTENNA_65 (.A(_04617_));
 sg13g2_antennanp ANTENNA_66 (.A(_04617_));
 sg13g2_antennanp ANTENNA_67 (.A(_04617_));
 sg13g2_antennanp ANTENNA_68 (.A(_04617_));
 sg13g2_antennanp ANTENNA_69 (.A(_04617_));
 sg13g2_antennanp ANTENNA_70 (.A(_04617_));
 sg13g2_antennanp ANTENNA_71 (.A(_04617_));
 sg13g2_antennanp ANTENNA_72 (.A(_04617_));
 sg13g2_antennanp ANTENNA_73 (.A(_04617_));
 sg13g2_antennanp ANTENNA_74 (.A(_04617_));
 sg13g2_antennanp ANTENNA_75 (.A(_04617_));
 sg13g2_antennanp ANTENNA_76 (.A(_04617_));
 sg13g2_antennanp ANTENNA_77 (.A(_04617_));
 sg13g2_antennanp ANTENNA_78 (.A(_04617_));
 sg13g2_antennanp ANTENNA_79 (.A(_04617_));
 sg13g2_antennanp ANTENNA_80 (.A(_04617_));
 sg13g2_antennanp ANTENNA_81 (.A(_04617_));
 sg13g2_antennanp ANTENNA_82 (.A(_04617_));
 sg13g2_antennanp ANTENNA_83 (.A(_04617_));
 sg13g2_antennanp ANTENNA_84 (.A(_04617_));
 sg13g2_antennanp ANTENNA_85 (.A(_04620_));
 sg13g2_antennanp ANTENNA_86 (.A(_04674_));
 sg13g2_antennanp ANTENNA_87 (.A(_04676_));
 sg13g2_antennanp ANTENNA_88 (.A(_05061_));
 sg13g2_antennanp ANTENNA_89 (.A(_05067_));
 sg13g2_antennanp ANTENNA_90 (.A(_05091_));
 sg13g2_antennanp ANTENNA_91 (.A(_05275_));
 sg13g2_antennanp ANTENNA_92 (.A(_05275_));
 sg13g2_antennanp ANTENNA_93 (.A(_05275_));
 sg13g2_antennanp ANTENNA_94 (.A(_05275_));
 sg13g2_antennanp ANTENNA_95 (.A(_05275_));
 sg13g2_antennanp ANTENNA_96 (.A(_05275_));
 sg13g2_antennanp ANTENNA_97 (.A(_05275_));
 sg13g2_antennanp ANTENNA_98 (.A(_05275_));
 sg13g2_antennanp ANTENNA_99 (.A(_05276_));
 sg13g2_antennanp ANTENNA_100 (.A(_05276_));
 sg13g2_antennanp ANTENNA_101 (.A(_05276_));
 sg13g2_antennanp ANTENNA_102 (.A(_05276_));
 sg13g2_antennanp ANTENNA_103 (.A(_05278_));
 sg13g2_antennanp ANTENNA_104 (.A(_05290_));
 sg13g2_antennanp ANTENNA_105 (.A(_05298_));
 sg13g2_antennanp ANTENNA_106 (.A(_05298_));
 sg13g2_antennanp ANTENNA_107 (.A(_05298_));
 sg13g2_antennanp ANTENNA_108 (.A(_05298_));
 sg13g2_antennanp ANTENNA_109 (.A(_05298_));
 sg13g2_antennanp ANTENNA_110 (.A(_05298_));
 sg13g2_antennanp ANTENNA_111 (.A(_05298_));
 sg13g2_antennanp ANTENNA_112 (.A(_05303_));
 sg13g2_antennanp ANTENNA_113 (.A(_05303_));
 sg13g2_antennanp ANTENNA_114 (.A(_05303_));
 sg13g2_antennanp ANTENNA_115 (.A(_05318_));
 sg13g2_antennanp ANTENNA_116 (.A(_05347_));
 sg13g2_antennanp ANTENNA_117 (.A(_05347_));
 sg13g2_antennanp ANTENNA_118 (.A(_05347_));
 sg13g2_antennanp ANTENNA_119 (.A(_05347_));
 sg13g2_antennanp ANTENNA_120 (.A(_05347_));
 sg13g2_antennanp ANTENNA_121 (.A(_05350_));
 sg13g2_antennanp ANTENNA_122 (.A(_05364_));
 sg13g2_antennanp ANTENNA_123 (.A(_05417_));
 sg13g2_antennanp ANTENNA_124 (.A(_05417_));
 sg13g2_antennanp ANTENNA_125 (.A(_05432_));
 sg13g2_antennanp ANTENNA_126 (.A(_05465_));
 sg13g2_antennanp ANTENNA_127 (.A(_05465_));
 sg13g2_antennanp ANTENNA_128 (.A(_05465_));
 sg13g2_antennanp ANTENNA_129 (.A(_05465_));
 sg13g2_antennanp ANTENNA_130 (.A(_05510_));
 sg13g2_antennanp ANTENNA_131 (.A(_05510_));
 sg13g2_antennanp ANTENNA_132 (.A(_05510_));
 sg13g2_antennanp ANTENNA_133 (.A(_05510_));
 sg13g2_antennanp ANTENNA_134 (.A(_05512_));
 sg13g2_antennanp ANTENNA_135 (.A(_05577_));
 sg13g2_antennanp ANTENNA_136 (.A(_05584_));
 sg13g2_antennanp ANTENNA_137 (.A(_05600_));
 sg13g2_antennanp ANTENNA_138 (.A(_05600_));
 sg13g2_antennanp ANTENNA_139 (.A(_05600_));
 sg13g2_antennanp ANTENNA_140 (.A(_05640_));
 sg13g2_antennanp ANTENNA_141 (.A(_05640_));
 sg13g2_antennanp ANTENNA_142 (.A(_05640_));
 sg13g2_antennanp ANTENNA_143 (.A(_05652_));
 sg13g2_antennanp ANTENNA_144 (.A(_05652_));
 sg13g2_antennanp ANTENNA_145 (.A(_05652_));
 sg13g2_antennanp ANTENNA_146 (.A(_05652_));
 sg13g2_antennanp ANTENNA_147 (.A(_05652_));
 sg13g2_antennanp ANTENNA_148 (.A(_05659_));
 sg13g2_antennanp ANTENNA_149 (.A(_05659_));
 sg13g2_antennanp ANTENNA_150 (.A(_05659_));
 sg13g2_antennanp ANTENNA_151 (.A(_05662_));
 sg13g2_antennanp ANTENNA_152 (.A(_05662_));
 sg13g2_antennanp ANTENNA_153 (.A(_05662_));
 sg13g2_antennanp ANTENNA_154 (.A(_05662_));
 sg13g2_antennanp ANTENNA_155 (.A(_05663_));
 sg13g2_antennanp ANTENNA_156 (.A(_05663_));
 sg13g2_antennanp ANTENNA_157 (.A(_05663_));
 sg13g2_antennanp ANTENNA_158 (.A(_05663_));
 sg13g2_antennanp ANTENNA_159 (.A(_05672_));
 sg13g2_antennanp ANTENNA_160 (.A(_05707_));
 sg13g2_antennanp ANTENNA_161 (.A(_05707_));
 sg13g2_antennanp ANTENNA_162 (.A(_05707_));
 sg13g2_antennanp ANTENNA_163 (.A(_05754_));
 sg13g2_antennanp ANTENNA_164 (.A(_05755_));
 sg13g2_antennanp ANTENNA_165 (.A(_05778_));
 sg13g2_antennanp ANTENNA_166 (.A(_05778_));
 sg13g2_antennanp ANTENNA_167 (.A(_05778_));
 sg13g2_antennanp ANTENNA_168 (.A(_05778_));
 sg13g2_antennanp ANTENNA_169 (.A(_05784_));
 sg13g2_antennanp ANTENNA_170 (.A(_05784_));
 sg13g2_antennanp ANTENNA_171 (.A(_05784_));
 sg13g2_antennanp ANTENNA_172 (.A(_05784_));
 sg13g2_antennanp ANTENNA_173 (.A(_05784_));
 sg13g2_antennanp ANTENNA_174 (.A(_05784_));
 sg13g2_antennanp ANTENNA_175 (.A(_05784_));
 sg13g2_antennanp ANTENNA_176 (.A(_05784_));
 sg13g2_antennanp ANTENNA_177 (.A(_05784_));
 sg13g2_antennanp ANTENNA_178 (.A(_05784_));
 sg13g2_antennanp ANTENNA_179 (.A(_05788_));
 sg13g2_antennanp ANTENNA_180 (.A(_05788_));
 sg13g2_antennanp ANTENNA_181 (.A(_05788_));
 sg13g2_antennanp ANTENNA_182 (.A(_05804_));
 sg13g2_antennanp ANTENNA_183 (.A(_05811_));
 sg13g2_antennanp ANTENNA_184 (.A(_05811_));
 sg13g2_antennanp ANTENNA_185 (.A(_05811_));
 sg13g2_antennanp ANTENNA_186 (.A(_05811_));
 sg13g2_antennanp ANTENNA_187 (.A(_05851_));
 sg13g2_antennanp ANTENNA_188 (.A(_05851_));
 sg13g2_antennanp ANTENNA_189 (.A(_05851_));
 sg13g2_antennanp ANTENNA_190 (.A(_05851_));
 sg13g2_antennanp ANTENNA_191 (.A(_05868_));
 sg13g2_antennanp ANTENNA_192 (.A(_05872_));
 sg13g2_antennanp ANTENNA_193 (.A(_05891_));
 sg13g2_antennanp ANTENNA_194 (.A(_05892_));
 sg13g2_antennanp ANTENNA_195 (.A(_05892_));
 sg13g2_antennanp ANTENNA_196 (.A(_05892_));
 sg13g2_antennanp ANTENNA_197 (.A(_05901_));
 sg13g2_antennanp ANTENNA_198 (.A(_05901_));
 sg13g2_antennanp ANTENNA_199 (.A(_05901_));
 sg13g2_antennanp ANTENNA_200 (.A(_05918_));
 sg13g2_antennanp ANTENNA_201 (.A(_05918_));
 sg13g2_antennanp ANTENNA_202 (.A(_05918_));
 sg13g2_antennanp ANTENNA_203 (.A(_05918_));
 sg13g2_antennanp ANTENNA_204 (.A(_05918_));
 sg13g2_antennanp ANTENNA_205 (.A(_05918_));
 sg13g2_antennanp ANTENNA_206 (.A(_05918_));
 sg13g2_antennanp ANTENNA_207 (.A(_05918_));
 sg13g2_antennanp ANTENNA_208 (.A(_05918_));
 sg13g2_antennanp ANTENNA_209 (.A(_05918_));
 sg13g2_antennanp ANTENNA_210 (.A(_05918_));
 sg13g2_antennanp ANTENNA_211 (.A(_05918_));
 sg13g2_antennanp ANTENNA_212 (.A(_05918_));
 sg13g2_antennanp ANTENNA_213 (.A(_05918_));
 sg13g2_antennanp ANTENNA_214 (.A(_05918_));
 sg13g2_antennanp ANTENNA_215 (.A(_05918_));
 sg13g2_antennanp ANTENNA_216 (.A(_05918_));
 sg13g2_antennanp ANTENNA_217 (.A(_05918_));
 sg13g2_antennanp ANTENNA_218 (.A(_05918_));
 sg13g2_antennanp ANTENNA_219 (.A(_05918_));
 sg13g2_antennanp ANTENNA_220 (.A(_05932_));
 sg13g2_antennanp ANTENNA_221 (.A(_05932_));
 sg13g2_antennanp ANTENNA_222 (.A(_05932_));
 sg13g2_antennanp ANTENNA_223 (.A(_05932_));
 sg13g2_antennanp ANTENNA_224 (.A(_05932_));
 sg13g2_antennanp ANTENNA_225 (.A(_05932_));
 sg13g2_antennanp ANTENNA_226 (.A(_05936_));
 sg13g2_antennanp ANTENNA_227 (.A(_05940_));
 sg13g2_antennanp ANTENNA_228 (.A(_05953_));
 sg13g2_antennanp ANTENNA_229 (.A(_05975_));
 sg13g2_antennanp ANTENNA_230 (.A(_05975_));
 sg13g2_antennanp ANTENNA_231 (.A(_05975_));
 sg13g2_antennanp ANTENNA_232 (.A(_05975_));
 sg13g2_antennanp ANTENNA_233 (.A(_06009_));
 sg13g2_antennanp ANTENNA_234 (.A(_06009_));
 sg13g2_antennanp ANTENNA_235 (.A(_06009_));
 sg13g2_antennanp ANTENNA_236 (.A(_06009_));
 sg13g2_antennanp ANTENNA_237 (.A(_06009_));
 sg13g2_antennanp ANTENNA_238 (.A(_06009_));
 sg13g2_antennanp ANTENNA_239 (.A(_06027_));
 sg13g2_antennanp ANTENNA_240 (.A(_06076_));
 sg13g2_antennanp ANTENNA_241 (.A(_06090_));
 sg13g2_antennanp ANTENNA_242 (.A(_06101_));
 sg13g2_antennanp ANTENNA_243 (.A(_06108_));
 sg13g2_antennanp ANTENNA_244 (.A(_06108_));
 sg13g2_antennanp ANTENNA_245 (.A(_06108_));
 sg13g2_antennanp ANTENNA_246 (.A(_06154_));
 sg13g2_antennanp ANTENNA_247 (.A(_06154_));
 sg13g2_antennanp ANTENNA_248 (.A(_06154_));
 sg13g2_antennanp ANTENNA_249 (.A(_06154_));
 sg13g2_antennanp ANTENNA_250 (.A(_06154_));
 sg13g2_antennanp ANTENNA_251 (.A(_06154_));
 sg13g2_antennanp ANTENNA_252 (.A(_06184_));
 sg13g2_antennanp ANTENNA_253 (.A(_06214_));
 sg13g2_antennanp ANTENNA_254 (.A(_06235_));
 sg13g2_antennanp ANTENNA_255 (.A(_06235_));
 sg13g2_antennanp ANTENNA_256 (.A(_06235_));
 sg13g2_antennanp ANTENNA_257 (.A(_06244_));
 sg13g2_antennanp ANTENNA_258 (.A(_06254_));
 sg13g2_antennanp ANTENNA_259 (.A(_06255_));
 sg13g2_antennanp ANTENNA_260 (.A(_06265_));
 sg13g2_antennanp ANTENNA_261 (.A(_06302_));
 sg13g2_antennanp ANTENNA_262 (.A(_06302_));
 sg13g2_antennanp ANTENNA_263 (.A(_06306_));
 sg13g2_antennanp ANTENNA_264 (.A(_06309_));
 sg13g2_antennanp ANTENNA_265 (.A(_06313_));
 sg13g2_antennanp ANTENNA_266 (.A(_06313_));
 sg13g2_antennanp ANTENNA_267 (.A(_06313_));
 sg13g2_antennanp ANTENNA_268 (.A(_06313_));
 sg13g2_antennanp ANTENNA_269 (.A(_06317_));
 sg13g2_antennanp ANTENNA_270 (.A(_06317_));
 sg13g2_antennanp ANTENNA_271 (.A(_06317_));
 sg13g2_antennanp ANTENNA_272 (.A(_06317_));
 sg13g2_antennanp ANTENNA_273 (.A(_06330_));
 sg13g2_antennanp ANTENNA_274 (.A(_06345_));
 sg13g2_antennanp ANTENNA_275 (.A(_06351_));
 sg13g2_antennanp ANTENNA_276 (.A(_06359_));
 sg13g2_antennanp ANTENNA_277 (.A(_06409_));
 sg13g2_antennanp ANTENNA_278 (.A(_06409_));
 sg13g2_antennanp ANTENNA_279 (.A(_06440_));
 sg13g2_antennanp ANTENNA_280 (.A(_06443_));
 sg13g2_antennanp ANTENNA_281 (.A(_06447_));
 sg13g2_antennanp ANTENNA_282 (.A(_06467_));
 sg13g2_antennanp ANTENNA_283 (.A(_06489_));
 sg13g2_antennanp ANTENNA_284 (.A(_06518_));
 sg13g2_antennanp ANTENNA_285 (.A(_06518_));
 sg13g2_antennanp ANTENNA_286 (.A(_06518_));
 sg13g2_antennanp ANTENNA_287 (.A(_06518_));
 sg13g2_antennanp ANTENNA_288 (.A(_06530_));
 sg13g2_antennanp ANTENNA_289 (.A(_06533_));
 sg13g2_antennanp ANTENNA_290 (.A(_06538_));
 sg13g2_antennanp ANTENNA_291 (.A(_06545_));
 sg13g2_antennanp ANTENNA_292 (.A(_06550_));
 sg13g2_antennanp ANTENNA_293 (.A(_06587_));
 sg13g2_antennanp ANTENNA_294 (.A(_06591_));
 sg13g2_antennanp ANTENNA_295 (.A(_06591_));
 sg13g2_antennanp ANTENNA_296 (.A(_06601_));
 sg13g2_antennanp ANTENNA_297 (.A(_06601_));
 sg13g2_antennanp ANTENNA_298 (.A(_06601_));
 sg13g2_antennanp ANTENNA_299 (.A(_06601_));
 sg13g2_antennanp ANTENNA_300 (.A(_06603_));
 sg13g2_antennanp ANTENNA_301 (.A(_06609_));
 sg13g2_antennanp ANTENNA_302 (.A(_06619_));
 sg13g2_antennanp ANTENNA_303 (.A(_06651_));
 sg13g2_antennanp ANTENNA_304 (.A(_06654_));
 sg13g2_antennanp ANTENNA_305 (.A(_06662_));
 sg13g2_antennanp ANTENNA_306 (.A(_06671_));
 sg13g2_antennanp ANTENNA_307 (.A(_06708_));
 sg13g2_antennanp ANTENNA_308 (.A(_06708_));
 sg13g2_antennanp ANTENNA_309 (.A(_06708_));
 sg13g2_antennanp ANTENNA_310 (.A(_06716_));
 sg13g2_antennanp ANTENNA_311 (.A(_06721_));
 sg13g2_antennanp ANTENNA_312 (.A(_06722_));
 sg13g2_antennanp ANTENNA_313 (.A(_06735_));
 sg13g2_antennanp ANTENNA_314 (.A(_06740_));
 sg13g2_antennanp ANTENNA_315 (.A(_06741_));
 sg13g2_antennanp ANTENNA_316 (.A(_06751_));
 sg13g2_antennanp ANTENNA_317 (.A(_06780_));
 sg13g2_antennanp ANTENNA_318 (.A(_06792_));
 sg13g2_antennanp ANTENNA_319 (.A(_06793_));
 sg13g2_antennanp ANTENNA_320 (.A(_06807_));
 sg13g2_antennanp ANTENNA_321 (.A(_06817_));
 sg13g2_antennanp ANTENNA_322 (.A(_06817_));
 sg13g2_antennanp ANTENNA_323 (.A(_06821_));
 sg13g2_antennanp ANTENNA_324 (.A(_06838_));
 sg13g2_antennanp ANTENNA_325 (.A(_06853_));
 sg13g2_antennanp ANTENNA_326 (.A(_06874_));
 sg13g2_antennanp ANTENNA_327 (.A(_06875_));
 sg13g2_antennanp ANTENNA_328 (.A(_06895_));
 sg13g2_antennanp ANTENNA_329 (.A(_06902_));
 sg13g2_antennanp ANTENNA_330 (.A(_06908_));
 sg13g2_antennanp ANTENNA_331 (.A(_06945_));
 sg13g2_antennanp ANTENNA_332 (.A(_06963_));
 sg13g2_antennanp ANTENNA_333 (.A(_06980_));
 sg13g2_antennanp ANTENNA_334 (.A(_06980_));
 sg13g2_antennanp ANTENNA_335 (.A(_06980_));
 sg13g2_antennanp ANTENNA_336 (.A(_06981_));
 sg13g2_antennanp ANTENNA_337 (.A(_06985_));
 sg13g2_antennanp ANTENNA_338 (.A(_07020_));
 sg13g2_antennanp ANTENNA_339 (.A(_07032_));
 sg13g2_antennanp ANTENNA_340 (.A(_07063_));
 sg13g2_antennanp ANTENNA_341 (.A(_07064_));
 sg13g2_antennanp ANTENNA_342 (.A(_07073_));
 sg13g2_antennanp ANTENNA_343 (.A(_07074_));
 sg13g2_antennanp ANTENNA_344 (.A(_07077_));
 sg13g2_antennanp ANTENNA_345 (.A(_07085_));
 sg13g2_antennanp ANTENNA_346 (.A(_07104_));
 sg13g2_antennanp ANTENNA_347 (.A(_07113_));
 sg13g2_antennanp ANTENNA_348 (.A(_07125_));
 sg13g2_antennanp ANTENNA_349 (.A(_07129_));
 sg13g2_antennanp ANTENNA_350 (.A(_07150_));
 sg13g2_antennanp ANTENNA_351 (.A(_07151_));
 sg13g2_antennanp ANTENNA_352 (.A(_07157_));
 sg13g2_antennanp ANTENNA_353 (.A(_07172_));
 sg13g2_antennanp ANTENNA_354 (.A(_07188_));
 sg13g2_antennanp ANTENNA_355 (.A(_07195_));
 sg13g2_antennanp ANTENNA_356 (.A(_07201_));
 sg13g2_antennanp ANTENNA_357 (.A(_07221_));
 sg13g2_antennanp ANTENNA_358 (.A(_07222_));
 sg13g2_antennanp ANTENNA_359 (.A(_07243_));
 sg13g2_antennanp ANTENNA_360 (.A(_07269_));
 sg13g2_antennanp ANTENNA_361 (.A(_07279_));
 sg13g2_antennanp ANTENNA_362 (.A(_07282_));
 sg13g2_antennanp ANTENNA_363 (.A(_07344_));
 sg13g2_antennanp ANTENNA_364 (.A(_07345_));
 sg13g2_antennanp ANTENNA_365 (.A(_07369_));
 sg13g2_antennanp ANTENNA_366 (.A(_07371_));
 sg13g2_antennanp ANTENNA_367 (.A(_07381_));
 sg13g2_antennanp ANTENNA_368 (.A(_07385_));
 sg13g2_antennanp ANTENNA_369 (.A(_07421_));
 sg13g2_antennanp ANTENNA_370 (.A(_07429_));
 sg13g2_antennanp ANTENNA_371 (.A(_07435_));
 sg13g2_antennanp ANTENNA_372 (.A(_07440_));
 sg13g2_antennanp ANTENNA_373 (.A(_07446_));
 sg13g2_antennanp ANTENNA_374 (.A(_07480_));
 sg13g2_antennanp ANTENNA_375 (.A(_07485_));
 sg13g2_antennanp ANTENNA_376 (.A(_07507_));
 sg13g2_antennanp ANTENNA_377 (.A(_07535_));
 sg13g2_antennanp ANTENNA_378 (.A(_07540_));
 sg13g2_antennanp ANTENNA_379 (.A(_07544_));
 sg13g2_antennanp ANTENNA_380 (.A(_07552_));
 sg13g2_antennanp ANTENNA_381 (.A(_07560_));
 sg13g2_antennanp ANTENNA_382 (.A(_07577_));
 sg13g2_antennanp ANTENNA_383 (.A(_07577_));
 sg13g2_antennanp ANTENNA_384 (.A(_07577_));
 sg13g2_antennanp ANTENNA_385 (.A(_07592_));
 sg13g2_antennanp ANTENNA_386 (.A(_07595_));
 sg13g2_antennanp ANTENNA_387 (.A(_07601_));
 sg13g2_antennanp ANTENNA_388 (.A(_07601_));
 sg13g2_antennanp ANTENNA_389 (.A(_07601_));
 sg13g2_antennanp ANTENNA_390 (.A(_07603_));
 sg13g2_antennanp ANTENNA_391 (.A(_07634_));
 sg13g2_antennanp ANTENNA_392 (.A(_07913_));
 sg13g2_antennanp ANTENNA_393 (.A(_07945_));
 sg13g2_antennanp ANTENNA_394 (.A(_07979_));
 sg13g2_antennanp ANTENNA_395 (.A(_08062_));
 sg13g2_antennanp ANTENNA_396 (.A(_08219_));
 sg13g2_antennanp ANTENNA_397 (.A(_08219_));
 sg13g2_antennanp ANTENNA_398 (.A(_08219_));
 sg13g2_antennanp ANTENNA_399 (.A(_08219_));
 sg13g2_antennanp ANTENNA_400 (.A(_08219_));
 sg13g2_antennanp ANTENNA_401 (.A(_08219_));
 sg13g2_antennanp ANTENNA_402 (.A(_08219_));
 sg13g2_antennanp ANTENNA_403 (.A(_08219_));
 sg13g2_antennanp ANTENNA_404 (.A(_08219_));
 sg13g2_antennanp ANTENNA_405 (.A(_08219_));
 sg13g2_antennanp ANTENNA_406 (.A(_08219_));
 sg13g2_antennanp ANTENNA_407 (.A(_08219_));
 sg13g2_antennanp ANTENNA_408 (.A(_08219_));
 sg13g2_antennanp ANTENNA_409 (.A(_08219_));
 sg13g2_antennanp ANTENNA_410 (.A(_08219_));
 sg13g2_antennanp ANTENNA_411 (.A(_08219_));
 sg13g2_antennanp ANTENNA_412 (.A(_08221_));
 sg13g2_antennanp ANTENNA_413 (.A(_08221_));
 sg13g2_antennanp ANTENNA_414 (.A(_08221_));
 sg13g2_antennanp ANTENNA_415 (.A(_08223_));
 sg13g2_antennanp ANTENNA_416 (.A(_08223_));
 sg13g2_antennanp ANTENNA_417 (.A(_08223_));
 sg13g2_antennanp ANTENNA_418 (.A(_08223_));
 sg13g2_antennanp ANTENNA_419 (.A(_08223_));
 sg13g2_antennanp ANTENNA_420 (.A(_08223_));
 sg13g2_antennanp ANTENNA_421 (.A(_08227_));
 sg13g2_antennanp ANTENNA_422 (.A(_08227_));
 sg13g2_antennanp ANTENNA_423 (.A(_08260_));
 sg13g2_antennanp ANTENNA_424 (.A(_08260_));
 sg13g2_antennanp ANTENNA_425 (.A(_08260_));
 sg13g2_antennanp ANTENNA_426 (.A(_08260_));
 sg13g2_antennanp ANTENNA_427 (.A(_08260_));
 sg13g2_antennanp ANTENNA_428 (.A(_08260_));
 sg13g2_antennanp ANTENNA_429 (.A(_08260_));
 sg13g2_antennanp ANTENNA_430 (.A(_08260_));
 sg13g2_antennanp ANTENNA_431 (.A(_08260_));
 sg13g2_antennanp ANTENNA_432 (.A(_08260_));
 sg13g2_antennanp ANTENNA_433 (.A(_08261_));
 sg13g2_antennanp ANTENNA_434 (.A(_08261_));
 sg13g2_antennanp ANTENNA_435 (.A(_08263_));
 sg13g2_antennanp ANTENNA_436 (.A(_08263_));
 sg13g2_antennanp ANTENNA_437 (.A(_08263_));
 sg13g2_antennanp ANTENNA_438 (.A(_08263_));
 sg13g2_antennanp ANTENNA_439 (.A(_08263_));
 sg13g2_antennanp ANTENNA_440 (.A(_08263_));
 sg13g2_antennanp ANTENNA_441 (.A(_08263_));
 sg13g2_antennanp ANTENNA_442 (.A(_08263_));
 sg13g2_antennanp ANTENNA_443 (.A(_08263_));
 sg13g2_antennanp ANTENNA_444 (.A(_08263_));
 sg13g2_antennanp ANTENNA_445 (.A(_08321_));
 sg13g2_antennanp ANTENNA_446 (.A(_08321_));
 sg13g2_antennanp ANTENNA_447 (.A(_08321_));
 sg13g2_antennanp ANTENNA_448 (.A(_08321_));
 sg13g2_antennanp ANTENNA_449 (.A(_08321_));
 sg13g2_antennanp ANTENNA_450 (.A(_08321_));
 sg13g2_antennanp ANTENNA_451 (.A(_08321_));
 sg13g2_antennanp ANTENNA_452 (.A(_08321_));
 sg13g2_antennanp ANTENNA_453 (.A(_08321_));
 sg13g2_antennanp ANTENNA_454 (.A(_08321_));
 sg13g2_antennanp ANTENNA_455 (.A(_08321_));
 sg13g2_antennanp ANTENNA_456 (.A(_08321_));
 sg13g2_antennanp ANTENNA_457 (.A(_08321_));
 sg13g2_antennanp ANTENNA_458 (.A(_08321_));
 sg13g2_antennanp ANTENNA_459 (.A(_08321_));
 sg13g2_antennanp ANTENNA_460 (.A(_08321_));
 sg13g2_antennanp ANTENNA_461 (.A(_08321_));
 sg13g2_antennanp ANTENNA_462 (.A(_08321_));
 sg13g2_antennanp ANTENNA_463 (.A(_08321_));
 sg13g2_antennanp ANTENNA_464 (.A(_08321_));
 sg13g2_antennanp ANTENNA_465 (.A(_08321_));
 sg13g2_antennanp ANTENNA_466 (.A(_08321_));
 sg13g2_antennanp ANTENNA_467 (.A(_08321_));
 sg13g2_antennanp ANTENNA_468 (.A(_08321_));
 sg13g2_antennanp ANTENNA_469 (.A(_08338_));
 sg13g2_antennanp ANTENNA_470 (.A(_08338_));
 sg13g2_antennanp ANTENNA_471 (.A(_08338_));
 sg13g2_antennanp ANTENNA_472 (.A(_08345_));
 sg13g2_antennanp ANTENNA_473 (.A(_08345_));
 sg13g2_antennanp ANTENNA_474 (.A(_08345_));
 sg13g2_antennanp ANTENNA_475 (.A(_08345_));
 sg13g2_antennanp ANTENNA_476 (.A(_08345_));
 sg13g2_antennanp ANTENNA_477 (.A(_08345_));
 sg13g2_antennanp ANTENNA_478 (.A(_08345_));
 sg13g2_antennanp ANTENNA_479 (.A(_08345_));
 sg13g2_antennanp ANTENNA_480 (.A(_08345_));
 sg13g2_antennanp ANTENNA_481 (.A(_08345_));
 sg13g2_antennanp ANTENNA_482 (.A(_08345_));
 sg13g2_antennanp ANTENNA_483 (.A(_08345_));
 sg13g2_antennanp ANTENNA_484 (.A(_08345_));
 sg13g2_antennanp ANTENNA_485 (.A(_08345_));
 sg13g2_antennanp ANTENNA_486 (.A(_08345_));
 sg13g2_antennanp ANTENNA_487 (.A(_08345_));
 sg13g2_antennanp ANTENNA_488 (.A(_08345_));
 sg13g2_antennanp ANTENNA_489 (.A(_08345_));
 sg13g2_antennanp ANTENNA_490 (.A(_08345_));
 sg13g2_antennanp ANTENNA_491 (.A(_08345_));
 sg13g2_antennanp ANTENNA_492 (.A(_08345_));
 sg13g2_antennanp ANTENNA_493 (.A(_08345_));
 sg13g2_antennanp ANTENNA_494 (.A(_08354_));
 sg13g2_antennanp ANTENNA_495 (.A(_08354_));
 sg13g2_antennanp ANTENNA_496 (.A(_08354_));
 sg13g2_antennanp ANTENNA_497 (.A(_08354_));
 sg13g2_antennanp ANTENNA_498 (.A(_08354_));
 sg13g2_antennanp ANTENNA_499 (.A(_08354_));
 sg13g2_antennanp ANTENNA_500 (.A(_08354_));
 sg13g2_antennanp ANTENNA_501 (.A(_08380_));
 sg13g2_antennanp ANTENNA_502 (.A(_08380_));
 sg13g2_antennanp ANTENNA_503 (.A(_08706_));
 sg13g2_antennanp ANTENNA_504 (.A(_08730_));
 sg13g2_antennanp ANTENNA_505 (.A(_08730_));
 sg13g2_antennanp ANTENNA_506 (.A(_08985_));
 sg13g2_antennanp ANTENNA_507 (.A(_08985_));
 sg13g2_antennanp ANTENNA_508 (.A(_08985_));
 sg13g2_antennanp ANTENNA_509 (.A(_08985_));
 sg13g2_antennanp ANTENNA_510 (.A(_08993_));
 sg13g2_antennanp ANTENNA_511 (.A(_08993_));
 sg13g2_antennanp ANTENNA_512 (.A(_08993_));
 sg13g2_antennanp ANTENNA_513 (.A(_08997_));
 sg13g2_antennanp ANTENNA_514 (.A(_08997_));
 sg13g2_antennanp ANTENNA_515 (.A(_08997_));
 sg13g2_antennanp ANTENNA_516 (.A(_08997_));
 sg13g2_antennanp ANTENNA_517 (.A(_09940_));
 sg13g2_antennanp ANTENNA_518 (.A(_10089_));
 sg13g2_antennanp ANTENNA_519 (.A(_10089_));
 sg13g2_antennanp ANTENNA_520 (.A(_10089_));
 sg13g2_antennanp ANTENNA_521 (.A(_10158_));
 sg13g2_antennanp ANTENNA_522 (.A(_10158_));
 sg13g2_antennanp ANTENNA_523 (.A(_10158_));
 sg13g2_antennanp ANTENNA_524 (.A(_10158_));
 sg13g2_antennanp ANTENNA_525 (.A(_10159_));
 sg13g2_antennanp ANTENNA_526 (.A(_10159_));
 sg13g2_antennanp ANTENNA_527 (.A(_10159_));
 sg13g2_antennanp ANTENNA_528 (.A(_10204_));
 sg13g2_antennanp ANTENNA_529 (.A(_10224_));
 sg13g2_antennanp ANTENNA_530 (.A(_10224_));
 sg13g2_antennanp ANTENNA_531 (.A(_10224_));
 sg13g2_antennanp ANTENNA_532 (.A(_10224_));
 sg13g2_antennanp ANTENNA_533 (.A(_10224_));
 sg13g2_antennanp ANTENNA_534 (.A(_10224_));
 sg13g2_antennanp ANTENNA_535 (.A(_10224_));
 sg13g2_antennanp ANTENNA_536 (.A(_10224_));
 sg13g2_antennanp ANTENNA_537 (.A(_10318_));
 sg13g2_antennanp ANTENNA_538 (.A(_10318_));
 sg13g2_antennanp ANTENNA_539 (.A(_10318_));
 sg13g2_antennanp ANTENNA_540 (.A(_10342_));
 sg13g2_antennanp ANTENNA_541 (.A(_10342_));
 sg13g2_antennanp ANTENNA_542 (.A(_10361_));
 sg13g2_antennanp ANTENNA_543 (.A(_10361_));
 sg13g2_antennanp ANTENNA_544 (.A(_10361_));
 sg13g2_antennanp ANTENNA_545 (.A(_10361_));
 sg13g2_antennanp ANTENNA_546 (.A(_10424_));
 sg13g2_antennanp ANTENNA_547 (.A(_10424_));
 sg13g2_antennanp ANTENNA_548 (.A(_10424_));
 sg13g2_antennanp ANTENNA_549 (.A(_10424_));
 sg13g2_antennanp ANTENNA_550 (.A(_10424_));
 sg13g2_antennanp ANTENNA_551 (.A(_10424_));
 sg13g2_antennanp ANTENNA_552 (.A(_10424_));
 sg13g2_antennanp ANTENNA_553 (.A(_10429_));
 sg13g2_antennanp ANTENNA_554 (.A(_10429_));
 sg13g2_antennanp ANTENNA_555 (.A(_10429_));
 sg13g2_antennanp ANTENNA_556 (.A(_10429_));
 sg13g2_antennanp ANTENNA_557 (.A(_10429_));
 sg13g2_antennanp ANTENNA_558 (.A(_10429_));
 sg13g2_antennanp ANTENNA_559 (.A(_10535_));
 sg13g2_antennanp ANTENNA_560 (.A(_10535_));
 sg13g2_antennanp ANTENNA_561 (.A(_10535_));
 sg13g2_antennanp ANTENNA_562 (.A(_10535_));
 sg13g2_antennanp ANTENNA_563 (.A(_10535_));
 sg13g2_antennanp ANTENNA_564 (.A(_10535_));
 sg13g2_antennanp ANTENNA_565 (.A(_10535_));
 sg13g2_antennanp ANTENNA_566 (.A(_10599_));
 sg13g2_antennanp ANTENNA_567 (.A(_10599_));
 sg13g2_antennanp ANTENNA_568 (.A(_10599_));
 sg13g2_antennanp ANTENNA_569 (.A(_10599_));
 sg13g2_antennanp ANTENNA_570 (.A(_10599_));
 sg13g2_antennanp ANTENNA_571 (.A(_10599_));
 sg13g2_antennanp ANTENNA_572 (.A(_10600_));
 sg13g2_antennanp ANTENNA_573 (.A(_10600_));
 sg13g2_antennanp ANTENNA_574 (.A(_10600_));
 sg13g2_antennanp ANTENNA_575 (.A(_10600_));
 sg13g2_antennanp ANTENNA_576 (.A(_10600_));
 sg13g2_antennanp ANTENNA_577 (.A(_10600_));
 sg13g2_antennanp ANTENNA_578 (.A(_10662_));
 sg13g2_antennanp ANTENNA_579 (.A(_10662_));
 sg13g2_antennanp ANTENNA_580 (.A(_10662_));
 sg13g2_antennanp ANTENNA_581 (.A(_10662_));
 sg13g2_antennanp ANTENNA_582 (.A(_10662_));
 sg13g2_antennanp ANTENNA_583 (.A(_10662_));
 sg13g2_antennanp ANTENNA_584 (.A(_10662_));
 sg13g2_antennanp ANTENNA_585 (.A(_10662_));
 sg13g2_antennanp ANTENNA_586 (.A(_10662_));
 sg13g2_antennanp ANTENNA_587 (.A(_10662_));
 sg13g2_antennanp ANTENNA_588 (.A(_10696_));
 sg13g2_antennanp ANTENNA_589 (.A(_10696_));
 sg13g2_antennanp ANTENNA_590 (.A(_10696_));
 sg13g2_antennanp ANTENNA_591 (.A(_10704_));
 sg13g2_antennanp ANTENNA_592 (.A(_10704_));
 sg13g2_antennanp ANTENNA_593 (.A(_10704_));
 sg13g2_antennanp ANTENNA_594 (.A(_10704_));
 sg13g2_antennanp ANTENNA_595 (.A(_10704_));
 sg13g2_antennanp ANTENNA_596 (.A(_10704_));
 sg13g2_antennanp ANTENNA_597 (.A(_10739_));
 sg13g2_antennanp ANTENNA_598 (.A(_10739_));
 sg13g2_antennanp ANTENNA_599 (.A(_10739_));
 sg13g2_antennanp ANTENNA_600 (.A(_10739_));
 sg13g2_antennanp ANTENNA_601 (.A(_10739_));
 sg13g2_antennanp ANTENNA_602 (.A(_10739_));
 sg13g2_antennanp ANTENNA_603 (.A(_10741_));
 sg13g2_antennanp ANTENNA_604 (.A(_10741_));
 sg13g2_antennanp ANTENNA_605 (.A(_10741_));
 sg13g2_antennanp ANTENNA_606 (.A(_10741_));
 sg13g2_antennanp ANTENNA_607 (.A(_10741_));
 sg13g2_antennanp ANTENNA_608 (.A(_10741_));
 sg13g2_antennanp ANTENNA_609 (.A(_10741_));
 sg13g2_antennanp ANTENNA_610 (.A(_10741_));
 sg13g2_antennanp ANTENNA_611 (.A(_10741_));
 sg13g2_antennanp ANTENNA_612 (.A(_10741_));
 sg13g2_antennanp ANTENNA_613 (.A(_10742_));
 sg13g2_antennanp ANTENNA_614 (.A(_10742_));
 sg13g2_antennanp ANTENNA_615 (.A(_10742_));
 sg13g2_antennanp ANTENNA_616 (.A(_10742_));
 sg13g2_antennanp ANTENNA_617 (.A(_10742_));
 sg13g2_antennanp ANTENNA_618 (.A(_10742_));
 sg13g2_antennanp ANTENNA_619 (.A(_10742_));
 sg13g2_antennanp ANTENNA_620 (.A(_10742_));
 sg13g2_antennanp ANTENNA_621 (.A(_10742_));
 sg13g2_antennanp ANTENNA_622 (.A(_10745_));
 sg13g2_antennanp ANTENNA_623 (.A(_10745_));
 sg13g2_antennanp ANTENNA_624 (.A(_10745_));
 sg13g2_antennanp ANTENNA_625 (.A(_10745_));
 sg13g2_antennanp ANTENNA_626 (.A(_10745_));
 sg13g2_antennanp ANTENNA_627 (.A(_10745_));
 sg13g2_antennanp ANTENNA_628 (.A(_10745_));
 sg13g2_antennanp ANTENNA_629 (.A(_10745_));
 sg13g2_antennanp ANTENNA_630 (.A(_10745_));
 sg13g2_antennanp ANTENNA_631 (.A(_10779_));
 sg13g2_antennanp ANTENNA_632 (.A(_10779_));
 sg13g2_antennanp ANTENNA_633 (.A(_10779_));
 sg13g2_antennanp ANTENNA_634 (.A(_10779_));
 sg13g2_antennanp ANTENNA_635 (.A(_10779_));
 sg13g2_antennanp ANTENNA_636 (.A(_10779_));
 sg13g2_antennanp ANTENNA_637 (.A(_10797_));
 sg13g2_antennanp ANTENNA_638 (.A(_10797_));
 sg13g2_antennanp ANTENNA_639 (.A(_10797_));
 sg13g2_antennanp ANTENNA_640 (.A(_10797_));
 sg13g2_antennanp ANTENNA_641 (.A(_10804_));
 sg13g2_antennanp ANTENNA_642 (.A(_10804_));
 sg13g2_antennanp ANTENNA_643 (.A(_10804_));
 sg13g2_antennanp ANTENNA_644 (.A(_10810_));
 sg13g2_antennanp ANTENNA_645 (.A(_10810_));
 sg13g2_antennanp ANTENNA_646 (.A(_10810_));
 sg13g2_antennanp ANTENNA_647 (.A(_10810_));
 sg13g2_antennanp ANTENNA_648 (.A(_10810_));
 sg13g2_antennanp ANTENNA_649 (.A(_10810_));
 sg13g2_antennanp ANTENNA_650 (.A(_10810_));
 sg13g2_antennanp ANTENNA_651 (.A(_10810_));
 sg13g2_antennanp ANTENNA_652 (.A(_10810_));
 sg13g2_antennanp ANTENNA_653 (.A(_10810_));
 sg13g2_antennanp ANTENNA_654 (.A(_10812_));
 sg13g2_antennanp ANTENNA_655 (.A(_10812_));
 sg13g2_antennanp ANTENNA_656 (.A(_10812_));
 sg13g2_antennanp ANTENNA_657 (.A(_10812_));
 sg13g2_antennanp ANTENNA_658 (.A(_10812_));
 sg13g2_antennanp ANTENNA_659 (.A(_10812_));
 sg13g2_antennanp ANTENNA_660 (.A(_10812_));
 sg13g2_antennanp ANTENNA_661 (.A(_10812_));
 sg13g2_antennanp ANTENNA_662 (.A(_10812_));
 sg13g2_antennanp ANTENNA_663 (.A(_10812_));
 sg13g2_antennanp ANTENNA_664 (.A(_10818_));
 sg13g2_antennanp ANTENNA_665 (.A(_10818_));
 sg13g2_antennanp ANTENNA_666 (.A(_10818_));
 sg13g2_antennanp ANTENNA_667 (.A(_10818_));
 sg13g2_antennanp ANTENNA_668 (.A(_10818_));
 sg13g2_antennanp ANTENNA_669 (.A(_10818_));
 sg13g2_antennanp ANTENNA_670 (.A(_10818_));
 sg13g2_antennanp ANTENNA_671 (.A(_10818_));
 sg13g2_antennanp ANTENNA_672 (.A(_10818_));
 sg13g2_antennanp ANTENNA_673 (.A(_10818_));
 sg13g2_antennanp ANTENNA_674 (.A(_10845_));
 sg13g2_antennanp ANTENNA_675 (.A(_10845_));
 sg13g2_antennanp ANTENNA_676 (.A(_10845_));
 sg13g2_antennanp ANTENNA_677 (.A(_10845_));
 sg13g2_antennanp ANTENNA_678 (.A(_10845_));
 sg13g2_antennanp ANTENNA_679 (.A(_10845_));
 sg13g2_antennanp ANTENNA_680 (.A(_10845_));
 sg13g2_antennanp ANTENNA_681 (.A(_10845_));
 sg13g2_antennanp ANTENNA_682 (.A(_10845_));
 sg13g2_antennanp ANTENNA_683 (.A(_10845_));
 sg13g2_antennanp ANTENNA_684 (.A(_10974_));
 sg13g2_antennanp ANTENNA_685 (.A(_10974_));
 sg13g2_antennanp ANTENNA_686 (.A(_10974_));
 sg13g2_antennanp ANTENNA_687 (.A(_10974_));
 sg13g2_antennanp ANTENNA_688 (.A(_10974_));
 sg13g2_antennanp ANTENNA_689 (.A(_10974_));
 sg13g2_antennanp ANTENNA_690 (.A(_10974_));
 sg13g2_antennanp ANTENNA_691 (.A(_10974_));
 sg13g2_antennanp ANTENNA_692 (.A(_10974_));
 sg13g2_antennanp ANTENNA_693 (.A(_10974_));
 sg13g2_antennanp ANTENNA_694 (.A(_11107_));
 sg13g2_antennanp ANTENNA_695 (.A(_11107_));
 sg13g2_antennanp ANTENNA_696 (.A(_11107_));
 sg13g2_antennanp ANTENNA_697 (.A(_11107_));
 sg13g2_antennanp ANTENNA_698 (.A(_11147_));
 sg13g2_antennanp ANTENNA_699 (.A(_11147_));
 sg13g2_antennanp ANTENNA_700 (.A(_11147_));
 sg13g2_antennanp ANTENNA_701 (.A(_11147_));
 sg13g2_antennanp ANTENNA_702 (.A(clk));
 sg13g2_antennanp ANTENNA_703 (.A(clk));
 sg13g2_antennanp ANTENNA_704 (.A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_antennanp ANTENNA_705 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_706 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_707 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_708 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_709 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_710 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_711 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_712 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_713 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_714 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_715 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_716 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_717 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_718 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_719 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_720 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_721 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_722 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_723 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_724 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_725 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_726 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_727 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_728 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_729 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_730 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_731 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_732 (.A(\top_ihp.oisc.regs[32][31] ));
 sg13g2_antennanp ANTENNA_733 (.A(\top_ihp.oisc.regs[32][31] ));
 sg13g2_antennanp ANTENNA_734 (.A(\top_ihp.oisc.regs[32][31] ));
 sg13g2_antennanp ANTENNA_735 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_736 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_737 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_738 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_739 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_740 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_741 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_742 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_743 (.A(\top_ihp.oisc.regs[50][16] ));
 sg13g2_antennanp ANTENNA_744 (.A(\top_ihp.oisc.regs[50][16] ));
 sg13g2_antennanp ANTENNA_745 (.A(\top_ihp.oisc.regs[50][16] ));
 sg13g2_antennanp ANTENNA_746 (.A(\top_ihp.oisc.regs[59][2] ));
 sg13g2_antennanp ANTENNA_747 (.A(\top_ihp.oisc.regs[59][2] ));
 sg13g2_antennanp ANTENNA_748 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_749 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_750 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_751 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_752 (.A(net54));
 sg13g2_antennanp ANTENNA_753 (.A(net54));
 sg13g2_antennanp ANTENNA_754 (.A(net54));
 sg13g2_antennanp ANTENNA_755 (.A(net54));
 sg13g2_antennanp ANTENNA_756 (.A(net54));
 sg13g2_antennanp ANTENNA_757 (.A(net54));
 sg13g2_antennanp ANTENNA_758 (.A(net54));
 sg13g2_antennanp ANTENNA_759 (.A(net54));
 sg13g2_antennanp ANTENNA_760 (.A(net54));
 sg13g2_antennanp ANTENNA_761 (.A(net56));
 sg13g2_antennanp ANTENNA_762 (.A(net56));
 sg13g2_antennanp ANTENNA_763 (.A(net56));
 sg13g2_antennanp ANTENNA_764 (.A(net56));
 sg13g2_antennanp ANTENNA_765 (.A(net56));
 sg13g2_antennanp ANTENNA_766 (.A(net56));
 sg13g2_antennanp ANTENNA_767 (.A(net56));
 sg13g2_antennanp ANTENNA_768 (.A(net56));
 sg13g2_antennanp ANTENNA_769 (.A(net56));
 sg13g2_antennanp ANTENNA_770 (.A(net90));
 sg13g2_antennanp ANTENNA_771 (.A(net90));
 sg13g2_antennanp ANTENNA_772 (.A(net90));
 sg13g2_antennanp ANTENNA_773 (.A(net90));
 sg13g2_antennanp ANTENNA_774 (.A(net90));
 sg13g2_antennanp ANTENNA_775 (.A(net90));
 sg13g2_antennanp ANTENNA_776 (.A(net90));
 sg13g2_antennanp ANTENNA_777 (.A(net90));
 sg13g2_antennanp ANTENNA_778 (.A(net117));
 sg13g2_antennanp ANTENNA_779 (.A(net117));
 sg13g2_antennanp ANTENNA_780 (.A(net117));
 sg13g2_antennanp ANTENNA_781 (.A(net117));
 sg13g2_antennanp ANTENNA_782 (.A(net117));
 sg13g2_antennanp ANTENNA_783 (.A(net117));
 sg13g2_antennanp ANTENNA_784 (.A(net117));
 sg13g2_antennanp ANTENNA_785 (.A(net117));
 sg13g2_antennanp ANTENNA_786 (.A(net117));
 sg13g2_antennanp ANTENNA_787 (.A(net117));
 sg13g2_antennanp ANTENNA_788 (.A(net117));
 sg13g2_antennanp ANTENNA_789 (.A(net117));
 sg13g2_antennanp ANTENNA_790 (.A(net117));
 sg13g2_antennanp ANTENNA_791 (.A(net117));
 sg13g2_antennanp ANTENNA_792 (.A(net117));
 sg13g2_antennanp ANTENNA_793 (.A(net117));
 sg13g2_antennanp ANTENNA_794 (.A(net117));
 sg13g2_antennanp ANTENNA_795 (.A(net117));
 sg13g2_antennanp ANTENNA_796 (.A(net117));
 sg13g2_antennanp ANTENNA_797 (.A(net117));
 sg13g2_antennanp ANTENNA_798 (.A(net118));
 sg13g2_antennanp ANTENNA_799 (.A(net118));
 sg13g2_antennanp ANTENNA_800 (.A(net118));
 sg13g2_antennanp ANTENNA_801 (.A(net118));
 sg13g2_antennanp ANTENNA_802 (.A(net118));
 sg13g2_antennanp ANTENNA_803 (.A(net118));
 sg13g2_antennanp ANTENNA_804 (.A(net118));
 sg13g2_antennanp ANTENNA_805 (.A(net118));
 sg13g2_antennanp ANTENNA_806 (.A(net118));
 sg13g2_antennanp ANTENNA_807 (.A(net121));
 sg13g2_antennanp ANTENNA_808 (.A(net121));
 sg13g2_antennanp ANTENNA_809 (.A(net121));
 sg13g2_antennanp ANTENNA_810 (.A(net121));
 sg13g2_antennanp ANTENNA_811 (.A(net121));
 sg13g2_antennanp ANTENNA_812 (.A(net121));
 sg13g2_antennanp ANTENNA_813 (.A(net121));
 sg13g2_antennanp ANTENNA_814 (.A(net121));
 sg13g2_antennanp ANTENNA_815 (.A(net121));
 sg13g2_antennanp ANTENNA_816 (.A(net121));
 sg13g2_antennanp ANTENNA_817 (.A(net121));
 sg13g2_antennanp ANTENNA_818 (.A(net121));
 sg13g2_antennanp ANTENNA_819 (.A(net121));
 sg13g2_antennanp ANTENNA_820 (.A(net123));
 sg13g2_antennanp ANTENNA_821 (.A(net123));
 sg13g2_antennanp ANTENNA_822 (.A(net123));
 sg13g2_antennanp ANTENNA_823 (.A(net123));
 sg13g2_antennanp ANTENNA_824 (.A(net123));
 sg13g2_antennanp ANTENNA_825 (.A(net123));
 sg13g2_antennanp ANTENNA_826 (.A(net123));
 sg13g2_antennanp ANTENNA_827 (.A(net123));
 sg13g2_antennanp ANTENNA_828 (.A(net123));
 sg13g2_antennanp ANTENNA_829 (.A(net123));
 sg13g2_antennanp ANTENNA_830 (.A(net123));
 sg13g2_antennanp ANTENNA_831 (.A(net123));
 sg13g2_antennanp ANTENNA_832 (.A(net123));
 sg13g2_antennanp ANTENNA_833 (.A(net123));
 sg13g2_antennanp ANTENNA_834 (.A(net124));
 sg13g2_antennanp ANTENNA_835 (.A(net124));
 sg13g2_antennanp ANTENNA_836 (.A(net124));
 sg13g2_antennanp ANTENNA_837 (.A(net124));
 sg13g2_antennanp ANTENNA_838 (.A(net124));
 sg13g2_antennanp ANTENNA_839 (.A(net124));
 sg13g2_antennanp ANTENNA_840 (.A(net124));
 sg13g2_antennanp ANTENNA_841 (.A(net124));
 sg13g2_antennanp ANTENNA_842 (.A(net124));
 sg13g2_antennanp ANTENNA_843 (.A(net126));
 sg13g2_antennanp ANTENNA_844 (.A(net126));
 sg13g2_antennanp ANTENNA_845 (.A(net126));
 sg13g2_antennanp ANTENNA_846 (.A(net126));
 sg13g2_antennanp ANTENNA_847 (.A(net126));
 sg13g2_antennanp ANTENNA_848 (.A(net126));
 sg13g2_antennanp ANTENNA_849 (.A(net126));
 sg13g2_antennanp ANTENNA_850 (.A(net126));
 sg13g2_antennanp ANTENNA_851 (.A(net127));
 sg13g2_antennanp ANTENNA_852 (.A(net127));
 sg13g2_antennanp ANTENNA_853 (.A(net127));
 sg13g2_antennanp ANTENNA_854 (.A(net127));
 sg13g2_antennanp ANTENNA_855 (.A(net127));
 sg13g2_antennanp ANTENNA_856 (.A(net127));
 sg13g2_antennanp ANTENNA_857 (.A(net127));
 sg13g2_antennanp ANTENNA_858 (.A(net127));
 sg13g2_antennanp ANTENNA_859 (.A(net127));
 sg13g2_antennanp ANTENNA_860 (.A(net127));
 sg13g2_antennanp ANTENNA_861 (.A(net127));
 sg13g2_antennanp ANTENNA_862 (.A(net127));
 sg13g2_antennanp ANTENNA_863 (.A(net127));
 sg13g2_antennanp ANTENNA_864 (.A(net127));
 sg13g2_antennanp ANTENNA_865 (.A(net127));
 sg13g2_antennanp ANTENNA_866 (.A(net127));
 sg13g2_antennanp ANTENNA_867 (.A(net127));
 sg13g2_antennanp ANTENNA_868 (.A(net127));
 sg13g2_antennanp ANTENNA_869 (.A(net127));
 sg13g2_antennanp ANTENNA_870 (.A(net127));
 sg13g2_antennanp ANTENNA_871 (.A(net127));
 sg13g2_antennanp ANTENNA_872 (.A(net127));
 sg13g2_antennanp ANTENNA_873 (.A(net127));
 sg13g2_antennanp ANTENNA_874 (.A(net127));
 sg13g2_antennanp ANTENNA_875 (.A(net127));
 sg13g2_antennanp ANTENNA_876 (.A(net127));
 sg13g2_antennanp ANTENNA_877 (.A(net127));
 sg13g2_antennanp ANTENNA_878 (.A(net127));
 sg13g2_antennanp ANTENNA_879 (.A(net130));
 sg13g2_antennanp ANTENNA_880 (.A(net130));
 sg13g2_antennanp ANTENNA_881 (.A(net130));
 sg13g2_antennanp ANTENNA_882 (.A(net130));
 sg13g2_antennanp ANTENNA_883 (.A(net130));
 sg13g2_antennanp ANTENNA_884 (.A(net130));
 sg13g2_antennanp ANTENNA_885 (.A(net130));
 sg13g2_antennanp ANTENNA_886 (.A(net130));
 sg13g2_antennanp ANTENNA_887 (.A(net132));
 sg13g2_antennanp ANTENNA_888 (.A(net132));
 sg13g2_antennanp ANTENNA_889 (.A(net132));
 sg13g2_antennanp ANTENNA_890 (.A(net132));
 sg13g2_antennanp ANTENNA_891 (.A(net132));
 sg13g2_antennanp ANTENNA_892 (.A(net132));
 sg13g2_antennanp ANTENNA_893 (.A(net132));
 sg13g2_antennanp ANTENNA_894 (.A(net132));
 sg13g2_antennanp ANTENNA_895 (.A(net132));
 sg13g2_antennanp ANTENNA_896 (.A(net134));
 sg13g2_antennanp ANTENNA_897 (.A(net134));
 sg13g2_antennanp ANTENNA_898 (.A(net134));
 sg13g2_antennanp ANTENNA_899 (.A(net134));
 sg13g2_antennanp ANTENNA_900 (.A(net134));
 sg13g2_antennanp ANTENNA_901 (.A(net134));
 sg13g2_antennanp ANTENNA_902 (.A(net134));
 sg13g2_antennanp ANTENNA_903 (.A(net134));
 sg13g2_antennanp ANTENNA_904 (.A(net134));
 sg13g2_antennanp ANTENNA_905 (.A(net134));
 sg13g2_antennanp ANTENNA_906 (.A(net134));
 sg13g2_antennanp ANTENNA_907 (.A(net134));
 sg13g2_antennanp ANTENNA_908 (.A(net134));
 sg13g2_antennanp ANTENNA_909 (.A(net134));
 sg13g2_antennanp ANTENNA_910 (.A(net134));
 sg13g2_antennanp ANTENNA_911 (.A(net134));
 sg13g2_antennanp ANTENNA_912 (.A(net134));
 sg13g2_antennanp ANTENNA_913 (.A(net134));
 sg13g2_antennanp ANTENNA_914 (.A(net134));
 sg13g2_antennanp ANTENNA_915 (.A(net134));
 sg13g2_antennanp ANTENNA_916 (.A(net134));
 sg13g2_antennanp ANTENNA_917 (.A(net134));
 sg13g2_antennanp ANTENNA_918 (.A(net134));
 sg13g2_antennanp ANTENNA_919 (.A(net134));
 sg13g2_antennanp ANTENNA_920 (.A(net134));
 sg13g2_antennanp ANTENNA_921 (.A(net134));
 sg13g2_antennanp ANTENNA_922 (.A(net134));
 sg13g2_antennanp ANTENNA_923 (.A(net134));
 sg13g2_antennanp ANTENNA_924 (.A(net134));
 sg13g2_antennanp ANTENNA_925 (.A(net134));
 sg13g2_antennanp ANTENNA_926 (.A(net134));
 sg13g2_antennanp ANTENNA_927 (.A(net134));
 sg13g2_antennanp ANTENNA_928 (.A(net134));
 sg13g2_antennanp ANTENNA_929 (.A(net134));
 sg13g2_antennanp ANTENNA_930 (.A(net143));
 sg13g2_antennanp ANTENNA_931 (.A(net143));
 sg13g2_antennanp ANTENNA_932 (.A(net143));
 sg13g2_antennanp ANTENNA_933 (.A(net143));
 sg13g2_antennanp ANTENNA_934 (.A(net143));
 sg13g2_antennanp ANTENNA_935 (.A(net143));
 sg13g2_antennanp ANTENNA_936 (.A(net143));
 sg13g2_antennanp ANTENNA_937 (.A(net143));
 sg13g2_antennanp ANTENNA_938 (.A(net143));
 sg13g2_antennanp ANTENNA_939 (.A(net159));
 sg13g2_antennanp ANTENNA_940 (.A(net159));
 sg13g2_antennanp ANTENNA_941 (.A(net159));
 sg13g2_antennanp ANTENNA_942 (.A(net159));
 sg13g2_antennanp ANTENNA_943 (.A(net159));
 sg13g2_antennanp ANTENNA_944 (.A(net159));
 sg13g2_antennanp ANTENNA_945 (.A(net159));
 sg13g2_antennanp ANTENNA_946 (.A(net159));
 sg13g2_antennanp ANTENNA_947 (.A(net159));
 sg13g2_antennanp ANTENNA_948 (.A(net173));
 sg13g2_antennanp ANTENNA_949 (.A(net173));
 sg13g2_antennanp ANTENNA_950 (.A(net173));
 sg13g2_antennanp ANTENNA_951 (.A(net173));
 sg13g2_antennanp ANTENNA_952 (.A(net173));
 sg13g2_antennanp ANTENNA_953 (.A(net173));
 sg13g2_antennanp ANTENNA_954 (.A(net173));
 sg13g2_antennanp ANTENNA_955 (.A(net173));
 sg13g2_antennanp ANTENNA_956 (.A(net177));
 sg13g2_antennanp ANTENNA_957 (.A(net177));
 sg13g2_antennanp ANTENNA_958 (.A(net177));
 sg13g2_antennanp ANTENNA_959 (.A(net177));
 sg13g2_antennanp ANTENNA_960 (.A(net177));
 sg13g2_antennanp ANTENNA_961 (.A(net177));
 sg13g2_antennanp ANTENNA_962 (.A(net177));
 sg13g2_antennanp ANTENNA_963 (.A(net177));
 sg13g2_antennanp ANTENNA_964 (.A(net177));
 sg13g2_antennanp ANTENNA_965 (.A(net177));
 sg13g2_antennanp ANTENNA_966 (.A(net177));
 sg13g2_antennanp ANTENNA_967 (.A(net188));
 sg13g2_antennanp ANTENNA_968 (.A(net188));
 sg13g2_antennanp ANTENNA_969 (.A(net188));
 sg13g2_antennanp ANTENNA_970 (.A(net188));
 sg13g2_antennanp ANTENNA_971 (.A(net188));
 sg13g2_antennanp ANTENNA_972 (.A(net188));
 sg13g2_antennanp ANTENNA_973 (.A(net188));
 sg13g2_antennanp ANTENNA_974 (.A(net188));
 sg13g2_antennanp ANTENNA_975 (.A(net231));
 sg13g2_antennanp ANTENNA_976 (.A(net231));
 sg13g2_antennanp ANTENNA_977 (.A(net231));
 sg13g2_antennanp ANTENNA_978 (.A(net231));
 sg13g2_antennanp ANTENNA_979 (.A(net231));
 sg13g2_antennanp ANTENNA_980 (.A(net231));
 sg13g2_antennanp ANTENNA_981 (.A(net231));
 sg13g2_antennanp ANTENNA_982 (.A(net231));
 sg13g2_antennanp ANTENNA_983 (.A(net231));
 sg13g2_antennanp ANTENNA_984 (.A(net255));
 sg13g2_antennanp ANTENNA_985 (.A(net255));
 sg13g2_antennanp ANTENNA_986 (.A(net255));
 sg13g2_antennanp ANTENNA_987 (.A(net255));
 sg13g2_antennanp ANTENNA_988 (.A(net255));
 sg13g2_antennanp ANTENNA_989 (.A(net255));
 sg13g2_antennanp ANTENNA_990 (.A(net255));
 sg13g2_antennanp ANTENNA_991 (.A(net255));
 sg13g2_antennanp ANTENNA_992 (.A(net255));
 sg13g2_antennanp ANTENNA_993 (.A(net255));
 sg13g2_antennanp ANTENNA_994 (.A(net255));
 sg13g2_antennanp ANTENNA_995 (.A(net263));
 sg13g2_antennanp ANTENNA_996 (.A(net263));
 sg13g2_antennanp ANTENNA_997 (.A(net263));
 sg13g2_antennanp ANTENNA_998 (.A(net263));
 sg13g2_antennanp ANTENNA_999 (.A(net263));
 sg13g2_antennanp ANTENNA_1000 (.A(net263));
 sg13g2_antennanp ANTENNA_1001 (.A(net263));
 sg13g2_antennanp ANTENNA_1002 (.A(net263));
 sg13g2_antennanp ANTENNA_1003 (.A(net264));
 sg13g2_antennanp ANTENNA_1004 (.A(net264));
 sg13g2_antennanp ANTENNA_1005 (.A(net264));
 sg13g2_antennanp ANTENNA_1006 (.A(net264));
 sg13g2_antennanp ANTENNA_1007 (.A(net264));
 sg13g2_antennanp ANTENNA_1008 (.A(net264));
 sg13g2_antennanp ANTENNA_1009 (.A(net264));
 sg13g2_antennanp ANTENNA_1010 (.A(net264));
 sg13g2_antennanp ANTENNA_1011 (.A(net264));
 sg13g2_antennanp ANTENNA_1012 (.A(net264));
 sg13g2_antennanp ANTENNA_1013 (.A(net264));
 sg13g2_antennanp ANTENNA_1014 (.A(net264));
 sg13g2_antennanp ANTENNA_1015 (.A(net264));
 sg13g2_antennanp ANTENNA_1016 (.A(net264));
 sg13g2_antennanp ANTENNA_1017 (.A(net264));
 sg13g2_antennanp ANTENNA_1018 (.A(net286));
 sg13g2_antennanp ANTENNA_1019 (.A(net286));
 sg13g2_antennanp ANTENNA_1020 (.A(net286));
 sg13g2_antennanp ANTENNA_1021 (.A(net286));
 sg13g2_antennanp ANTENNA_1022 (.A(net286));
 sg13g2_antennanp ANTENNA_1023 (.A(net286));
 sg13g2_antennanp ANTENNA_1024 (.A(net286));
 sg13g2_antennanp ANTENNA_1025 (.A(net286));
 sg13g2_antennanp ANTENNA_1026 (.A(net286));
 sg13g2_antennanp ANTENNA_1027 (.A(net286));
 sg13g2_antennanp ANTENNA_1028 (.A(net286));
 sg13g2_antennanp ANTENNA_1029 (.A(net286));
 sg13g2_antennanp ANTENNA_1030 (.A(net286));
 sg13g2_antennanp ANTENNA_1031 (.A(net286));
 sg13g2_antennanp ANTENNA_1032 (.A(net286));
 sg13g2_antennanp ANTENNA_1033 (.A(net286));
 sg13g2_antennanp ANTENNA_1034 (.A(net286));
 sg13g2_antennanp ANTENNA_1035 (.A(net286));
 sg13g2_antennanp ANTENNA_1036 (.A(net286));
 sg13g2_antennanp ANTENNA_1037 (.A(net286));
 sg13g2_antennanp ANTENNA_1038 (.A(net286));
 sg13g2_antennanp ANTENNA_1039 (.A(net286));
 sg13g2_antennanp ANTENNA_1040 (.A(net286));
 sg13g2_antennanp ANTENNA_1041 (.A(net286));
 sg13g2_antennanp ANTENNA_1042 (.A(net286));
 sg13g2_antennanp ANTENNA_1043 (.A(net286));
 sg13g2_antennanp ANTENNA_1044 (.A(net286));
 sg13g2_antennanp ANTENNA_1045 (.A(net286));
 sg13g2_antennanp ANTENNA_1046 (.A(net286));
 sg13g2_antennanp ANTENNA_1047 (.A(net286));
 sg13g2_antennanp ANTENNA_1048 (.A(net286));
 sg13g2_antennanp ANTENNA_1049 (.A(net286));
 sg13g2_antennanp ANTENNA_1050 (.A(net286));
 sg13g2_antennanp ANTENNA_1051 (.A(net286));
 sg13g2_antennanp ANTENNA_1052 (.A(net286));
 sg13g2_antennanp ANTENNA_1053 (.A(net286));
 sg13g2_antennanp ANTENNA_1054 (.A(net286));
 sg13g2_antennanp ANTENNA_1055 (.A(net286));
 sg13g2_antennanp ANTENNA_1056 (.A(net286));
 sg13g2_antennanp ANTENNA_1057 (.A(net286));
 sg13g2_antennanp ANTENNA_1058 (.A(net286));
 sg13g2_antennanp ANTENNA_1059 (.A(net286));
 sg13g2_antennanp ANTENNA_1060 (.A(net286));
 sg13g2_antennanp ANTENNA_1061 (.A(net286));
 sg13g2_antennanp ANTENNA_1062 (.A(net293));
 sg13g2_antennanp ANTENNA_1063 (.A(net293));
 sg13g2_antennanp ANTENNA_1064 (.A(net293));
 sg13g2_antennanp ANTENNA_1065 (.A(net293));
 sg13g2_antennanp ANTENNA_1066 (.A(net293));
 sg13g2_antennanp ANTENNA_1067 (.A(net293));
 sg13g2_antennanp ANTENNA_1068 (.A(net293));
 sg13g2_antennanp ANTENNA_1069 (.A(net293));
 sg13g2_antennanp ANTENNA_1070 (.A(net293));
 sg13g2_antennanp ANTENNA_1071 (.A(net293));
 sg13g2_antennanp ANTENNA_1072 (.A(net293));
 sg13g2_antennanp ANTENNA_1073 (.A(net293));
 sg13g2_antennanp ANTENNA_1074 (.A(net293));
 sg13g2_antennanp ANTENNA_1075 (.A(net293));
 sg13g2_antennanp ANTENNA_1076 (.A(net293));
 sg13g2_antennanp ANTENNA_1077 (.A(net293));
 sg13g2_antennanp ANTENNA_1078 (.A(net293));
 sg13g2_antennanp ANTENNA_1079 (.A(net293));
 sg13g2_antennanp ANTENNA_1080 (.A(net293));
 sg13g2_antennanp ANTENNA_1081 (.A(net293));
 sg13g2_antennanp ANTENNA_1082 (.A(net300));
 sg13g2_antennanp ANTENNA_1083 (.A(net300));
 sg13g2_antennanp ANTENNA_1084 (.A(net300));
 sg13g2_antennanp ANTENNA_1085 (.A(net300));
 sg13g2_antennanp ANTENNA_1086 (.A(net300));
 sg13g2_antennanp ANTENNA_1087 (.A(net300));
 sg13g2_antennanp ANTENNA_1088 (.A(net300));
 sg13g2_antennanp ANTENNA_1089 (.A(net300));
 sg13g2_antennanp ANTENNA_1090 (.A(net316));
 sg13g2_antennanp ANTENNA_1091 (.A(net316));
 sg13g2_antennanp ANTENNA_1092 (.A(net316));
 sg13g2_antennanp ANTENNA_1093 (.A(net316));
 sg13g2_antennanp ANTENNA_1094 (.A(net316));
 sg13g2_antennanp ANTENNA_1095 (.A(net316));
 sg13g2_antennanp ANTENNA_1096 (.A(net316));
 sg13g2_antennanp ANTENNA_1097 (.A(net316));
 sg13g2_antennanp ANTENNA_1098 (.A(net316));
 sg13g2_antennanp ANTENNA_1099 (.A(net316));
 sg13g2_antennanp ANTENNA_1100 (.A(net316));
 sg13g2_antennanp ANTENNA_1101 (.A(net316));
 sg13g2_antennanp ANTENNA_1102 (.A(net316));
 sg13g2_antennanp ANTENNA_1103 (.A(net323));
 sg13g2_antennanp ANTENNA_1104 (.A(net323));
 sg13g2_antennanp ANTENNA_1105 (.A(net323));
 sg13g2_antennanp ANTENNA_1106 (.A(net323));
 sg13g2_antennanp ANTENNA_1107 (.A(net323));
 sg13g2_antennanp ANTENNA_1108 (.A(net323));
 sg13g2_antennanp ANTENNA_1109 (.A(net323));
 sg13g2_antennanp ANTENNA_1110 (.A(net323));
 sg13g2_antennanp ANTENNA_1111 (.A(net323));
 sg13g2_antennanp ANTENNA_1112 (.A(net323));
 sg13g2_antennanp ANTENNA_1113 (.A(net323));
 sg13g2_antennanp ANTENNA_1114 (.A(net323));
 sg13g2_antennanp ANTENNA_1115 (.A(net323));
 sg13g2_antennanp ANTENNA_1116 (.A(net323));
 sg13g2_antennanp ANTENNA_1117 (.A(net323));
 sg13g2_antennanp ANTENNA_1118 (.A(net323));
 sg13g2_antennanp ANTENNA_1119 (.A(net323));
 sg13g2_antennanp ANTENNA_1120 (.A(net326));
 sg13g2_antennanp ANTENNA_1121 (.A(net326));
 sg13g2_antennanp ANTENNA_1122 (.A(net326));
 sg13g2_antennanp ANTENNA_1123 (.A(net326));
 sg13g2_antennanp ANTENNA_1124 (.A(net326));
 sg13g2_antennanp ANTENNA_1125 (.A(net326));
 sg13g2_antennanp ANTENNA_1126 (.A(net326));
 sg13g2_antennanp ANTENNA_1127 (.A(net326));
 sg13g2_antennanp ANTENNA_1128 (.A(net326));
 sg13g2_antennanp ANTENNA_1129 (.A(net326));
 sg13g2_antennanp ANTENNA_1130 (.A(net326));
 sg13g2_antennanp ANTENNA_1131 (.A(net326));
 sg13g2_antennanp ANTENNA_1132 (.A(net326));
 sg13g2_antennanp ANTENNA_1133 (.A(net326));
 sg13g2_antennanp ANTENNA_1134 (.A(net372));
 sg13g2_antennanp ANTENNA_1135 (.A(net372));
 sg13g2_antennanp ANTENNA_1136 (.A(net372));
 sg13g2_antennanp ANTENNA_1137 (.A(net372));
 sg13g2_antennanp ANTENNA_1138 (.A(net372));
 sg13g2_antennanp ANTENNA_1139 (.A(net372));
 sg13g2_antennanp ANTENNA_1140 (.A(net372));
 sg13g2_antennanp ANTENNA_1141 (.A(net372));
 sg13g2_antennanp ANTENNA_1142 (.A(net396));
 sg13g2_antennanp ANTENNA_1143 (.A(net396));
 sg13g2_antennanp ANTENNA_1144 (.A(net396));
 sg13g2_antennanp ANTENNA_1145 (.A(net396));
 sg13g2_antennanp ANTENNA_1146 (.A(net396));
 sg13g2_antennanp ANTENNA_1147 (.A(net396));
 sg13g2_antennanp ANTENNA_1148 (.A(net396));
 sg13g2_antennanp ANTENNA_1149 (.A(net396));
 sg13g2_antennanp ANTENNA_1150 (.A(net396));
 sg13g2_antennanp ANTENNA_1151 (.A(net396));
 sg13g2_antennanp ANTENNA_1152 (.A(net396));
 sg13g2_antennanp ANTENNA_1153 (.A(net396));
 sg13g2_antennanp ANTENNA_1154 (.A(net396));
 sg13g2_antennanp ANTENNA_1155 (.A(net396));
 sg13g2_antennanp ANTENNA_1156 (.A(net396));
 sg13g2_antennanp ANTENNA_1157 (.A(net403));
 sg13g2_antennanp ANTENNA_1158 (.A(net403));
 sg13g2_antennanp ANTENNA_1159 (.A(net403));
 sg13g2_antennanp ANTENNA_1160 (.A(net403));
 sg13g2_antennanp ANTENNA_1161 (.A(net403));
 sg13g2_antennanp ANTENNA_1162 (.A(net403));
 sg13g2_antennanp ANTENNA_1163 (.A(net403));
 sg13g2_antennanp ANTENNA_1164 (.A(net403));
 sg13g2_antennanp ANTENNA_1165 (.A(net403));
 sg13g2_antennanp ANTENNA_1166 (.A(net423));
 sg13g2_antennanp ANTENNA_1167 (.A(net423));
 sg13g2_antennanp ANTENNA_1168 (.A(net423));
 sg13g2_antennanp ANTENNA_1169 (.A(net423));
 sg13g2_antennanp ANTENNA_1170 (.A(net423));
 sg13g2_antennanp ANTENNA_1171 (.A(net423));
 sg13g2_antennanp ANTENNA_1172 (.A(net423));
 sg13g2_antennanp ANTENNA_1173 (.A(net423));
 sg13g2_antennanp ANTENNA_1174 (.A(net435));
 sg13g2_antennanp ANTENNA_1175 (.A(net435));
 sg13g2_antennanp ANTENNA_1176 (.A(net435));
 sg13g2_antennanp ANTENNA_1177 (.A(net435));
 sg13g2_antennanp ANTENNA_1178 (.A(net435));
 sg13g2_antennanp ANTENNA_1179 (.A(net435));
 sg13g2_antennanp ANTENNA_1180 (.A(net435));
 sg13g2_antennanp ANTENNA_1181 (.A(net435));
 sg13g2_antennanp ANTENNA_1182 (.A(net435));
 sg13g2_antennanp ANTENNA_1183 (.A(net440));
 sg13g2_antennanp ANTENNA_1184 (.A(net440));
 sg13g2_antennanp ANTENNA_1185 (.A(net440));
 sg13g2_antennanp ANTENNA_1186 (.A(net440));
 sg13g2_antennanp ANTENNA_1187 (.A(net440));
 sg13g2_antennanp ANTENNA_1188 (.A(net440));
 sg13g2_antennanp ANTENNA_1189 (.A(net440));
 sg13g2_antennanp ANTENNA_1190 (.A(net440));
 sg13g2_antennanp ANTENNA_1191 (.A(net440));
 sg13g2_antennanp ANTENNA_1192 (.A(net440));
 sg13g2_antennanp ANTENNA_1193 (.A(net440));
 sg13g2_antennanp ANTENNA_1194 (.A(net440));
 sg13g2_antennanp ANTENNA_1195 (.A(net441));
 sg13g2_antennanp ANTENNA_1196 (.A(net441));
 sg13g2_antennanp ANTENNA_1197 (.A(net441));
 sg13g2_antennanp ANTENNA_1198 (.A(net441));
 sg13g2_antennanp ANTENNA_1199 (.A(net441));
 sg13g2_antennanp ANTENNA_1200 (.A(net441));
 sg13g2_antennanp ANTENNA_1201 (.A(net441));
 sg13g2_antennanp ANTENNA_1202 (.A(net441));
 sg13g2_antennanp ANTENNA_1203 (.A(net441));
 sg13g2_antennanp ANTENNA_1204 (.A(net444));
 sg13g2_antennanp ANTENNA_1205 (.A(net444));
 sg13g2_antennanp ANTENNA_1206 (.A(net444));
 sg13g2_antennanp ANTENNA_1207 (.A(net444));
 sg13g2_antennanp ANTENNA_1208 (.A(net444));
 sg13g2_antennanp ANTENNA_1209 (.A(net444));
 sg13g2_antennanp ANTENNA_1210 (.A(net444));
 sg13g2_antennanp ANTENNA_1211 (.A(net444));
 sg13g2_antennanp ANTENNA_1212 (.A(net444));
 sg13g2_antennanp ANTENNA_1213 (.A(net444));
 sg13g2_antennanp ANTENNA_1214 (.A(net444));
 sg13g2_antennanp ANTENNA_1215 (.A(net444));
 sg13g2_antennanp ANTENNA_1216 (.A(net444));
 sg13g2_antennanp ANTENNA_1217 (.A(net444));
 sg13g2_antennanp ANTENNA_1218 (.A(net444));
 sg13g2_antennanp ANTENNA_1219 (.A(net444));
 sg13g2_antennanp ANTENNA_1220 (.A(net444));
 sg13g2_antennanp ANTENNA_1221 (.A(net444));
 sg13g2_antennanp ANTENNA_1222 (.A(net444));
 sg13g2_antennanp ANTENNA_1223 (.A(net444));
 sg13g2_antennanp ANTENNA_1224 (.A(net444));
 sg13g2_antennanp ANTENNA_1225 (.A(net444));
 sg13g2_antennanp ANTENNA_1226 (.A(net444));
 sg13g2_antennanp ANTENNA_1227 (.A(net449));
 sg13g2_antennanp ANTENNA_1228 (.A(net449));
 sg13g2_antennanp ANTENNA_1229 (.A(net449));
 sg13g2_antennanp ANTENNA_1230 (.A(net449));
 sg13g2_antennanp ANTENNA_1231 (.A(net449));
 sg13g2_antennanp ANTENNA_1232 (.A(net449));
 sg13g2_antennanp ANTENNA_1233 (.A(net449));
 sg13g2_antennanp ANTENNA_1234 (.A(net449));
 sg13g2_antennanp ANTENNA_1235 (.A(net487));
 sg13g2_antennanp ANTENNA_1236 (.A(net487));
 sg13g2_antennanp ANTENNA_1237 (.A(net487));
 sg13g2_antennanp ANTENNA_1238 (.A(net487));
 sg13g2_antennanp ANTENNA_1239 (.A(net487));
 sg13g2_antennanp ANTENNA_1240 (.A(net487));
 sg13g2_antennanp ANTENNA_1241 (.A(net487));
 sg13g2_antennanp ANTENNA_1242 (.A(net487));
 sg13g2_antennanp ANTENNA_1243 (.A(net487));
 sg13g2_antennanp ANTENNA_1244 (.A(net595));
 sg13g2_antennanp ANTENNA_1245 (.A(net595));
 sg13g2_antennanp ANTENNA_1246 (.A(net595));
 sg13g2_antennanp ANTENNA_1247 (.A(net595));
 sg13g2_antennanp ANTENNA_1248 (.A(net595));
 sg13g2_antennanp ANTENNA_1249 (.A(net595));
 sg13g2_antennanp ANTENNA_1250 (.A(net595));
 sg13g2_antennanp ANTENNA_1251 (.A(net595));
 sg13g2_antennanp ANTENNA_1252 (.A(net595));
 sg13g2_antennanp ANTENNA_1253 (.A(net595));
 sg13g2_antennanp ANTENNA_1254 (.A(net595));
 sg13g2_antennanp ANTENNA_1255 (.A(net595));
 sg13g2_antennanp ANTENNA_1256 (.A(net595));
 sg13g2_antennanp ANTENNA_1257 (.A(net595));
 sg13g2_antennanp ANTENNA_1258 (.A(net595));
 sg13g2_antennanp ANTENNA_1259 (.A(net595));
 sg13g2_antennanp ANTENNA_1260 (.A(net595));
 sg13g2_antennanp ANTENNA_1261 (.A(net595));
 sg13g2_antennanp ANTENNA_1262 (.A(net595));
 sg13g2_antennanp ANTENNA_1263 (.A(net603));
 sg13g2_antennanp ANTENNA_1264 (.A(net603));
 sg13g2_antennanp ANTENNA_1265 (.A(net603));
 sg13g2_antennanp ANTENNA_1266 (.A(net603));
 sg13g2_antennanp ANTENNA_1267 (.A(net603));
 sg13g2_antennanp ANTENNA_1268 (.A(net603));
 sg13g2_antennanp ANTENNA_1269 (.A(net603));
 sg13g2_antennanp ANTENNA_1270 (.A(net603));
 sg13g2_antennanp ANTENNA_1271 (.A(net603));
 sg13g2_antennanp ANTENNA_1272 (.A(net603));
 sg13g2_antennanp ANTENNA_1273 (.A(net603));
 sg13g2_antennanp ANTENNA_1274 (.A(net603));
 sg13g2_antennanp ANTENNA_1275 (.A(net603));
 sg13g2_antennanp ANTENNA_1276 (.A(net672));
 sg13g2_antennanp ANTENNA_1277 (.A(net672));
 sg13g2_antennanp ANTENNA_1278 (.A(net672));
 sg13g2_antennanp ANTENNA_1279 (.A(net672));
 sg13g2_antennanp ANTENNA_1280 (.A(net672));
 sg13g2_antennanp ANTENNA_1281 (.A(net672));
 sg13g2_antennanp ANTENNA_1282 (.A(net672));
 sg13g2_antennanp ANTENNA_1283 (.A(net672));
 sg13g2_antennanp ANTENNA_1284 (.A(net672));
 sg13g2_antennanp ANTENNA_1285 (.A(net672));
 sg13g2_antennanp ANTENNA_1286 (.A(net672));
 sg13g2_antennanp ANTENNA_1287 (.A(net672));
 sg13g2_antennanp ANTENNA_1288 (.A(net672));
 sg13g2_antennanp ANTENNA_1289 (.A(net692));
 sg13g2_antennanp ANTENNA_1290 (.A(net692));
 sg13g2_antennanp ANTENNA_1291 (.A(net692));
 sg13g2_antennanp ANTENNA_1292 (.A(net692));
 sg13g2_antennanp ANTENNA_1293 (.A(net692));
 sg13g2_antennanp ANTENNA_1294 (.A(net692));
 sg13g2_antennanp ANTENNA_1295 (.A(net692));
 sg13g2_antennanp ANTENNA_1296 (.A(net692));
 sg13g2_antennanp ANTENNA_1297 (.A(net692));
 sg13g2_antennanp ANTENNA_1298 (.A(net718));
 sg13g2_antennanp ANTENNA_1299 (.A(net718));
 sg13g2_antennanp ANTENNA_1300 (.A(net718));
 sg13g2_antennanp ANTENNA_1301 (.A(net718));
 sg13g2_antennanp ANTENNA_1302 (.A(net718));
 sg13g2_antennanp ANTENNA_1303 (.A(net718));
 sg13g2_antennanp ANTENNA_1304 (.A(net718));
 sg13g2_antennanp ANTENNA_1305 (.A(net718));
 sg13g2_antennanp ANTENNA_1306 (.A(net718));
 sg13g2_antennanp ANTENNA_1307 (.A(net718));
 sg13g2_antennanp ANTENNA_1308 (.A(net718));
 sg13g2_antennanp ANTENNA_1309 (.A(net718));
 sg13g2_antennanp ANTENNA_1310 (.A(net748));
 sg13g2_antennanp ANTENNA_1311 (.A(net748));
 sg13g2_antennanp ANTENNA_1312 (.A(net748));
 sg13g2_antennanp ANTENNA_1313 (.A(net748));
 sg13g2_antennanp ANTENNA_1314 (.A(net748));
 sg13g2_antennanp ANTENNA_1315 (.A(net748));
 sg13g2_antennanp ANTENNA_1316 (.A(net748));
 sg13g2_antennanp ANTENNA_1317 (.A(net748));
 sg13g2_antennanp ANTENNA_1318 (.A(net748));
 sg13g2_antennanp ANTENNA_1319 (.A(net748));
 sg13g2_antennanp ANTENNA_1320 (.A(net748));
 sg13g2_antennanp ANTENNA_1321 (.A(net748));
 sg13g2_antennanp ANTENNA_1322 (.A(net748));
 sg13g2_antennanp ANTENNA_1323 (.A(net748));
 sg13g2_antennanp ANTENNA_1324 (.A(net748));
 sg13g2_antennanp ANTENNA_1325 (.A(net748));
 sg13g2_antennanp ANTENNA_1326 (.A(net1046));
 sg13g2_antennanp ANTENNA_1327 (.A(net1046));
 sg13g2_antennanp ANTENNA_1328 (.A(net1046));
 sg13g2_antennanp ANTENNA_1329 (.A(net1046));
 sg13g2_antennanp ANTENNA_1330 (.A(net1046));
 sg13g2_antennanp ANTENNA_1331 (.A(net1046));
 sg13g2_antennanp ANTENNA_1332 (.A(net1046));
 sg13g2_antennanp ANTENNA_1333 (.A(net1046));
 sg13g2_antennanp ANTENNA_1334 (.A(net1053));
 sg13g2_antennanp ANTENNA_1335 (.A(net1053));
 sg13g2_antennanp ANTENNA_1336 (.A(net1053));
 sg13g2_antennanp ANTENNA_1337 (.A(net1053));
 sg13g2_antennanp ANTENNA_1338 (.A(net1053));
 sg13g2_antennanp ANTENNA_1339 (.A(net1053));
 sg13g2_antennanp ANTENNA_1340 (.A(net1053));
 sg13g2_antennanp ANTENNA_1341 (.A(net1053));
 sg13g2_antennanp ANTENNA_1342 (.A(net1053));
 sg13g2_antennanp ANTENNA_1343 (.A(net1053));
 sg13g2_antennanp ANTENNA_1344 (.A(net1053));
 sg13g2_antennanp ANTENNA_1345 (.A(net1053));
 sg13g2_antennanp ANTENNA_1346 (.A(net1053));
 sg13g2_antennanp ANTENNA_1347 (.A(net1053));
 sg13g2_antennanp ANTENNA_1348 (.A(net1053));
 sg13g2_antennanp ANTENNA_1349 (.A(net1053));
 sg13g2_antennanp ANTENNA_1350 (.A(net1053));
 sg13g2_antennanp ANTENNA_1351 (.A(net1053));
 sg13g2_antennanp ANTENNA_1352 (.A(net1053));
 sg13g2_antennanp ANTENNA_1353 (.A(net1053));
 sg13g2_antennanp ANTENNA_1354 (.A(net1421));
 sg13g2_antennanp ANTENNA_1355 (.A(net1421));
 sg13g2_antennanp ANTENNA_1356 (.A(net1421));
 sg13g2_antennanp ANTENNA_1357 (.A(net1421));
 sg13g2_antennanp ANTENNA_1358 (.A(net1421));
 sg13g2_antennanp ANTENNA_1359 (.A(net1421));
 sg13g2_antennanp ANTENNA_1360 (.A(net1421));
 sg13g2_antennanp ANTENNA_1361 (.A(net1421));
 sg13g2_antennanp ANTENNA_1362 (.A(net1421));
 sg13g2_antennanp ANTENNA_1363 (.A(net1421));
 sg13g2_antennanp ANTENNA_1364 (.A(net1421));
 sg13g2_antennanp ANTENNA_1365 (.A(net1421));
 sg13g2_antennanp ANTENNA_1366 (.A(net1421));
 sg13g2_antennanp ANTENNA_1367 (.A(net1421));
 sg13g2_antennanp ANTENNA_1368 (.A(net1421));
 sg13g2_antennanp ANTENNA_1369 (.A(net1421));
 sg13g2_antennanp ANTENNA_1370 (.A(net1421));
 sg13g2_antennanp ANTENNA_1371 (.A(net1421));
 sg13g2_antennanp ANTENNA_1372 (.A(net1421));
 sg13g2_antennanp ANTENNA_1373 (.A(net1421));
 sg13g2_antennanp ANTENNA_1374 (.A(net1421));
 sg13g2_antennanp ANTENNA_1375 (.A(net1421));
 sg13g2_antennanp ANTENNA_1376 (.A(net1421));
 sg13g2_antennanp ANTENNA_1377 (.A(net1421));
 sg13g2_antennanp ANTENNA_1378 (.A(net1421));
 sg13g2_antennanp ANTENNA_1379 (.A(net1421));
 sg13g2_antennanp ANTENNA_1380 (.A(net1421));
 sg13g2_antennanp ANTENNA_1381 (.A(net1421));
 sg13g2_antennanp ANTENNA_1382 (.A(net1421));
 sg13g2_antennanp ANTENNA_1383 (.A(net1421));
 sg13g2_antennanp ANTENNA_1384 (.A(net1421));
 sg13g2_antennanp ANTENNA_1385 (.A(net1421));
 sg13g2_antennanp ANTENNA_1386 (.A(net1421));
 sg13g2_antennanp ANTENNA_1387 (.A(net1421));
 sg13g2_antennanp ANTENNA_1388 (.A(net1421));
 sg13g2_antennanp ANTENNA_1389 (.A(net1421));
 sg13g2_antennanp ANTENNA_1390 (.A(net1421));
 sg13g2_antennanp ANTENNA_1391 (.A(net1421));
 sg13g2_antennanp ANTENNA_1392 (.A(net1421));
 sg13g2_antennanp ANTENNA_1393 (.A(net1421));
 sg13g2_antennanp ANTENNA_1394 (.A(net1421));
 sg13g2_antennanp ANTENNA_1395 (.A(net1421));
 sg13g2_antennanp ANTENNA_1396 (.A(net1421));
 sg13g2_antennanp ANTENNA_1397 (.A(net1421));
 sg13g2_antennanp ANTENNA_1398 (.A(net1421));
 sg13g2_antennanp ANTENNA_1399 (.A(net1421));
 sg13g2_antennanp ANTENNA_1400 (.A(net1421));
 sg13g2_antennanp ANTENNA_1401 (.A(net1421));
 sg13g2_antennanp ANTENNA_1402 (.A(net1421));
 sg13g2_antennanp ANTENNA_1403 (.A(net1421));
 sg13g2_antennanp ANTENNA_1404 (.A(net1421));
 sg13g2_antennanp ANTENNA_1405 (.A(_00356_));
 sg13g2_antennanp ANTENNA_1406 (.A(_00410_));
 sg13g2_antennanp ANTENNA_1407 (.A(_00422_));
 sg13g2_antennanp ANTENNA_1408 (.A(_00425_));
 sg13g2_antennanp ANTENNA_1409 (.A(_00432_));
 sg13g2_antennanp ANTENNA_1410 (.A(_00443_));
 sg13g2_antennanp ANTENNA_1411 (.A(_02799_));
 sg13g2_antennanp ANTENNA_1412 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1413 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1414 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1415 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1416 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1417 (.A(_02946_));
 sg13g2_antennanp ANTENNA_1418 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1419 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1420 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1421 (.A(_03019_));
 sg13g2_antennanp ANTENNA_1422 (.A(_03060_));
 sg13g2_antennanp ANTENNA_1423 (.A(_03060_));
 sg13g2_antennanp ANTENNA_1424 (.A(_03060_));
 sg13g2_antennanp ANTENNA_1425 (.A(_03079_));
 sg13g2_antennanp ANTENNA_1426 (.A(_03079_));
 sg13g2_antennanp ANTENNA_1427 (.A(_03268_));
 sg13g2_antennanp ANTENNA_1428 (.A(_03268_));
 sg13g2_antennanp ANTENNA_1429 (.A(_03268_));
 sg13g2_antennanp ANTENNA_1430 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1431 (.A(_03684_));
 sg13g2_antennanp ANTENNA_1432 (.A(_03714_));
 sg13g2_antennanp ANTENNA_1433 (.A(_03714_));
 sg13g2_antennanp ANTENNA_1434 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1435 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1436 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1437 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1438 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1439 (.A(_03760_));
 sg13g2_antennanp ANTENNA_1440 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1441 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1442 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1443 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1444 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1445 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1446 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1447 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1448 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1449 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1450 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1451 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1452 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1453 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1454 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1455 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1456 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1457 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1458 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1459 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1460 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1461 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1462 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1463 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1464 (.A(_04617_));
 sg13g2_antennanp ANTENNA_1465 (.A(_04620_));
 sg13g2_antennanp ANTENNA_1466 (.A(_04674_));
 sg13g2_antennanp ANTENNA_1467 (.A(_04676_));
 sg13g2_antennanp ANTENNA_1468 (.A(_04676_));
 sg13g2_antennanp ANTENNA_1469 (.A(_05061_));
 sg13g2_antennanp ANTENNA_1470 (.A(_05061_));
 sg13g2_antennanp ANTENNA_1471 (.A(_05067_));
 sg13g2_antennanp ANTENNA_1472 (.A(_05067_));
 sg13g2_antennanp ANTENNA_1473 (.A(_05091_));
 sg13g2_antennanp ANTENNA_1474 (.A(_05091_));
 sg13g2_antennanp ANTENNA_1475 (.A(_05091_));
 sg13g2_antennanp ANTENNA_1476 (.A(_05276_));
 sg13g2_antennanp ANTENNA_1477 (.A(_05276_));
 sg13g2_antennanp ANTENNA_1478 (.A(_05276_));
 sg13g2_antennanp ANTENNA_1479 (.A(_05276_));
 sg13g2_antennanp ANTENNA_1480 (.A(_05278_));
 sg13g2_antennanp ANTENNA_1481 (.A(_05290_));
 sg13g2_antennanp ANTENNA_1482 (.A(_05303_));
 sg13g2_antennanp ANTENNA_1483 (.A(_05303_));
 sg13g2_antennanp ANTENNA_1484 (.A(_05303_));
 sg13g2_antennanp ANTENNA_1485 (.A(_05318_));
 sg13g2_antennanp ANTENNA_1486 (.A(_05347_));
 sg13g2_antennanp ANTENNA_1487 (.A(_05347_));
 sg13g2_antennanp ANTENNA_1488 (.A(_05347_));
 sg13g2_antennanp ANTENNA_1489 (.A(_05347_));
 sg13g2_antennanp ANTENNA_1490 (.A(_05347_));
 sg13g2_antennanp ANTENNA_1491 (.A(_05350_));
 sg13g2_antennanp ANTENNA_1492 (.A(_05364_));
 sg13g2_antennanp ANTENNA_1493 (.A(_05432_));
 sg13g2_antennanp ANTENNA_1494 (.A(_05465_));
 sg13g2_antennanp ANTENNA_1495 (.A(_05465_));
 sg13g2_antennanp ANTENNA_1496 (.A(_05465_));
 sg13g2_antennanp ANTENNA_1497 (.A(_05465_));
 sg13g2_antennanp ANTENNA_1498 (.A(_05512_));
 sg13g2_antennanp ANTENNA_1499 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1500 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1501 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1502 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1503 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1504 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1505 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1506 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1507 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1508 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1509 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1510 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1511 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1512 (.A(_05525_));
 sg13g2_antennanp ANTENNA_1513 (.A(_05577_));
 sg13g2_antennanp ANTENNA_1514 (.A(_05584_));
 sg13g2_antennanp ANTENNA_1515 (.A(_05640_));
 sg13g2_antennanp ANTENNA_1516 (.A(_05640_));
 sg13g2_antennanp ANTENNA_1517 (.A(_05640_));
 sg13g2_antennanp ANTENNA_1518 (.A(_05652_));
 sg13g2_antennanp ANTENNA_1519 (.A(_05652_));
 sg13g2_antennanp ANTENNA_1520 (.A(_05652_));
 sg13g2_antennanp ANTENNA_1521 (.A(_05663_));
 sg13g2_antennanp ANTENNA_1522 (.A(_05663_));
 sg13g2_antennanp ANTENNA_1523 (.A(_05663_));
 sg13g2_antennanp ANTENNA_1524 (.A(_05663_));
 sg13g2_antennanp ANTENNA_1525 (.A(_05672_));
 sg13g2_antennanp ANTENNA_1526 (.A(_05707_));
 sg13g2_antennanp ANTENNA_1527 (.A(_05707_));
 sg13g2_antennanp ANTENNA_1528 (.A(_05707_));
 sg13g2_antennanp ANTENNA_1529 (.A(_05754_));
 sg13g2_antennanp ANTENNA_1530 (.A(_05788_));
 sg13g2_antennanp ANTENNA_1531 (.A(_05788_));
 sg13g2_antennanp ANTENNA_1532 (.A(_05788_));
 sg13g2_antennanp ANTENNA_1533 (.A(_05788_));
 sg13g2_antennanp ANTENNA_1534 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1535 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1536 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1537 (.A(_05811_));
 sg13g2_antennanp ANTENNA_1538 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1539 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1540 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1541 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1542 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1543 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1544 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1545 (.A(_05851_));
 sg13g2_antennanp ANTENNA_1546 (.A(_05868_));
 sg13g2_antennanp ANTENNA_1547 (.A(_05872_));
 sg13g2_antennanp ANTENNA_1548 (.A(_05892_));
 sg13g2_antennanp ANTENNA_1549 (.A(_05892_));
 sg13g2_antennanp ANTENNA_1550 (.A(_05892_));
 sg13g2_antennanp ANTENNA_1551 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1552 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1553 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1554 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1555 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1556 (.A(_05901_));
 sg13g2_antennanp ANTENNA_1557 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1558 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1559 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1560 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1561 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1562 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1563 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1564 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1565 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1566 (.A(_05932_));
 sg13g2_antennanp ANTENNA_1567 (.A(_05936_));
 sg13g2_antennanp ANTENNA_1568 (.A(_05940_));
 sg13g2_antennanp ANTENNA_1569 (.A(_05953_));
 sg13g2_antennanp ANTENNA_1570 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1571 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1572 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1573 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1574 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1575 (.A(_06009_));
 sg13g2_antennanp ANTENNA_1576 (.A(_06027_));
 sg13g2_antennanp ANTENNA_1577 (.A(_06076_));
 sg13g2_antennanp ANTENNA_1578 (.A(_06090_));
 sg13g2_antennanp ANTENNA_1579 (.A(_06090_));
 sg13g2_antennanp ANTENNA_1580 (.A(_06101_));
 sg13g2_antennanp ANTENNA_1581 (.A(_06184_));
 sg13g2_antennanp ANTENNA_1582 (.A(_06214_));
 sg13g2_antennanp ANTENNA_1583 (.A(_06244_));
 sg13g2_antennanp ANTENNA_1584 (.A(_06254_));
 sg13g2_antennanp ANTENNA_1585 (.A(_06255_));
 sg13g2_antennanp ANTENNA_1586 (.A(_06265_));
 sg13g2_antennanp ANTENNA_1587 (.A(_06302_));
 sg13g2_antennanp ANTENNA_1588 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1589 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1590 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1591 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1592 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1593 (.A(_06313_));
 sg13g2_antennanp ANTENNA_1594 (.A(_06345_));
 sg13g2_antennanp ANTENNA_1595 (.A(_06351_));
 sg13g2_antennanp ANTENNA_1596 (.A(_06359_));
 sg13g2_antennanp ANTENNA_1597 (.A(_06440_));
 sg13g2_antennanp ANTENNA_1598 (.A(_06440_));
 sg13g2_antennanp ANTENNA_1599 (.A(_06443_));
 sg13g2_antennanp ANTENNA_1600 (.A(_06447_));
 sg13g2_antennanp ANTENNA_1601 (.A(_06467_));
 sg13g2_antennanp ANTENNA_1602 (.A(_06489_));
 sg13g2_antennanp ANTENNA_1603 (.A(_06530_));
 sg13g2_antennanp ANTENNA_1604 (.A(_06533_));
 sg13g2_antennanp ANTENNA_1605 (.A(_06538_));
 sg13g2_antennanp ANTENNA_1606 (.A(_06545_));
 sg13g2_antennanp ANTENNA_1607 (.A(_06587_));
 sg13g2_antennanp ANTENNA_1608 (.A(_06591_));
 sg13g2_antennanp ANTENNA_1609 (.A(_06591_));
 sg13g2_antennanp ANTENNA_1610 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1611 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1612 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1613 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1614 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1615 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1616 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1617 (.A(_06601_));
 sg13g2_antennanp ANTENNA_1618 (.A(_06603_));
 sg13g2_antennanp ANTENNA_1619 (.A(_06603_));
 sg13g2_antennanp ANTENNA_1620 (.A(_06609_));
 sg13g2_antennanp ANTENNA_1621 (.A(_06619_));
 sg13g2_antennanp ANTENNA_1622 (.A(_06651_));
 sg13g2_antennanp ANTENNA_1623 (.A(_06654_));
 sg13g2_antennanp ANTENNA_1624 (.A(_06662_));
 sg13g2_antennanp ANTENNA_1625 (.A(_06671_));
 sg13g2_antennanp ANTENNA_1626 (.A(_06708_));
 sg13g2_antennanp ANTENNA_1627 (.A(_06708_));
 sg13g2_antennanp ANTENNA_1628 (.A(_06708_));
 sg13g2_antennanp ANTENNA_1629 (.A(_06716_));
 sg13g2_antennanp ANTENNA_1630 (.A(_06721_));
 sg13g2_antennanp ANTENNA_1631 (.A(_06722_));
 sg13g2_antennanp ANTENNA_1632 (.A(_06735_));
 sg13g2_antennanp ANTENNA_1633 (.A(_06740_));
 sg13g2_antennanp ANTENNA_1634 (.A(_06741_));
 sg13g2_antennanp ANTENNA_1635 (.A(_06751_));
 sg13g2_antennanp ANTENNA_1636 (.A(_06780_));
 sg13g2_antennanp ANTENNA_1637 (.A(_06792_));
 sg13g2_antennanp ANTENNA_1638 (.A(_06793_));
 sg13g2_antennanp ANTENNA_1639 (.A(_06807_));
 sg13g2_antennanp ANTENNA_1640 (.A(_06838_));
 sg13g2_antennanp ANTENNA_1641 (.A(_06853_));
 sg13g2_antennanp ANTENNA_1642 (.A(_06874_));
 sg13g2_antennanp ANTENNA_1643 (.A(_06875_));
 sg13g2_antennanp ANTENNA_1644 (.A(_06895_));
 sg13g2_antennanp ANTENNA_1645 (.A(_06902_));
 sg13g2_antennanp ANTENNA_1646 (.A(_06945_));
 sg13g2_antennanp ANTENNA_1647 (.A(_06963_));
 sg13g2_antennanp ANTENNA_1648 (.A(_06980_));
 sg13g2_antennanp ANTENNA_1649 (.A(_06980_));
 sg13g2_antennanp ANTENNA_1650 (.A(_06980_));
 sg13g2_antennanp ANTENNA_1651 (.A(_06980_));
 sg13g2_antennanp ANTENNA_1652 (.A(_06981_));
 sg13g2_antennanp ANTENNA_1653 (.A(_06985_));
 sg13g2_antennanp ANTENNA_1654 (.A(_07020_));
 sg13g2_antennanp ANTENNA_1655 (.A(_07032_));
 sg13g2_antennanp ANTENNA_1656 (.A(_07063_));
 sg13g2_antennanp ANTENNA_1657 (.A(_07064_));
 sg13g2_antennanp ANTENNA_1658 (.A(_07064_));
 sg13g2_antennanp ANTENNA_1659 (.A(_07073_));
 sg13g2_antennanp ANTENNA_1660 (.A(_07074_));
 sg13g2_antennanp ANTENNA_1661 (.A(_07077_));
 sg13g2_antennanp ANTENNA_1662 (.A(_07085_));
 sg13g2_antennanp ANTENNA_1663 (.A(_07104_));
 sg13g2_antennanp ANTENNA_1664 (.A(_07113_));
 sg13g2_antennanp ANTENNA_1665 (.A(_07125_));
 sg13g2_antennanp ANTENNA_1666 (.A(_07129_));
 sg13g2_antennanp ANTENNA_1667 (.A(_07150_));
 sg13g2_antennanp ANTENNA_1668 (.A(_07151_));
 sg13g2_antennanp ANTENNA_1669 (.A(_07157_));
 sg13g2_antennanp ANTENNA_1670 (.A(_07157_));
 sg13g2_antennanp ANTENNA_1671 (.A(_07157_));
 sg13g2_antennanp ANTENNA_1672 (.A(_07172_));
 sg13g2_antennanp ANTENNA_1673 (.A(_07188_));
 sg13g2_antennanp ANTENNA_1674 (.A(_07195_));
 sg13g2_antennanp ANTENNA_1675 (.A(_07201_));
 sg13g2_antennanp ANTENNA_1676 (.A(_07221_));
 sg13g2_antennanp ANTENNA_1677 (.A(_07222_));
 sg13g2_antennanp ANTENNA_1678 (.A(_07243_));
 sg13g2_antennanp ANTENNA_1679 (.A(_07243_));
 sg13g2_antennanp ANTENNA_1680 (.A(_07269_));
 sg13g2_antennanp ANTENNA_1681 (.A(_07279_));
 sg13g2_antennanp ANTENNA_1682 (.A(_07282_));
 sg13g2_antennanp ANTENNA_1683 (.A(_07344_));
 sg13g2_antennanp ANTENNA_1684 (.A(_07345_));
 sg13g2_antennanp ANTENNA_1685 (.A(_07371_));
 sg13g2_antennanp ANTENNA_1686 (.A(_07381_));
 sg13g2_antennanp ANTENNA_1687 (.A(_07385_));
 sg13g2_antennanp ANTENNA_1688 (.A(_07421_));
 sg13g2_antennanp ANTENNA_1689 (.A(_07429_));
 sg13g2_antennanp ANTENNA_1690 (.A(_07435_));
 sg13g2_antennanp ANTENNA_1691 (.A(_07440_));
 sg13g2_antennanp ANTENNA_1692 (.A(_07446_));
 sg13g2_antennanp ANTENNA_1693 (.A(_07480_));
 sg13g2_antennanp ANTENNA_1694 (.A(_07485_));
 sg13g2_antennanp ANTENNA_1695 (.A(_07507_));
 sg13g2_antennanp ANTENNA_1696 (.A(_07535_));
 sg13g2_antennanp ANTENNA_1697 (.A(_07540_));
 sg13g2_antennanp ANTENNA_1698 (.A(_07544_));
 sg13g2_antennanp ANTENNA_1699 (.A(_07552_));
 sg13g2_antennanp ANTENNA_1700 (.A(_07560_));
 sg13g2_antennanp ANTENNA_1701 (.A(_07592_));
 sg13g2_antennanp ANTENNA_1702 (.A(_07595_));
 sg13g2_antennanp ANTENNA_1703 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1704 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1705 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1706 (.A(_07601_));
 sg13g2_antennanp ANTENNA_1707 (.A(_07603_));
 sg13g2_antennanp ANTENNA_1708 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1709 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1710 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1711 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1712 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1713 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1714 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1715 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1716 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1717 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1718 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1719 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1720 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1721 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1722 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1723 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1724 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1725 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1726 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1727 (.A(_07633_));
 sg13g2_antennanp ANTENNA_1728 (.A(_07634_));
 sg13g2_antennanp ANTENNA_1729 (.A(_07913_));
 sg13g2_antennanp ANTENNA_1730 (.A(_07945_));
 sg13g2_antennanp ANTENNA_1731 (.A(_07979_));
 sg13g2_antennanp ANTENNA_1732 (.A(_08062_));
 sg13g2_antennanp ANTENNA_1733 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1734 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1735 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1736 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1737 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1738 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1739 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1740 (.A(_08219_));
 sg13g2_antennanp ANTENNA_1741 (.A(_08221_));
 sg13g2_antennanp ANTENNA_1742 (.A(_08221_));
 sg13g2_antennanp ANTENNA_1743 (.A(_08221_));
 sg13g2_antennanp ANTENNA_1744 (.A(_08223_));
 sg13g2_antennanp ANTENNA_1745 (.A(_08223_));
 sg13g2_antennanp ANTENNA_1746 (.A(_08223_));
 sg13g2_antennanp ANTENNA_1747 (.A(_08223_));
 sg13g2_antennanp ANTENNA_1748 (.A(_08227_));
 sg13g2_antennanp ANTENNA_1749 (.A(_08227_));
 sg13g2_antennanp ANTENNA_1750 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1751 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1752 (.A(_08260_));
 sg13g2_antennanp ANTENNA_1753 (.A(_08261_));
 sg13g2_antennanp ANTENNA_1754 (.A(_08261_));
 sg13g2_antennanp ANTENNA_1755 (.A(_08261_));
 sg13g2_antennanp ANTENNA_1756 (.A(_08261_));
 sg13g2_antennanp ANTENNA_1757 (.A(_08261_));
 sg13g2_antennanp ANTENNA_1758 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1759 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1760 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1761 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1762 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1763 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1764 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1765 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1766 (.A(_08263_));
 sg13g2_antennanp ANTENNA_1767 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1768 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1769 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1770 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1771 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1772 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1773 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1774 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1775 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1776 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1777 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1778 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1779 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1780 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1781 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1782 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1783 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1784 (.A(_08321_));
 sg13g2_antennanp ANTENNA_1785 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1786 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1787 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1788 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1789 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1790 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1791 (.A(_08354_));
 sg13g2_antennanp ANTENNA_1792 (.A(_08380_));
 sg13g2_antennanp ANTENNA_1793 (.A(_08380_));
 sg13g2_antennanp ANTENNA_1794 (.A(_08380_));
 sg13g2_antennanp ANTENNA_1795 (.A(_08380_));
 sg13g2_antennanp ANTENNA_1796 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1797 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1798 (.A(_08706_));
 sg13g2_antennanp ANTENNA_1799 (.A(_08730_));
 sg13g2_antennanp ANTENNA_1800 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1801 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1802 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1803 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1804 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1805 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1806 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1807 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1808 (.A(_08985_));
 sg13g2_antennanp ANTENNA_1809 (.A(_08993_));
 sg13g2_antennanp ANTENNA_1810 (.A(_08993_));
 sg13g2_antennanp ANTENNA_1811 (.A(_08993_));
 sg13g2_antennanp ANTENNA_1812 (.A(_09940_));
 sg13g2_antennanp ANTENNA_1813 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1814 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1815 (.A(_10089_));
 sg13g2_antennanp ANTENNA_1816 (.A(_10158_));
 sg13g2_antennanp ANTENNA_1817 (.A(_10158_));
 sg13g2_antennanp ANTENNA_1818 (.A(_10158_));
 sg13g2_antennanp ANTENNA_1819 (.A(_10158_));
 sg13g2_antennanp ANTENNA_1820 (.A(_10159_));
 sg13g2_antennanp ANTENNA_1821 (.A(_10159_));
 sg13g2_antennanp ANTENNA_1822 (.A(_10159_));
 sg13g2_antennanp ANTENNA_1823 (.A(_10204_));
 sg13g2_antennanp ANTENNA_1824 (.A(_10318_));
 sg13g2_antennanp ANTENNA_1825 (.A(_10318_));
 sg13g2_antennanp ANTENNA_1826 (.A(_10318_));
 sg13g2_antennanp ANTENNA_1827 (.A(_10342_));
 sg13g2_antennanp ANTENNA_1828 (.A(_10342_));
 sg13g2_antennanp ANTENNA_1829 (.A(_10361_));
 sg13g2_antennanp ANTENNA_1830 (.A(_10361_));
 sg13g2_antennanp ANTENNA_1831 (.A(_10361_));
 sg13g2_antennanp ANTENNA_1832 (.A(_10361_));
 sg13g2_antennanp ANTENNA_1833 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1834 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1835 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1836 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1837 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1838 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1839 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1840 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1841 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1842 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1843 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1844 (.A(_10424_));
 sg13g2_antennanp ANTENNA_1845 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1846 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1847 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1848 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1849 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1850 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1851 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1852 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1853 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1854 (.A(_10429_));
 sg13g2_antennanp ANTENNA_1855 (.A(_10450_));
 sg13g2_antennanp ANTENNA_1856 (.A(_10450_));
 sg13g2_antennanp ANTENNA_1857 (.A(_10450_));
 sg13g2_antennanp ANTENNA_1858 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1859 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1860 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1861 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1862 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1863 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1864 (.A(_10535_));
 sg13g2_antennanp ANTENNA_1865 (.A(_10599_));
 sg13g2_antennanp ANTENNA_1866 (.A(_10599_));
 sg13g2_antennanp ANTENNA_1867 (.A(_10599_));
 sg13g2_antennanp ANTENNA_1868 (.A(_10600_));
 sg13g2_antennanp ANTENNA_1869 (.A(_10600_));
 sg13g2_antennanp ANTENNA_1870 (.A(_10600_));
 sg13g2_antennanp ANTENNA_1871 (.A(_10600_));
 sg13g2_antennanp ANTENNA_1872 (.A(_10704_));
 sg13g2_antennanp ANTENNA_1873 (.A(_10704_));
 sg13g2_antennanp ANTENNA_1874 (.A(_10704_));
 sg13g2_antennanp ANTENNA_1875 (.A(_10726_));
 sg13g2_antennanp ANTENNA_1876 (.A(_10726_));
 sg13g2_antennanp ANTENNA_1877 (.A(_10726_));
 sg13g2_antennanp ANTENNA_1878 (.A(_10739_));
 sg13g2_antennanp ANTENNA_1879 (.A(_10739_));
 sg13g2_antennanp ANTENNA_1880 (.A(_10739_));
 sg13g2_antennanp ANTENNA_1881 (.A(_10739_));
 sg13g2_antennanp ANTENNA_1882 (.A(_10740_));
 sg13g2_antennanp ANTENNA_1883 (.A(_10740_));
 sg13g2_antennanp ANTENNA_1884 (.A(_10740_));
 sg13g2_antennanp ANTENNA_1885 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1886 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1887 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1888 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1889 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1890 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1891 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1892 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1893 (.A(_10742_));
 sg13g2_antennanp ANTENNA_1894 (.A(_10745_));
 sg13g2_antennanp ANTENNA_1895 (.A(_10745_));
 sg13g2_antennanp ANTENNA_1896 (.A(_10745_));
 sg13g2_antennanp ANTENNA_1897 (.A(_10779_));
 sg13g2_antennanp ANTENNA_1898 (.A(_10779_));
 sg13g2_antennanp ANTENNA_1899 (.A(_10779_));
 sg13g2_antennanp ANTENNA_1900 (.A(_10797_));
 sg13g2_antennanp ANTENNA_1901 (.A(_10797_));
 sg13g2_antennanp ANTENNA_1902 (.A(_10797_));
 sg13g2_antennanp ANTENNA_1903 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1904 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1905 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1906 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1907 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1908 (.A(_10812_));
 sg13g2_antennanp ANTENNA_1909 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1910 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1911 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1912 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1913 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1914 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1915 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1916 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1917 (.A(_10845_));
 sg13g2_antennanp ANTENNA_1918 (.A(clk));
 sg13g2_antennanp ANTENNA_1919 (.A(clk));
 sg13g2_antennanp ANTENNA_1920 (.A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_antennanp ANTENNA_1921 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_1922 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_1923 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_1924 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1925 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1926 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1927 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1928 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1929 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1930 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1931 (.A(\top_ihp.oisc.reg_rb[2] ));
 sg13g2_antennanp ANTENNA_1932 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_1933 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_1934 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_1935 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_1936 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1937 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1938 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_1939 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_1940 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_1941 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_1942 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1943 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1944 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_1945 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_1946 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_1947 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_1948 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1949 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1950 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1951 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_1952 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1953 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1954 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1955 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_1956 (.A(\top_ihp.oisc.regs[59][23] ));
 sg13g2_antennanp ANTENNA_1957 (.A(\top_ihp.oisc.regs[59][23] ));
 sg13g2_antennanp ANTENNA_1958 (.A(\top_ihp.oisc.regs[59][23] ));
 sg13g2_antennanp ANTENNA_1959 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_1960 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_1961 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_1962 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_1963 (.A(net54));
 sg13g2_antennanp ANTENNA_1964 (.A(net54));
 sg13g2_antennanp ANTENNA_1965 (.A(net54));
 sg13g2_antennanp ANTENNA_1966 (.A(net54));
 sg13g2_antennanp ANTENNA_1967 (.A(net54));
 sg13g2_antennanp ANTENNA_1968 (.A(net54));
 sg13g2_antennanp ANTENNA_1969 (.A(net54));
 sg13g2_antennanp ANTENNA_1970 (.A(net54));
 sg13g2_antennanp ANTENNA_1971 (.A(net56));
 sg13g2_antennanp ANTENNA_1972 (.A(net56));
 sg13g2_antennanp ANTENNA_1973 (.A(net56));
 sg13g2_antennanp ANTENNA_1974 (.A(net56));
 sg13g2_antennanp ANTENNA_1975 (.A(net56));
 sg13g2_antennanp ANTENNA_1976 (.A(net56));
 sg13g2_antennanp ANTENNA_1977 (.A(net56));
 sg13g2_antennanp ANTENNA_1978 (.A(net56));
 sg13g2_antennanp ANTENNA_1979 (.A(net56));
 sg13g2_antennanp ANTENNA_1980 (.A(net59));
 sg13g2_antennanp ANTENNA_1981 (.A(net59));
 sg13g2_antennanp ANTENNA_1982 (.A(net59));
 sg13g2_antennanp ANTENNA_1983 (.A(net59));
 sg13g2_antennanp ANTENNA_1984 (.A(net59));
 sg13g2_antennanp ANTENNA_1985 (.A(net59));
 sg13g2_antennanp ANTENNA_1986 (.A(net59));
 sg13g2_antennanp ANTENNA_1987 (.A(net59));
 sg13g2_antennanp ANTENNA_1988 (.A(net69));
 sg13g2_antennanp ANTENNA_1989 (.A(net69));
 sg13g2_antennanp ANTENNA_1990 (.A(net69));
 sg13g2_antennanp ANTENNA_1991 (.A(net69));
 sg13g2_antennanp ANTENNA_1992 (.A(net69));
 sg13g2_antennanp ANTENNA_1993 (.A(net69));
 sg13g2_antennanp ANTENNA_1994 (.A(net69));
 sg13g2_antennanp ANTENNA_1995 (.A(net69));
 sg13g2_antennanp ANTENNA_1996 (.A(net90));
 sg13g2_antennanp ANTENNA_1997 (.A(net90));
 sg13g2_antennanp ANTENNA_1998 (.A(net90));
 sg13g2_antennanp ANTENNA_1999 (.A(net90));
 sg13g2_antennanp ANTENNA_2000 (.A(net90));
 sg13g2_antennanp ANTENNA_2001 (.A(net90));
 sg13g2_antennanp ANTENNA_2002 (.A(net90));
 sg13g2_antennanp ANTENNA_2003 (.A(net90));
 sg13g2_antennanp ANTENNA_2004 (.A(net90));
 sg13g2_antennanp ANTENNA_2005 (.A(net117));
 sg13g2_antennanp ANTENNA_2006 (.A(net117));
 sg13g2_antennanp ANTENNA_2007 (.A(net117));
 sg13g2_antennanp ANTENNA_2008 (.A(net117));
 sg13g2_antennanp ANTENNA_2009 (.A(net117));
 sg13g2_antennanp ANTENNA_2010 (.A(net117));
 sg13g2_antennanp ANTENNA_2011 (.A(net117));
 sg13g2_antennanp ANTENNA_2012 (.A(net117));
 sg13g2_antennanp ANTENNA_2013 (.A(net117));
 sg13g2_antennanp ANTENNA_2014 (.A(net117));
 sg13g2_antennanp ANTENNA_2015 (.A(net117));
 sg13g2_antennanp ANTENNA_2016 (.A(net117));
 sg13g2_antennanp ANTENNA_2017 (.A(net117));
 sg13g2_antennanp ANTENNA_2018 (.A(net117));
 sg13g2_antennanp ANTENNA_2019 (.A(net117));
 sg13g2_antennanp ANTENNA_2020 (.A(net117));
 sg13g2_antennanp ANTENNA_2021 (.A(net117));
 sg13g2_antennanp ANTENNA_2022 (.A(net117));
 sg13g2_antennanp ANTENNA_2023 (.A(net117));
 sg13g2_antennanp ANTENNA_2024 (.A(net117));
 sg13g2_antennanp ANTENNA_2025 (.A(net121));
 sg13g2_antennanp ANTENNA_2026 (.A(net121));
 sg13g2_antennanp ANTENNA_2027 (.A(net121));
 sg13g2_antennanp ANTENNA_2028 (.A(net121));
 sg13g2_antennanp ANTENNA_2029 (.A(net121));
 sg13g2_antennanp ANTENNA_2030 (.A(net121));
 sg13g2_antennanp ANTENNA_2031 (.A(net121));
 sg13g2_antennanp ANTENNA_2032 (.A(net121));
 sg13g2_antennanp ANTENNA_2033 (.A(net123));
 sg13g2_antennanp ANTENNA_2034 (.A(net123));
 sg13g2_antennanp ANTENNA_2035 (.A(net123));
 sg13g2_antennanp ANTENNA_2036 (.A(net123));
 sg13g2_antennanp ANTENNA_2037 (.A(net123));
 sg13g2_antennanp ANTENNA_2038 (.A(net123));
 sg13g2_antennanp ANTENNA_2039 (.A(net123));
 sg13g2_antennanp ANTENNA_2040 (.A(net123));
 sg13g2_antennanp ANTENNA_2041 (.A(net123));
 sg13g2_antennanp ANTENNA_2042 (.A(net125));
 sg13g2_antennanp ANTENNA_2043 (.A(net125));
 sg13g2_antennanp ANTENNA_2044 (.A(net125));
 sg13g2_antennanp ANTENNA_2045 (.A(net125));
 sg13g2_antennanp ANTENNA_2046 (.A(net125));
 sg13g2_antennanp ANTENNA_2047 (.A(net125));
 sg13g2_antennanp ANTENNA_2048 (.A(net125));
 sg13g2_antennanp ANTENNA_2049 (.A(net125));
 sg13g2_antennanp ANTENNA_2050 (.A(net126));
 sg13g2_antennanp ANTENNA_2051 (.A(net126));
 sg13g2_antennanp ANTENNA_2052 (.A(net126));
 sg13g2_antennanp ANTENNA_2053 (.A(net126));
 sg13g2_antennanp ANTENNA_2054 (.A(net126));
 sg13g2_antennanp ANTENNA_2055 (.A(net126));
 sg13g2_antennanp ANTENNA_2056 (.A(net126));
 sg13g2_antennanp ANTENNA_2057 (.A(net126));
 sg13g2_antennanp ANTENNA_2058 (.A(net127));
 sg13g2_antennanp ANTENNA_2059 (.A(net127));
 sg13g2_antennanp ANTENNA_2060 (.A(net127));
 sg13g2_antennanp ANTENNA_2061 (.A(net127));
 sg13g2_antennanp ANTENNA_2062 (.A(net127));
 sg13g2_antennanp ANTENNA_2063 (.A(net127));
 sg13g2_antennanp ANTENNA_2064 (.A(net127));
 sg13g2_antennanp ANTENNA_2065 (.A(net127));
 sg13g2_antennanp ANTENNA_2066 (.A(net127));
 sg13g2_antennanp ANTENNA_2067 (.A(net127));
 sg13g2_antennanp ANTENNA_2068 (.A(net127));
 sg13g2_antennanp ANTENNA_2069 (.A(net127));
 sg13g2_antennanp ANTENNA_2070 (.A(net127));
 sg13g2_antennanp ANTENNA_2071 (.A(net127));
 sg13g2_antennanp ANTENNA_2072 (.A(net127));
 sg13g2_antennanp ANTENNA_2073 (.A(net127));
 sg13g2_antennanp ANTENNA_2074 (.A(net127));
 sg13g2_antennanp ANTENNA_2075 (.A(net127));
 sg13g2_antennanp ANTENNA_2076 (.A(net127));
 sg13g2_antennanp ANTENNA_2077 (.A(net127));
 sg13g2_antennanp ANTENNA_2078 (.A(net130));
 sg13g2_antennanp ANTENNA_2079 (.A(net130));
 sg13g2_antennanp ANTENNA_2080 (.A(net130));
 sg13g2_antennanp ANTENNA_2081 (.A(net130));
 sg13g2_antennanp ANTENNA_2082 (.A(net130));
 sg13g2_antennanp ANTENNA_2083 (.A(net130));
 sg13g2_antennanp ANTENNA_2084 (.A(net130));
 sg13g2_antennanp ANTENNA_2085 (.A(net130));
 sg13g2_antennanp ANTENNA_2086 (.A(net130));
 sg13g2_antennanp ANTENNA_2087 (.A(net130));
 sg13g2_antennanp ANTENNA_2088 (.A(net130));
 sg13g2_antennanp ANTENNA_2089 (.A(net130));
 sg13g2_antennanp ANTENNA_2090 (.A(net130));
 sg13g2_antennanp ANTENNA_2091 (.A(net130));
 sg13g2_antennanp ANTENNA_2092 (.A(net130));
 sg13g2_antennanp ANTENNA_2093 (.A(net130));
 sg13g2_antennanp ANTENNA_2094 (.A(net130));
 sg13g2_antennanp ANTENNA_2095 (.A(net130));
 sg13g2_antennanp ANTENNA_2096 (.A(net130));
 sg13g2_antennanp ANTENNA_2097 (.A(net130));
 sg13g2_antennanp ANTENNA_2098 (.A(net130));
 sg13g2_antennanp ANTENNA_2099 (.A(net130));
 sg13g2_antennanp ANTENNA_2100 (.A(net130));
 sg13g2_antennanp ANTENNA_2101 (.A(net132));
 sg13g2_antennanp ANTENNA_2102 (.A(net132));
 sg13g2_antennanp ANTENNA_2103 (.A(net132));
 sg13g2_antennanp ANTENNA_2104 (.A(net132));
 sg13g2_antennanp ANTENNA_2105 (.A(net132));
 sg13g2_antennanp ANTENNA_2106 (.A(net132));
 sg13g2_antennanp ANTENNA_2107 (.A(net132));
 sg13g2_antennanp ANTENNA_2108 (.A(net132));
 sg13g2_antennanp ANTENNA_2109 (.A(net132));
 sg13g2_antennanp ANTENNA_2110 (.A(net134));
 sg13g2_antennanp ANTENNA_2111 (.A(net134));
 sg13g2_antennanp ANTENNA_2112 (.A(net134));
 sg13g2_antennanp ANTENNA_2113 (.A(net134));
 sg13g2_antennanp ANTENNA_2114 (.A(net134));
 sg13g2_antennanp ANTENNA_2115 (.A(net134));
 sg13g2_antennanp ANTENNA_2116 (.A(net134));
 sg13g2_antennanp ANTENNA_2117 (.A(net134));
 sg13g2_antennanp ANTENNA_2118 (.A(net134));
 sg13g2_antennanp ANTENNA_2119 (.A(net134));
 sg13g2_antennanp ANTENNA_2120 (.A(net134));
 sg13g2_antennanp ANTENNA_2121 (.A(net134));
 sg13g2_antennanp ANTENNA_2122 (.A(net134));
 sg13g2_antennanp ANTENNA_2123 (.A(net134));
 sg13g2_antennanp ANTENNA_2124 (.A(net134));
 sg13g2_antennanp ANTENNA_2125 (.A(net134));
 sg13g2_antennanp ANTENNA_2126 (.A(net134));
 sg13g2_antennanp ANTENNA_2127 (.A(net134));
 sg13g2_antennanp ANTENNA_2128 (.A(net134));
 sg13g2_antennanp ANTENNA_2129 (.A(net134));
 sg13g2_antennanp ANTENNA_2130 (.A(net143));
 sg13g2_antennanp ANTENNA_2131 (.A(net143));
 sg13g2_antennanp ANTENNA_2132 (.A(net143));
 sg13g2_antennanp ANTENNA_2133 (.A(net143));
 sg13g2_antennanp ANTENNA_2134 (.A(net143));
 sg13g2_antennanp ANTENNA_2135 (.A(net143));
 sg13g2_antennanp ANTENNA_2136 (.A(net143));
 sg13g2_antennanp ANTENNA_2137 (.A(net143));
 sg13g2_antennanp ANTENNA_2138 (.A(net143));
 sg13g2_antennanp ANTENNA_2139 (.A(net159));
 sg13g2_antennanp ANTENNA_2140 (.A(net159));
 sg13g2_antennanp ANTENNA_2141 (.A(net159));
 sg13g2_antennanp ANTENNA_2142 (.A(net159));
 sg13g2_antennanp ANTENNA_2143 (.A(net159));
 sg13g2_antennanp ANTENNA_2144 (.A(net159));
 sg13g2_antennanp ANTENNA_2145 (.A(net159));
 sg13g2_antennanp ANTENNA_2146 (.A(net159));
 sg13g2_antennanp ANTENNA_2147 (.A(net177));
 sg13g2_antennanp ANTENNA_2148 (.A(net177));
 sg13g2_antennanp ANTENNA_2149 (.A(net177));
 sg13g2_antennanp ANTENNA_2150 (.A(net177));
 sg13g2_antennanp ANTENNA_2151 (.A(net177));
 sg13g2_antennanp ANTENNA_2152 (.A(net177));
 sg13g2_antennanp ANTENNA_2153 (.A(net177));
 sg13g2_antennanp ANTENNA_2154 (.A(net177));
 sg13g2_antennanp ANTENNA_2155 (.A(net177));
 sg13g2_antennanp ANTENNA_2156 (.A(net177));
 sg13g2_antennanp ANTENNA_2157 (.A(net177));
 sg13g2_antennanp ANTENNA_2158 (.A(net177));
 sg13g2_antennanp ANTENNA_2159 (.A(net177));
 sg13g2_antennanp ANTENNA_2160 (.A(net177));
 sg13g2_antennanp ANTENNA_2161 (.A(net188));
 sg13g2_antennanp ANTENNA_2162 (.A(net188));
 sg13g2_antennanp ANTENNA_2163 (.A(net188));
 sg13g2_antennanp ANTENNA_2164 (.A(net188));
 sg13g2_antennanp ANTENNA_2165 (.A(net188));
 sg13g2_antennanp ANTENNA_2166 (.A(net188));
 sg13g2_antennanp ANTENNA_2167 (.A(net188));
 sg13g2_antennanp ANTENNA_2168 (.A(net188));
 sg13g2_antennanp ANTENNA_2169 (.A(net264));
 sg13g2_antennanp ANTENNA_2170 (.A(net264));
 sg13g2_antennanp ANTENNA_2171 (.A(net264));
 sg13g2_antennanp ANTENNA_2172 (.A(net264));
 sg13g2_antennanp ANTENNA_2173 (.A(net264));
 sg13g2_antennanp ANTENNA_2174 (.A(net264));
 sg13g2_antennanp ANTENNA_2175 (.A(net264));
 sg13g2_antennanp ANTENNA_2176 (.A(net264));
 sg13g2_antennanp ANTENNA_2177 (.A(net264));
 sg13g2_antennanp ANTENNA_2178 (.A(net323));
 sg13g2_antennanp ANTENNA_2179 (.A(net323));
 sg13g2_antennanp ANTENNA_2180 (.A(net323));
 sg13g2_antennanp ANTENNA_2181 (.A(net323));
 sg13g2_antennanp ANTENNA_2182 (.A(net323));
 sg13g2_antennanp ANTENNA_2183 (.A(net323));
 sg13g2_antennanp ANTENNA_2184 (.A(net323));
 sg13g2_antennanp ANTENNA_2185 (.A(net323));
 sg13g2_antennanp ANTENNA_2186 (.A(net323));
 sg13g2_antennanp ANTENNA_2187 (.A(net326));
 sg13g2_antennanp ANTENNA_2188 (.A(net326));
 sg13g2_antennanp ANTENNA_2189 (.A(net326));
 sg13g2_antennanp ANTENNA_2190 (.A(net326));
 sg13g2_antennanp ANTENNA_2191 (.A(net326));
 sg13g2_antennanp ANTENNA_2192 (.A(net326));
 sg13g2_antennanp ANTENNA_2193 (.A(net326));
 sg13g2_antennanp ANTENNA_2194 (.A(net326));
 sg13g2_antennanp ANTENNA_2195 (.A(net345));
 sg13g2_antennanp ANTENNA_2196 (.A(net345));
 sg13g2_antennanp ANTENNA_2197 (.A(net345));
 sg13g2_antennanp ANTENNA_2198 (.A(net345));
 sg13g2_antennanp ANTENNA_2199 (.A(net345));
 sg13g2_antennanp ANTENNA_2200 (.A(net345));
 sg13g2_antennanp ANTENNA_2201 (.A(net345));
 sg13g2_antennanp ANTENNA_2202 (.A(net345));
 sg13g2_antennanp ANTENNA_2203 (.A(net372));
 sg13g2_antennanp ANTENNA_2204 (.A(net372));
 sg13g2_antennanp ANTENNA_2205 (.A(net372));
 sg13g2_antennanp ANTENNA_2206 (.A(net372));
 sg13g2_antennanp ANTENNA_2207 (.A(net372));
 sg13g2_antennanp ANTENNA_2208 (.A(net372));
 sg13g2_antennanp ANTENNA_2209 (.A(net372));
 sg13g2_antennanp ANTENNA_2210 (.A(net372));
 sg13g2_antennanp ANTENNA_2211 (.A(net403));
 sg13g2_antennanp ANTENNA_2212 (.A(net403));
 sg13g2_antennanp ANTENNA_2213 (.A(net403));
 sg13g2_antennanp ANTENNA_2214 (.A(net403));
 sg13g2_antennanp ANTENNA_2215 (.A(net403));
 sg13g2_antennanp ANTENNA_2216 (.A(net403));
 sg13g2_antennanp ANTENNA_2217 (.A(net403));
 sg13g2_antennanp ANTENNA_2218 (.A(net403));
 sg13g2_antennanp ANTENNA_2219 (.A(net403));
 sg13g2_antennanp ANTENNA_2220 (.A(net435));
 sg13g2_antennanp ANTENNA_2221 (.A(net435));
 sg13g2_antennanp ANTENNA_2222 (.A(net435));
 sg13g2_antennanp ANTENNA_2223 (.A(net435));
 sg13g2_antennanp ANTENNA_2224 (.A(net435));
 sg13g2_antennanp ANTENNA_2225 (.A(net435));
 sg13g2_antennanp ANTENNA_2226 (.A(net435));
 sg13g2_antennanp ANTENNA_2227 (.A(net435));
 sg13g2_antennanp ANTENNA_2228 (.A(net435));
 sg13g2_antennanp ANTENNA_2229 (.A(net444));
 sg13g2_antennanp ANTENNA_2230 (.A(net444));
 sg13g2_antennanp ANTENNA_2231 (.A(net444));
 sg13g2_antennanp ANTENNA_2232 (.A(net444));
 sg13g2_antennanp ANTENNA_2233 (.A(net444));
 sg13g2_antennanp ANTENNA_2234 (.A(net444));
 sg13g2_antennanp ANTENNA_2235 (.A(net444));
 sg13g2_antennanp ANTENNA_2236 (.A(net444));
 sg13g2_antennanp ANTENNA_2237 (.A(net444));
 sg13g2_antennanp ANTENNA_2238 (.A(net446));
 sg13g2_antennanp ANTENNA_2239 (.A(net446));
 sg13g2_antennanp ANTENNA_2240 (.A(net446));
 sg13g2_antennanp ANTENNA_2241 (.A(net446));
 sg13g2_antennanp ANTENNA_2242 (.A(net446));
 sg13g2_antennanp ANTENNA_2243 (.A(net446));
 sg13g2_antennanp ANTENNA_2244 (.A(net446));
 sg13g2_antennanp ANTENNA_2245 (.A(net446));
 sg13g2_antennanp ANTENNA_2246 (.A(net449));
 sg13g2_antennanp ANTENNA_2247 (.A(net449));
 sg13g2_antennanp ANTENNA_2248 (.A(net449));
 sg13g2_antennanp ANTENNA_2249 (.A(net449));
 sg13g2_antennanp ANTENNA_2250 (.A(net449));
 sg13g2_antennanp ANTENNA_2251 (.A(net449));
 sg13g2_antennanp ANTENNA_2252 (.A(net449));
 sg13g2_antennanp ANTENNA_2253 (.A(net449));
 sg13g2_antennanp ANTENNA_2254 (.A(net449));
 sg13g2_antennanp ANTENNA_2255 (.A(net449));
 sg13g2_antennanp ANTENNA_2256 (.A(net449));
 sg13g2_antennanp ANTENNA_2257 (.A(net449));
 sg13g2_antennanp ANTENNA_2258 (.A(net449));
 sg13g2_antennanp ANTENNA_2259 (.A(net449));
 sg13g2_antennanp ANTENNA_2260 (.A(net449));
 sg13g2_antennanp ANTENNA_2261 (.A(net487));
 sg13g2_antennanp ANTENNA_2262 (.A(net487));
 sg13g2_antennanp ANTENNA_2263 (.A(net487));
 sg13g2_antennanp ANTENNA_2264 (.A(net487));
 sg13g2_antennanp ANTENNA_2265 (.A(net487));
 sg13g2_antennanp ANTENNA_2266 (.A(net487));
 sg13g2_antennanp ANTENNA_2267 (.A(net487));
 sg13g2_antennanp ANTENNA_2268 (.A(net487));
 sg13g2_antennanp ANTENNA_2269 (.A(net487));
 sg13g2_antennanp ANTENNA_2270 (.A(net598));
 sg13g2_antennanp ANTENNA_2271 (.A(net598));
 sg13g2_antennanp ANTENNA_2272 (.A(net598));
 sg13g2_antennanp ANTENNA_2273 (.A(net598));
 sg13g2_antennanp ANTENNA_2274 (.A(net598));
 sg13g2_antennanp ANTENNA_2275 (.A(net598));
 sg13g2_antennanp ANTENNA_2276 (.A(net598));
 sg13g2_antennanp ANTENNA_2277 (.A(net598));
 sg13g2_antennanp ANTENNA_2278 (.A(net605));
 sg13g2_antennanp ANTENNA_2279 (.A(net605));
 sg13g2_antennanp ANTENNA_2280 (.A(net605));
 sg13g2_antennanp ANTENNA_2281 (.A(net605));
 sg13g2_antennanp ANTENNA_2282 (.A(net605));
 sg13g2_antennanp ANTENNA_2283 (.A(net605));
 sg13g2_antennanp ANTENNA_2284 (.A(net605));
 sg13g2_antennanp ANTENNA_2285 (.A(net605));
 sg13g2_antennanp ANTENNA_2286 (.A(net672));
 sg13g2_antennanp ANTENNA_2287 (.A(net672));
 sg13g2_antennanp ANTENNA_2288 (.A(net672));
 sg13g2_antennanp ANTENNA_2289 (.A(net672));
 sg13g2_antennanp ANTENNA_2290 (.A(net672));
 sg13g2_antennanp ANTENNA_2291 (.A(net672));
 sg13g2_antennanp ANTENNA_2292 (.A(net672));
 sg13g2_antennanp ANTENNA_2293 (.A(net672));
 sg13g2_antennanp ANTENNA_2294 (.A(net748));
 sg13g2_antennanp ANTENNA_2295 (.A(net748));
 sg13g2_antennanp ANTENNA_2296 (.A(net748));
 sg13g2_antennanp ANTENNA_2297 (.A(net748));
 sg13g2_antennanp ANTENNA_2298 (.A(net748));
 sg13g2_antennanp ANTENNA_2299 (.A(net748));
 sg13g2_antennanp ANTENNA_2300 (.A(net748));
 sg13g2_antennanp ANTENNA_2301 (.A(net748));
 sg13g2_antennanp ANTENNA_2302 (.A(net748));
 sg13g2_antennanp ANTENNA_2303 (.A(net1421));
 sg13g2_antennanp ANTENNA_2304 (.A(net1421));
 sg13g2_antennanp ANTENNA_2305 (.A(net1421));
 sg13g2_antennanp ANTENNA_2306 (.A(net1421));
 sg13g2_antennanp ANTENNA_2307 (.A(net1421));
 sg13g2_antennanp ANTENNA_2308 (.A(net1421));
 sg13g2_antennanp ANTENNA_2309 (.A(net1421));
 sg13g2_antennanp ANTENNA_2310 (.A(net1421));
 sg13g2_antennanp ANTENNA_2311 (.A(net1421));
 sg13g2_antennanp ANTENNA_2312 (.A(net1421));
 sg13g2_antennanp ANTENNA_2313 (.A(net1421));
 sg13g2_antennanp ANTENNA_2314 (.A(net1421));
 sg13g2_antennanp ANTENNA_2315 (.A(net1421));
 sg13g2_antennanp ANTENNA_2316 (.A(net1421));
 sg13g2_antennanp ANTENNA_2317 (.A(net1421));
 sg13g2_antennanp ANTENNA_2318 (.A(net1421));
 sg13g2_antennanp ANTENNA_2319 (.A(net1421));
 sg13g2_antennanp ANTENNA_2320 (.A(net1421));
 sg13g2_antennanp ANTENNA_2321 (.A(net1421));
 sg13g2_antennanp ANTENNA_2322 (.A(net1421));
 sg13g2_antennanp ANTENNA_2323 (.A(net1421));
 sg13g2_antennanp ANTENNA_2324 (.A(net1421));
 sg13g2_antennanp ANTENNA_2325 (.A(net1421));
 sg13g2_antennanp ANTENNA_2326 (.A(_00356_));
 sg13g2_antennanp ANTENNA_2327 (.A(_00410_));
 sg13g2_antennanp ANTENNA_2328 (.A(_00422_));
 sg13g2_antennanp ANTENNA_2329 (.A(_00425_));
 sg13g2_antennanp ANTENNA_2330 (.A(_00432_));
 sg13g2_antennanp ANTENNA_2331 (.A(_02799_));
 sg13g2_antennanp ANTENNA_2332 (.A(_03060_));
 sg13g2_antennanp ANTENNA_2333 (.A(_03060_));
 sg13g2_antennanp ANTENNA_2334 (.A(_03060_));
 sg13g2_antennanp ANTENNA_2335 (.A(_03268_));
 sg13g2_antennanp ANTENNA_2336 (.A(_03268_));
 sg13g2_antennanp ANTENNA_2337 (.A(_03268_));
 sg13g2_antennanp ANTENNA_2338 (.A(_03268_));
 sg13g2_antennanp ANTENNA_2339 (.A(_03684_));
 sg13g2_antennanp ANTENNA_2340 (.A(_03684_));
 sg13g2_antennanp ANTENNA_2341 (.A(_03714_));
 sg13g2_antennanp ANTENNA_2342 (.A(_03714_));
 sg13g2_antennanp ANTENNA_2343 (.A(_03714_));
 sg13g2_antennanp ANTENNA_2344 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2345 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2346 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2347 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2348 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2349 (.A(_03760_));
 sg13g2_antennanp ANTENNA_2350 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2351 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2352 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2353 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2354 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2355 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2356 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2357 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2358 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2359 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2360 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2361 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2362 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2363 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2364 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2365 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2366 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2367 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2368 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2369 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2370 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2371 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2372 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2373 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2374 (.A(_04617_));
 sg13g2_antennanp ANTENNA_2375 (.A(_04620_));
 sg13g2_antennanp ANTENNA_2376 (.A(_04674_));
 sg13g2_antennanp ANTENNA_2377 (.A(_04676_));
 sg13g2_antennanp ANTENNA_2378 (.A(_05061_));
 sg13g2_antennanp ANTENNA_2379 (.A(_05067_));
 sg13g2_antennanp ANTENNA_2380 (.A(_05091_));
 sg13g2_antennanp ANTENNA_2381 (.A(_05276_));
 sg13g2_antennanp ANTENNA_2382 (.A(_05276_));
 sg13g2_antennanp ANTENNA_2383 (.A(_05276_));
 sg13g2_antennanp ANTENNA_2384 (.A(_05276_));
 sg13g2_antennanp ANTENNA_2385 (.A(_05278_));
 sg13g2_antennanp ANTENNA_2386 (.A(_05290_));
 sg13g2_antennanp ANTENNA_2387 (.A(_05303_));
 sg13g2_antennanp ANTENNA_2388 (.A(_05303_));
 sg13g2_antennanp ANTENNA_2389 (.A(_05303_));
 sg13g2_antennanp ANTENNA_2390 (.A(_05303_));
 sg13g2_antennanp ANTENNA_2391 (.A(_05318_));
 sg13g2_antennanp ANTENNA_2392 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2393 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2394 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2395 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2396 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2397 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2398 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2399 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2400 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2401 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2402 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2403 (.A(_05347_));
 sg13g2_antennanp ANTENNA_2404 (.A(_05350_));
 sg13g2_antennanp ANTENNA_2405 (.A(_05364_));
 sg13g2_antennanp ANTENNA_2406 (.A(_05432_));
 sg13g2_antennanp ANTENNA_2407 (.A(_05465_));
 sg13g2_antennanp ANTENNA_2408 (.A(_05465_));
 sg13g2_antennanp ANTENNA_2409 (.A(_05465_));
 sg13g2_antennanp ANTENNA_2410 (.A(_05465_));
 sg13g2_antennanp ANTENNA_2411 (.A(_05512_));
 sg13g2_antennanp ANTENNA_2412 (.A(_05577_));
 sg13g2_antennanp ANTENNA_2413 (.A(_05584_));
 sg13g2_antennanp ANTENNA_2414 (.A(_05652_));
 sg13g2_antennanp ANTENNA_2415 (.A(_05652_));
 sg13g2_antennanp ANTENNA_2416 (.A(_05652_));
 sg13g2_antennanp ANTENNA_2417 (.A(_05652_));
 sg13g2_antennanp ANTENNA_2418 (.A(_05672_));
 sg13g2_antennanp ANTENNA_2419 (.A(_05754_));
 sg13g2_antennanp ANTENNA_2420 (.A(_05788_));
 sg13g2_antennanp ANTENNA_2421 (.A(_05788_));
 sg13g2_antennanp ANTENNA_2422 (.A(_05788_));
 sg13g2_antennanp ANTENNA_2423 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2424 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2425 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2426 (.A(_05811_));
 sg13g2_antennanp ANTENNA_2427 (.A(_05868_));
 sg13g2_antennanp ANTENNA_2428 (.A(_05872_));
 sg13g2_antennanp ANTENNA_2429 (.A(_05892_));
 sg13g2_antennanp ANTENNA_2430 (.A(_05892_));
 sg13g2_antennanp ANTENNA_2431 (.A(_05892_));
 sg13g2_antennanp ANTENNA_2432 (.A(_05892_));
 sg13g2_antennanp ANTENNA_2433 (.A(_05892_));
 sg13g2_antennanp ANTENNA_2434 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2435 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2436 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2437 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2438 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2439 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2440 (.A(_05901_));
 sg13g2_antennanp ANTENNA_2441 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2442 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2443 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2444 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2445 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2446 (.A(_05932_));
 sg13g2_antennanp ANTENNA_2447 (.A(_05936_));
 sg13g2_antennanp ANTENNA_2448 (.A(_05940_));
 sg13g2_antennanp ANTENNA_2449 (.A(_05953_));
 sg13g2_antennanp ANTENNA_2450 (.A(_06009_));
 sg13g2_antennanp ANTENNA_2451 (.A(_06009_));
 sg13g2_antennanp ANTENNA_2452 (.A(_06027_));
 sg13g2_antennanp ANTENNA_2453 (.A(_06076_));
 sg13g2_antennanp ANTENNA_2454 (.A(_06090_));
 sg13g2_antennanp ANTENNA_2455 (.A(_06101_));
 sg13g2_antennanp ANTENNA_2456 (.A(_06167_));
 sg13g2_antennanp ANTENNA_2457 (.A(_06184_));
 sg13g2_antennanp ANTENNA_2458 (.A(_06214_));
 sg13g2_antennanp ANTENNA_2459 (.A(_06244_));
 sg13g2_antennanp ANTENNA_2460 (.A(_06254_));
 sg13g2_antennanp ANTENNA_2461 (.A(_06255_));
 sg13g2_antennanp ANTENNA_2462 (.A(_06265_));
 sg13g2_antennanp ANTENNA_2463 (.A(_06302_));
 sg13g2_antennanp ANTENNA_2464 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2465 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2466 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2467 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2468 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2469 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2470 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2471 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2472 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2473 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2474 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2475 (.A(_06313_));
 sg13g2_antennanp ANTENNA_2476 (.A(_06330_));
 sg13g2_antennanp ANTENNA_2477 (.A(_06345_));
 sg13g2_antennanp ANTENNA_2478 (.A(_06351_));
 sg13g2_antennanp ANTENNA_2479 (.A(_06359_));
 sg13g2_antennanp ANTENNA_2480 (.A(_06440_));
 sg13g2_antennanp ANTENNA_2481 (.A(_06440_));
 sg13g2_antennanp ANTENNA_2482 (.A(_06443_));
 sg13g2_antennanp ANTENNA_2483 (.A(_06447_));
 sg13g2_antennanp ANTENNA_2484 (.A(_06489_));
 sg13g2_antennanp ANTENNA_2485 (.A(_06489_));
 sg13g2_antennanp ANTENNA_2486 (.A(_06530_));
 sg13g2_antennanp ANTENNA_2487 (.A(_06533_));
 sg13g2_antennanp ANTENNA_2488 (.A(_06538_));
 sg13g2_antennanp ANTENNA_2489 (.A(_06545_));
 sg13g2_antennanp ANTENNA_2490 (.A(_06587_));
 sg13g2_antennanp ANTENNA_2491 (.A(_06591_));
 sg13g2_antennanp ANTENNA_2492 (.A(_06591_));
 sg13g2_antennanp ANTENNA_2493 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2494 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2495 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2496 (.A(_06601_));
 sg13g2_antennanp ANTENNA_2497 (.A(_06603_));
 sg13g2_antennanp ANTENNA_2498 (.A(_06609_));
 sg13g2_antennanp ANTENNA_2499 (.A(_06619_));
 sg13g2_antennanp ANTENNA_2500 (.A(_06651_));
 sg13g2_antennanp ANTENNA_2501 (.A(_06654_));
 sg13g2_antennanp ANTENNA_2502 (.A(_06654_));
 sg13g2_antennanp ANTENNA_2503 (.A(_06662_));
 sg13g2_antennanp ANTENNA_2504 (.A(_06671_));
 sg13g2_antennanp ANTENNA_2505 (.A(_06708_));
 sg13g2_antennanp ANTENNA_2506 (.A(_06708_));
 sg13g2_antennanp ANTENNA_2507 (.A(_06708_));
 sg13g2_antennanp ANTENNA_2508 (.A(_06716_));
 sg13g2_antennanp ANTENNA_2509 (.A(_06721_));
 sg13g2_antennanp ANTENNA_2510 (.A(_06722_));
 sg13g2_antennanp ANTENNA_2511 (.A(_06735_));
 sg13g2_antennanp ANTENNA_2512 (.A(_06740_));
 sg13g2_antennanp ANTENNA_2513 (.A(_06741_));
 sg13g2_antennanp ANTENNA_2514 (.A(_06751_));
 sg13g2_antennanp ANTENNA_2515 (.A(_06780_));
 sg13g2_antennanp ANTENNA_2516 (.A(_06792_));
 sg13g2_antennanp ANTENNA_2517 (.A(_06793_));
 sg13g2_antennanp ANTENNA_2518 (.A(_06807_));
 sg13g2_antennanp ANTENNA_2519 (.A(_06838_));
 sg13g2_antennanp ANTENNA_2520 (.A(_06853_));
 sg13g2_antennanp ANTENNA_2521 (.A(_06874_));
 sg13g2_antennanp ANTENNA_2522 (.A(_06875_));
 sg13g2_antennanp ANTENNA_2523 (.A(_06902_));
 sg13g2_antennanp ANTENNA_2524 (.A(_06945_));
 sg13g2_antennanp ANTENNA_2525 (.A(_06963_));
 sg13g2_antennanp ANTENNA_2526 (.A(_06980_));
 sg13g2_antennanp ANTENNA_2527 (.A(_06980_));
 sg13g2_antennanp ANTENNA_2528 (.A(_06980_));
 sg13g2_antennanp ANTENNA_2529 (.A(_06980_));
 sg13g2_antennanp ANTENNA_2530 (.A(_06981_));
 sg13g2_antennanp ANTENNA_2531 (.A(_06985_));
 sg13g2_antennanp ANTENNA_2532 (.A(_07020_));
 sg13g2_antennanp ANTENNA_2533 (.A(_07032_));
 sg13g2_antennanp ANTENNA_2534 (.A(_07063_));
 sg13g2_antennanp ANTENNA_2535 (.A(_07064_));
 sg13g2_antennanp ANTENNA_2536 (.A(_07064_));
 sg13g2_antennanp ANTENNA_2537 (.A(_07073_));
 sg13g2_antennanp ANTENNA_2538 (.A(_07074_));
 sg13g2_antennanp ANTENNA_2539 (.A(_07077_));
 sg13g2_antennanp ANTENNA_2540 (.A(_07085_));
 sg13g2_antennanp ANTENNA_2541 (.A(_07104_));
 sg13g2_antennanp ANTENNA_2542 (.A(_07113_));
 sg13g2_antennanp ANTENNA_2543 (.A(_07125_));
 sg13g2_antennanp ANTENNA_2544 (.A(_07129_));
 sg13g2_antennanp ANTENNA_2545 (.A(_07150_));
 sg13g2_antennanp ANTENNA_2546 (.A(_07151_));
 sg13g2_antennanp ANTENNA_2547 (.A(_07157_));
 sg13g2_antennanp ANTENNA_2548 (.A(_07172_));
 sg13g2_antennanp ANTENNA_2549 (.A(_07188_));
 sg13g2_antennanp ANTENNA_2550 (.A(_07195_));
 sg13g2_antennanp ANTENNA_2551 (.A(_07201_));
 sg13g2_antennanp ANTENNA_2552 (.A(_07221_));
 sg13g2_antennanp ANTENNA_2553 (.A(_07222_));
 sg13g2_antennanp ANTENNA_2554 (.A(_07243_));
 sg13g2_antennanp ANTENNA_2555 (.A(_07269_));
 sg13g2_antennanp ANTENNA_2556 (.A(_07282_));
 sg13g2_antennanp ANTENNA_2557 (.A(_07344_));
 sg13g2_antennanp ANTENNA_2558 (.A(_07345_));
 sg13g2_antennanp ANTENNA_2559 (.A(_07371_));
 sg13g2_antennanp ANTENNA_2560 (.A(_07381_));
 sg13g2_antennanp ANTENNA_2561 (.A(_07385_));
 sg13g2_antennanp ANTENNA_2562 (.A(_07421_));
 sg13g2_antennanp ANTENNA_2563 (.A(_07429_));
 sg13g2_antennanp ANTENNA_2564 (.A(_07435_));
 sg13g2_antennanp ANTENNA_2565 (.A(_07440_));
 sg13g2_antennanp ANTENNA_2566 (.A(_07446_));
 sg13g2_antennanp ANTENNA_2567 (.A(_07480_));
 sg13g2_antennanp ANTENNA_2568 (.A(_07485_));
 sg13g2_antennanp ANTENNA_2569 (.A(_07507_));
 sg13g2_antennanp ANTENNA_2570 (.A(_07535_));
 sg13g2_antennanp ANTENNA_2571 (.A(_07540_));
 sg13g2_antennanp ANTENNA_2572 (.A(_07552_));
 sg13g2_antennanp ANTENNA_2573 (.A(_07560_));
 sg13g2_antennanp ANTENNA_2574 (.A(_07592_));
 sg13g2_antennanp ANTENNA_2575 (.A(_07592_));
 sg13g2_antennanp ANTENNA_2576 (.A(_07595_));
 sg13g2_antennanp ANTENNA_2577 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2578 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2579 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2580 (.A(_07601_));
 sg13g2_antennanp ANTENNA_2581 (.A(_07603_));
 sg13g2_antennanp ANTENNA_2582 (.A(_07634_));
 sg13g2_antennanp ANTENNA_2583 (.A(_07913_));
 sg13g2_antennanp ANTENNA_2584 (.A(_07945_));
 sg13g2_antennanp ANTENNA_2585 (.A(_07979_));
 sg13g2_antennanp ANTENNA_2586 (.A(_08062_));
 sg13g2_antennanp ANTENNA_2587 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2588 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2589 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2590 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2591 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2592 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2593 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2594 (.A(_08219_));
 sg13g2_antennanp ANTENNA_2595 (.A(_08223_));
 sg13g2_antennanp ANTENNA_2596 (.A(_08223_));
 sg13g2_antennanp ANTENNA_2597 (.A(_08223_));
 sg13g2_antennanp ANTENNA_2598 (.A(_08223_));
 sg13g2_antennanp ANTENNA_2599 (.A(_08227_));
 sg13g2_antennanp ANTENNA_2600 (.A(_08227_));
 sg13g2_antennanp ANTENNA_2601 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2602 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2603 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2604 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2605 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2606 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2607 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2608 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2609 (.A(_08260_));
 sg13g2_antennanp ANTENNA_2610 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2611 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2612 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2613 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2614 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2615 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2616 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2617 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2618 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2619 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2620 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2621 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2622 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2623 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2624 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2625 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2626 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2627 (.A(_08321_));
 sg13g2_antennanp ANTENNA_2628 (.A(_08380_));
 sg13g2_antennanp ANTENNA_2629 (.A(_08380_));
 sg13g2_antennanp ANTENNA_2630 (.A(_08380_));
 sg13g2_antennanp ANTENNA_2631 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2632 (.A(_08706_));
 sg13g2_antennanp ANTENNA_2633 (.A(_08730_));
 sg13g2_antennanp ANTENNA_2634 (.A(_08985_));
 sg13g2_antennanp ANTENNA_2635 (.A(_08985_));
 sg13g2_antennanp ANTENNA_2636 (.A(_08985_));
 sg13g2_antennanp ANTENNA_2637 (.A(_08985_));
 sg13g2_antennanp ANTENNA_2638 (.A(_08993_));
 sg13g2_antennanp ANTENNA_2639 (.A(_08993_));
 sg13g2_antennanp ANTENNA_2640 (.A(_08993_));
 sg13g2_antennanp ANTENNA_2641 (.A(_09940_));
 sg13g2_antennanp ANTENNA_2642 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2643 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2644 (.A(_10089_));
 sg13g2_antennanp ANTENNA_2645 (.A(_10158_));
 sg13g2_antennanp ANTENNA_2646 (.A(_10158_));
 sg13g2_antennanp ANTENNA_2647 (.A(_10158_));
 sg13g2_antennanp ANTENNA_2648 (.A(_10158_));
 sg13g2_antennanp ANTENNA_2649 (.A(_10159_));
 sg13g2_antennanp ANTENNA_2650 (.A(_10159_));
 sg13g2_antennanp ANTENNA_2651 (.A(_10159_));
 sg13g2_antennanp ANTENNA_2652 (.A(_10204_));
 sg13g2_antennanp ANTENNA_2653 (.A(_10318_));
 sg13g2_antennanp ANTENNA_2654 (.A(_10318_));
 sg13g2_antennanp ANTENNA_2655 (.A(_10318_));
 sg13g2_antennanp ANTENNA_2656 (.A(_10342_));
 sg13g2_antennanp ANTENNA_2657 (.A(_10342_));
 sg13g2_antennanp ANTENNA_2658 (.A(_10361_));
 sg13g2_antennanp ANTENNA_2659 (.A(_10361_));
 sg13g2_antennanp ANTENNA_2660 (.A(_10361_));
 sg13g2_antennanp ANTENNA_2661 (.A(_10361_));
 sg13g2_antennanp ANTENNA_2662 (.A(_10424_));
 sg13g2_antennanp ANTENNA_2663 (.A(_10424_));
 sg13g2_antennanp ANTENNA_2664 (.A(_10424_));
 sg13g2_antennanp ANTENNA_2665 (.A(_10424_));
 sg13g2_antennanp ANTENNA_2666 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2667 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2668 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2669 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2670 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2671 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2672 (.A(_10429_));
 sg13g2_antennanp ANTENNA_2673 (.A(_10450_));
 sg13g2_antennanp ANTENNA_2674 (.A(_10450_));
 sg13g2_antennanp ANTENNA_2675 (.A(_10450_));
 sg13g2_antennanp ANTENNA_2676 (.A(_10450_));
 sg13g2_antennanp ANTENNA_2677 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2678 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2679 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2680 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2681 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2682 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2683 (.A(_10535_));
 sg13g2_antennanp ANTENNA_2684 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2685 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2686 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2687 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2688 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2689 (.A(_10599_));
 sg13g2_antennanp ANTENNA_2690 (.A(_10600_));
 sg13g2_antennanp ANTENNA_2691 (.A(_10600_));
 sg13g2_antennanp ANTENNA_2692 (.A(_10600_));
 sg13g2_antennanp ANTENNA_2693 (.A(_10600_));
 sg13g2_antennanp ANTENNA_2694 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2695 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2696 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2697 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2698 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2699 (.A(_10704_));
 sg13g2_antennanp ANTENNA_2700 (.A(_10726_));
 sg13g2_antennanp ANTENNA_2701 (.A(_10726_));
 sg13g2_antennanp ANTENNA_2702 (.A(_10726_));
 sg13g2_antennanp ANTENNA_2703 (.A(_10739_));
 sg13g2_antennanp ANTENNA_2704 (.A(_10739_));
 sg13g2_antennanp ANTENNA_2705 (.A(_10739_));
 sg13g2_antennanp ANTENNA_2706 (.A(_10739_));
 sg13g2_antennanp ANTENNA_2707 (.A(_10740_));
 sg13g2_antennanp ANTENNA_2708 (.A(_10740_));
 sg13g2_antennanp ANTENNA_2709 (.A(_10740_));
 sg13g2_antennanp ANTENNA_2710 (.A(_10741_));
 sg13g2_antennanp ANTENNA_2711 (.A(_10741_));
 sg13g2_antennanp ANTENNA_2712 (.A(_10741_));
 sg13g2_antennanp ANTENNA_2713 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2714 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2715 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2716 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2717 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2718 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2719 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2720 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2721 (.A(_10742_));
 sg13g2_antennanp ANTENNA_2722 (.A(_10745_));
 sg13g2_antennanp ANTENNA_2723 (.A(_10745_));
 sg13g2_antennanp ANTENNA_2724 (.A(_10745_));
 sg13g2_antennanp ANTENNA_2725 (.A(_10779_));
 sg13g2_antennanp ANTENNA_2726 (.A(_10779_));
 sg13g2_antennanp ANTENNA_2727 (.A(_10779_));
 sg13g2_antennanp ANTENNA_2728 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2729 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2730 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2731 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2732 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2733 (.A(_10810_));
 sg13g2_antennanp ANTENNA_2734 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2735 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2736 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2737 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2738 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2739 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2740 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2741 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2742 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2743 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2744 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2745 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2746 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2747 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2748 (.A(_10812_));
 sg13g2_antennanp ANTENNA_2749 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2750 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2751 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2752 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2753 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2754 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2755 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2756 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2757 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2758 (.A(_10818_));
 sg13g2_antennanp ANTENNA_2759 (.A(_10845_));
 sg13g2_antennanp ANTENNA_2760 (.A(_10845_));
 sg13g2_antennanp ANTENNA_2761 (.A(_10845_));
 sg13g2_antennanp ANTENNA_2762 (.A(clk));
 sg13g2_antennanp ANTENNA_2763 (.A(clk));
 sg13g2_antennanp ANTENNA_2764 (.A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_antennanp ANTENNA_2765 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_2766 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_2767 (.A(\top_ihp.oisc.op_b[27] ));
 sg13g2_antennanp ANTENNA_2768 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_2769 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_2770 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_2771 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_2772 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2773 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2774 (.A(\top_ihp.oisc.regs[32][20] ));
 sg13g2_antennanp ANTENNA_2775 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_2776 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_2777 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_2778 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_2779 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_2780 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2781 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2782 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_2783 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_2784 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_2785 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_2786 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2787 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2788 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2789 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_2790 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2791 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2792 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2793 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_2794 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_2795 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_2796 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_2797 (.A(\top_ihp.oisc.regs[8][15] ));
 sg13g2_antennanp ANTENNA_2798 (.A(net56));
 sg13g2_antennanp ANTENNA_2799 (.A(net56));
 sg13g2_antennanp ANTENNA_2800 (.A(net56));
 sg13g2_antennanp ANTENNA_2801 (.A(net56));
 sg13g2_antennanp ANTENNA_2802 (.A(net56));
 sg13g2_antennanp ANTENNA_2803 (.A(net56));
 sg13g2_antennanp ANTENNA_2804 (.A(net56));
 sg13g2_antennanp ANTENNA_2805 (.A(net56));
 sg13g2_antennanp ANTENNA_2806 (.A(net56));
 sg13g2_antennanp ANTENNA_2807 (.A(net69));
 sg13g2_antennanp ANTENNA_2808 (.A(net69));
 sg13g2_antennanp ANTENNA_2809 (.A(net69));
 sg13g2_antennanp ANTENNA_2810 (.A(net69));
 sg13g2_antennanp ANTENNA_2811 (.A(net69));
 sg13g2_antennanp ANTENNA_2812 (.A(net69));
 sg13g2_antennanp ANTENNA_2813 (.A(net69));
 sg13g2_antennanp ANTENNA_2814 (.A(net69));
 sg13g2_antennanp ANTENNA_2815 (.A(net74));
 sg13g2_antennanp ANTENNA_2816 (.A(net74));
 sg13g2_antennanp ANTENNA_2817 (.A(net74));
 sg13g2_antennanp ANTENNA_2818 (.A(net74));
 sg13g2_antennanp ANTENNA_2819 (.A(net74));
 sg13g2_antennanp ANTENNA_2820 (.A(net74));
 sg13g2_antennanp ANTENNA_2821 (.A(net74));
 sg13g2_antennanp ANTENNA_2822 (.A(net74));
 sg13g2_antennanp ANTENNA_2823 (.A(net74));
 sg13g2_antennanp ANTENNA_2824 (.A(net74));
 sg13g2_antennanp ANTENNA_2825 (.A(net74));
 sg13g2_antennanp ANTENNA_2826 (.A(net74));
 sg13g2_antennanp ANTENNA_2827 (.A(net123));
 sg13g2_antennanp ANTENNA_2828 (.A(net123));
 sg13g2_antennanp ANTENNA_2829 (.A(net123));
 sg13g2_antennanp ANTENNA_2830 (.A(net123));
 sg13g2_antennanp ANTENNA_2831 (.A(net123));
 sg13g2_antennanp ANTENNA_2832 (.A(net123));
 sg13g2_antennanp ANTENNA_2833 (.A(net123));
 sg13g2_antennanp ANTENNA_2834 (.A(net123));
 sg13g2_antennanp ANTENNA_2835 (.A(net123));
 sg13g2_antennanp ANTENNA_2836 (.A(net127));
 sg13g2_antennanp ANTENNA_2837 (.A(net127));
 sg13g2_antennanp ANTENNA_2838 (.A(net127));
 sg13g2_antennanp ANTENNA_2839 (.A(net127));
 sg13g2_antennanp ANTENNA_2840 (.A(net127));
 sg13g2_antennanp ANTENNA_2841 (.A(net127));
 sg13g2_antennanp ANTENNA_2842 (.A(net127));
 sg13g2_antennanp ANTENNA_2843 (.A(net127));
 sg13g2_antennanp ANTENNA_2844 (.A(net127));
 sg13g2_antennanp ANTENNA_2845 (.A(net127));
 sg13g2_antennanp ANTENNA_2846 (.A(net127));
 sg13g2_antennanp ANTENNA_2847 (.A(net127));
 sg13g2_antennanp ANTENNA_2848 (.A(net127));
 sg13g2_antennanp ANTENNA_2849 (.A(net127));
 sg13g2_antennanp ANTENNA_2850 (.A(net127));
 sg13g2_antennanp ANTENNA_2851 (.A(net127));
 sg13g2_antennanp ANTENNA_2852 (.A(net127));
 sg13g2_antennanp ANTENNA_2853 (.A(net127));
 sg13g2_antennanp ANTENNA_2854 (.A(net127));
 sg13g2_antennanp ANTENNA_2855 (.A(net127));
 sg13g2_antennanp ANTENNA_2856 (.A(net127));
 sg13g2_antennanp ANTENNA_2857 (.A(net127));
 sg13g2_antennanp ANTENNA_2858 (.A(net127));
 sg13g2_antennanp ANTENNA_2859 (.A(net127));
 sg13g2_antennanp ANTENNA_2860 (.A(net127));
 sg13g2_antennanp ANTENNA_2861 (.A(net127));
 sg13g2_antennanp ANTENNA_2862 (.A(net127));
 sg13g2_antennanp ANTENNA_2863 (.A(net127));
 sg13g2_antennanp ANTENNA_2864 (.A(net127));
 sg13g2_antennanp ANTENNA_2865 (.A(net127));
 sg13g2_antennanp ANTENNA_2866 (.A(net127));
 sg13g2_antennanp ANTENNA_2867 (.A(net127));
 sg13g2_antennanp ANTENNA_2868 (.A(net127));
 sg13g2_antennanp ANTENNA_2869 (.A(net127));
 sg13g2_antennanp ANTENNA_2870 (.A(net127));
 sg13g2_antennanp ANTENNA_2871 (.A(net127));
 sg13g2_antennanp ANTENNA_2872 (.A(net127));
 sg13g2_antennanp ANTENNA_2873 (.A(net127));
 sg13g2_antennanp ANTENNA_2874 (.A(net127));
 sg13g2_antennanp ANTENNA_2875 (.A(net127));
 sg13g2_antennanp ANTENNA_2876 (.A(net127));
 sg13g2_antennanp ANTENNA_2877 (.A(net127));
 sg13g2_antennanp ANTENNA_2878 (.A(net127));
 sg13g2_antennanp ANTENNA_2879 (.A(net127));
 sg13g2_antennanp ANTENNA_2880 (.A(net127));
 sg13g2_antennanp ANTENNA_2881 (.A(net127));
 sg13g2_antennanp ANTENNA_2882 (.A(net127));
 sg13g2_antennanp ANTENNA_2883 (.A(net127));
 sg13g2_antennanp ANTENNA_2884 (.A(net127));
 sg13g2_antennanp ANTENNA_2885 (.A(net127));
 sg13g2_antennanp ANTENNA_2886 (.A(net127));
 sg13g2_antennanp ANTENNA_2887 (.A(net127));
 sg13g2_antennanp ANTENNA_2888 (.A(net127));
 sg13g2_antennanp ANTENNA_2889 (.A(net127));
 sg13g2_antennanp ANTENNA_2890 (.A(net127));
 sg13g2_antennanp ANTENNA_2891 (.A(net127));
 sg13g2_antennanp ANTENNA_2892 (.A(net127));
 sg13g2_antennanp ANTENNA_2893 (.A(net127));
 sg13g2_antennanp ANTENNA_2894 (.A(net127));
 sg13g2_antennanp ANTENNA_2895 (.A(net127));
 sg13g2_antennanp ANTENNA_2896 (.A(net127));
 sg13g2_antennanp ANTENNA_2897 (.A(net127));
 sg13g2_antennanp ANTENNA_2898 (.A(net127));
 sg13g2_antennanp ANTENNA_2899 (.A(net127));
 sg13g2_antennanp ANTENNA_2900 (.A(net127));
 sg13g2_antennanp ANTENNA_2901 (.A(net127));
 sg13g2_antennanp ANTENNA_2902 (.A(net127));
 sg13g2_antennanp ANTENNA_2903 (.A(net127));
 sg13g2_antennanp ANTENNA_2904 (.A(net127));
 sg13g2_antennanp ANTENNA_2905 (.A(net127));
 sg13g2_antennanp ANTENNA_2906 (.A(net127));
 sg13g2_antennanp ANTENNA_2907 (.A(net127));
 sg13g2_antennanp ANTENNA_2908 (.A(net127));
 sg13g2_antennanp ANTENNA_2909 (.A(net127));
 sg13g2_antennanp ANTENNA_2910 (.A(net127));
 sg13g2_antennanp ANTENNA_2911 (.A(net130));
 sg13g2_antennanp ANTENNA_2912 (.A(net130));
 sg13g2_antennanp ANTENNA_2913 (.A(net130));
 sg13g2_antennanp ANTENNA_2914 (.A(net130));
 sg13g2_antennanp ANTENNA_2915 (.A(net130));
 sg13g2_antennanp ANTENNA_2916 (.A(net130));
 sg13g2_antennanp ANTENNA_2917 (.A(net130));
 sg13g2_antennanp ANTENNA_2918 (.A(net130));
 sg13g2_antennanp ANTENNA_2919 (.A(net130));
 sg13g2_antennanp ANTENNA_2920 (.A(net130));
 sg13g2_antennanp ANTENNA_2921 (.A(net130));
 sg13g2_antennanp ANTENNA_2922 (.A(net130));
 sg13g2_antennanp ANTENNA_2923 (.A(net130));
 sg13g2_antennanp ANTENNA_2924 (.A(net130));
 sg13g2_antennanp ANTENNA_2925 (.A(net130));
 sg13g2_antennanp ANTENNA_2926 (.A(net130));
 sg13g2_antennanp ANTENNA_2927 (.A(net130));
 sg13g2_antennanp ANTENNA_2928 (.A(net130));
 sg13g2_antennanp ANTENNA_2929 (.A(net130));
 sg13g2_antennanp ANTENNA_2930 (.A(net130));
 sg13g2_antennanp ANTENNA_2931 (.A(net130));
 sg13g2_antennanp ANTENNA_2932 (.A(net130));
 sg13g2_antennanp ANTENNA_2933 (.A(net130));
 sg13g2_antennanp ANTENNA_2934 (.A(net132));
 sg13g2_antennanp ANTENNA_2935 (.A(net132));
 sg13g2_antennanp ANTENNA_2936 (.A(net132));
 sg13g2_antennanp ANTENNA_2937 (.A(net132));
 sg13g2_antennanp ANTENNA_2938 (.A(net132));
 sg13g2_antennanp ANTENNA_2939 (.A(net132));
 sg13g2_antennanp ANTENNA_2940 (.A(net132));
 sg13g2_antennanp ANTENNA_2941 (.A(net132));
 sg13g2_antennanp ANTENNA_2942 (.A(net132));
 sg13g2_antennanp ANTENNA_2943 (.A(net134));
 sg13g2_antennanp ANTENNA_2944 (.A(net134));
 sg13g2_antennanp ANTENNA_2945 (.A(net134));
 sg13g2_antennanp ANTENNA_2946 (.A(net134));
 sg13g2_antennanp ANTENNA_2947 (.A(net134));
 sg13g2_antennanp ANTENNA_2948 (.A(net134));
 sg13g2_antennanp ANTENNA_2949 (.A(net134));
 sg13g2_antennanp ANTENNA_2950 (.A(net134));
 sg13g2_antennanp ANTENNA_2951 (.A(net134));
 sg13g2_antennanp ANTENNA_2952 (.A(net134));
 sg13g2_antennanp ANTENNA_2953 (.A(net134));
 sg13g2_antennanp ANTENNA_2954 (.A(net134));
 sg13g2_antennanp ANTENNA_2955 (.A(net134));
 sg13g2_antennanp ANTENNA_2956 (.A(net134));
 sg13g2_antennanp ANTENNA_2957 (.A(net134));
 sg13g2_antennanp ANTENNA_2958 (.A(net134));
 sg13g2_antennanp ANTENNA_2959 (.A(net134));
 sg13g2_antennanp ANTENNA_2960 (.A(net134));
 sg13g2_antennanp ANTENNA_2961 (.A(net134));
 sg13g2_antennanp ANTENNA_2962 (.A(net134));
 sg13g2_antennanp ANTENNA_2963 (.A(net143));
 sg13g2_antennanp ANTENNA_2964 (.A(net143));
 sg13g2_antennanp ANTENNA_2965 (.A(net143));
 sg13g2_antennanp ANTENNA_2966 (.A(net143));
 sg13g2_antennanp ANTENNA_2967 (.A(net143));
 sg13g2_antennanp ANTENNA_2968 (.A(net143));
 sg13g2_antennanp ANTENNA_2969 (.A(net143));
 sg13g2_antennanp ANTENNA_2970 (.A(net143));
 sg13g2_antennanp ANTENNA_2971 (.A(net143));
 sg13g2_antennanp ANTENNA_2972 (.A(net159));
 sg13g2_antennanp ANTENNA_2973 (.A(net159));
 sg13g2_antennanp ANTENNA_2974 (.A(net159));
 sg13g2_antennanp ANTENNA_2975 (.A(net159));
 sg13g2_antennanp ANTENNA_2976 (.A(net159));
 sg13g2_antennanp ANTENNA_2977 (.A(net159));
 sg13g2_antennanp ANTENNA_2978 (.A(net159));
 sg13g2_antennanp ANTENNA_2979 (.A(net159));
 sg13g2_antennanp ANTENNA_2980 (.A(net159));
 sg13g2_antennanp ANTENNA_2981 (.A(net177));
 sg13g2_antennanp ANTENNA_2982 (.A(net177));
 sg13g2_antennanp ANTENNA_2983 (.A(net177));
 sg13g2_antennanp ANTENNA_2984 (.A(net177));
 sg13g2_antennanp ANTENNA_2985 (.A(net177));
 sg13g2_antennanp ANTENNA_2986 (.A(net177));
 sg13g2_antennanp ANTENNA_2987 (.A(net177));
 sg13g2_antennanp ANTENNA_2988 (.A(net177));
 sg13g2_antennanp ANTENNA_2989 (.A(net177));
 sg13g2_antennanp ANTENNA_2990 (.A(net263));
 sg13g2_antennanp ANTENNA_2991 (.A(net263));
 sg13g2_antennanp ANTENNA_2992 (.A(net263));
 sg13g2_antennanp ANTENNA_2993 (.A(net263));
 sg13g2_antennanp ANTENNA_2994 (.A(net263));
 sg13g2_antennanp ANTENNA_2995 (.A(net263));
 sg13g2_antennanp ANTENNA_2996 (.A(net263));
 sg13g2_antennanp ANTENNA_2997 (.A(net263));
 sg13g2_antennanp ANTENNA_2998 (.A(net264));
 sg13g2_antennanp ANTENNA_2999 (.A(net264));
 sg13g2_antennanp ANTENNA_3000 (.A(net264));
 sg13g2_antennanp ANTENNA_3001 (.A(net264));
 sg13g2_antennanp ANTENNA_3002 (.A(net264));
 sg13g2_antennanp ANTENNA_3003 (.A(net264));
 sg13g2_antennanp ANTENNA_3004 (.A(net264));
 sg13g2_antennanp ANTENNA_3005 (.A(net264));
 sg13g2_antennanp ANTENNA_3006 (.A(net264));
 sg13g2_antennanp ANTENNA_3007 (.A(net314));
 sg13g2_antennanp ANTENNA_3008 (.A(net314));
 sg13g2_antennanp ANTENNA_3009 (.A(net314));
 sg13g2_antennanp ANTENNA_3010 (.A(net314));
 sg13g2_antennanp ANTENNA_3011 (.A(net314));
 sg13g2_antennanp ANTENNA_3012 (.A(net314));
 sg13g2_antennanp ANTENNA_3013 (.A(net314));
 sg13g2_antennanp ANTENNA_3014 (.A(net314));
 sg13g2_antennanp ANTENNA_3015 (.A(net323));
 sg13g2_antennanp ANTENNA_3016 (.A(net323));
 sg13g2_antennanp ANTENNA_3017 (.A(net323));
 sg13g2_antennanp ANTENNA_3018 (.A(net323));
 sg13g2_antennanp ANTENNA_3019 (.A(net323));
 sg13g2_antennanp ANTENNA_3020 (.A(net323));
 sg13g2_antennanp ANTENNA_3021 (.A(net323));
 sg13g2_antennanp ANTENNA_3022 (.A(net323));
 sg13g2_antennanp ANTENNA_3023 (.A(net323));
 sg13g2_antennanp ANTENNA_3024 (.A(net326));
 sg13g2_antennanp ANTENNA_3025 (.A(net326));
 sg13g2_antennanp ANTENNA_3026 (.A(net326));
 sg13g2_antennanp ANTENNA_3027 (.A(net326));
 sg13g2_antennanp ANTENNA_3028 (.A(net326));
 sg13g2_antennanp ANTENNA_3029 (.A(net326));
 sg13g2_antennanp ANTENNA_3030 (.A(net326));
 sg13g2_antennanp ANTENNA_3031 (.A(net326));
 sg13g2_antennanp ANTENNA_3032 (.A(net372));
 sg13g2_antennanp ANTENNA_3033 (.A(net372));
 sg13g2_antennanp ANTENNA_3034 (.A(net372));
 sg13g2_antennanp ANTENNA_3035 (.A(net372));
 sg13g2_antennanp ANTENNA_3036 (.A(net372));
 sg13g2_antennanp ANTENNA_3037 (.A(net372));
 sg13g2_antennanp ANTENNA_3038 (.A(net372));
 sg13g2_antennanp ANTENNA_3039 (.A(net372));
 sg13g2_antennanp ANTENNA_3040 (.A(net403));
 sg13g2_antennanp ANTENNA_3041 (.A(net403));
 sg13g2_antennanp ANTENNA_3042 (.A(net403));
 sg13g2_antennanp ANTENNA_3043 (.A(net403));
 sg13g2_antennanp ANTENNA_3044 (.A(net403));
 sg13g2_antennanp ANTENNA_3045 (.A(net403));
 sg13g2_antennanp ANTENNA_3046 (.A(net403));
 sg13g2_antennanp ANTENNA_3047 (.A(net403));
 sg13g2_antennanp ANTENNA_3048 (.A(net403));
 sg13g2_antennanp ANTENNA_3049 (.A(net435));
 sg13g2_antennanp ANTENNA_3050 (.A(net435));
 sg13g2_antennanp ANTENNA_3051 (.A(net435));
 sg13g2_antennanp ANTENNA_3052 (.A(net435));
 sg13g2_antennanp ANTENNA_3053 (.A(net435));
 sg13g2_antennanp ANTENNA_3054 (.A(net435));
 sg13g2_antennanp ANTENNA_3055 (.A(net435));
 sg13g2_antennanp ANTENNA_3056 (.A(net435));
 sg13g2_antennanp ANTENNA_3057 (.A(net435));
 sg13g2_antennanp ANTENNA_3058 (.A(net444));
 sg13g2_antennanp ANTENNA_3059 (.A(net444));
 sg13g2_antennanp ANTENNA_3060 (.A(net444));
 sg13g2_antennanp ANTENNA_3061 (.A(net444));
 sg13g2_antennanp ANTENNA_3062 (.A(net444));
 sg13g2_antennanp ANTENNA_3063 (.A(net444));
 sg13g2_antennanp ANTENNA_3064 (.A(net444));
 sg13g2_antennanp ANTENNA_3065 (.A(net444));
 sg13g2_antennanp ANTENNA_3066 (.A(net444));
 sg13g2_antennanp ANTENNA_3067 (.A(net444));
 sg13g2_antennanp ANTENNA_3068 (.A(net444));
 sg13g2_antennanp ANTENNA_3069 (.A(net444));
 sg13g2_antennanp ANTENNA_3070 (.A(net444));
 sg13g2_antennanp ANTENNA_3071 (.A(net444));
 sg13g2_antennanp ANTENNA_3072 (.A(net444));
 sg13g2_antennanp ANTENNA_3073 (.A(net444));
 sg13g2_antennanp ANTENNA_3074 (.A(net444));
 sg13g2_antennanp ANTENNA_3075 (.A(net444));
 sg13g2_antennanp ANTENNA_3076 (.A(net444));
 sg13g2_antennanp ANTENNA_3077 (.A(net444));
 sg13g2_antennanp ANTENNA_3078 (.A(net444));
 sg13g2_antennanp ANTENNA_3079 (.A(net444));
 sg13g2_antennanp ANTENNA_3080 (.A(net444));
 sg13g2_antennanp ANTENNA_3081 (.A(net449));
 sg13g2_antennanp ANTENNA_3082 (.A(net449));
 sg13g2_antennanp ANTENNA_3083 (.A(net449));
 sg13g2_antennanp ANTENNA_3084 (.A(net449));
 sg13g2_antennanp ANTENNA_3085 (.A(net449));
 sg13g2_antennanp ANTENNA_3086 (.A(net449));
 sg13g2_antennanp ANTENNA_3087 (.A(net449));
 sg13g2_antennanp ANTENNA_3088 (.A(net449));
 sg13g2_antennanp ANTENNA_3089 (.A(net487));
 sg13g2_antennanp ANTENNA_3090 (.A(net487));
 sg13g2_antennanp ANTENNA_3091 (.A(net487));
 sg13g2_antennanp ANTENNA_3092 (.A(net487));
 sg13g2_antennanp ANTENNA_3093 (.A(net487));
 sg13g2_antennanp ANTENNA_3094 (.A(net487));
 sg13g2_antennanp ANTENNA_3095 (.A(net487));
 sg13g2_antennanp ANTENNA_3096 (.A(net487));
 sg13g2_antennanp ANTENNA_3097 (.A(net487));
 sg13g2_antennanp ANTENNA_3098 (.A(net1421));
 sg13g2_antennanp ANTENNA_3099 (.A(net1421));
 sg13g2_antennanp ANTENNA_3100 (.A(net1421));
 sg13g2_antennanp ANTENNA_3101 (.A(net1421));
 sg13g2_antennanp ANTENNA_3102 (.A(net1421));
 sg13g2_antennanp ANTENNA_3103 (.A(net1421));
 sg13g2_antennanp ANTENNA_3104 (.A(net1421));
 sg13g2_antennanp ANTENNA_3105 (.A(net1421));
 sg13g2_antennanp ANTENNA_3106 (.A(net1421));
 sg13g2_antennanp ANTENNA_3107 (.A(net1421));
 sg13g2_antennanp ANTENNA_3108 (.A(net1421));
 sg13g2_antennanp ANTENNA_3109 (.A(net1421));
 sg13g2_antennanp ANTENNA_3110 (.A(net1421));
 sg13g2_antennanp ANTENNA_3111 (.A(net1421));
 sg13g2_antennanp ANTENNA_3112 (.A(net1421));
 sg13g2_antennanp ANTENNA_3113 (.A(net1421));
 sg13g2_antennanp ANTENNA_3114 (.A(net1421));
 sg13g2_antennanp ANTENNA_3115 (.A(net1421));
 sg13g2_antennanp ANTENNA_3116 (.A(net1421));
 sg13g2_antennanp ANTENNA_3117 (.A(net1421));
 sg13g2_antennanp ANTENNA_3118 (.A(net1421));
 sg13g2_antennanp ANTENNA_3119 (.A(net1421));
 sg13g2_antennanp ANTENNA_3120 (.A(net1421));
 sg13g2_antennanp ANTENNA_3121 (.A(_00356_));
 sg13g2_antennanp ANTENNA_3122 (.A(_00410_));
 sg13g2_antennanp ANTENNA_3123 (.A(_00422_));
 sg13g2_antennanp ANTENNA_3124 (.A(_00425_));
 sg13g2_antennanp ANTENNA_3125 (.A(_00432_));
 sg13g2_antennanp ANTENNA_3126 (.A(_02799_));
 sg13g2_antennanp ANTENNA_3127 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3128 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3129 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3130 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3131 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3132 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3133 (.A(_03714_));
 sg13g2_antennanp ANTENNA_3134 (.A(_03714_));
 sg13g2_antennanp ANTENNA_3135 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3136 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3137 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3138 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3139 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3140 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3141 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3142 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3143 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3144 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3145 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3146 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3147 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3148 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3149 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3150 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3151 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3152 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3153 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3154 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3155 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3156 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3157 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3158 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3159 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3160 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3161 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3162 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3163 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3164 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3165 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3166 (.A(_04620_));
 sg13g2_antennanp ANTENNA_3167 (.A(_04674_));
 sg13g2_antennanp ANTENNA_3168 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3169 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3170 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3171 (.A(_05061_));
 sg13g2_antennanp ANTENNA_3172 (.A(_05067_));
 sg13g2_antennanp ANTENNA_3173 (.A(_05091_));
 sg13g2_antennanp ANTENNA_3174 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3175 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3176 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3177 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3178 (.A(_05278_));
 sg13g2_antennanp ANTENNA_3179 (.A(_05290_));
 sg13g2_antennanp ANTENNA_3180 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3181 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3182 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3183 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3184 (.A(_05318_));
 sg13g2_antennanp ANTENNA_3185 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3186 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3187 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3188 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3189 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3190 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3191 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3192 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3193 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3194 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3195 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3196 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3197 (.A(_05350_));
 sg13g2_antennanp ANTENNA_3198 (.A(_05364_));
 sg13g2_antennanp ANTENNA_3199 (.A(_05432_));
 sg13g2_antennanp ANTENNA_3200 (.A(_05512_));
 sg13g2_antennanp ANTENNA_3201 (.A(_05577_));
 sg13g2_antennanp ANTENNA_3202 (.A(_05584_));
 sg13g2_antennanp ANTENNA_3203 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3204 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3205 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3206 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3207 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3208 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3209 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3210 (.A(_05672_));
 sg13g2_antennanp ANTENNA_3211 (.A(_05754_));
 sg13g2_antennanp ANTENNA_3212 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3213 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3214 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3215 (.A(_05788_));
 sg13g2_antennanp ANTENNA_3216 (.A(_05788_));
 sg13g2_antennanp ANTENNA_3217 (.A(_05788_));
 sg13g2_antennanp ANTENNA_3218 (.A(_05788_));
 sg13g2_antennanp ANTENNA_3219 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3220 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3221 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3222 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3223 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3224 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3225 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3226 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3227 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3228 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3229 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3230 (.A(_05851_));
 sg13g2_antennanp ANTENNA_3231 (.A(_05868_));
 sg13g2_antennanp ANTENNA_3232 (.A(_05872_));
 sg13g2_antennanp ANTENNA_3233 (.A(_05892_));
 sg13g2_antennanp ANTENNA_3234 (.A(_05892_));
 sg13g2_antennanp ANTENNA_3235 (.A(_05892_));
 sg13g2_antennanp ANTENNA_3236 (.A(_05892_));
 sg13g2_antennanp ANTENNA_3237 (.A(_05892_));
 sg13g2_antennanp ANTENNA_3238 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3239 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3240 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3241 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3242 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3243 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3244 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3245 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3246 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3247 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3248 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3249 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3250 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3251 (.A(_05936_));
 sg13g2_antennanp ANTENNA_3252 (.A(_05940_));
 sg13g2_antennanp ANTENNA_3253 (.A(_05953_));
 sg13g2_antennanp ANTENNA_3254 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3255 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3256 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3257 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3258 (.A(_06027_));
 sg13g2_antennanp ANTENNA_3259 (.A(_06090_));
 sg13g2_antennanp ANTENNA_3260 (.A(_06101_));
 sg13g2_antennanp ANTENNA_3261 (.A(_06167_));
 sg13g2_antennanp ANTENNA_3262 (.A(_06184_));
 sg13g2_antennanp ANTENNA_3263 (.A(_06214_));
 sg13g2_antennanp ANTENNA_3264 (.A(_06244_));
 sg13g2_antennanp ANTENNA_3265 (.A(_06254_));
 sg13g2_antennanp ANTENNA_3266 (.A(_06255_));
 sg13g2_antennanp ANTENNA_3267 (.A(_06265_));
 sg13g2_antennanp ANTENNA_3268 (.A(_06302_));
 sg13g2_antennanp ANTENNA_3269 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3270 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3271 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3272 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3273 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3274 (.A(_06330_));
 sg13g2_antennanp ANTENNA_3275 (.A(_06345_));
 sg13g2_antennanp ANTENNA_3276 (.A(_06345_));
 sg13g2_antennanp ANTENNA_3277 (.A(_06351_));
 sg13g2_antennanp ANTENNA_3278 (.A(_06351_));
 sg13g2_antennanp ANTENNA_3279 (.A(_06351_));
 sg13g2_antennanp ANTENNA_3280 (.A(_06359_));
 sg13g2_antennanp ANTENNA_3281 (.A(_06359_));
 sg13g2_antennanp ANTENNA_3282 (.A(_06440_));
 sg13g2_antennanp ANTENNA_3283 (.A(_06443_));
 sg13g2_antennanp ANTENNA_3284 (.A(_06447_));
 sg13g2_antennanp ANTENNA_3285 (.A(_06489_));
 sg13g2_antennanp ANTENNA_3286 (.A(_06489_));
 sg13g2_antennanp ANTENNA_3287 (.A(_06530_));
 sg13g2_antennanp ANTENNA_3288 (.A(_06533_));
 sg13g2_antennanp ANTENNA_3289 (.A(_06538_));
 sg13g2_antennanp ANTENNA_3290 (.A(_06545_));
 sg13g2_antennanp ANTENNA_3291 (.A(_06587_));
 sg13g2_antennanp ANTENNA_3292 (.A(_06591_));
 sg13g2_antennanp ANTENNA_3293 (.A(_06591_));
 sg13g2_antennanp ANTENNA_3294 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3295 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3296 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3297 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3298 (.A(_06603_));
 sg13g2_antennanp ANTENNA_3299 (.A(_06603_));
 sg13g2_antennanp ANTENNA_3300 (.A(_06609_));
 sg13g2_antennanp ANTENNA_3301 (.A(_06619_));
 sg13g2_antennanp ANTENNA_3302 (.A(_06651_));
 sg13g2_antennanp ANTENNA_3303 (.A(_06654_));
 sg13g2_antennanp ANTENNA_3304 (.A(_06662_));
 sg13g2_antennanp ANTENNA_3305 (.A(_06671_));
 sg13g2_antennanp ANTENNA_3306 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3307 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3308 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3309 (.A(_06716_));
 sg13g2_antennanp ANTENNA_3310 (.A(_06721_));
 sg13g2_antennanp ANTENNA_3311 (.A(_06722_));
 sg13g2_antennanp ANTENNA_3312 (.A(_06735_));
 sg13g2_antennanp ANTENNA_3313 (.A(_06740_));
 sg13g2_antennanp ANTENNA_3314 (.A(_06741_));
 sg13g2_antennanp ANTENNA_3315 (.A(_06751_));
 sg13g2_antennanp ANTENNA_3316 (.A(_06780_));
 sg13g2_antennanp ANTENNA_3317 (.A(_06792_));
 sg13g2_antennanp ANTENNA_3318 (.A(_06793_));
 sg13g2_antennanp ANTENNA_3319 (.A(_06807_));
 sg13g2_antennanp ANTENNA_3320 (.A(_06838_));
 sg13g2_antennanp ANTENNA_3321 (.A(_06853_));
 sg13g2_antennanp ANTENNA_3322 (.A(_06874_));
 sg13g2_antennanp ANTENNA_3323 (.A(_06875_));
 sg13g2_antennanp ANTENNA_3324 (.A(_06902_));
 sg13g2_antennanp ANTENNA_3325 (.A(_06945_));
 sg13g2_antennanp ANTENNA_3326 (.A(_06963_));
 sg13g2_antennanp ANTENNA_3327 (.A(_06980_));
 sg13g2_antennanp ANTENNA_3328 (.A(_06980_));
 sg13g2_antennanp ANTENNA_3329 (.A(_06980_));
 sg13g2_antennanp ANTENNA_3330 (.A(_06981_));
 sg13g2_antennanp ANTENNA_3331 (.A(_06985_));
 sg13g2_antennanp ANTENNA_3332 (.A(_07020_));
 sg13g2_antennanp ANTENNA_3333 (.A(_07032_));
 sg13g2_antennanp ANTENNA_3334 (.A(_07063_));
 sg13g2_antennanp ANTENNA_3335 (.A(_07064_));
 sg13g2_antennanp ANTENNA_3336 (.A(_07064_));
 sg13g2_antennanp ANTENNA_3337 (.A(_07073_));
 sg13g2_antennanp ANTENNA_3338 (.A(_07074_));
 sg13g2_antennanp ANTENNA_3339 (.A(_07077_));
 sg13g2_antennanp ANTENNA_3340 (.A(_07085_));
 sg13g2_antennanp ANTENNA_3341 (.A(_07104_));
 sg13g2_antennanp ANTENNA_3342 (.A(_07113_));
 sg13g2_antennanp ANTENNA_3343 (.A(_07125_));
 sg13g2_antennanp ANTENNA_3344 (.A(_07129_));
 sg13g2_antennanp ANTENNA_3345 (.A(_07150_));
 sg13g2_antennanp ANTENNA_3346 (.A(_07151_));
 sg13g2_antennanp ANTENNA_3347 (.A(_07157_));
 sg13g2_antennanp ANTENNA_3348 (.A(_07172_));
 sg13g2_antennanp ANTENNA_3349 (.A(_07188_));
 sg13g2_antennanp ANTENNA_3350 (.A(_07195_));
 sg13g2_antennanp ANTENNA_3351 (.A(_07201_));
 sg13g2_antennanp ANTENNA_3352 (.A(_07221_));
 sg13g2_antennanp ANTENNA_3353 (.A(_07222_));
 sg13g2_antennanp ANTENNA_3354 (.A(_07243_));
 sg13g2_antennanp ANTENNA_3355 (.A(_07269_));
 sg13g2_antennanp ANTENNA_3356 (.A(_07279_));
 sg13g2_antennanp ANTENNA_3357 (.A(_07282_));
 sg13g2_antennanp ANTENNA_3358 (.A(_07344_));
 sg13g2_antennanp ANTENNA_3359 (.A(_07345_));
 sg13g2_antennanp ANTENNA_3360 (.A(_07371_));
 sg13g2_antennanp ANTENNA_3361 (.A(_07381_));
 sg13g2_antennanp ANTENNA_3362 (.A(_07385_));
 sg13g2_antennanp ANTENNA_3363 (.A(_07429_));
 sg13g2_antennanp ANTENNA_3364 (.A(_07435_));
 sg13g2_antennanp ANTENNA_3365 (.A(_07440_));
 sg13g2_antennanp ANTENNA_3366 (.A(_07446_));
 sg13g2_antennanp ANTENNA_3367 (.A(_07485_));
 sg13g2_antennanp ANTENNA_3368 (.A(_07507_));
 sg13g2_antennanp ANTENNA_3369 (.A(_07535_));
 sg13g2_antennanp ANTENNA_3370 (.A(_07540_));
 sg13g2_antennanp ANTENNA_3371 (.A(_07544_));
 sg13g2_antennanp ANTENNA_3372 (.A(_07552_));
 sg13g2_antennanp ANTENNA_3373 (.A(_07560_));
 sg13g2_antennanp ANTENNA_3374 (.A(_07592_));
 sg13g2_antennanp ANTENNA_3375 (.A(_07595_));
 sg13g2_antennanp ANTENNA_3376 (.A(_07601_));
 sg13g2_antennanp ANTENNA_3377 (.A(_07601_));
 sg13g2_antennanp ANTENNA_3378 (.A(_07601_));
 sg13g2_antennanp ANTENNA_3379 (.A(_07601_));
 sg13g2_antennanp ANTENNA_3380 (.A(_07603_));
 sg13g2_antennanp ANTENNA_3381 (.A(_07634_));
 sg13g2_antennanp ANTENNA_3382 (.A(_07913_));
 sg13g2_antennanp ANTENNA_3383 (.A(_07945_));
 sg13g2_antennanp ANTENNA_3384 (.A(_07979_));
 sg13g2_antennanp ANTENNA_3385 (.A(_08062_));
 sg13g2_antennanp ANTENNA_3386 (.A(_08227_));
 sg13g2_antennanp ANTENNA_3387 (.A(_08227_));
 sg13g2_antennanp ANTENNA_3388 (.A(_08227_));
 sg13g2_antennanp ANTENNA_3389 (.A(_08227_));
 sg13g2_antennanp ANTENNA_3390 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3391 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3392 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3393 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3394 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3395 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3396 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3397 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3398 (.A(_08260_));
 sg13g2_antennanp ANTENNA_3399 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3400 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3401 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3402 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3403 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3404 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3405 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3406 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3407 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3408 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3409 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3410 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3411 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3412 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3413 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3414 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3415 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3416 (.A(_08321_));
 sg13g2_antennanp ANTENNA_3417 (.A(_08380_));
 sg13g2_antennanp ANTENNA_3418 (.A(_08380_));
 sg13g2_antennanp ANTENNA_3419 (.A(_08380_));
 sg13g2_antennanp ANTENNA_3420 (.A(_08380_));
 sg13g2_antennanp ANTENNA_3421 (.A(_08706_));
 sg13g2_antennanp ANTENNA_3422 (.A(_08706_));
 sg13g2_antennanp ANTENNA_3423 (.A(_08730_));
 sg13g2_antennanp ANTENNA_3424 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3425 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3426 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3427 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3428 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3429 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3430 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3431 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3432 (.A(_08985_));
 sg13g2_antennanp ANTENNA_3433 (.A(_08993_));
 sg13g2_antennanp ANTENNA_3434 (.A(_08993_));
 sg13g2_antennanp ANTENNA_3435 (.A(_08993_));
 sg13g2_antennanp ANTENNA_3436 (.A(_09940_));
 sg13g2_antennanp ANTENNA_3437 (.A(_10089_));
 sg13g2_antennanp ANTENNA_3438 (.A(_10089_));
 sg13g2_antennanp ANTENNA_3439 (.A(_10089_));
 sg13g2_antennanp ANTENNA_3440 (.A(_10158_));
 sg13g2_antennanp ANTENNA_3441 (.A(_10158_));
 sg13g2_antennanp ANTENNA_3442 (.A(_10158_));
 sg13g2_antennanp ANTENNA_3443 (.A(_10158_));
 sg13g2_antennanp ANTENNA_3444 (.A(_10204_));
 sg13g2_antennanp ANTENNA_3445 (.A(_10342_));
 sg13g2_antennanp ANTENNA_3446 (.A(_10342_));
 sg13g2_antennanp ANTENNA_3447 (.A(_10361_));
 sg13g2_antennanp ANTENNA_3448 (.A(_10361_));
 sg13g2_antennanp ANTENNA_3449 (.A(_10361_));
 sg13g2_antennanp ANTENNA_3450 (.A(_10361_));
 sg13g2_antennanp ANTENNA_3451 (.A(_10361_));
 sg13g2_antennanp ANTENNA_3452 (.A(_10424_));
 sg13g2_antennanp ANTENNA_3453 (.A(_10424_));
 sg13g2_antennanp ANTENNA_3454 (.A(_10424_));
 sg13g2_antennanp ANTENNA_3455 (.A(_10424_));
 sg13g2_antennanp ANTENNA_3456 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3457 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3458 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3459 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3460 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3461 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3462 (.A(_10429_));
 sg13g2_antennanp ANTENNA_3463 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3464 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3465 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3466 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3467 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3468 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3469 (.A(_10535_));
 sg13g2_antennanp ANTENNA_3470 (.A(_10600_));
 sg13g2_antennanp ANTENNA_3471 (.A(_10600_));
 sg13g2_antennanp ANTENNA_3472 (.A(_10600_));
 sg13g2_antennanp ANTENNA_3473 (.A(_10600_));
 sg13g2_antennanp ANTENNA_3474 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3475 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3476 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3477 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3478 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3479 (.A(_10704_));
 sg13g2_antennanp ANTENNA_3480 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3481 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3482 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3483 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3484 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3485 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3486 (.A(_10739_));
 sg13g2_antennanp ANTENNA_3487 (.A(_10740_));
 sg13g2_antennanp ANTENNA_3488 (.A(_10740_));
 sg13g2_antennanp ANTENNA_3489 (.A(_10740_));
 sg13g2_antennanp ANTENNA_3490 (.A(_10741_));
 sg13g2_antennanp ANTENNA_3491 (.A(_10741_));
 sg13g2_antennanp ANTENNA_3492 (.A(_10741_));
 sg13g2_antennanp ANTENNA_3493 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3494 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3495 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3496 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3497 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3498 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3499 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3500 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3501 (.A(_10742_));
 sg13g2_antennanp ANTENNA_3502 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3503 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3504 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3505 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3506 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3507 (.A(_10745_));
 sg13g2_antennanp ANTENNA_3508 (.A(_10779_));
 sg13g2_antennanp ANTENNA_3509 (.A(_10779_));
 sg13g2_antennanp ANTENNA_3510 (.A(_10779_));
 sg13g2_antennanp ANTENNA_3511 (.A(_10804_));
 sg13g2_antennanp ANTENNA_3512 (.A(_10804_));
 sg13g2_antennanp ANTENNA_3513 (.A(_10804_));
 sg13g2_antennanp ANTENNA_3514 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3515 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3516 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3517 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3518 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3519 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3520 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3521 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3522 (.A(_10810_));
 sg13g2_antennanp ANTENNA_3523 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3524 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3525 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3526 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3527 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3528 (.A(_10812_));
 sg13g2_antennanp ANTENNA_3529 (.A(_10818_));
 sg13g2_antennanp ANTENNA_3530 (.A(_10818_));
 sg13g2_antennanp ANTENNA_3531 (.A(_10818_));
 sg13g2_antennanp ANTENNA_3532 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3533 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3534 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3535 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3536 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3537 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3538 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3539 (.A(_10845_));
 sg13g2_antennanp ANTENNA_3540 (.A(clk));
 sg13g2_antennanp ANTENNA_3541 (.A(clk));
 sg13g2_antennanp ANTENNA_3542 (.A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_antennanp ANTENNA_3543 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_3544 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_3545 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_3546 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_3547 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_3548 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_3549 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_3550 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_3551 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_3552 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_3553 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_3554 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_3555 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_3556 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_3557 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3558 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3559 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3560 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_3561 (.A(net54));
 sg13g2_antennanp ANTENNA_3562 (.A(net54));
 sg13g2_antennanp ANTENNA_3563 (.A(net54));
 sg13g2_antennanp ANTENNA_3564 (.A(net54));
 sg13g2_antennanp ANTENNA_3565 (.A(net54));
 sg13g2_antennanp ANTENNA_3566 (.A(net54));
 sg13g2_antennanp ANTENNA_3567 (.A(net54));
 sg13g2_antennanp ANTENNA_3568 (.A(net54));
 sg13g2_antennanp ANTENNA_3569 (.A(net54));
 sg13g2_antennanp ANTENNA_3570 (.A(net56));
 sg13g2_antennanp ANTENNA_3571 (.A(net56));
 sg13g2_antennanp ANTENNA_3572 (.A(net56));
 sg13g2_antennanp ANTENNA_3573 (.A(net56));
 sg13g2_antennanp ANTENNA_3574 (.A(net56));
 sg13g2_antennanp ANTENNA_3575 (.A(net56));
 sg13g2_antennanp ANTENNA_3576 (.A(net56));
 sg13g2_antennanp ANTENNA_3577 (.A(net56));
 sg13g2_antennanp ANTENNA_3578 (.A(net56));
 sg13g2_antennanp ANTENNA_3579 (.A(net117));
 sg13g2_antennanp ANTENNA_3580 (.A(net117));
 sg13g2_antennanp ANTENNA_3581 (.A(net117));
 sg13g2_antennanp ANTENNA_3582 (.A(net117));
 sg13g2_antennanp ANTENNA_3583 (.A(net117));
 sg13g2_antennanp ANTENNA_3584 (.A(net117));
 sg13g2_antennanp ANTENNA_3585 (.A(net117));
 sg13g2_antennanp ANTENNA_3586 (.A(net117));
 sg13g2_antennanp ANTENNA_3587 (.A(net117));
 sg13g2_antennanp ANTENNA_3588 (.A(net117));
 sg13g2_antennanp ANTENNA_3589 (.A(net117));
 sg13g2_antennanp ANTENNA_3590 (.A(net117));
 sg13g2_antennanp ANTENNA_3591 (.A(net117));
 sg13g2_antennanp ANTENNA_3592 (.A(net117));
 sg13g2_antennanp ANTENNA_3593 (.A(net117));
 sg13g2_antennanp ANTENNA_3594 (.A(net117));
 sg13g2_antennanp ANTENNA_3595 (.A(net117));
 sg13g2_antennanp ANTENNA_3596 (.A(net117));
 sg13g2_antennanp ANTENNA_3597 (.A(net117));
 sg13g2_antennanp ANTENNA_3598 (.A(net117));
 sg13g2_antennanp ANTENNA_3599 (.A(net123));
 sg13g2_antennanp ANTENNA_3600 (.A(net123));
 sg13g2_antennanp ANTENNA_3601 (.A(net123));
 sg13g2_antennanp ANTENNA_3602 (.A(net123));
 sg13g2_antennanp ANTENNA_3603 (.A(net123));
 sg13g2_antennanp ANTENNA_3604 (.A(net123));
 sg13g2_antennanp ANTENNA_3605 (.A(net123));
 sg13g2_antennanp ANTENNA_3606 (.A(net123));
 sg13g2_antennanp ANTENNA_3607 (.A(net123));
 sg13g2_antennanp ANTENNA_3608 (.A(net127));
 sg13g2_antennanp ANTENNA_3609 (.A(net127));
 sg13g2_antennanp ANTENNA_3610 (.A(net127));
 sg13g2_antennanp ANTENNA_3611 (.A(net127));
 sg13g2_antennanp ANTENNA_3612 (.A(net127));
 sg13g2_antennanp ANTENNA_3613 (.A(net127));
 sg13g2_antennanp ANTENNA_3614 (.A(net127));
 sg13g2_antennanp ANTENNA_3615 (.A(net127));
 sg13g2_antennanp ANTENNA_3616 (.A(net130));
 sg13g2_antennanp ANTENNA_3617 (.A(net130));
 sg13g2_antennanp ANTENNA_3618 (.A(net130));
 sg13g2_antennanp ANTENNA_3619 (.A(net130));
 sg13g2_antennanp ANTENNA_3620 (.A(net130));
 sg13g2_antennanp ANTENNA_3621 (.A(net130));
 sg13g2_antennanp ANTENNA_3622 (.A(net130));
 sg13g2_antennanp ANTENNA_3623 (.A(net130));
 sg13g2_antennanp ANTENNA_3624 (.A(net130));
 sg13g2_antennanp ANTENNA_3625 (.A(net130));
 sg13g2_antennanp ANTENNA_3626 (.A(net130));
 sg13g2_antennanp ANTENNA_3627 (.A(net130));
 sg13g2_antennanp ANTENNA_3628 (.A(net130));
 sg13g2_antennanp ANTENNA_3629 (.A(net130));
 sg13g2_antennanp ANTENNA_3630 (.A(net130));
 sg13g2_antennanp ANTENNA_3631 (.A(net130));
 sg13g2_antennanp ANTENNA_3632 (.A(net130));
 sg13g2_antennanp ANTENNA_3633 (.A(net130));
 sg13g2_antennanp ANTENNA_3634 (.A(net130));
 sg13g2_antennanp ANTENNA_3635 (.A(net130));
 sg13g2_antennanp ANTENNA_3636 (.A(net130));
 sg13g2_antennanp ANTENNA_3637 (.A(net130));
 sg13g2_antennanp ANTENNA_3638 (.A(net130));
 sg13g2_antennanp ANTENNA_3639 (.A(net130));
 sg13g2_antennanp ANTENNA_3640 (.A(net132));
 sg13g2_antennanp ANTENNA_3641 (.A(net132));
 sg13g2_antennanp ANTENNA_3642 (.A(net132));
 sg13g2_antennanp ANTENNA_3643 (.A(net132));
 sg13g2_antennanp ANTENNA_3644 (.A(net132));
 sg13g2_antennanp ANTENNA_3645 (.A(net132));
 sg13g2_antennanp ANTENNA_3646 (.A(net132));
 sg13g2_antennanp ANTENNA_3647 (.A(net132));
 sg13g2_antennanp ANTENNA_3648 (.A(net132));
 sg13g2_antennanp ANTENNA_3649 (.A(net134));
 sg13g2_antennanp ANTENNA_3650 (.A(net134));
 sg13g2_antennanp ANTENNA_3651 (.A(net134));
 sg13g2_antennanp ANTENNA_3652 (.A(net134));
 sg13g2_antennanp ANTENNA_3653 (.A(net134));
 sg13g2_antennanp ANTENNA_3654 (.A(net134));
 sg13g2_antennanp ANTENNA_3655 (.A(net134));
 sg13g2_antennanp ANTENNA_3656 (.A(net134));
 sg13g2_antennanp ANTENNA_3657 (.A(net134));
 sg13g2_antennanp ANTENNA_3658 (.A(net134));
 sg13g2_antennanp ANTENNA_3659 (.A(net134));
 sg13g2_antennanp ANTENNA_3660 (.A(net134));
 sg13g2_antennanp ANTENNA_3661 (.A(net134));
 sg13g2_antennanp ANTENNA_3662 (.A(net134));
 sg13g2_antennanp ANTENNA_3663 (.A(net134));
 sg13g2_antennanp ANTENNA_3664 (.A(net134));
 sg13g2_antennanp ANTENNA_3665 (.A(net134));
 sg13g2_antennanp ANTENNA_3666 (.A(net134));
 sg13g2_antennanp ANTENNA_3667 (.A(net134));
 sg13g2_antennanp ANTENNA_3668 (.A(net134));
 sg13g2_antennanp ANTENNA_3669 (.A(net143));
 sg13g2_antennanp ANTENNA_3670 (.A(net143));
 sg13g2_antennanp ANTENNA_3671 (.A(net143));
 sg13g2_antennanp ANTENNA_3672 (.A(net143));
 sg13g2_antennanp ANTENNA_3673 (.A(net143));
 sg13g2_antennanp ANTENNA_3674 (.A(net143));
 sg13g2_antennanp ANTENNA_3675 (.A(net143));
 sg13g2_antennanp ANTENNA_3676 (.A(net143));
 sg13g2_antennanp ANTENNA_3677 (.A(net143));
 sg13g2_antennanp ANTENNA_3678 (.A(net159));
 sg13g2_antennanp ANTENNA_3679 (.A(net159));
 sg13g2_antennanp ANTENNA_3680 (.A(net159));
 sg13g2_antennanp ANTENNA_3681 (.A(net159));
 sg13g2_antennanp ANTENNA_3682 (.A(net159));
 sg13g2_antennanp ANTENNA_3683 (.A(net159));
 sg13g2_antennanp ANTENNA_3684 (.A(net159));
 sg13g2_antennanp ANTENNA_3685 (.A(net159));
 sg13g2_antennanp ANTENNA_3686 (.A(net177));
 sg13g2_antennanp ANTENNA_3687 (.A(net177));
 sg13g2_antennanp ANTENNA_3688 (.A(net177));
 sg13g2_antennanp ANTENNA_3689 (.A(net177));
 sg13g2_antennanp ANTENNA_3690 (.A(net177));
 sg13g2_antennanp ANTENNA_3691 (.A(net177));
 sg13g2_antennanp ANTENNA_3692 (.A(net177));
 sg13g2_antennanp ANTENNA_3693 (.A(net177));
 sg13g2_antennanp ANTENNA_3694 (.A(net177));
 sg13g2_antennanp ANTENNA_3695 (.A(net264));
 sg13g2_antennanp ANTENNA_3696 (.A(net264));
 sg13g2_antennanp ANTENNA_3697 (.A(net264));
 sg13g2_antennanp ANTENNA_3698 (.A(net264));
 sg13g2_antennanp ANTENNA_3699 (.A(net264));
 sg13g2_antennanp ANTENNA_3700 (.A(net264));
 sg13g2_antennanp ANTENNA_3701 (.A(net264));
 sg13g2_antennanp ANTENNA_3702 (.A(net264));
 sg13g2_antennanp ANTENNA_3703 (.A(net264));
 sg13g2_antennanp ANTENNA_3704 (.A(net274));
 sg13g2_antennanp ANTENNA_3705 (.A(net274));
 sg13g2_antennanp ANTENNA_3706 (.A(net274));
 sg13g2_antennanp ANTENNA_3707 (.A(net274));
 sg13g2_antennanp ANTENNA_3708 (.A(net274));
 sg13g2_antennanp ANTENNA_3709 (.A(net274));
 sg13g2_antennanp ANTENNA_3710 (.A(net274));
 sg13g2_antennanp ANTENNA_3711 (.A(net274));
 sg13g2_antennanp ANTENNA_3712 (.A(net274));
 sg13g2_antennanp ANTENNA_3713 (.A(net274));
 sg13g2_antennanp ANTENNA_3714 (.A(net314));
 sg13g2_antennanp ANTENNA_3715 (.A(net314));
 sg13g2_antennanp ANTENNA_3716 (.A(net314));
 sg13g2_antennanp ANTENNA_3717 (.A(net314));
 sg13g2_antennanp ANTENNA_3718 (.A(net314));
 sg13g2_antennanp ANTENNA_3719 (.A(net314));
 sg13g2_antennanp ANTENNA_3720 (.A(net314));
 sg13g2_antennanp ANTENNA_3721 (.A(net314));
 sg13g2_antennanp ANTENNA_3722 (.A(net323));
 sg13g2_antennanp ANTENNA_3723 (.A(net323));
 sg13g2_antennanp ANTENNA_3724 (.A(net323));
 sg13g2_antennanp ANTENNA_3725 (.A(net323));
 sg13g2_antennanp ANTENNA_3726 (.A(net323));
 sg13g2_antennanp ANTENNA_3727 (.A(net323));
 sg13g2_antennanp ANTENNA_3728 (.A(net323));
 sg13g2_antennanp ANTENNA_3729 (.A(net323));
 sg13g2_antennanp ANTENNA_3730 (.A(net323));
 sg13g2_antennanp ANTENNA_3731 (.A(net323));
 sg13g2_antennanp ANTENNA_3732 (.A(net323));
 sg13g2_antennanp ANTENNA_3733 (.A(net323));
 sg13g2_antennanp ANTENNA_3734 (.A(net323));
 sg13g2_antennanp ANTENNA_3735 (.A(net323));
 sg13g2_antennanp ANTENNA_3736 (.A(net323));
 sg13g2_antennanp ANTENNA_3737 (.A(net323));
 sg13g2_antennanp ANTENNA_3738 (.A(net326));
 sg13g2_antennanp ANTENNA_3739 (.A(net326));
 sg13g2_antennanp ANTENNA_3740 (.A(net326));
 sg13g2_antennanp ANTENNA_3741 (.A(net326));
 sg13g2_antennanp ANTENNA_3742 (.A(net326));
 sg13g2_antennanp ANTENNA_3743 (.A(net326));
 sg13g2_antennanp ANTENNA_3744 (.A(net326));
 sg13g2_antennanp ANTENNA_3745 (.A(net326));
 sg13g2_antennanp ANTENNA_3746 (.A(net403));
 sg13g2_antennanp ANTENNA_3747 (.A(net403));
 sg13g2_antennanp ANTENNA_3748 (.A(net403));
 sg13g2_antennanp ANTENNA_3749 (.A(net403));
 sg13g2_antennanp ANTENNA_3750 (.A(net403));
 sg13g2_antennanp ANTENNA_3751 (.A(net403));
 sg13g2_antennanp ANTENNA_3752 (.A(net403));
 sg13g2_antennanp ANTENNA_3753 (.A(net403));
 sg13g2_antennanp ANTENNA_3754 (.A(net403));
 sg13g2_antennanp ANTENNA_3755 (.A(net403));
 sg13g2_antennanp ANTENNA_3756 (.A(net403));
 sg13g2_antennanp ANTENNA_3757 (.A(net403));
 sg13g2_antennanp ANTENNA_3758 (.A(net403));
 sg13g2_antennanp ANTENNA_3759 (.A(net403));
 sg13g2_antennanp ANTENNA_3760 (.A(net403));
 sg13g2_antennanp ANTENNA_3761 (.A(net403));
 sg13g2_antennanp ANTENNA_3762 (.A(net403));
 sg13g2_antennanp ANTENNA_3763 (.A(net403));
 sg13g2_antennanp ANTENNA_3764 (.A(net403));
 sg13g2_antennanp ANTENNA_3765 (.A(net403));
 sg13g2_antennanp ANTENNA_3766 (.A(net435));
 sg13g2_antennanp ANTENNA_3767 (.A(net435));
 sg13g2_antennanp ANTENNA_3768 (.A(net435));
 sg13g2_antennanp ANTENNA_3769 (.A(net435));
 sg13g2_antennanp ANTENNA_3770 (.A(net435));
 sg13g2_antennanp ANTENNA_3771 (.A(net435));
 sg13g2_antennanp ANTENNA_3772 (.A(net435));
 sg13g2_antennanp ANTENNA_3773 (.A(net435));
 sg13g2_antennanp ANTENNA_3774 (.A(net435));
 sg13g2_antennanp ANTENNA_3775 (.A(net444));
 sg13g2_antennanp ANTENNA_3776 (.A(net444));
 sg13g2_antennanp ANTENNA_3777 (.A(net444));
 sg13g2_antennanp ANTENNA_3778 (.A(net444));
 sg13g2_antennanp ANTENNA_3779 (.A(net444));
 sg13g2_antennanp ANTENNA_3780 (.A(net444));
 sg13g2_antennanp ANTENNA_3781 (.A(net444));
 sg13g2_antennanp ANTENNA_3782 (.A(net444));
 sg13g2_antennanp ANTENNA_3783 (.A(net444));
 sg13g2_antennanp ANTENNA_3784 (.A(net605));
 sg13g2_antennanp ANTENNA_3785 (.A(net605));
 sg13g2_antennanp ANTENNA_3786 (.A(net605));
 sg13g2_antennanp ANTENNA_3787 (.A(net605));
 sg13g2_antennanp ANTENNA_3788 (.A(net605));
 sg13g2_antennanp ANTENNA_3789 (.A(net605));
 sg13g2_antennanp ANTENNA_3790 (.A(net605));
 sg13g2_antennanp ANTENNA_3791 (.A(net605));
 sg13g2_antennanp ANTENNA_3792 (.A(net1421));
 sg13g2_antennanp ANTENNA_3793 (.A(net1421));
 sg13g2_antennanp ANTENNA_3794 (.A(net1421));
 sg13g2_antennanp ANTENNA_3795 (.A(net1421));
 sg13g2_antennanp ANTENNA_3796 (.A(net1421));
 sg13g2_antennanp ANTENNA_3797 (.A(net1421));
 sg13g2_antennanp ANTENNA_3798 (.A(net1421));
 sg13g2_antennanp ANTENNA_3799 (.A(net1421));
 sg13g2_antennanp ANTENNA_3800 (.A(net1421));
 sg13g2_antennanp ANTENNA_3801 (.A(net1421));
 sg13g2_antennanp ANTENNA_3802 (.A(net1421));
 sg13g2_antennanp ANTENNA_3803 (.A(net1421));
 sg13g2_antennanp ANTENNA_3804 (.A(net1421));
 sg13g2_antennanp ANTENNA_3805 (.A(net1421));
 sg13g2_antennanp ANTENNA_3806 (.A(net1421));
 sg13g2_antennanp ANTENNA_3807 (.A(net1421));
 sg13g2_antennanp ANTENNA_3808 (.A(net1421));
 sg13g2_antennanp ANTENNA_3809 (.A(net1421));
 sg13g2_antennanp ANTENNA_3810 (.A(net1421));
 sg13g2_antennanp ANTENNA_3811 (.A(net1421));
 sg13g2_antennanp ANTENNA_3812 (.A(net1421));
 sg13g2_antennanp ANTENNA_3813 (.A(net1421));
 sg13g2_antennanp ANTENNA_3814 (.A(net1421));
 sg13g2_antennanp ANTENNA_3815 (.A(net1421));
 sg13g2_antennanp ANTENNA_3816 (.A(net1421));
 sg13g2_antennanp ANTENNA_3817 (.A(net1421));
 sg13g2_antennanp ANTENNA_3818 (.A(net1421));
 sg13g2_antennanp ANTENNA_3819 (.A(_00356_));
 sg13g2_antennanp ANTENNA_3820 (.A(_00410_));
 sg13g2_antennanp ANTENNA_3821 (.A(_00422_));
 sg13g2_antennanp ANTENNA_3822 (.A(_00425_));
 sg13g2_antennanp ANTENNA_3823 (.A(_00432_));
 sg13g2_antennanp ANTENNA_3824 (.A(_02799_));
 sg13g2_antennanp ANTENNA_3825 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3826 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3827 (.A(_03060_));
 sg13g2_antennanp ANTENNA_3828 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3829 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3830 (.A(_03268_));
 sg13g2_antennanp ANTENNA_3831 (.A(_03714_));
 sg13g2_antennanp ANTENNA_3832 (.A(_03714_));
 sg13g2_antennanp ANTENNA_3833 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3834 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3835 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3836 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3837 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3838 (.A(_03760_));
 sg13g2_antennanp ANTENNA_3839 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3840 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3841 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3842 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3843 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3844 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3845 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3846 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3847 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3848 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3849 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3850 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3851 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3852 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3853 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3854 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3855 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3856 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3857 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3858 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3859 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3860 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3861 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3862 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3863 (.A(_04617_));
 sg13g2_antennanp ANTENNA_3864 (.A(_04620_));
 sg13g2_antennanp ANTENNA_3865 (.A(_04674_));
 sg13g2_antennanp ANTENNA_3866 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3867 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3868 (.A(_04676_));
 sg13g2_antennanp ANTENNA_3869 (.A(_05061_));
 sg13g2_antennanp ANTENNA_3870 (.A(_05067_));
 sg13g2_antennanp ANTENNA_3871 (.A(_05091_));
 sg13g2_antennanp ANTENNA_3872 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3873 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3874 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3875 (.A(_05276_));
 sg13g2_antennanp ANTENNA_3876 (.A(_05278_));
 sg13g2_antennanp ANTENNA_3877 (.A(_05290_));
 sg13g2_antennanp ANTENNA_3878 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3879 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3880 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3881 (.A(_05303_));
 sg13g2_antennanp ANTENNA_3882 (.A(_05318_));
 sg13g2_antennanp ANTENNA_3883 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3884 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3885 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3886 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3887 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3888 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3889 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3890 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3891 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3892 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3893 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3894 (.A(_05347_));
 sg13g2_antennanp ANTENNA_3895 (.A(_05350_));
 sg13g2_antennanp ANTENNA_3896 (.A(_05364_));
 sg13g2_antennanp ANTENNA_3897 (.A(_05432_));
 sg13g2_antennanp ANTENNA_3898 (.A(_05512_));
 sg13g2_antennanp ANTENNA_3899 (.A(_05577_));
 sg13g2_antennanp ANTENNA_3900 (.A(_05584_));
 sg13g2_antennanp ANTENNA_3901 (.A(_05600_));
 sg13g2_antennanp ANTENNA_3902 (.A(_05600_));
 sg13g2_antennanp ANTENNA_3903 (.A(_05600_));
 sg13g2_antennanp ANTENNA_3904 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3905 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3906 (.A(_05652_));
 sg13g2_antennanp ANTENNA_3907 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3908 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3909 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3910 (.A(_05662_));
 sg13g2_antennanp ANTENNA_3911 (.A(_05672_));
 sg13g2_antennanp ANTENNA_3912 (.A(_05754_));
 sg13g2_antennanp ANTENNA_3913 (.A(_05778_));
 sg13g2_antennanp ANTENNA_3914 (.A(_05778_));
 sg13g2_antennanp ANTENNA_3915 (.A(_05778_));
 sg13g2_antennanp ANTENNA_3916 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3917 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3918 (.A(_05784_));
 sg13g2_antennanp ANTENNA_3919 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3920 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3921 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3922 (.A(_05811_));
 sg13g2_antennanp ANTENNA_3923 (.A(_05868_));
 sg13g2_antennanp ANTENNA_3924 (.A(_05872_));
 sg13g2_antennanp ANTENNA_3925 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3926 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3927 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3928 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3929 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3930 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3931 (.A(_05901_));
 sg13g2_antennanp ANTENNA_3932 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3933 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3934 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3935 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3936 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3937 (.A(_05932_));
 sg13g2_antennanp ANTENNA_3938 (.A(_05936_));
 sg13g2_antennanp ANTENNA_3939 (.A(_05940_));
 sg13g2_antennanp ANTENNA_3940 (.A(_05953_));
 sg13g2_antennanp ANTENNA_3941 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3942 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3943 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3944 (.A(_06009_));
 sg13g2_antennanp ANTENNA_3945 (.A(_06027_));
 sg13g2_antennanp ANTENNA_3946 (.A(_06076_));
 sg13g2_antennanp ANTENNA_3947 (.A(_06101_));
 sg13g2_antennanp ANTENNA_3948 (.A(_06167_));
 sg13g2_antennanp ANTENNA_3949 (.A(_06184_));
 sg13g2_antennanp ANTENNA_3950 (.A(_06214_));
 sg13g2_antennanp ANTENNA_3951 (.A(_06244_));
 sg13g2_antennanp ANTENNA_3952 (.A(_06254_));
 sg13g2_antennanp ANTENNA_3953 (.A(_06255_));
 sg13g2_antennanp ANTENNA_3954 (.A(_06265_));
 sg13g2_antennanp ANTENNA_3955 (.A(_06302_));
 sg13g2_antennanp ANTENNA_3956 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3957 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3958 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3959 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3960 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3961 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3962 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3963 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3964 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3965 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3966 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3967 (.A(_06313_));
 sg13g2_antennanp ANTENNA_3968 (.A(_06330_));
 sg13g2_antennanp ANTENNA_3969 (.A(_06345_));
 sg13g2_antennanp ANTENNA_3970 (.A(_06351_));
 sg13g2_antennanp ANTENNA_3971 (.A(_06359_));
 sg13g2_antennanp ANTENNA_3972 (.A(_06440_));
 sg13g2_antennanp ANTENNA_3973 (.A(_06443_));
 sg13g2_antennanp ANTENNA_3974 (.A(_06447_));
 sg13g2_antennanp ANTENNA_3975 (.A(_06489_));
 sg13g2_antennanp ANTENNA_3976 (.A(_06530_));
 sg13g2_antennanp ANTENNA_3977 (.A(_06533_));
 sg13g2_antennanp ANTENNA_3978 (.A(_06538_));
 sg13g2_antennanp ANTENNA_3979 (.A(_06545_));
 sg13g2_antennanp ANTENNA_3980 (.A(_06545_));
 sg13g2_antennanp ANTENNA_3981 (.A(_06587_));
 sg13g2_antennanp ANTENNA_3982 (.A(_06591_));
 sg13g2_antennanp ANTENNA_3983 (.A(_06591_));
 sg13g2_antennanp ANTENNA_3984 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3985 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3986 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3987 (.A(_06601_));
 sg13g2_antennanp ANTENNA_3988 (.A(_06603_));
 sg13g2_antennanp ANTENNA_3989 (.A(_06609_));
 sg13g2_antennanp ANTENNA_3990 (.A(_06619_));
 sg13g2_antennanp ANTENNA_3991 (.A(_06651_));
 sg13g2_antennanp ANTENNA_3992 (.A(_06654_));
 sg13g2_antennanp ANTENNA_3993 (.A(_06662_));
 sg13g2_antennanp ANTENNA_3994 (.A(_06671_));
 sg13g2_antennanp ANTENNA_3995 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3996 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3997 (.A(_06708_));
 sg13g2_antennanp ANTENNA_3998 (.A(_06716_));
 sg13g2_antennanp ANTENNA_3999 (.A(_06721_));
 sg13g2_antennanp ANTENNA_4000 (.A(_06722_));
 sg13g2_antennanp ANTENNA_4001 (.A(_06735_));
 sg13g2_antennanp ANTENNA_4002 (.A(_06740_));
 sg13g2_antennanp ANTENNA_4003 (.A(_06741_));
 sg13g2_antennanp ANTENNA_4004 (.A(_06751_));
 sg13g2_antennanp ANTENNA_4005 (.A(_06780_));
 sg13g2_antennanp ANTENNA_4006 (.A(_06792_));
 sg13g2_antennanp ANTENNA_4007 (.A(_06793_));
 sg13g2_antennanp ANTENNA_4008 (.A(_06807_));
 sg13g2_antennanp ANTENNA_4009 (.A(_06838_));
 sg13g2_antennanp ANTENNA_4010 (.A(_06853_));
 sg13g2_antennanp ANTENNA_4011 (.A(_06874_));
 sg13g2_antennanp ANTENNA_4012 (.A(_06875_));
 sg13g2_antennanp ANTENNA_4013 (.A(_06902_));
 sg13g2_antennanp ANTENNA_4014 (.A(_06945_));
 sg13g2_antennanp ANTENNA_4015 (.A(_06963_));
 sg13g2_antennanp ANTENNA_4016 (.A(_06980_));
 sg13g2_antennanp ANTENNA_4017 (.A(_06980_));
 sg13g2_antennanp ANTENNA_4018 (.A(_06980_));
 sg13g2_antennanp ANTENNA_4019 (.A(_06980_));
 sg13g2_antennanp ANTENNA_4020 (.A(_06981_));
 sg13g2_antennanp ANTENNA_4021 (.A(_06985_));
 sg13g2_antennanp ANTENNA_4022 (.A(_07020_));
 sg13g2_antennanp ANTENNA_4023 (.A(_07032_));
 sg13g2_antennanp ANTENNA_4024 (.A(_07063_));
 sg13g2_antennanp ANTENNA_4025 (.A(_07064_));
 sg13g2_antennanp ANTENNA_4026 (.A(_07064_));
 sg13g2_antennanp ANTENNA_4027 (.A(_07073_));
 sg13g2_antennanp ANTENNA_4028 (.A(_07074_));
 sg13g2_antennanp ANTENNA_4029 (.A(_07077_));
 sg13g2_antennanp ANTENNA_4030 (.A(_07085_));
 sg13g2_antennanp ANTENNA_4031 (.A(_07104_));
 sg13g2_antennanp ANTENNA_4032 (.A(_07113_));
 sg13g2_antennanp ANTENNA_4033 (.A(_07125_));
 sg13g2_antennanp ANTENNA_4034 (.A(_07129_));
 sg13g2_antennanp ANTENNA_4035 (.A(_07150_));
 sg13g2_antennanp ANTENNA_4036 (.A(_07151_));
 sg13g2_antennanp ANTENNA_4037 (.A(_07151_));
 sg13g2_antennanp ANTENNA_4038 (.A(_07157_));
 sg13g2_antennanp ANTENNA_4039 (.A(_07172_));
 sg13g2_antennanp ANTENNA_4040 (.A(_07188_));
 sg13g2_antennanp ANTENNA_4041 (.A(_07195_));
 sg13g2_antennanp ANTENNA_4042 (.A(_07201_));
 sg13g2_antennanp ANTENNA_4043 (.A(_07221_));
 sg13g2_antennanp ANTENNA_4044 (.A(_07222_));
 sg13g2_antennanp ANTENNA_4045 (.A(_07243_));
 sg13g2_antennanp ANTENNA_4046 (.A(_07243_));
 sg13g2_antennanp ANTENNA_4047 (.A(_07269_));
 sg13g2_antennanp ANTENNA_4048 (.A(_07282_));
 sg13g2_antennanp ANTENNA_4049 (.A(_07344_));
 sg13g2_antennanp ANTENNA_4050 (.A(_07371_));
 sg13g2_antennanp ANTENNA_4051 (.A(_07381_));
 sg13g2_antennanp ANTENNA_4052 (.A(_07385_));
 sg13g2_antennanp ANTENNA_4053 (.A(_07421_));
 sg13g2_antennanp ANTENNA_4054 (.A(_07429_));
 sg13g2_antennanp ANTENNA_4055 (.A(_07429_));
 sg13g2_antennanp ANTENNA_4056 (.A(_07435_));
 sg13g2_antennanp ANTENNA_4057 (.A(_07435_));
 sg13g2_antennanp ANTENNA_4058 (.A(_07440_));
 sg13g2_antennanp ANTENNA_4059 (.A(_07446_));
 sg13g2_antennanp ANTENNA_4060 (.A(_07485_));
 sg13g2_antennanp ANTENNA_4061 (.A(_07507_));
 sg13g2_antennanp ANTENNA_4062 (.A(_07535_));
 sg13g2_antennanp ANTENNA_4063 (.A(_07535_));
 sg13g2_antennanp ANTENNA_4064 (.A(_07540_));
 sg13g2_antennanp ANTENNA_4065 (.A(_07552_));
 sg13g2_antennanp ANTENNA_4066 (.A(_07560_));
 sg13g2_antennanp ANTENNA_4067 (.A(_07592_));
 sg13g2_antennanp ANTENNA_4068 (.A(_07595_));
 sg13g2_antennanp ANTENNA_4069 (.A(_07601_));
 sg13g2_antennanp ANTENNA_4070 (.A(_07601_));
 sg13g2_antennanp ANTENNA_4071 (.A(_07601_));
 sg13g2_antennanp ANTENNA_4072 (.A(_07601_));
 sg13g2_antennanp ANTENNA_4073 (.A(_07603_));
 sg13g2_antennanp ANTENNA_4074 (.A(_07634_));
 sg13g2_antennanp ANTENNA_4075 (.A(_07913_));
 sg13g2_antennanp ANTENNA_4076 (.A(_07945_));
 sg13g2_antennanp ANTENNA_4077 (.A(_07945_));
 sg13g2_antennanp ANTENNA_4078 (.A(_07979_));
 sg13g2_antennanp ANTENNA_4079 (.A(_08062_));
 sg13g2_antennanp ANTENNA_4080 (.A(_08227_));
 sg13g2_antennanp ANTENNA_4081 (.A(_08227_));
 sg13g2_antennanp ANTENNA_4082 (.A(_08227_));
 sg13g2_antennanp ANTENNA_4083 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4084 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4085 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4086 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4087 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4088 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4089 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4090 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4091 (.A(_08260_));
 sg13g2_antennanp ANTENNA_4092 (.A(_08261_));
 sg13g2_antennanp ANTENNA_4093 (.A(_08261_));
 sg13g2_antennanp ANTENNA_4094 (.A(_08261_));
 sg13g2_antennanp ANTENNA_4095 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4096 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4097 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4098 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4099 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4100 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4101 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4102 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4103 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4104 (.A(_08263_));
 sg13g2_antennanp ANTENNA_4105 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4106 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4107 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4108 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4109 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4110 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4111 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4112 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4113 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4114 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4115 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4116 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4117 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4118 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4119 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4120 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4121 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4122 (.A(_08321_));
 sg13g2_antennanp ANTENNA_4123 (.A(_08380_));
 sg13g2_antennanp ANTENNA_4124 (.A(_08380_));
 sg13g2_antennanp ANTENNA_4125 (.A(_08380_));
 sg13g2_antennanp ANTENNA_4126 (.A(_08380_));
 sg13g2_antennanp ANTENNA_4127 (.A(_08706_));
 sg13g2_antennanp ANTENNA_4128 (.A(_08730_));
 sg13g2_antennanp ANTENNA_4129 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4130 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4131 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4132 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4133 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4134 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4135 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4136 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4137 (.A(_08985_));
 sg13g2_antennanp ANTENNA_4138 (.A(_08993_));
 sg13g2_antennanp ANTENNA_4139 (.A(_08993_));
 sg13g2_antennanp ANTENNA_4140 (.A(_08993_));
 sg13g2_antennanp ANTENNA_4141 (.A(_09940_));
 sg13g2_antennanp ANTENNA_4142 (.A(_10089_));
 sg13g2_antennanp ANTENNA_4143 (.A(_10089_));
 sg13g2_antennanp ANTENNA_4144 (.A(_10089_));
 sg13g2_antennanp ANTENNA_4145 (.A(_10158_));
 sg13g2_antennanp ANTENNA_4146 (.A(_10158_));
 sg13g2_antennanp ANTENNA_4147 (.A(_10158_));
 sg13g2_antennanp ANTENNA_4148 (.A(_10158_));
 sg13g2_antennanp ANTENNA_4149 (.A(_10204_));
 sg13g2_antennanp ANTENNA_4150 (.A(_10342_));
 sg13g2_antennanp ANTENNA_4151 (.A(_10342_));
 sg13g2_antennanp ANTENNA_4152 (.A(_10361_));
 sg13g2_antennanp ANTENNA_4153 (.A(_10361_));
 sg13g2_antennanp ANTENNA_4154 (.A(_10361_));
 sg13g2_antennanp ANTENNA_4155 (.A(_10361_));
 sg13g2_antennanp ANTENNA_4156 (.A(_10361_));
 sg13g2_antennanp ANTENNA_4157 (.A(_10424_));
 sg13g2_antennanp ANTENNA_4158 (.A(_10424_));
 sg13g2_antennanp ANTENNA_4159 (.A(_10424_));
 sg13g2_antennanp ANTENNA_4160 (.A(_10424_));
 sg13g2_antennanp ANTENNA_4161 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4162 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4163 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4164 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4165 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4166 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4167 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4168 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4169 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4170 (.A(_10429_));
 sg13g2_antennanp ANTENNA_4171 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4172 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4173 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4174 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4175 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4176 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4177 (.A(_10535_));
 sg13g2_antennanp ANTENNA_4178 (.A(_10599_));
 sg13g2_antennanp ANTENNA_4179 (.A(_10599_));
 sg13g2_antennanp ANTENNA_4180 (.A(_10599_));
 sg13g2_antennanp ANTENNA_4181 (.A(_10600_));
 sg13g2_antennanp ANTENNA_4182 (.A(_10600_));
 sg13g2_antennanp ANTENNA_4183 (.A(_10600_));
 sg13g2_antennanp ANTENNA_4184 (.A(_10600_));
 sg13g2_antennanp ANTENNA_4185 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4186 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4187 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4188 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4189 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4190 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4191 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4192 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4193 (.A(_10704_));
 sg13g2_antennanp ANTENNA_4194 (.A(_10739_));
 sg13g2_antennanp ANTENNA_4195 (.A(_10739_));
 sg13g2_antennanp ANTENNA_4196 (.A(_10739_));
 sg13g2_antennanp ANTENNA_4197 (.A(_10739_));
 sg13g2_antennanp ANTENNA_4198 (.A(_10740_));
 sg13g2_antennanp ANTENNA_4199 (.A(_10740_));
 sg13g2_antennanp ANTENNA_4200 (.A(_10740_));
 sg13g2_antennanp ANTENNA_4201 (.A(_10741_));
 sg13g2_antennanp ANTENNA_4202 (.A(_10741_));
 sg13g2_antennanp ANTENNA_4203 (.A(_10741_));
 sg13g2_antennanp ANTENNA_4204 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4205 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4206 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4207 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4208 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4209 (.A(_10742_));
 sg13g2_antennanp ANTENNA_4210 (.A(_10779_));
 sg13g2_antennanp ANTENNA_4211 (.A(_10779_));
 sg13g2_antennanp ANTENNA_4212 (.A(_10779_));
 sg13g2_antennanp ANTENNA_4213 (.A(_10804_));
 sg13g2_antennanp ANTENNA_4214 (.A(_10804_));
 sg13g2_antennanp ANTENNA_4215 (.A(_10804_));
 sg13g2_antennanp ANTENNA_4216 (.A(_10810_));
 sg13g2_antennanp ANTENNA_4217 (.A(_10810_));
 sg13g2_antennanp ANTENNA_4218 (.A(_10810_));
 sg13g2_antennanp ANTENNA_4219 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4220 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4221 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4222 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4223 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4224 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4225 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4226 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4227 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4228 (.A(_10812_));
 sg13g2_antennanp ANTENNA_4229 (.A(_10818_));
 sg13g2_antennanp ANTENNA_4230 (.A(_10818_));
 sg13g2_antennanp ANTENNA_4231 (.A(_10818_));
 sg13g2_antennanp ANTENNA_4232 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4233 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4234 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4235 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4236 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4237 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4238 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4239 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4240 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4241 (.A(_10845_));
 sg13g2_antennanp ANTENNA_4242 (.A(clk));
 sg13g2_antennanp ANTENNA_4243 (.A(clk));
 sg13g2_antennanp ANTENNA_4244 (.A(\top_ihp.oisc.micro_res_addr[2] ));
 sg13g2_antennanp ANTENNA_4245 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_4246 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_4247 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_4248 (.A(\top_ihp.oisc.regs[32][10] ));
 sg13g2_antennanp ANTENNA_4249 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_4250 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_4251 (.A(\top_ihp.oisc.regs[32][11] ));
 sg13g2_antennanp ANTENNA_4252 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_4253 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_4254 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_4255 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_4256 (.A(\top_ihp.oisc.regs[32][25] ));
 sg13g2_antennanp ANTENNA_4257 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_4258 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_4259 (.A(\top_ihp.oisc.regs[32][27] ));
 sg13g2_antennanp ANTENNA_4260 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_4261 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_4262 (.A(\top_ihp.oisc.regs[32][2] ));
 sg13g2_antennanp ANTENNA_4263 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_4264 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_4265 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_4266 (.A(\top_ihp.oisc.regs[32][5] ));
 sg13g2_antennanp ANTENNA_4267 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_4268 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_4269 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_4270 (.A(\top_ihp.oisc.regs[32][6] ));
 sg13g2_antennanp ANTENNA_4271 (.A(net54));
 sg13g2_antennanp ANTENNA_4272 (.A(net54));
 sg13g2_antennanp ANTENNA_4273 (.A(net54));
 sg13g2_antennanp ANTENNA_4274 (.A(net54));
 sg13g2_antennanp ANTENNA_4275 (.A(net54));
 sg13g2_antennanp ANTENNA_4276 (.A(net54));
 sg13g2_antennanp ANTENNA_4277 (.A(net54));
 sg13g2_antennanp ANTENNA_4278 (.A(net54));
 sg13g2_antennanp ANTENNA_4279 (.A(net54));
 sg13g2_antennanp ANTENNA_4280 (.A(net56));
 sg13g2_antennanp ANTENNA_4281 (.A(net56));
 sg13g2_antennanp ANTENNA_4282 (.A(net56));
 sg13g2_antennanp ANTENNA_4283 (.A(net56));
 sg13g2_antennanp ANTENNA_4284 (.A(net56));
 sg13g2_antennanp ANTENNA_4285 (.A(net56));
 sg13g2_antennanp ANTENNA_4286 (.A(net56));
 sg13g2_antennanp ANTENNA_4287 (.A(net56));
 sg13g2_antennanp ANTENNA_4288 (.A(net56));
 sg13g2_antennanp ANTENNA_4289 (.A(net90));
 sg13g2_antennanp ANTENNA_4290 (.A(net90));
 sg13g2_antennanp ANTENNA_4291 (.A(net90));
 sg13g2_antennanp ANTENNA_4292 (.A(net90));
 sg13g2_antennanp ANTENNA_4293 (.A(net90));
 sg13g2_antennanp ANTENNA_4294 (.A(net90));
 sg13g2_antennanp ANTENNA_4295 (.A(net90));
 sg13g2_antennanp ANTENNA_4296 (.A(net90));
 sg13g2_antennanp ANTENNA_4297 (.A(net90));
 sg13g2_antennanp ANTENNA_4298 (.A(net117));
 sg13g2_antennanp ANTENNA_4299 (.A(net117));
 sg13g2_antennanp ANTENNA_4300 (.A(net117));
 sg13g2_antennanp ANTENNA_4301 (.A(net117));
 sg13g2_antennanp ANTENNA_4302 (.A(net117));
 sg13g2_antennanp ANTENNA_4303 (.A(net117));
 sg13g2_antennanp ANTENNA_4304 (.A(net117));
 sg13g2_antennanp ANTENNA_4305 (.A(net117));
 sg13g2_antennanp ANTENNA_4306 (.A(net117));
 sg13g2_antennanp ANTENNA_4307 (.A(net117));
 sg13g2_antennanp ANTENNA_4308 (.A(net117));
 sg13g2_antennanp ANTENNA_4309 (.A(net117));
 sg13g2_antennanp ANTENNA_4310 (.A(net117));
 sg13g2_antennanp ANTENNA_4311 (.A(net117));
 sg13g2_antennanp ANTENNA_4312 (.A(net117));
 sg13g2_antennanp ANTENNA_4313 (.A(net117));
 sg13g2_antennanp ANTENNA_4314 (.A(net117));
 sg13g2_antennanp ANTENNA_4315 (.A(net117));
 sg13g2_antennanp ANTENNA_4316 (.A(net117));
 sg13g2_antennanp ANTENNA_4317 (.A(net117));
 sg13g2_antennanp ANTENNA_4318 (.A(net125));
 sg13g2_antennanp ANTENNA_4319 (.A(net125));
 sg13g2_antennanp ANTENNA_4320 (.A(net125));
 sg13g2_antennanp ANTENNA_4321 (.A(net125));
 sg13g2_antennanp ANTENNA_4322 (.A(net125));
 sg13g2_antennanp ANTENNA_4323 (.A(net125));
 sg13g2_antennanp ANTENNA_4324 (.A(net125));
 sg13g2_antennanp ANTENNA_4325 (.A(net125));
 sg13g2_antennanp ANTENNA_4326 (.A(net125));
 sg13g2_antennanp ANTENNA_4327 (.A(net125));
 sg13g2_antennanp ANTENNA_4328 (.A(net125));
 sg13g2_antennanp ANTENNA_4329 (.A(net125));
 sg13g2_antennanp ANTENNA_4330 (.A(net125));
 sg13g2_antennanp ANTENNA_4331 (.A(net125));
 sg13g2_antennanp ANTENNA_4332 (.A(net125));
 sg13g2_antennanp ANTENNA_4333 (.A(net125));
 sg13g2_antennanp ANTENNA_4334 (.A(net125));
 sg13g2_antennanp ANTENNA_4335 (.A(net125));
 sg13g2_antennanp ANTENNA_4336 (.A(net125));
 sg13g2_antennanp ANTENNA_4337 (.A(net127));
 sg13g2_antennanp ANTENNA_4338 (.A(net127));
 sg13g2_antennanp ANTENNA_4339 (.A(net127));
 sg13g2_antennanp ANTENNA_4340 (.A(net127));
 sg13g2_antennanp ANTENNA_4341 (.A(net127));
 sg13g2_antennanp ANTENNA_4342 (.A(net127));
 sg13g2_antennanp ANTENNA_4343 (.A(net127));
 sg13g2_antennanp ANTENNA_4344 (.A(net127));
 sg13g2_antennanp ANTENNA_4345 (.A(net127));
 sg13g2_antennanp ANTENNA_4346 (.A(net127));
 sg13g2_antennanp ANTENNA_4347 (.A(net127));
 sg13g2_antennanp ANTENNA_4348 (.A(net127));
 sg13g2_antennanp ANTENNA_4349 (.A(net127));
 sg13g2_antennanp ANTENNA_4350 (.A(net127));
 sg13g2_antennanp ANTENNA_4351 (.A(net127));
 sg13g2_antennanp ANTENNA_4352 (.A(net127));
 sg13g2_antennanp ANTENNA_4353 (.A(net130));
 sg13g2_antennanp ANTENNA_4354 (.A(net130));
 sg13g2_antennanp ANTENNA_4355 (.A(net130));
 sg13g2_antennanp ANTENNA_4356 (.A(net130));
 sg13g2_antennanp ANTENNA_4357 (.A(net130));
 sg13g2_antennanp ANTENNA_4358 (.A(net130));
 sg13g2_antennanp ANTENNA_4359 (.A(net130));
 sg13g2_antennanp ANTENNA_4360 (.A(net130));
 sg13g2_antennanp ANTENNA_4361 (.A(net130));
 sg13g2_antennanp ANTENNA_4362 (.A(net130));
 sg13g2_antennanp ANTENNA_4363 (.A(net130));
 sg13g2_antennanp ANTENNA_4364 (.A(net130));
 sg13g2_antennanp ANTENNA_4365 (.A(net130));
 sg13g2_antennanp ANTENNA_4366 (.A(net130));
 sg13g2_antennanp ANTENNA_4367 (.A(net130));
 sg13g2_antennanp ANTENNA_4368 (.A(net130));
 sg13g2_antennanp ANTENNA_4369 (.A(net130));
 sg13g2_antennanp ANTENNA_4370 (.A(net130));
 sg13g2_antennanp ANTENNA_4371 (.A(net130));
 sg13g2_antennanp ANTENNA_4372 (.A(net130));
 sg13g2_antennanp ANTENNA_4373 (.A(net130));
 sg13g2_antennanp ANTENNA_4374 (.A(net130));
 sg13g2_antennanp ANTENNA_4375 (.A(net130));
 sg13g2_antennanp ANTENNA_4376 (.A(net132));
 sg13g2_antennanp ANTENNA_4377 (.A(net132));
 sg13g2_antennanp ANTENNA_4378 (.A(net132));
 sg13g2_antennanp ANTENNA_4379 (.A(net132));
 sg13g2_antennanp ANTENNA_4380 (.A(net132));
 sg13g2_antennanp ANTENNA_4381 (.A(net132));
 sg13g2_antennanp ANTENNA_4382 (.A(net132));
 sg13g2_antennanp ANTENNA_4383 (.A(net132));
 sg13g2_antennanp ANTENNA_4384 (.A(net132));
 sg13g2_antennanp ANTENNA_4385 (.A(net134));
 sg13g2_antennanp ANTENNA_4386 (.A(net134));
 sg13g2_antennanp ANTENNA_4387 (.A(net134));
 sg13g2_antennanp ANTENNA_4388 (.A(net134));
 sg13g2_antennanp ANTENNA_4389 (.A(net134));
 sg13g2_antennanp ANTENNA_4390 (.A(net134));
 sg13g2_antennanp ANTENNA_4391 (.A(net134));
 sg13g2_antennanp ANTENNA_4392 (.A(net134));
 sg13g2_antennanp ANTENNA_4393 (.A(net134));
 sg13g2_antennanp ANTENNA_4394 (.A(net134));
 sg13g2_antennanp ANTENNA_4395 (.A(net134));
 sg13g2_antennanp ANTENNA_4396 (.A(net134));
 sg13g2_antennanp ANTENNA_4397 (.A(net134));
 sg13g2_antennanp ANTENNA_4398 (.A(net134));
 sg13g2_antennanp ANTENNA_4399 (.A(net134));
 sg13g2_antennanp ANTENNA_4400 (.A(net134));
 sg13g2_antennanp ANTENNA_4401 (.A(net134));
 sg13g2_antennanp ANTENNA_4402 (.A(net134));
 sg13g2_antennanp ANTENNA_4403 (.A(net134));
 sg13g2_antennanp ANTENNA_4404 (.A(net134));
 sg13g2_antennanp ANTENNA_4405 (.A(net138));
 sg13g2_antennanp ANTENNA_4406 (.A(net138));
 sg13g2_antennanp ANTENNA_4407 (.A(net138));
 sg13g2_antennanp ANTENNA_4408 (.A(net138));
 sg13g2_antennanp ANTENNA_4409 (.A(net138));
 sg13g2_antennanp ANTENNA_4410 (.A(net138));
 sg13g2_antennanp ANTENNA_4411 (.A(net138));
 sg13g2_antennanp ANTENNA_4412 (.A(net138));
 sg13g2_antennanp ANTENNA_4413 (.A(net138));
 sg13g2_antennanp ANTENNA_4414 (.A(net138));
 sg13g2_antennanp ANTENNA_4415 (.A(net138));
 sg13g2_antennanp ANTENNA_4416 (.A(net138));
 sg13g2_antennanp ANTENNA_4417 (.A(net177));
 sg13g2_antennanp ANTENNA_4418 (.A(net177));
 sg13g2_antennanp ANTENNA_4419 (.A(net177));
 sg13g2_antennanp ANTENNA_4420 (.A(net177));
 sg13g2_antennanp ANTENNA_4421 (.A(net177));
 sg13g2_antennanp ANTENNA_4422 (.A(net177));
 sg13g2_antennanp ANTENNA_4423 (.A(net177));
 sg13g2_antennanp ANTENNA_4424 (.A(net177));
 sg13g2_antennanp ANTENNA_4425 (.A(net177));
 sg13g2_antennanp ANTENNA_4426 (.A(net177));
 sg13g2_antennanp ANTENNA_4427 (.A(net177));
 sg13g2_antennanp ANTENNA_4428 (.A(net177));
 sg13g2_antennanp ANTENNA_4429 (.A(net177));
 sg13g2_antennanp ANTENNA_4430 (.A(net177));
 sg13g2_antennanp ANTENNA_4431 (.A(net177));
 sg13g2_antennanp ANTENNA_4432 (.A(net177));
 sg13g2_antennanp ANTENNA_4433 (.A(net177));
 sg13g2_antennanp ANTENNA_4434 (.A(net264));
 sg13g2_antennanp ANTENNA_4435 (.A(net264));
 sg13g2_antennanp ANTENNA_4436 (.A(net264));
 sg13g2_antennanp ANTENNA_4437 (.A(net264));
 sg13g2_antennanp ANTENNA_4438 (.A(net264));
 sg13g2_antennanp ANTENNA_4439 (.A(net264));
 sg13g2_antennanp ANTENNA_4440 (.A(net264));
 sg13g2_antennanp ANTENNA_4441 (.A(net264));
 sg13g2_antennanp ANTENNA_4442 (.A(net264));
 sg13g2_antennanp ANTENNA_4443 (.A(net274));
 sg13g2_antennanp ANTENNA_4444 (.A(net274));
 sg13g2_antennanp ANTENNA_4445 (.A(net274));
 sg13g2_antennanp ANTENNA_4446 (.A(net274));
 sg13g2_antennanp ANTENNA_4447 (.A(net274));
 sg13g2_antennanp ANTENNA_4448 (.A(net274));
 sg13g2_antennanp ANTENNA_4449 (.A(net274));
 sg13g2_antennanp ANTENNA_4450 (.A(net274));
 sg13g2_antennanp ANTENNA_4451 (.A(net274));
 sg13g2_antennanp ANTENNA_4452 (.A(net274));
 sg13g2_antennanp ANTENNA_4453 (.A(net274));
 sg13g2_antennanp ANTENNA_4454 (.A(net274));
 sg13g2_antennanp ANTENNA_4455 (.A(net274));
 sg13g2_antennanp ANTENNA_4456 (.A(net293));
 sg13g2_antennanp ANTENNA_4457 (.A(net293));
 sg13g2_antennanp ANTENNA_4458 (.A(net293));
 sg13g2_antennanp ANTENNA_4459 (.A(net293));
 sg13g2_antennanp ANTENNA_4460 (.A(net293));
 sg13g2_antennanp ANTENNA_4461 (.A(net293));
 sg13g2_antennanp ANTENNA_4462 (.A(net293));
 sg13g2_antennanp ANTENNA_4463 (.A(net293));
 sg13g2_antennanp ANTENNA_4464 (.A(net314));
 sg13g2_antennanp ANTENNA_4465 (.A(net314));
 sg13g2_antennanp ANTENNA_4466 (.A(net314));
 sg13g2_antennanp ANTENNA_4467 (.A(net314));
 sg13g2_antennanp ANTENNA_4468 (.A(net314));
 sg13g2_antennanp ANTENNA_4469 (.A(net314));
 sg13g2_antennanp ANTENNA_4470 (.A(net314));
 sg13g2_antennanp ANTENNA_4471 (.A(net314));
 sg13g2_antennanp ANTENNA_4472 (.A(net314));
 sg13g2_antennanp ANTENNA_4473 (.A(net314));
 sg13g2_antennanp ANTENNA_4474 (.A(net314));
 sg13g2_antennanp ANTENNA_4475 (.A(net314));
 sg13g2_antennanp ANTENNA_4476 (.A(net314));
 sg13g2_antennanp ANTENNA_4477 (.A(net314));
 sg13g2_antennanp ANTENNA_4478 (.A(net314));
 sg13g2_antennanp ANTENNA_4479 (.A(net314));
 sg13g2_antennanp ANTENNA_4480 (.A(net314));
 sg13g2_antennanp ANTENNA_4481 (.A(net314));
 sg13g2_antennanp ANTENNA_4482 (.A(net314));
 sg13g2_antennanp ANTENNA_4483 (.A(net314));
 sg13g2_antennanp ANTENNA_4484 (.A(net314));
 sg13g2_antennanp ANTENNA_4485 (.A(net314));
 sg13g2_antennanp ANTENNA_4486 (.A(net323));
 sg13g2_antennanp ANTENNA_4487 (.A(net323));
 sg13g2_antennanp ANTENNA_4488 (.A(net323));
 sg13g2_antennanp ANTENNA_4489 (.A(net323));
 sg13g2_antennanp ANTENNA_4490 (.A(net323));
 sg13g2_antennanp ANTENNA_4491 (.A(net323));
 sg13g2_antennanp ANTENNA_4492 (.A(net323));
 sg13g2_antennanp ANTENNA_4493 (.A(net323));
 sg13g2_antennanp ANTENNA_4494 (.A(net323));
 sg13g2_antennanp ANTENNA_4495 (.A(net326));
 sg13g2_antennanp ANTENNA_4496 (.A(net326));
 sg13g2_antennanp ANTENNA_4497 (.A(net326));
 sg13g2_antennanp ANTENNA_4498 (.A(net326));
 sg13g2_antennanp ANTENNA_4499 (.A(net326));
 sg13g2_antennanp ANTENNA_4500 (.A(net326));
 sg13g2_antennanp ANTENNA_4501 (.A(net326));
 sg13g2_antennanp ANTENNA_4502 (.A(net326));
 sg13g2_antennanp ANTENNA_4503 (.A(net403));
 sg13g2_antennanp ANTENNA_4504 (.A(net403));
 sg13g2_antennanp ANTENNA_4505 (.A(net403));
 sg13g2_antennanp ANTENNA_4506 (.A(net403));
 sg13g2_antennanp ANTENNA_4507 (.A(net403));
 sg13g2_antennanp ANTENNA_4508 (.A(net403));
 sg13g2_antennanp ANTENNA_4509 (.A(net403));
 sg13g2_antennanp ANTENNA_4510 (.A(net403));
 sg13g2_antennanp ANTENNA_4511 (.A(net403));
 sg13g2_antennanp ANTENNA_4512 (.A(net435));
 sg13g2_antennanp ANTENNA_4513 (.A(net435));
 sg13g2_antennanp ANTENNA_4514 (.A(net435));
 sg13g2_antennanp ANTENNA_4515 (.A(net435));
 sg13g2_antennanp ANTENNA_4516 (.A(net435));
 sg13g2_antennanp ANTENNA_4517 (.A(net435));
 sg13g2_antennanp ANTENNA_4518 (.A(net435));
 sg13g2_antennanp ANTENNA_4519 (.A(net435));
 sg13g2_antennanp ANTENNA_4520 (.A(net435));
 sg13g2_antennanp ANTENNA_4521 (.A(net444));
 sg13g2_antennanp ANTENNA_4522 (.A(net444));
 sg13g2_antennanp ANTENNA_4523 (.A(net444));
 sg13g2_antennanp ANTENNA_4524 (.A(net444));
 sg13g2_antennanp ANTENNA_4525 (.A(net444));
 sg13g2_antennanp ANTENNA_4526 (.A(net444));
 sg13g2_antennanp ANTENNA_4527 (.A(net444));
 sg13g2_antennanp ANTENNA_4528 (.A(net444));
 sg13g2_antennanp ANTENNA_4529 (.A(net444));
 sg13g2_antennanp ANTENNA_4530 (.A(net444));
 sg13g2_antennanp ANTENNA_4531 (.A(net444));
 sg13g2_antennanp ANTENNA_4532 (.A(net444));
 sg13g2_antennanp ANTENNA_4533 (.A(net444));
 sg13g2_antennanp ANTENNA_4534 (.A(net444));
 sg13g2_antennanp ANTENNA_4535 (.A(net444));
 sg13g2_antennanp ANTENNA_4536 (.A(net444));
 sg13g2_antennanp ANTENNA_4537 (.A(net444));
 sg13g2_antennanp ANTENNA_4538 (.A(net444));
 sg13g2_antennanp ANTENNA_4539 (.A(net444));
 sg13g2_antennanp ANTENNA_4540 (.A(net444));
 sg13g2_antennanp ANTENNA_4541 (.A(net444));
 sg13g2_antennanp ANTENNA_4542 (.A(net444));
 sg13g2_antennanp ANTENNA_4543 (.A(net444));
 sg13g2_antennanp ANTENNA_4544 (.A(net449));
 sg13g2_antennanp ANTENNA_4545 (.A(net449));
 sg13g2_antennanp ANTENNA_4546 (.A(net449));
 sg13g2_antennanp ANTENNA_4547 (.A(net449));
 sg13g2_antennanp ANTENNA_4548 (.A(net449));
 sg13g2_antennanp ANTENNA_4549 (.A(net449));
 sg13g2_antennanp ANTENNA_4550 (.A(net449));
 sg13g2_antennanp ANTENNA_4551 (.A(net449));
 sg13g2_antennanp ANTENNA_4552 (.A(net672));
 sg13g2_antennanp ANTENNA_4553 (.A(net672));
 sg13g2_antennanp ANTENNA_4554 (.A(net672));
 sg13g2_antennanp ANTENNA_4555 (.A(net672));
 sg13g2_antennanp ANTENNA_4556 (.A(net672));
 sg13g2_antennanp ANTENNA_4557 (.A(net672));
 sg13g2_antennanp ANTENNA_4558 (.A(net672));
 sg13g2_antennanp ANTENNA_4559 (.A(net672));
 sg13g2_antennanp ANTENNA_4560 (.A(net1421));
 sg13g2_antennanp ANTENNA_4561 (.A(net1421));
 sg13g2_antennanp ANTENNA_4562 (.A(net1421));
 sg13g2_antennanp ANTENNA_4563 (.A(net1421));
 sg13g2_antennanp ANTENNA_4564 (.A(net1421));
 sg13g2_antennanp ANTENNA_4565 (.A(net1421));
 sg13g2_antennanp ANTENNA_4566 (.A(net1421));
 sg13g2_antennanp ANTENNA_4567 (.A(net1421));
 sg13g2_antennanp ANTENNA_4568 (.A(net1421));
 sg13g2_antennanp ANTENNA_4569 (.A(net1421));
 sg13g2_antennanp ANTENNA_4570 (.A(net1421));
 sg13g2_antennanp ANTENNA_4571 (.A(net1421));
 sg13g2_antennanp ANTENNA_4572 (.A(net1421));
 sg13g2_antennanp ANTENNA_4573 (.A(net1421));
 sg13g2_antennanp ANTENNA_4574 (.A(net1421));
 sg13g2_antennanp ANTENNA_4575 (.A(net1421));
 sg13g2_antennanp ANTENNA_4576 (.A(net1421));
 sg13g2_antennanp ANTENNA_4577 (.A(net1421));
 sg13g2_antennanp ANTENNA_4578 (.A(net1421));
 sg13g2_antennanp ANTENNA_4579 (.A(net1421));
 sg13g2_antennanp ANTENNA_4580 (.A(net1421));
 sg13g2_antennanp ANTENNA_4581 (.A(net1421));
 sg13g2_antennanp ANTENNA_4582 (.A(net1421));
 sg13g2_antennanp ANTENNA_4583 (.A(net1421));
 sg13g2_antennanp ANTENNA_4584 (.A(net1421));
 sg13g2_antennanp ANTENNA_4585 (.A(net1421));
 sg13g2_antennanp ANTENNA_4586 (.A(net1421));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_fill_2 FILLER_0_21 ();
 sg13g2_fill_1 FILLER_0_23 ();
 sg13g2_fill_1 FILLER_0_28 ();
 sg13g2_fill_1 FILLER_0_33 ();
 sg13g2_decap_8 FILLER_0_38 ();
 sg13g2_decap_8 FILLER_0_45 ();
 sg13g2_decap_8 FILLER_0_52 ();
 sg13g2_decap_8 FILLER_0_59 ();
 sg13g2_decap_8 FILLER_0_66 ();
 sg13g2_decap_8 FILLER_0_73 ();
 sg13g2_decap_8 FILLER_0_80 ();
 sg13g2_decap_8 FILLER_0_87 ();
 sg13g2_decap_8 FILLER_0_94 ();
 sg13g2_decap_8 FILLER_0_101 ();
 sg13g2_decap_8 FILLER_0_108 ();
 sg13g2_decap_8 FILLER_0_115 ();
 sg13g2_decap_8 FILLER_0_122 ();
 sg13g2_decap_8 FILLER_0_129 ();
 sg13g2_decap_8 FILLER_0_136 ();
 sg13g2_decap_8 FILLER_0_143 ();
 sg13g2_decap_8 FILLER_0_150 ();
 sg13g2_fill_1 FILLER_0_157 ();
 sg13g2_decap_8 FILLER_0_165 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_0_200 ();
 sg13g2_decap_8 FILLER_0_207 ();
 sg13g2_decap_8 FILLER_0_214 ();
 sg13g2_decap_8 FILLER_0_221 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_4 FILLER_0_284 ();
 sg13g2_fill_2 FILLER_0_288 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_4 FILLER_0_319 ();
 sg13g2_fill_1 FILLER_0_323 ();
 sg13g2_decap_8 FILLER_0_328 ();
 sg13g2_decap_8 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_342 ();
 sg13g2_decap_8 FILLER_0_349 ();
 sg13g2_decap_8 FILLER_0_356 ();
 sg13g2_decap_8 FILLER_0_363 ();
 sg13g2_decap_8 FILLER_0_370 ();
 sg13g2_decap_8 FILLER_0_377 ();
 sg13g2_decap_8 FILLER_0_384 ();
 sg13g2_decap_8 FILLER_0_391 ();
 sg13g2_decap_8 FILLER_0_398 ();
 sg13g2_decap_8 FILLER_0_405 ();
 sg13g2_decap_8 FILLER_0_412 ();
 sg13g2_decap_8 FILLER_0_419 ();
 sg13g2_decap_8 FILLER_0_426 ();
 sg13g2_decap_8 FILLER_0_433 ();
 sg13g2_decap_8 FILLER_0_440 ();
 sg13g2_decap_8 FILLER_0_447 ();
 sg13g2_decap_8 FILLER_0_454 ();
 sg13g2_decap_8 FILLER_0_461 ();
 sg13g2_decap_8 FILLER_0_468 ();
 sg13g2_decap_8 FILLER_0_475 ();
 sg13g2_decap_8 FILLER_0_482 ();
 sg13g2_decap_8 FILLER_0_489 ();
 sg13g2_decap_8 FILLER_0_496 ();
 sg13g2_decap_8 FILLER_0_503 ();
 sg13g2_decap_8 FILLER_0_510 ();
 sg13g2_decap_8 FILLER_0_517 ();
 sg13g2_decap_8 FILLER_0_524 ();
 sg13g2_decap_8 FILLER_0_531 ();
 sg13g2_decap_8 FILLER_0_538 ();
 sg13g2_decap_8 FILLER_0_545 ();
 sg13g2_decap_8 FILLER_0_552 ();
 sg13g2_decap_8 FILLER_0_559 ();
 sg13g2_decap_8 FILLER_0_566 ();
 sg13g2_decap_8 FILLER_0_573 ();
 sg13g2_decap_8 FILLER_0_580 ();
 sg13g2_decap_8 FILLER_0_587 ();
 sg13g2_decap_8 FILLER_0_594 ();
 sg13g2_decap_8 FILLER_0_601 ();
 sg13g2_decap_8 FILLER_0_608 ();
 sg13g2_decap_8 FILLER_0_615 ();
 sg13g2_decap_8 FILLER_0_622 ();
 sg13g2_decap_8 FILLER_0_629 ();
 sg13g2_decap_8 FILLER_0_636 ();
 sg13g2_decap_8 FILLER_0_643 ();
 sg13g2_decap_8 FILLER_0_650 ();
 sg13g2_decap_8 FILLER_0_657 ();
 sg13g2_decap_8 FILLER_0_664 ();
 sg13g2_decap_8 FILLER_0_671 ();
 sg13g2_decap_4 FILLER_0_678 ();
 sg13g2_fill_2 FILLER_0_682 ();
 sg13g2_decap_8 FILLER_0_710 ();
 sg13g2_decap_8 FILLER_0_717 ();
 sg13g2_decap_8 FILLER_0_724 ();
 sg13g2_decap_8 FILLER_0_731 ();
 sg13g2_decap_8 FILLER_0_738 ();
 sg13g2_fill_1 FILLER_0_745 ();
 sg13g2_decap_8 FILLER_0_808 ();
 sg13g2_decap_8 FILLER_0_815 ();
 sg13g2_decap_8 FILLER_0_822 ();
 sg13g2_decap_8 FILLER_0_829 ();
 sg13g2_decap_8 FILLER_0_836 ();
 sg13g2_decap_8 FILLER_0_843 ();
 sg13g2_decap_8 FILLER_0_850 ();
 sg13g2_decap_8 FILLER_0_857 ();
 sg13g2_decap_8 FILLER_0_864 ();
 sg13g2_decap_8 FILLER_0_871 ();
 sg13g2_decap_8 FILLER_0_878 ();
 sg13g2_decap_8 FILLER_0_885 ();
 sg13g2_decap_8 FILLER_0_892 ();
 sg13g2_decap_4 FILLER_0_899 ();
 sg13g2_fill_2 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_1009 ();
 sg13g2_decap_8 FILLER_0_1016 ();
 sg13g2_decap_8 FILLER_0_1023 ();
 sg13g2_decap_8 FILLER_0_1030 ();
 sg13g2_decap_4 FILLER_0_1037 ();
 sg13g2_fill_2 FILLER_0_1041 ();
 sg13g2_fill_1 FILLER_0_1053 ();
 sg13g2_fill_2 FILLER_0_1080 ();
 sg13g2_fill_1 FILLER_0_1082 ();
 sg13g2_decap_8 FILLER_0_1098 ();
 sg13g2_decap_8 FILLER_0_1105 ();
 sg13g2_decap_8 FILLER_0_1112 ();
 sg13g2_decap_8 FILLER_0_1119 ();
 sg13g2_decap_8 FILLER_0_1126 ();
 sg13g2_decap_8 FILLER_0_1133 ();
 sg13g2_decap_8 FILLER_0_1140 ();
 sg13g2_decap_8 FILLER_0_1147 ();
 sg13g2_decap_8 FILLER_0_1154 ();
 sg13g2_decap_8 FILLER_0_1161 ();
 sg13g2_decap_8 FILLER_0_1168 ();
 sg13g2_decap_4 FILLER_0_1175 ();
 sg13g2_fill_1 FILLER_0_1179 ();
 sg13g2_decap_8 FILLER_0_1183 ();
 sg13g2_fill_2 FILLER_0_1190 ();
 sg13g2_fill_1 FILLER_0_1192 ();
 sg13g2_decap_8 FILLER_0_1208 ();
 sg13g2_decap_8 FILLER_0_1215 ();
 sg13g2_decap_8 FILLER_0_1222 ();
 sg13g2_decap_8 FILLER_0_1229 ();
 sg13g2_decap_8 FILLER_0_1236 ();
 sg13g2_decap_8 FILLER_0_1243 ();
 sg13g2_decap_8 FILLER_0_1250 ();
 sg13g2_decap_8 FILLER_0_1257 ();
 sg13g2_decap_8 FILLER_0_1264 ();
 sg13g2_decap_8 FILLER_0_1271 ();
 sg13g2_decap_8 FILLER_0_1278 ();
 sg13g2_decap_8 FILLER_0_1285 ();
 sg13g2_decap_8 FILLER_0_1292 ();
 sg13g2_decap_8 FILLER_0_1299 ();
 sg13g2_decap_8 FILLER_0_1306 ();
 sg13g2_decap_8 FILLER_0_1313 ();
 sg13g2_decap_8 FILLER_0_1320 ();
 sg13g2_decap_8 FILLER_0_1327 ();
 sg13g2_decap_8 FILLER_0_1334 ();
 sg13g2_decap_8 FILLER_0_1341 ();
 sg13g2_decap_8 FILLER_0_1348 ();
 sg13g2_decap_8 FILLER_0_1355 ();
 sg13g2_decap_8 FILLER_0_1362 ();
 sg13g2_decap_8 FILLER_0_1369 ();
 sg13g2_decap_8 FILLER_0_1376 ();
 sg13g2_decap_8 FILLER_0_1383 ();
 sg13g2_fill_1 FILLER_0_1390 ();
 sg13g2_decap_4 FILLER_0_1417 ();
 sg13g2_fill_1 FILLER_0_1421 ();
 sg13g2_decap_8 FILLER_0_1461 ();
 sg13g2_decap_8 FILLER_0_1468 ();
 sg13g2_decap_8 FILLER_0_1475 ();
 sg13g2_decap_8 FILLER_0_1482 ();
 sg13g2_decap_8 FILLER_0_1489 ();
 sg13g2_decap_8 FILLER_0_1496 ();
 sg13g2_decap_8 FILLER_0_1503 ();
 sg13g2_decap_8 FILLER_0_1510 ();
 sg13g2_decap_8 FILLER_0_1517 ();
 sg13g2_decap_4 FILLER_0_1524 ();
 sg13g2_fill_2 FILLER_0_1528 ();
 sg13g2_decap_8 FILLER_0_1542 ();
 sg13g2_decap_8 FILLER_0_1549 ();
 sg13g2_decap_8 FILLER_0_1556 ();
 sg13g2_fill_2 FILLER_0_1563 ();
 sg13g2_fill_1 FILLER_0_1565 ();
 sg13g2_decap_8 FILLER_0_1596 ();
 sg13g2_decap_8 FILLER_0_1633 ();
 sg13g2_decap_8 FILLER_0_1640 ();
 sg13g2_fill_2 FILLER_0_1647 ();
 sg13g2_decap_8 FILLER_0_1679 ();
 sg13g2_decap_8 FILLER_0_1686 ();
 sg13g2_decap_8 FILLER_0_1693 ();
 sg13g2_decap_8 FILLER_0_1700 ();
 sg13g2_decap_8 FILLER_0_1707 ();
 sg13g2_decap_8 FILLER_0_1714 ();
 sg13g2_decap_8 FILLER_0_1721 ();
 sg13g2_decap_8 FILLER_0_1728 ();
 sg13g2_fill_2 FILLER_0_1735 ();
 sg13g2_decap_8 FILLER_0_1741 ();
 sg13g2_decap_8 FILLER_0_1748 ();
 sg13g2_decap_8 FILLER_0_1755 ();
 sg13g2_fill_2 FILLER_0_1762 ();
 sg13g2_fill_1 FILLER_0_1764 ();
 sg13g2_decap_4 FILLER_0_1799 ();
 sg13g2_fill_1 FILLER_0_1803 ();
 sg13g2_decap_8 FILLER_0_1830 ();
 sg13g2_decap_8 FILLER_0_1837 ();
 sg13g2_decap_8 FILLER_0_1844 ();
 sg13g2_decap_8 FILLER_0_1851 ();
 sg13g2_decap_8 FILLER_0_1858 ();
 sg13g2_decap_8 FILLER_0_1865 ();
 sg13g2_decap_8 FILLER_0_1872 ();
 sg13g2_decap_8 FILLER_0_1879 ();
 sg13g2_fill_1 FILLER_0_1886 ();
 sg13g2_decap_8 FILLER_0_1917 ();
 sg13g2_decap_8 FILLER_0_1924 ();
 sg13g2_decap_8 FILLER_0_1931 ();
 sg13g2_decap_8 FILLER_0_1938 ();
 sg13g2_decap_8 FILLER_0_1945 ();
 sg13g2_decap_4 FILLER_0_1952 ();
 sg13g2_fill_1 FILLER_0_1960 ();
 sg13g2_decap_8 FILLER_0_1987 ();
 sg13g2_fill_2 FILLER_0_1994 ();
 sg13g2_fill_2 FILLER_0_2011 ();
 sg13g2_decap_8 FILLER_0_2023 ();
 sg13g2_decap_8 FILLER_0_2030 ();
 sg13g2_fill_2 FILLER_0_2037 ();
 sg13g2_fill_1 FILLER_0_2039 ();
 sg13g2_decap_8 FILLER_0_2043 ();
 sg13g2_fill_2 FILLER_0_2050 ();
 sg13g2_decap_8 FILLER_0_2078 ();
 sg13g2_decap_8 FILLER_0_2085 ();
 sg13g2_fill_2 FILLER_0_2092 ();
 sg13g2_decap_8 FILLER_0_2098 ();
 sg13g2_decap_4 FILLER_0_2105 ();
 sg13g2_decap_8 FILLER_0_2139 ();
 sg13g2_decap_8 FILLER_0_2146 ();
 sg13g2_decap_8 FILLER_0_2153 ();
 sg13g2_decap_8 FILLER_0_2160 ();
 sg13g2_decap_8 FILLER_0_2167 ();
 sg13g2_decap_8 FILLER_0_2174 ();
 sg13g2_decap_4 FILLER_0_2181 ();
 sg13g2_fill_1 FILLER_0_2185 ();
 sg13g2_decap_8 FILLER_0_2201 ();
 sg13g2_decap_4 FILLER_0_2208 ();
 sg13g2_fill_1 FILLER_0_2212 ();
 sg13g2_decap_8 FILLER_0_2265 ();
 sg13g2_decap_8 FILLER_0_2272 ();
 sg13g2_decap_8 FILLER_0_2279 ();
 sg13g2_decap_8 FILLER_0_2286 ();
 sg13g2_decap_4 FILLER_0_2293 ();
 sg13g2_fill_2 FILLER_0_2297 ();
 sg13g2_decap_8 FILLER_0_2303 ();
 sg13g2_decap_4 FILLER_0_2310 ();
 sg13g2_fill_2 FILLER_0_2314 ();
 sg13g2_fill_2 FILLER_0_2320 ();
 sg13g2_fill_1 FILLER_0_2322 ();
 sg13g2_decap_8 FILLER_0_2327 ();
 sg13g2_decap_8 FILLER_0_2334 ();
 sg13g2_decap_8 FILLER_0_2341 ();
 sg13g2_decap_8 FILLER_0_2348 ();
 sg13g2_decap_8 FILLER_0_2355 ();
 sg13g2_decap_8 FILLER_0_2362 ();
 sg13g2_decap_8 FILLER_0_2369 ();
 sg13g2_decap_8 FILLER_0_2376 ();
 sg13g2_decap_8 FILLER_0_2383 ();
 sg13g2_decap_8 FILLER_0_2390 ();
 sg13g2_decap_8 FILLER_0_2397 ();
 sg13g2_decap_8 FILLER_0_2404 ();
 sg13g2_fill_2 FILLER_0_2411 ();
 sg13g2_fill_1 FILLER_0_2413 ();
 sg13g2_decap_8 FILLER_0_2480 ();
 sg13g2_decap_8 FILLER_0_2487 ();
 sg13g2_decap_8 FILLER_0_2494 ();
 sg13g2_decap_8 FILLER_0_2501 ();
 sg13g2_decap_8 FILLER_0_2508 ();
 sg13g2_decap_8 FILLER_0_2515 ();
 sg13g2_decap_8 FILLER_0_2522 ();
 sg13g2_decap_8 FILLER_0_2529 ();
 sg13g2_decap_8 FILLER_0_2536 ();
 sg13g2_decap_8 FILLER_0_2543 ();
 sg13g2_decap_8 FILLER_0_2550 ();
 sg13g2_decap_8 FILLER_0_2557 ();
 sg13g2_decap_8 FILLER_0_2564 ();
 sg13g2_decap_8 FILLER_0_2571 ();
 sg13g2_decap_8 FILLER_0_2578 ();
 sg13g2_decap_8 FILLER_0_2585 ();
 sg13g2_decap_8 FILLER_0_2592 ();
 sg13g2_decap_8 FILLER_0_2599 ();
 sg13g2_decap_8 FILLER_0_2606 ();
 sg13g2_decap_8 FILLER_0_2613 ();
 sg13g2_decap_8 FILLER_0_2620 ();
 sg13g2_decap_8 FILLER_0_2627 ();
 sg13g2_decap_8 FILLER_0_2634 ();
 sg13g2_decap_8 FILLER_0_2641 ();
 sg13g2_decap_8 FILLER_0_2648 ();
 sg13g2_decap_8 FILLER_0_2655 ();
 sg13g2_decap_8 FILLER_0_2662 ();
 sg13g2_fill_1 FILLER_0_2669 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_4 FILLER_1_7 ();
 sg13g2_fill_1 FILLER_1_11 ();
 sg13g2_fill_2 FILLER_1_50 ();
 sg13g2_fill_2 FILLER_1_60 ();
 sg13g2_fill_1 FILLER_1_62 ();
 sg13g2_fill_2 FILLER_1_67 ();
 sg13g2_decap_8 FILLER_1_95 ();
 sg13g2_decap_4 FILLER_1_102 ();
 sg13g2_fill_1 FILLER_1_110 ();
 sg13g2_fill_1 FILLER_1_115 ();
 sg13g2_decap_4 FILLER_1_120 ();
 sg13g2_fill_1 FILLER_1_124 ();
 sg13g2_fill_1 FILLER_1_166 ();
 sg13g2_fill_1 FILLER_1_171 ();
 sg13g2_fill_1 FILLER_1_176 ();
 sg13g2_fill_2 FILLER_1_181 ();
 sg13g2_fill_1 FILLER_1_191 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_fill_2 FILLER_1_203 ();
 sg13g2_fill_1 FILLER_1_205 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_4 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_246 ();
 sg13g2_decap_8 FILLER_1_253 ();
 sg13g2_decap_8 FILLER_1_260 ();
 sg13g2_fill_1 FILLER_1_267 ();
 sg13g2_fill_2 FILLER_1_324 ();
 sg13g2_fill_1 FILLER_1_364 ();
 sg13g2_fill_1 FILLER_1_369 ();
 sg13g2_decap_8 FILLER_1_374 ();
 sg13g2_decap_4 FILLER_1_381 ();
 sg13g2_decap_8 FILLER_1_415 ();
 sg13g2_decap_8 FILLER_1_422 ();
 sg13g2_decap_8 FILLER_1_429 ();
 sg13g2_fill_2 FILLER_1_436 ();
 sg13g2_decap_8 FILLER_1_516 ();
 sg13g2_decap_4 FILLER_1_523 ();
 sg13g2_fill_1 FILLER_1_527 ();
 sg13g2_decap_8 FILLER_1_559 ();
 sg13g2_decap_8 FILLER_1_566 ();
 sg13g2_decap_4 FILLER_1_573 ();
 sg13g2_decap_8 FILLER_1_603 ();
 sg13g2_decap_4 FILLER_1_610 ();
 sg13g2_decap_8 FILLER_1_640 ();
 sg13g2_decap_8 FILLER_1_647 ();
 sg13g2_decap_8 FILLER_1_654 ();
 sg13g2_decap_8 FILLER_1_661 ();
 sg13g2_decap_4 FILLER_1_668 ();
 sg13g2_fill_2 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_684 ();
 sg13g2_decap_4 FILLER_1_691 ();
 sg13g2_fill_1 FILLER_1_695 ();
 sg13g2_decap_4 FILLER_1_748 ();
 sg13g2_fill_2 FILLER_1_752 ();
 sg13g2_decap_4 FILLER_1_790 ();
 sg13g2_fill_1 FILLER_1_820 ();
 sg13g2_fill_2 FILLER_1_860 ();
 sg13g2_fill_1 FILLER_1_862 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_fill_2 FILLER_1_899 ();
 sg13g2_fill_2 FILLER_1_927 ();
 sg13g2_fill_2 FILLER_1_990 ();
 sg13g2_decap_8 FILLER_1_1018 ();
 sg13g2_fill_2 FILLER_1_1025 ();
 sg13g2_fill_1 FILLER_1_1027 ();
 sg13g2_decap_8 FILLER_1_1054 ();
 sg13g2_decap_8 FILLER_1_1061 ();
 sg13g2_decap_8 FILLER_1_1078 ();
 sg13g2_fill_1 FILLER_1_1085 ();
 sg13g2_decap_4 FILLER_1_1122 ();
 sg13g2_fill_2 FILLER_1_1126 ();
 sg13g2_decap_8 FILLER_1_1154 ();
 sg13g2_decap_4 FILLER_1_1161 ();
 sg13g2_decap_4 FILLER_1_1191 ();
 sg13g2_fill_1 FILLER_1_1195 ();
 sg13g2_decap_8 FILLER_1_1206 ();
 sg13g2_decap_4 FILLER_1_1213 ();
 sg13g2_decap_4 FILLER_1_1279 ();
 sg13g2_fill_2 FILLER_1_1283 ();
 sg13g2_fill_1 FILLER_1_1295 ();
 sg13g2_decap_8 FILLER_1_1328 ();
 sg13g2_decap_8 FILLER_1_1335 ();
 sg13g2_decap_8 FILLER_1_1342 ();
 sg13g2_decap_8 FILLER_1_1349 ();
 sg13g2_decap_4 FILLER_1_1356 ();
 sg13g2_decap_4 FILLER_1_1386 ();
 sg13g2_fill_1 FILLER_1_1390 ();
 sg13g2_decap_8 FILLER_1_1401 ();
 sg13g2_decap_8 FILLER_1_1408 ();
 sg13g2_fill_1 FILLER_1_1415 ();
 sg13g2_decap_4 FILLER_1_1467 ();
 sg13g2_decap_8 FILLER_1_1497 ();
 sg13g2_fill_2 FILLER_1_1504 ();
 sg13g2_fill_1 FILLER_1_1506 ();
 sg13g2_decap_8 FILLER_1_1543 ();
 sg13g2_decap_4 FILLER_1_1550 ();
 sg13g2_fill_1 FILLER_1_1554 ();
 sg13g2_fill_2 FILLER_1_1560 ();
 sg13g2_fill_1 FILLER_1_1562 ();
 sg13g2_decap_8 FILLER_1_1593 ();
 sg13g2_decap_4 FILLER_1_1600 ();
 sg13g2_fill_1 FILLER_1_1604 ();
 sg13g2_decap_4 FILLER_1_1639 ();
 sg13g2_fill_1 FILLER_1_1643 ();
 sg13g2_decap_8 FILLER_1_1674 ();
 sg13g2_decap_8 FILLER_1_1681 ();
 sg13g2_decap_8 FILLER_1_1702 ();
 sg13g2_fill_2 FILLER_1_1709 ();
 sg13g2_decap_4 FILLER_1_1721 ();
 sg13g2_fill_1 FILLER_1_1725 ();
 sg13g2_decap_4 FILLER_1_1838 ();
 sg13g2_fill_1 FILLER_1_1842 ();
 sg13g2_decap_8 FILLER_1_1905 ();
 sg13g2_decap_4 FILLER_1_1912 ();
 sg13g2_fill_2 FILLER_1_1916 ();
 sg13g2_fill_2 FILLER_1_1922 ();
 sg13g2_decap_8 FILLER_1_1950 ();
 sg13g2_decap_8 FILLER_1_1957 ();
 sg13g2_decap_8 FILLER_1_1964 ();
 sg13g2_decap_8 FILLER_1_1971 ();
 sg13g2_decap_8 FILLER_1_1978 ();
 sg13g2_decap_8 FILLER_1_1985 ();
 sg13g2_fill_1 FILLER_1_1992 ();
 sg13g2_fill_1 FILLER_1_2036 ();
 sg13g2_fill_1 FILLER_1_2075 ();
 sg13g2_decap_8 FILLER_1_2132 ();
 sg13g2_decap_8 FILLER_1_2139 ();
 sg13g2_fill_2 FILLER_1_2146 ();
 sg13g2_decap_8 FILLER_1_2178 ();
 sg13g2_fill_1 FILLER_1_2185 ();
 sg13g2_decap_8 FILLER_1_2222 ();
 sg13g2_fill_2 FILLER_1_2233 ();
 sg13g2_fill_1 FILLER_1_2235 ();
 sg13g2_fill_2 FILLER_1_2281 ();
 sg13g2_decap_4 FILLER_1_2351 ();
 sg13g2_fill_1 FILLER_1_2355 ();
 sg13g2_fill_2 FILLER_1_2386 ();
 sg13g2_fill_2 FILLER_1_2414 ();
 sg13g2_fill_1 FILLER_1_2416 ();
 sg13g2_fill_1 FILLER_1_2450 ();
 sg13g2_decap_8 FILLER_1_2484 ();
 sg13g2_fill_2 FILLER_1_2521 ();
 sg13g2_fill_1 FILLER_1_2523 ();
 sg13g2_decap_8 FILLER_1_2532 ();
 sg13g2_decap_8 FILLER_1_2539 ();
 sg13g2_decap_8 FILLER_1_2546 ();
 sg13g2_decap_8 FILLER_1_2553 ();
 sg13g2_decap_8 FILLER_1_2560 ();
 sg13g2_decap_8 FILLER_1_2567 ();
 sg13g2_decap_8 FILLER_1_2574 ();
 sg13g2_decap_8 FILLER_1_2581 ();
 sg13g2_decap_8 FILLER_1_2588 ();
 sg13g2_decap_8 FILLER_1_2595 ();
 sg13g2_decap_8 FILLER_1_2602 ();
 sg13g2_decap_8 FILLER_1_2609 ();
 sg13g2_decap_8 FILLER_1_2616 ();
 sg13g2_decap_8 FILLER_1_2623 ();
 sg13g2_decap_8 FILLER_1_2630 ();
 sg13g2_decap_8 FILLER_1_2637 ();
 sg13g2_decap_8 FILLER_1_2644 ();
 sg13g2_decap_8 FILLER_1_2651 ();
 sg13g2_decap_8 FILLER_1_2658 ();
 sg13g2_decap_4 FILLER_1_2665 ();
 sg13g2_fill_1 FILLER_1_2669 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_62 ();
 sg13g2_fill_1 FILLER_2_67 ();
 sg13g2_fill_2 FILLER_2_75 ();
 sg13g2_fill_2 FILLER_2_85 ();
 sg13g2_fill_1 FILLER_2_87 ();
 sg13g2_fill_1 FILLER_2_92 ();
 sg13g2_fill_1 FILLER_2_97 ();
 sg13g2_fill_1 FILLER_2_107 ();
 sg13g2_fill_1 FILLER_2_117 ();
 sg13g2_fill_1 FILLER_2_122 ();
 sg13g2_fill_1 FILLER_2_160 ();
 sg13g2_fill_2 FILLER_2_180 ();
 sg13g2_fill_1 FILLER_2_182 ();
 sg13g2_fill_1 FILLER_2_188 ();
 sg13g2_fill_1 FILLER_2_205 ();
 sg13g2_fill_1 FILLER_2_219 ();
 sg13g2_fill_2 FILLER_2_237 ();
 sg13g2_decap_8 FILLER_2_255 ();
 sg13g2_fill_1 FILLER_2_267 ();
 sg13g2_fill_2 FILLER_2_272 ();
 sg13g2_decap_4 FILLER_2_282 ();
 sg13g2_fill_1 FILLER_2_286 ();
 sg13g2_fill_2 FILLER_2_300 ();
 sg13g2_fill_1 FILLER_2_302 ();
 sg13g2_fill_1 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_fill_1 FILLER_2_354 ();
 sg13g2_fill_1 FILLER_2_363 ();
 sg13g2_fill_1 FILLER_2_369 ();
 sg13g2_fill_1 FILLER_2_395 ();
 sg13g2_decap_4 FILLER_2_422 ();
 sg13g2_fill_2 FILLER_2_426 ();
 sg13g2_fill_2 FILLER_2_454 ();
 sg13g2_fill_1 FILLER_2_456 ();
 sg13g2_fill_1 FILLER_2_460 ();
 sg13g2_fill_1 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_483 ();
 sg13g2_decap_8 FILLER_2_490 ();
 sg13g2_decap_4 FILLER_2_497 ();
 sg13g2_fill_2 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_602 ();
 sg13g2_decap_4 FILLER_2_609 ();
 sg13g2_fill_2 FILLER_2_618 ();
 sg13g2_decap_8 FILLER_2_625 ();
 sg13g2_decap_8 FILLER_2_632 ();
 sg13g2_fill_2 FILLER_2_639 ();
 sg13g2_fill_1 FILLER_2_641 ();
 sg13g2_fill_1 FILLER_2_668 ();
 sg13g2_decap_8 FILLER_2_695 ();
 sg13g2_decap_4 FILLER_2_702 ();
 sg13g2_fill_1 FILLER_2_738 ();
 sg13g2_fill_1 FILLER_2_764 ();
 sg13g2_fill_2 FILLER_2_780 ();
 sg13g2_fill_1 FILLER_2_808 ();
 sg13g2_fill_2 FILLER_2_835 ();
 sg13g2_fill_2 FILLER_2_863 ();
 sg13g2_fill_2 FILLER_2_908 ();
 sg13g2_decap_4 FILLER_2_920 ();
 sg13g2_fill_2 FILLER_2_924 ();
 sg13g2_fill_1 FILLER_2_973 ();
 sg13g2_fill_2 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_1054 ();
 sg13g2_fill_2 FILLER_2_1061 ();
 sg13g2_fill_1 FILLER_2_1063 ();
 sg13g2_decap_4 FILLER_2_1126 ();
 sg13g2_fill_2 FILLER_2_1130 ();
 sg13g2_fill_2 FILLER_2_1178 ();
 sg13g2_fill_1 FILLER_2_1186 ();
 sg13g2_decap_8 FILLER_2_1275 ();
 sg13g2_decap_8 FILLER_2_1282 ();
 sg13g2_fill_1 FILLER_2_1328 ();
 sg13g2_decap_8 FILLER_2_1355 ();
 sg13g2_decap_4 FILLER_2_1388 ();
 sg13g2_fill_1 FILLER_2_1418 ();
 sg13g2_fill_1 FILLER_2_1431 ();
 sg13g2_fill_1 FILLER_2_1458 ();
 sg13g2_decap_4 FILLER_2_1498 ();
 sg13g2_fill_2 FILLER_2_1502 ();
 sg13g2_fill_1 FILLER_2_1533 ();
 sg13g2_fill_1 FILLER_2_1573 ();
 sg13g2_fill_1 FILLER_2_1582 ();
 sg13g2_decap_8 FILLER_2_1589 ();
 sg13g2_decap_8 FILLER_2_1596 ();
 sg13g2_decap_8 FILLER_2_1603 ();
 sg13g2_decap_8 FILLER_2_1610 ();
 sg13g2_decap_4 FILLER_2_1627 ();
 sg13g2_fill_2 FILLER_2_1631 ();
 sg13g2_decap_8 FILLER_2_1638 ();
 sg13g2_decap_8 FILLER_2_1645 ();
 sg13g2_fill_2 FILLER_2_1652 ();
 sg13g2_fill_2 FILLER_2_1658 ();
 sg13g2_fill_1 FILLER_2_1667 ();
 sg13g2_decap_4 FILLER_2_1680 ();
 sg13g2_fill_2 FILLER_2_1694 ();
 sg13g2_fill_2 FILLER_2_1748 ();
 sg13g2_decap_8 FILLER_2_1792 ();
 sg13g2_fill_1 FILLER_2_1816 ();
 sg13g2_decap_8 FILLER_2_1869 ();
 sg13g2_decap_4 FILLER_2_1876 ();
 sg13g2_fill_1 FILLER_2_1884 ();
 sg13g2_fill_2 FILLER_2_1889 ();
 sg13g2_fill_2 FILLER_2_1895 ();
 sg13g2_decap_4 FILLER_2_1926 ();
 sg13g2_fill_2 FILLER_2_1934 ();
 sg13g2_fill_1 FILLER_2_1936 ();
 sg13g2_fill_1 FILLER_2_1941 ();
 sg13g2_fill_1 FILLER_2_1968 ();
 sg13g2_decap_8 FILLER_2_1995 ();
 sg13g2_decap_8 FILLER_2_2002 ();
 sg13g2_decap_8 FILLER_2_2009 ();
 sg13g2_fill_1 FILLER_2_2049 ();
 sg13g2_fill_2 FILLER_2_2054 ();
 sg13g2_fill_2 FILLER_2_2106 ();
 sg13g2_fill_2 FILLER_2_2115 ();
 sg13g2_decap_8 FILLER_2_2146 ();
 sg13g2_fill_1 FILLER_2_2153 ();
 sg13g2_decap_8 FILLER_2_2158 ();
 sg13g2_fill_2 FILLER_2_2165 ();
 sg13g2_fill_1 FILLER_2_2167 ();
 sg13g2_decap_8 FILLER_2_2224 ();
 sg13g2_fill_2 FILLER_2_2231 ();
 sg13g2_fill_1 FILLER_2_2233 ();
 sg13g2_fill_2 FILLER_2_2240 ();
 sg13g2_fill_1 FILLER_2_2251 ();
 sg13g2_fill_1 FILLER_2_2278 ();
 sg13g2_fill_1 FILLER_2_2305 ();
 sg13g2_fill_1 FILLER_2_2310 ();
 sg13g2_fill_1 FILLER_2_2337 ();
 sg13g2_decap_4 FILLER_2_2394 ();
 sg13g2_decap_4 FILLER_2_2402 ();
 sg13g2_fill_2 FILLER_2_2406 ();
 sg13g2_fill_2 FILLER_2_2439 ();
 sg13g2_fill_1 FILLER_2_2459 ();
 sg13g2_fill_1 FILLER_2_2497 ();
 sg13g2_decap_8 FILLER_2_2554 ();
 sg13g2_decap_8 FILLER_2_2561 ();
 sg13g2_decap_8 FILLER_2_2568 ();
 sg13g2_decap_8 FILLER_2_2575 ();
 sg13g2_decap_8 FILLER_2_2582 ();
 sg13g2_decap_8 FILLER_2_2589 ();
 sg13g2_decap_8 FILLER_2_2596 ();
 sg13g2_decap_8 FILLER_2_2603 ();
 sg13g2_decap_8 FILLER_2_2610 ();
 sg13g2_decap_8 FILLER_2_2617 ();
 sg13g2_decap_8 FILLER_2_2624 ();
 sg13g2_decap_8 FILLER_2_2631 ();
 sg13g2_decap_8 FILLER_2_2638 ();
 sg13g2_decap_8 FILLER_2_2645 ();
 sg13g2_decap_8 FILLER_2_2652 ();
 sg13g2_decap_8 FILLER_2_2659 ();
 sg13g2_decap_4 FILLER_2_2666 ();
 sg13g2_fill_2 FILLER_3_0 ();
 sg13g2_fill_2 FILLER_3_36 ();
 sg13g2_fill_1 FILLER_3_38 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_54 ();
 sg13g2_fill_1 FILLER_3_58 ();
 sg13g2_fill_1 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_76 ();
 sg13g2_decap_8 FILLER_3_83 ();
 sg13g2_fill_2 FILLER_3_107 ();
 sg13g2_fill_2 FILLER_3_113 ();
 sg13g2_fill_1 FILLER_3_127 ();
 sg13g2_fill_1 FILLER_3_138 ();
 sg13g2_fill_1 FILLER_3_148 ();
 sg13g2_fill_1 FILLER_3_160 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_fill_2 FILLER_3_176 ();
 sg13g2_fill_2 FILLER_3_182 ();
 sg13g2_fill_2 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_231 ();
 sg13g2_fill_1 FILLER_3_244 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_2 FILLER_3_279 ();
 sg13g2_fill_2 FILLER_3_289 ();
 sg13g2_fill_1 FILLER_3_304 ();
 sg13g2_fill_2 FILLER_3_337 ();
 sg13g2_fill_1 FILLER_3_339 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_fill_1 FILLER_3_379 ();
 sg13g2_fill_1 FILLER_3_405 ();
 sg13g2_decap_8 FILLER_3_411 ();
 sg13g2_fill_2 FILLER_3_418 ();
 sg13g2_decap_8 FILLER_3_459 ();
 sg13g2_decap_8 FILLER_3_466 ();
 sg13g2_decap_8 FILLER_3_473 ();
 sg13g2_decap_8 FILLER_3_480 ();
 sg13g2_decap_8 FILLER_3_487 ();
 sg13g2_fill_2 FILLER_3_494 ();
 sg13g2_fill_1 FILLER_3_496 ();
 sg13g2_decap_8 FILLER_3_500 ();
 sg13g2_decap_8 FILLER_3_507 ();
 sg13g2_decap_8 FILLER_3_514 ();
 sg13g2_fill_2 FILLER_3_521 ();
 sg13g2_fill_2 FILLER_3_537 ();
 sg13g2_decap_8 FILLER_3_569 ();
 sg13g2_fill_2 FILLER_3_576 ();
 sg13g2_fill_1 FILLER_3_598 ();
 sg13g2_fill_1 FILLER_3_603 ();
 sg13g2_decap_4 FILLER_3_635 ();
 sg13g2_fill_1 FILLER_3_639 ();
 sg13g2_fill_2 FILLER_3_645 ();
 sg13g2_fill_1 FILLER_3_647 ();
 sg13g2_fill_1 FILLER_3_674 ();
 sg13g2_decap_4 FILLER_3_685 ();
 sg13g2_fill_1 FILLER_3_689 ();
 sg13g2_fill_2 FILLER_3_708 ();
 sg13g2_fill_1 FILLER_3_734 ();
 sg13g2_decap_4 FILLER_3_786 ();
 sg13g2_fill_1 FILLER_3_810 ();
 sg13g2_fill_1 FILLER_3_817 ();
 sg13g2_decap_4 FILLER_3_906 ();
 sg13g2_fill_2 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_1012 ();
 sg13g2_decap_8 FILLER_3_1019 ();
 sg13g2_decap_4 FILLER_3_1026 ();
 sg13g2_fill_2 FILLER_3_1030 ();
 sg13g2_decap_4 FILLER_3_1040 ();
 sg13g2_fill_2 FILLER_3_1077 ();
 sg13g2_decap_8 FILLER_3_1095 ();
 sg13g2_decap_8 FILLER_3_1102 ();
 sg13g2_fill_1 FILLER_3_1109 ();
 sg13g2_decap_8 FILLER_3_1145 ();
 sg13g2_fill_2 FILLER_3_1152 ();
 sg13g2_fill_2 FILLER_3_1183 ();
 sg13g2_decap_4 FILLER_3_1221 ();
 sg13g2_fill_1 FILLER_3_1225 ();
 sg13g2_decap_8 FILLER_3_1245 ();
 sg13g2_fill_1 FILLER_3_1258 ();
 sg13g2_decap_8 FILLER_3_1295 ();
 sg13g2_fill_2 FILLER_3_1302 ();
 sg13g2_fill_1 FILLER_3_1304 ();
 sg13g2_decap_4 FILLER_3_1351 ();
 sg13g2_fill_1 FILLER_3_1355 ();
 sg13g2_decap_8 FILLER_3_1366 ();
 sg13g2_fill_2 FILLER_3_1373 ();
 sg13g2_fill_1 FILLER_3_1375 ();
 sg13g2_decap_8 FILLER_3_1386 ();
 sg13g2_fill_2 FILLER_3_1393 ();
 sg13g2_fill_1 FILLER_3_1421 ();
 sg13g2_fill_2 FILLER_3_1455 ();
 sg13g2_fill_2 FILLER_3_1463 ();
 sg13g2_fill_1 FILLER_3_1575 ();
 sg13g2_decap_8 FILLER_3_1605 ();
 sg13g2_decap_4 FILLER_3_1633 ();
 sg13g2_fill_2 FILLER_3_1722 ();
 sg13g2_decap_8 FILLER_3_1747 ();
 sg13g2_fill_2 FILLER_3_1754 ();
 sg13g2_fill_1 FILLER_3_1768 ();
 sg13g2_decap_8 FILLER_3_1795 ();
 sg13g2_fill_2 FILLER_3_1802 ();
 sg13g2_fill_1 FILLER_3_1804 ();
 sg13g2_fill_2 FILLER_3_1813 ();
 sg13g2_fill_1 FILLER_3_1815 ();
 sg13g2_decap_8 FILLER_3_1826 ();
 sg13g2_fill_2 FILLER_3_1833 ();
 sg13g2_fill_1 FILLER_3_1835 ();
 sg13g2_decap_8 FILLER_3_1846 ();
 sg13g2_decap_8 FILLER_3_1853 ();
 sg13g2_fill_2 FILLER_3_1860 ();
 sg13g2_decap_4 FILLER_3_1888 ();
 sg13g2_fill_2 FILLER_3_1892 ();
 sg13g2_fill_1 FILLER_3_1919 ();
 sg13g2_fill_1 FILLER_3_1925 ();
 sg13g2_fill_1 FILLER_3_1956 ();
 sg13g2_fill_1 FILLER_3_1961 ();
 sg13g2_decap_8 FILLER_3_2014 ();
 sg13g2_decap_8 FILLER_3_2021 ();
 sg13g2_decap_8 FILLER_3_2028 ();
 sg13g2_decap_8 FILLER_3_2035 ();
 sg13g2_fill_1 FILLER_3_2042 ();
 sg13g2_fill_2 FILLER_3_2059 ();
 sg13g2_fill_1 FILLER_3_2072 ();
 sg13g2_fill_1 FILLER_3_2119 ();
 sg13g2_fill_1 FILLER_3_2125 ();
 sg13g2_fill_2 FILLER_3_2152 ();
 sg13g2_decap_8 FILLER_3_2196 ();
 sg13g2_decap_8 FILLER_3_2203 ();
 sg13g2_fill_2 FILLER_3_2210 ();
 sg13g2_fill_2 FILLER_3_2222 ();
 sg13g2_fill_1 FILLER_3_2224 ();
 sg13g2_decap_4 FILLER_3_2251 ();
 sg13g2_fill_2 FILLER_3_2255 ();
 sg13g2_decap_4 FILLER_3_2283 ();
 sg13g2_fill_1 FILLER_3_2287 ();
 sg13g2_decap_8 FILLER_3_2292 ();
 sg13g2_decap_8 FILLER_3_2299 ();
 sg13g2_decap_8 FILLER_3_2306 ();
 sg13g2_fill_1 FILLER_3_2313 ();
 sg13g2_decap_8 FILLER_3_2344 ();
 sg13g2_fill_1 FILLER_3_2351 ();
 sg13g2_decap_8 FILLER_3_2356 ();
 sg13g2_fill_2 FILLER_3_2405 ();
 sg13g2_decap_8 FILLER_3_2415 ();
 sg13g2_decap_8 FILLER_3_2422 ();
 sg13g2_decap_8 FILLER_3_2429 ();
 sg13g2_fill_1 FILLER_3_2446 ();
 sg13g2_fill_2 FILLER_3_2480 ();
 sg13g2_decap_4 FILLER_3_2486 ();
 sg13g2_decap_4 FILLER_3_2500 ();
 sg13g2_decap_4 FILLER_3_2508 ();
 sg13g2_fill_2 FILLER_3_2512 ();
 sg13g2_fill_1 FILLER_3_2518 ();
 sg13g2_decap_8 FILLER_3_2549 ();
 sg13g2_decap_8 FILLER_3_2556 ();
 sg13g2_decap_8 FILLER_3_2563 ();
 sg13g2_decap_8 FILLER_3_2570 ();
 sg13g2_decap_8 FILLER_3_2577 ();
 sg13g2_decap_8 FILLER_3_2584 ();
 sg13g2_decap_8 FILLER_3_2591 ();
 sg13g2_decap_8 FILLER_3_2598 ();
 sg13g2_decap_8 FILLER_3_2605 ();
 sg13g2_decap_8 FILLER_3_2612 ();
 sg13g2_decap_8 FILLER_3_2619 ();
 sg13g2_decap_8 FILLER_3_2626 ();
 sg13g2_decap_8 FILLER_3_2633 ();
 sg13g2_decap_8 FILLER_3_2640 ();
 sg13g2_decap_8 FILLER_3_2647 ();
 sg13g2_decap_8 FILLER_3_2654 ();
 sg13g2_decap_8 FILLER_3_2661 ();
 sg13g2_fill_2 FILLER_3_2668 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_decap_4 FILLER_4_9 ();
 sg13g2_fill_2 FILLER_4_30 ();
 sg13g2_decap_8 FILLER_4_78 ();
 sg13g2_decap_4 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_89 ();
 sg13g2_fill_1 FILLER_4_103 ();
 sg13g2_fill_1 FILLER_4_113 ();
 sg13g2_fill_1 FILLER_4_157 ();
 sg13g2_fill_2 FILLER_4_163 ();
 sg13g2_fill_2 FILLER_4_170 ();
 sg13g2_fill_1 FILLER_4_172 ();
 sg13g2_fill_2 FILLER_4_178 ();
 sg13g2_fill_1 FILLER_4_225 ();
 sg13g2_fill_2 FILLER_4_236 ();
 sg13g2_fill_2 FILLER_4_247 ();
 sg13g2_fill_1 FILLER_4_260 ();
 sg13g2_decap_8 FILLER_4_289 ();
 sg13g2_decap_8 FILLER_4_300 ();
 sg13g2_decap_8 FILLER_4_307 ();
 sg13g2_decap_4 FILLER_4_314 ();
 sg13g2_decap_4 FILLER_4_335 ();
 sg13g2_fill_1 FILLER_4_355 ();
 sg13g2_fill_2 FILLER_4_361 ();
 sg13g2_fill_2 FILLER_4_384 ();
 sg13g2_decap_8 FILLER_4_390 ();
 sg13g2_decap_8 FILLER_4_397 ();
 sg13g2_decap_4 FILLER_4_430 ();
 sg13g2_fill_1 FILLER_4_444 ();
 sg13g2_fill_2 FILLER_4_455 ();
 sg13g2_decap_4 FILLER_4_461 ();
 sg13g2_fill_1 FILLER_4_465 ();
 sg13g2_fill_1 FILLER_4_471 ();
 sg13g2_fill_1 FILLER_4_477 ();
 sg13g2_decap_4 FILLER_4_482 ();
 sg13g2_fill_2 FILLER_4_486 ();
 sg13g2_fill_2 FILLER_4_492 ();
 sg13g2_fill_1 FILLER_4_494 ();
 sg13g2_fill_1 FILLER_4_503 ();
 sg13g2_fill_1 FILLER_4_509 ();
 sg13g2_fill_2 FILLER_4_514 ();
 sg13g2_fill_2 FILLER_4_521 ();
 sg13g2_fill_2 FILLER_4_528 ();
 sg13g2_decap_8 FILLER_4_536 ();
 sg13g2_decap_8 FILLER_4_543 ();
 sg13g2_decap_8 FILLER_4_550 ();
 sg13g2_decap_4 FILLER_4_561 ();
 sg13g2_decap_8 FILLER_4_569 ();
 sg13g2_decap_8 FILLER_4_576 ();
 sg13g2_decap_4 FILLER_4_583 ();
 sg13g2_fill_1 FILLER_4_587 ();
 sg13g2_decap_8 FILLER_4_648 ();
 sg13g2_decap_8 FILLER_4_655 ();
 sg13g2_fill_1 FILLER_4_662 ();
 sg13g2_decap_4 FILLER_4_683 ();
 sg13g2_decap_8 FILLER_4_696 ();
 sg13g2_decap_8 FILLER_4_703 ();
 sg13g2_fill_2 FILLER_4_726 ();
 sg13g2_decap_8 FILLER_4_796 ();
 sg13g2_fill_2 FILLER_4_803 ();
 sg13g2_fill_1 FILLER_4_805 ();
 sg13g2_decap_4 FILLER_4_818 ();
 sg13g2_fill_2 FILLER_4_822 ();
 sg13g2_decap_8 FILLER_4_865 ();
 sg13g2_fill_2 FILLER_4_872 ();
 sg13g2_fill_2 FILLER_4_879 ();
 sg13g2_fill_1 FILLER_4_973 ();
 sg13g2_fill_2 FILLER_4_977 ();
 sg13g2_fill_1 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1035 ();
 sg13g2_fill_2 FILLER_4_1042 ();
 sg13g2_decap_8 FILLER_4_1049 ();
 sg13g2_fill_2 FILLER_4_1056 ();
 sg13g2_fill_1 FILLER_4_1128 ();
 sg13g2_fill_2 FILLER_4_1139 ();
 sg13g2_fill_1 FILLER_4_1141 ();
 sg13g2_fill_2 FILLER_4_1178 ();
 sg13g2_fill_2 FILLER_4_1190 ();
 sg13g2_fill_1 FILLER_4_1192 ();
 sg13g2_fill_2 FILLER_4_1199 ();
 sg13g2_fill_2 FILLER_4_1204 ();
 sg13g2_fill_1 FILLER_4_1206 ();
 sg13g2_fill_1 FILLER_4_1213 ();
 sg13g2_fill_1 FILLER_4_1234 ();
 sg13g2_decap_8 FILLER_4_1245 ();
 sg13g2_fill_1 FILLER_4_1281 ();
 sg13g2_fill_2 FILLER_4_1318 ();
 sg13g2_fill_2 FILLER_4_1325 ();
 sg13g2_decap_4 FILLER_4_1395 ();
 sg13g2_fill_1 FILLER_4_1409 ();
 sg13g2_decap_8 FILLER_4_1413 ();
 sg13g2_fill_1 FILLER_4_1420 ();
 sg13g2_decap_4 FILLER_4_1431 ();
 sg13g2_decap_4 FILLER_4_1477 ();
 sg13g2_fill_2 FILLER_4_1500 ();
 sg13g2_fill_1 FILLER_4_1502 ();
 sg13g2_decap_8 FILLER_4_1513 ();
 sg13g2_decap_4 FILLER_4_1520 ();
 sg13g2_fill_2 FILLER_4_1524 ();
 sg13g2_fill_1 FILLER_4_1536 ();
 sg13g2_fill_2 FILLER_4_1553 ();
 sg13g2_fill_1 FILLER_4_1610 ();
 sg13g2_decap_4 FILLER_4_1637 ();
 sg13g2_fill_1 FILLER_4_1671 ();
 sg13g2_decap_8 FILLER_4_1750 ();
 sg13g2_decap_8 FILLER_4_1757 ();
 sg13g2_fill_1 FILLER_4_1764 ();
 sg13g2_decap_8 FILLER_4_1772 ();
 sg13g2_decap_8 FILLER_4_1779 ();
 sg13g2_fill_2 FILLER_4_1786 ();
 sg13g2_fill_2 FILLER_4_1791 ();
 sg13g2_fill_1 FILLER_4_1806 ();
 sg13g2_decap_4 FILLER_4_1842 ();
 sg13g2_decap_4 FILLER_4_1882 ();
 sg13g2_fill_1 FILLER_4_1906 ();
 sg13g2_fill_2 FILLER_4_1942 ();
 sg13g2_decap_8 FILLER_4_1970 ();
 sg13g2_decap_4 FILLER_4_1977 ();
 sg13g2_fill_1 FILLER_4_1981 ();
 sg13g2_decap_8 FILLER_4_1998 ();
 sg13g2_decap_4 FILLER_4_2015 ();
 sg13g2_decap_8 FILLER_4_2045 ();
 sg13g2_decap_4 FILLER_4_2052 ();
 sg13g2_fill_1 FILLER_4_2080 ();
 sg13g2_fill_1 FILLER_4_2090 ();
 sg13g2_decap_4 FILLER_4_2117 ();
 sg13g2_fill_1 FILLER_4_2121 ();
 sg13g2_decap_8 FILLER_4_2127 ();
 sg13g2_decap_4 FILLER_4_2134 ();
 sg13g2_decap_4 FILLER_4_2142 ();
 sg13g2_fill_1 FILLER_4_2146 ();
 sg13g2_fill_1 FILLER_4_2159 ();
 sg13g2_fill_1 FILLER_4_2170 ();
 sg13g2_fill_1 FILLER_4_2199 ();
 sg13g2_fill_1 FILLER_4_2210 ();
 sg13g2_decap_4 FILLER_4_2260 ();
 sg13g2_fill_2 FILLER_4_2277 ();
 sg13g2_decap_8 FILLER_4_2309 ();
 sg13g2_decap_4 FILLER_4_2320 ();
 sg13g2_fill_1 FILLER_4_2324 ();
 sg13g2_decap_8 FILLER_4_2329 ();
 sg13g2_decap_4 FILLER_4_2336 ();
 sg13g2_fill_1 FILLER_4_2340 ();
 sg13g2_fill_1 FILLER_4_2371 ();
 sg13g2_fill_2 FILLER_4_2394 ();
 sg13g2_fill_2 FILLER_4_2400 ();
 sg13g2_decap_8 FILLER_4_2432 ();
 sg13g2_decap_4 FILLER_4_2439 ();
 sg13g2_fill_2 FILLER_4_2443 ();
 sg13g2_decap_8 FILLER_4_2475 ();
 sg13g2_decap_8 FILLER_4_2482 ();
 sg13g2_decap_8 FILLER_4_2489 ();
 sg13g2_decap_8 FILLER_4_2496 ();
 sg13g2_decap_8 FILLER_4_2503 ();
 sg13g2_decap_4 FILLER_4_2510 ();
 sg13g2_fill_2 FILLER_4_2514 ();
 sg13g2_decap_8 FILLER_4_2537 ();
 sg13g2_decap_8 FILLER_4_2544 ();
 sg13g2_decap_8 FILLER_4_2551 ();
 sg13g2_decap_8 FILLER_4_2558 ();
 sg13g2_decap_8 FILLER_4_2565 ();
 sg13g2_decap_8 FILLER_4_2572 ();
 sg13g2_decap_8 FILLER_4_2579 ();
 sg13g2_decap_8 FILLER_4_2586 ();
 sg13g2_decap_8 FILLER_4_2593 ();
 sg13g2_decap_8 FILLER_4_2600 ();
 sg13g2_decap_8 FILLER_4_2607 ();
 sg13g2_decap_8 FILLER_4_2614 ();
 sg13g2_decap_8 FILLER_4_2621 ();
 sg13g2_decap_8 FILLER_4_2628 ();
 sg13g2_decap_8 FILLER_4_2635 ();
 sg13g2_decap_8 FILLER_4_2642 ();
 sg13g2_decap_8 FILLER_4_2649 ();
 sg13g2_decap_8 FILLER_4_2656 ();
 sg13g2_decap_8 FILLER_4_2663 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_fill_2 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_34 ();
 sg13g2_decap_8 FILLER_5_41 ();
 sg13g2_decap_8 FILLER_5_48 ();
 sg13g2_decap_8 FILLER_5_55 ();
 sg13g2_fill_1 FILLER_5_62 ();
 sg13g2_fill_1 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_85 ();
 sg13g2_decap_4 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_96 ();
 sg13g2_fill_2 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_117 ();
 sg13g2_fill_1 FILLER_5_127 ();
 sg13g2_fill_1 FILLER_5_132 ();
 sg13g2_fill_1 FILLER_5_147 ();
 sg13g2_fill_1 FILLER_5_191 ();
 sg13g2_fill_1 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_221 ();
 sg13g2_fill_1 FILLER_5_227 ();
 sg13g2_fill_1 FILLER_5_233 ();
 sg13g2_fill_1 FILLER_5_239 ();
 sg13g2_fill_1 FILLER_5_272 ();
 sg13g2_decap_8 FILLER_5_288 ();
 sg13g2_fill_1 FILLER_5_295 ();
 sg13g2_decap_8 FILLER_5_299 ();
 sg13g2_decap_4 FILLER_5_306 ();
 sg13g2_fill_1 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_316 ();
 sg13g2_fill_1 FILLER_5_323 ();
 sg13g2_decap_8 FILLER_5_328 ();
 sg13g2_decap_4 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_344 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_fill_1 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_fill_1 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_fill_2 FILLER_5_408 ();
 sg13g2_fill_1 FILLER_5_410 ();
 sg13g2_fill_1 FILLER_5_415 ();
 sg13g2_decap_4 FILLER_5_446 ();
 sg13g2_decap_4 FILLER_5_455 ();
 sg13g2_fill_1 FILLER_5_488 ();
 sg13g2_fill_2 FILLER_5_529 ();
 sg13g2_fill_1 FILLER_5_531 ();
 sg13g2_fill_2 FILLER_5_572 ();
 sg13g2_fill_1 FILLER_5_574 ();
 sg13g2_decap_8 FILLER_5_579 ();
 sg13g2_fill_2 FILLER_5_586 ();
 sg13g2_fill_1 FILLER_5_603 ();
 sg13g2_fill_1 FILLER_5_609 ();
 sg13g2_decap_4 FILLER_5_615 ();
 sg13g2_fill_2 FILLER_5_619 ();
 sg13g2_fill_2 FILLER_5_626 ();
 sg13g2_fill_1 FILLER_5_628 ();
 sg13g2_decap_8 FILLER_5_637 ();
 sg13g2_decap_8 FILLER_5_644 ();
 sg13g2_decap_8 FILLER_5_651 ();
 sg13g2_decap_8 FILLER_5_658 ();
 sg13g2_decap_8 FILLER_5_665 ();
 sg13g2_decap_4 FILLER_5_672 ();
 sg13g2_fill_2 FILLER_5_676 ();
 sg13g2_fill_1 FILLER_5_689 ();
 sg13g2_fill_2 FILLER_5_719 ();
 sg13g2_fill_2 FILLER_5_785 ();
 sg13g2_fill_1 FILLER_5_787 ();
 sg13g2_decap_4 FILLER_5_802 ();
 sg13g2_fill_2 FILLER_5_806 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_857 ();
 sg13g2_decap_4 FILLER_5_864 ();
 sg13g2_fill_2 FILLER_5_868 ();
 sg13g2_decap_8 FILLER_5_874 ();
 sg13g2_fill_2 FILLER_5_881 ();
 sg13g2_fill_1 FILLER_5_883 ();
 sg13g2_fill_2 FILLER_5_894 ();
 sg13g2_fill_2 FILLER_5_914 ();
 sg13g2_fill_2 FILLER_5_930 ();
 sg13g2_fill_2 FILLER_5_958 ();
 sg13g2_fill_1 FILLER_5_1006 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_decap_8 FILLER_5_1026 ();
 sg13g2_decap_8 FILLER_5_1033 ();
 sg13g2_decap_8 FILLER_5_1040 ();
 sg13g2_decap_8 FILLER_5_1047 ();
 sg13g2_decap_8 FILLER_5_1054 ();
 sg13g2_decap_8 FILLER_5_1061 ();
 sg13g2_decap_8 FILLER_5_1068 ();
 sg13g2_decap_8 FILLER_5_1075 ();
 sg13g2_decap_8 FILLER_5_1082 ();
 sg13g2_decap_8 FILLER_5_1089 ();
 sg13g2_decap_8 FILLER_5_1096 ();
 sg13g2_decap_8 FILLER_5_1103 ();
 sg13g2_decap_4 FILLER_5_1110 ();
 sg13g2_fill_2 FILLER_5_1114 ();
 sg13g2_decap_8 FILLER_5_1121 ();
 sg13g2_decap_8 FILLER_5_1128 ();
 sg13g2_decap_4 FILLER_5_1135 ();
 sg13g2_fill_1 FILLER_5_1139 ();
 sg13g2_decap_8 FILLER_5_1150 ();
 sg13g2_decap_4 FILLER_5_1157 ();
 sg13g2_fill_1 FILLER_5_1161 ();
 sg13g2_decap_4 FILLER_5_1193 ();
 sg13g2_fill_1 FILLER_5_1197 ();
 sg13g2_decap_8 FILLER_5_1216 ();
 sg13g2_decap_8 FILLER_5_1223 ();
 sg13g2_fill_2 FILLER_5_1230 ();
 sg13g2_fill_1 FILLER_5_1232 ();
 sg13g2_decap_8 FILLER_5_1238 ();
 sg13g2_decap_4 FILLER_5_1245 ();
 sg13g2_fill_2 FILLER_5_1260 ();
 sg13g2_fill_1 FILLER_5_1262 ();
 sg13g2_fill_2 FILLER_5_1269 ();
 sg13g2_decap_8 FILLER_5_1281 ();
 sg13g2_fill_1 FILLER_5_1301 ();
 sg13g2_decap_4 FILLER_5_1328 ();
 sg13g2_decap_4 FILLER_5_1342 ();
 sg13g2_fill_1 FILLER_5_1346 ();
 sg13g2_fill_1 FILLER_5_1353 ();
 sg13g2_fill_2 FILLER_5_1364 ();
 sg13g2_decap_8 FILLER_5_1398 ();
 sg13g2_fill_2 FILLER_5_1405 ();
 sg13g2_fill_1 FILLER_5_1416 ();
 sg13g2_fill_1 FILLER_5_1430 ();
 sg13g2_fill_1 FILLER_5_1460 ();
 sg13g2_fill_1 FILLER_5_1467 ();
 sg13g2_decap_8 FILLER_5_1496 ();
 sg13g2_fill_2 FILLER_5_1503 ();
 sg13g2_decap_8 FILLER_5_1541 ();
 sg13g2_fill_1 FILLER_5_1548 ();
 sg13g2_decap_8 FILLER_5_1591 ();
 sg13g2_decap_8 FILLER_5_1598 ();
 sg13g2_decap_8 FILLER_5_1605 ();
 sg13g2_decap_8 FILLER_5_1612 ();
 sg13g2_decap_8 FILLER_5_1619 ();
 sg13g2_fill_1 FILLER_5_1626 ();
 sg13g2_fill_1 FILLER_5_1666 ();
 sg13g2_fill_1 FILLER_5_1714 ();
 sg13g2_decap_8 FILLER_5_1734 ();
 sg13g2_decap_8 FILLER_5_1741 ();
 sg13g2_decap_8 FILLER_5_1748 ();
 sg13g2_decap_8 FILLER_5_1755 ();
 sg13g2_fill_2 FILLER_5_1762 ();
 sg13g2_fill_1 FILLER_5_1764 ();
 sg13g2_fill_2 FILLER_5_1768 ();
 sg13g2_fill_1 FILLER_5_1770 ();
 sg13g2_decap_4 FILLER_5_1776 ();
 sg13g2_fill_2 FILLER_5_1780 ();
 sg13g2_fill_2 FILLER_5_1791 ();
 sg13g2_decap_4 FILLER_5_1798 ();
 sg13g2_fill_1 FILLER_5_1802 ();
 sg13g2_decap_8 FILLER_5_1812 ();
 sg13g2_fill_1 FILLER_5_1819 ();
 sg13g2_decap_8 FILLER_5_1830 ();
 sg13g2_fill_1 FILLER_5_1837 ();
 sg13g2_decap_8 FILLER_5_1873 ();
 sg13g2_fill_2 FILLER_5_1880 ();
 sg13g2_fill_2 FILLER_5_1895 ();
 sg13g2_fill_1 FILLER_5_1897 ();
 sg13g2_fill_2 FILLER_5_1933 ();
 sg13g2_decap_4 FILLER_5_1963 ();
 sg13g2_fill_2 FILLER_5_1977 ();
 sg13g2_decap_8 FILLER_5_2011 ();
 sg13g2_decap_4 FILLER_5_2018 ();
 sg13g2_fill_2 FILLER_5_2067 ();
 sg13g2_fill_2 FILLER_5_2091 ();
 sg13g2_fill_1 FILLER_5_2099 ();
 sg13g2_decap_4 FILLER_5_2117 ();
 sg13g2_fill_2 FILLER_5_2121 ();
 sg13g2_fill_1 FILLER_5_2164 ();
 sg13g2_fill_1 FILLER_5_2217 ();
 sg13g2_fill_1 FILLER_5_2224 ();
 sg13g2_fill_1 FILLER_5_2272 ();
 sg13g2_decap_8 FILLER_5_2276 ();
 sg13g2_decap_8 FILLER_5_2283 ();
 sg13g2_decap_8 FILLER_5_2290 ();
 sg13g2_decap_8 FILLER_5_2297 ();
 sg13g2_fill_2 FILLER_5_2304 ();
 sg13g2_fill_1 FILLER_5_2306 ();
 sg13g2_fill_1 FILLER_5_2310 ();
 sg13g2_decap_8 FILLER_5_2315 ();
 sg13g2_decap_8 FILLER_5_2322 ();
 sg13g2_decap_8 FILLER_5_2329 ();
 sg13g2_decap_8 FILLER_5_2336 ();
 sg13g2_decap_8 FILLER_5_2343 ();
 sg13g2_fill_2 FILLER_5_2354 ();
 sg13g2_decap_8 FILLER_5_2359 ();
 sg13g2_fill_2 FILLER_5_2366 ();
 sg13g2_fill_1 FILLER_5_2368 ();
 sg13g2_fill_2 FILLER_5_2381 ();
 sg13g2_decap_8 FILLER_5_2443 ();
 sg13g2_decap_8 FILLER_5_2467 ();
 sg13g2_decap_8 FILLER_5_2474 ();
 sg13g2_decap_8 FILLER_5_2481 ();
 sg13g2_decap_4 FILLER_5_2488 ();
 sg13g2_fill_2 FILLER_5_2492 ();
 sg13g2_decap_8 FILLER_5_2498 ();
 sg13g2_decap_8 FILLER_5_2505 ();
 sg13g2_decap_4 FILLER_5_2512 ();
 sg13g2_fill_2 FILLER_5_2516 ();
 sg13g2_fill_1 FILLER_5_2532 ();
 sg13g2_decap_8 FILLER_5_2563 ();
 sg13g2_decap_8 FILLER_5_2570 ();
 sg13g2_decap_8 FILLER_5_2577 ();
 sg13g2_decap_8 FILLER_5_2584 ();
 sg13g2_decap_4 FILLER_5_2591 ();
 sg13g2_fill_1 FILLER_5_2595 ();
 sg13g2_decap_8 FILLER_5_2600 ();
 sg13g2_decap_8 FILLER_5_2607 ();
 sg13g2_decap_8 FILLER_5_2614 ();
 sg13g2_decap_8 FILLER_5_2621 ();
 sg13g2_decap_8 FILLER_5_2628 ();
 sg13g2_decap_8 FILLER_5_2635 ();
 sg13g2_decap_8 FILLER_5_2642 ();
 sg13g2_decap_8 FILLER_5_2649 ();
 sg13g2_decap_8 FILLER_5_2656 ();
 sg13g2_decap_8 FILLER_5_2663 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_4 FILLER_6_7 ();
 sg13g2_fill_1 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_38 ();
 sg13g2_decap_8 FILLER_6_45 ();
 sg13g2_fill_1 FILLER_6_52 ();
 sg13g2_decap_8 FILLER_6_83 ();
 sg13g2_decap_4 FILLER_6_90 ();
 sg13g2_fill_2 FILLER_6_94 ();
 sg13g2_fill_1 FILLER_6_100 ();
 sg13g2_fill_1 FILLER_6_114 ();
 sg13g2_fill_2 FILLER_6_119 ();
 sg13g2_fill_2 FILLER_6_141 ();
 sg13g2_fill_2 FILLER_6_166 ();
 sg13g2_fill_1 FILLER_6_177 ();
 sg13g2_fill_2 FILLER_6_186 ();
 sg13g2_fill_1 FILLER_6_188 ();
 sg13g2_fill_1 FILLER_6_195 ();
 sg13g2_fill_2 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_209 ();
 sg13g2_fill_1 FILLER_6_222 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_267 ();
 sg13g2_fill_1 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_decap_8 FILLER_6_298 ();
 sg13g2_decap_8 FILLER_6_305 ();
 sg13g2_decap_8 FILLER_6_312 ();
 sg13g2_decap_4 FILLER_6_319 ();
 sg13g2_fill_1 FILLER_6_323 ();
 sg13g2_fill_1 FILLER_6_328 ();
 sg13g2_decap_8 FILLER_6_334 ();
 sg13g2_decap_4 FILLER_6_341 ();
 sg13g2_fill_1 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_362 ();
 sg13g2_decap_4 FILLER_6_369 ();
 sg13g2_fill_1 FILLER_6_373 ();
 sg13g2_fill_1 FILLER_6_379 ();
 sg13g2_decap_4 FILLER_6_398 ();
 sg13g2_fill_2 FILLER_6_402 ();
 sg13g2_decap_8 FILLER_6_415 ();
 sg13g2_decap_8 FILLER_6_422 ();
 sg13g2_decap_4 FILLER_6_429 ();
 sg13g2_fill_1 FILLER_6_433 ();
 sg13g2_fill_1 FILLER_6_444 ();
 sg13g2_fill_1 FILLER_6_464 ();
 sg13g2_fill_1 FILLER_6_483 ();
 sg13g2_fill_1 FILLER_6_489 ();
 sg13g2_fill_1 FILLER_6_494 ();
 sg13g2_fill_1 FILLER_6_498 ();
 sg13g2_fill_1 FILLER_6_508 ();
 sg13g2_fill_1 FILLER_6_518 ();
 sg13g2_fill_1 FILLER_6_523 ();
 sg13g2_fill_1 FILLER_6_529 ();
 sg13g2_fill_2 FILLER_6_534 ();
 sg13g2_decap_4 FILLER_6_546 ();
 sg13g2_fill_1 FILLER_6_550 ();
 sg13g2_decap_8 FILLER_6_559 ();
 sg13g2_decap_8 FILLER_6_566 ();
 sg13g2_decap_8 FILLER_6_573 ();
 sg13g2_fill_1 FILLER_6_580 ();
 sg13g2_fill_2 FILLER_6_625 ();
 sg13g2_decap_4 FILLER_6_635 ();
 sg13g2_fill_2 FILLER_6_639 ();
 sg13g2_fill_2 FILLER_6_667 ();
 sg13g2_fill_1 FILLER_6_696 ();
 sg13g2_fill_1 FILLER_6_744 ();
 sg13g2_fill_2 FILLER_6_761 ();
 sg13g2_decap_8 FILLER_6_810 ();
 sg13g2_decap_8 FILLER_6_817 ();
 sg13g2_fill_2 FILLER_6_824 ();
 sg13g2_fill_1 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_fill_2 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_862 ();
 sg13g2_decap_4 FILLER_6_869 ();
 sg13g2_fill_2 FILLER_6_873 ();
 sg13g2_fill_1 FILLER_6_910 ();
 sg13g2_fill_1 FILLER_6_922 ();
 sg13g2_fill_2 FILLER_6_929 ();
 sg13g2_fill_1 FILLER_6_941 ();
 sg13g2_fill_2 FILLER_6_948 ();
 sg13g2_fill_1 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_1030 ();
 sg13g2_decap_8 FILLER_6_1037 ();
 sg13g2_decap_8 FILLER_6_1044 ();
 sg13g2_decap_8 FILLER_6_1051 ();
 sg13g2_decap_4 FILLER_6_1058 ();
 sg13g2_fill_1 FILLER_6_1062 ();
 sg13g2_decap_8 FILLER_6_1076 ();
 sg13g2_fill_2 FILLER_6_1104 ();
 sg13g2_fill_1 FILLER_6_1109 ();
 sg13g2_fill_2 FILLER_6_1117 ();
 sg13g2_decap_8 FILLER_6_1156 ();
 sg13g2_decap_8 FILLER_6_1163 ();
 sg13g2_decap_8 FILLER_6_1170 ();
 sg13g2_decap_4 FILLER_6_1177 ();
 sg13g2_decap_4 FILLER_6_1200 ();
 sg13g2_decap_4 FILLER_6_1236 ();
 sg13g2_fill_2 FILLER_6_1240 ();
 sg13g2_decap_8 FILLER_6_1299 ();
 sg13g2_decap_8 FILLER_6_1306 ();
 sg13g2_fill_1 FILLER_6_1313 ();
 sg13g2_decap_8 FILLER_6_1320 ();
 sg13g2_decap_8 FILLER_6_1327 ();
 sg13g2_decap_4 FILLER_6_1366 ();
 sg13g2_decap_4 FILLER_6_1380 ();
 sg13g2_decap_8 FILLER_6_1425 ();
 sg13g2_decap_8 FILLER_6_1432 ();
 sg13g2_fill_2 FILLER_6_1439 ();
 sg13g2_fill_1 FILLER_6_1441 ();
 sg13g2_fill_1 FILLER_6_1480 ();
 sg13g2_decap_8 FILLER_6_1492 ();
 sg13g2_decap_4 FILLER_6_1499 ();
 sg13g2_fill_2 FILLER_6_1503 ();
 sg13g2_fill_1 FILLER_6_1541 ();
 sg13g2_fill_1 FILLER_6_1557 ();
 sg13g2_fill_2 FILLER_6_1561 ();
 sg13g2_fill_1 FILLER_6_1563 ();
 sg13g2_decap_4 FILLER_6_1570 ();
 sg13g2_decap_8 FILLER_6_1604 ();
 sg13g2_decap_8 FILLER_6_1611 ();
 sg13g2_fill_1 FILLER_6_1618 ();
 sg13g2_fill_1 FILLER_6_1634 ();
 sg13g2_fill_1 FILLER_6_1638 ();
 sg13g2_fill_2 FILLER_6_1662 ();
 sg13g2_fill_2 FILLER_6_1680 ();
 sg13g2_fill_2 FILLER_6_1706 ();
 sg13g2_decap_8 FILLER_6_1747 ();
 sg13g2_decap_8 FILLER_6_1754 ();
 sg13g2_decap_8 FILLER_6_1761 ();
 sg13g2_decap_4 FILLER_6_1768 ();
 sg13g2_decap_4 FILLER_6_1780 ();
 sg13g2_fill_1 FILLER_6_1784 ();
 sg13g2_decap_8 FILLER_6_1839 ();
 sg13g2_decap_4 FILLER_6_1846 ();
 sg13g2_decap_8 FILLER_6_1854 ();
 sg13g2_decap_4 FILLER_6_1861 ();
 sg13g2_fill_1 FILLER_6_1865 ();
 sg13g2_decap_8 FILLER_6_1874 ();
 sg13g2_decap_8 FILLER_6_1881 ();
 sg13g2_fill_1 FILLER_6_1888 ();
 sg13g2_fill_2 FILLER_6_1948 ();
 sg13g2_fill_2 FILLER_6_1986 ();
 sg13g2_fill_2 FILLER_6_1998 ();
 sg13g2_fill_1 FILLER_6_2005 ();
 sg13g2_decap_8 FILLER_6_2043 ();
 sg13g2_decap_8 FILLER_6_2050 ();
 sg13g2_fill_1 FILLER_6_2057 ();
 sg13g2_fill_2 FILLER_6_2133 ();
 sg13g2_fill_1 FILLER_6_2159 ();
 sg13g2_fill_1 FILLER_6_2195 ();
 sg13g2_fill_1 FILLER_6_2213 ();
 sg13g2_fill_2 FILLER_6_2235 ();
 sg13g2_fill_2 FILLER_6_2246 ();
 sg13g2_decap_4 FILLER_6_2340 ();
 sg13g2_fill_2 FILLER_6_2344 ();
 sg13g2_fill_2 FILLER_6_2384 ();
 sg13g2_decap_8 FILLER_6_2425 ();
 sg13g2_decap_8 FILLER_6_2432 ();
 sg13g2_decap_8 FILLER_6_2439 ();
 sg13g2_fill_2 FILLER_6_2446 ();
 sg13g2_fill_1 FILLER_6_2466 ();
 sg13g2_fill_1 FILLER_6_2475 ();
 sg13g2_fill_2 FILLER_6_2484 ();
 sg13g2_fill_2 FILLER_6_2546 ();
 sg13g2_decap_8 FILLER_6_2574 ();
 sg13g2_decap_4 FILLER_6_2581 ();
 sg13g2_decap_8 FILLER_6_2615 ();
 sg13g2_decap_8 FILLER_6_2622 ();
 sg13g2_decap_8 FILLER_6_2629 ();
 sg13g2_decap_8 FILLER_6_2636 ();
 sg13g2_decap_8 FILLER_6_2643 ();
 sg13g2_decap_8 FILLER_6_2650 ();
 sg13g2_decap_8 FILLER_6_2657 ();
 sg13g2_decap_4 FILLER_6_2664 ();
 sg13g2_fill_2 FILLER_6_2668 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_7 ();
 sg13g2_fill_1 FILLER_7_9 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_4 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_36 ();
 sg13g2_decap_4 FILLER_7_43 ();
 sg13g2_fill_2 FILLER_7_47 ();
 sg13g2_decap_8 FILLER_7_78 ();
 sg13g2_decap_8 FILLER_7_85 ();
 sg13g2_fill_1 FILLER_7_92 ();
 sg13g2_fill_1 FILLER_7_114 ();
 sg13g2_fill_2 FILLER_7_127 ();
 sg13g2_fill_2 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_2 FILLER_7_162 ();
 sg13g2_fill_2 FILLER_7_173 ();
 sg13g2_fill_1 FILLER_7_175 ();
 sg13g2_fill_2 FILLER_7_180 ();
 sg13g2_fill_1 FILLER_7_182 ();
 sg13g2_decap_4 FILLER_7_188 ();
 sg13g2_fill_1 FILLER_7_192 ();
 sg13g2_decap_8 FILLER_7_202 ();
 sg13g2_fill_2 FILLER_7_209 ();
 sg13g2_fill_1 FILLER_7_211 ();
 sg13g2_fill_2 FILLER_7_232 ();
 sg13g2_fill_1 FILLER_7_234 ();
 sg13g2_fill_2 FILLER_7_244 ();
 sg13g2_fill_1 FILLER_7_246 ();
 sg13g2_decap_4 FILLER_7_253 ();
 sg13g2_fill_1 FILLER_7_257 ();
 sg13g2_fill_1 FILLER_7_267 ();
 sg13g2_fill_1 FILLER_7_273 ();
 sg13g2_fill_1 FILLER_7_279 ();
 sg13g2_fill_1 FILLER_7_283 ();
 sg13g2_fill_1 FILLER_7_290 ();
 sg13g2_fill_1 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_335 ();
 sg13g2_fill_2 FILLER_7_342 ();
 sg13g2_fill_1 FILLER_7_344 ();
 sg13g2_fill_2 FILLER_7_353 ();
 sg13g2_decap_4 FILLER_7_398 ();
 sg13g2_fill_1 FILLER_7_402 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_decap_8 FILLER_7_427 ();
 sg13g2_decap_8 FILLER_7_434 ();
 sg13g2_decap_8 FILLER_7_441 ();
 sg13g2_fill_2 FILLER_7_448 ();
 sg13g2_fill_1 FILLER_7_450 ();
 sg13g2_fill_1 FILLER_7_477 ();
 sg13g2_fill_1 FILLER_7_488 ();
 sg13g2_fill_1 FILLER_7_517 ();
 sg13g2_decap_8 FILLER_7_532 ();
 sg13g2_decap_8 FILLER_7_539 ();
 sg13g2_decap_8 FILLER_7_546 ();
 sg13g2_decap_8 FILLER_7_557 ();
 sg13g2_decap_4 FILLER_7_564 ();
 sg13g2_fill_2 FILLER_7_568 ();
 sg13g2_decap_8 FILLER_7_574 ();
 sg13g2_decap_4 FILLER_7_581 ();
 sg13g2_fill_1 FILLER_7_585 ();
 sg13g2_fill_2 FILLER_7_622 ();
 sg13g2_fill_1 FILLER_7_624 ();
 sg13g2_decap_8 FILLER_7_651 ();
 sg13g2_fill_2 FILLER_7_658 ();
 sg13g2_fill_1 FILLER_7_660 ();
 sg13g2_fill_1 FILLER_7_683 ();
 sg13g2_decap_4 FILLER_7_735 ();
 sg13g2_decap_8 FILLER_7_785 ();
 sg13g2_fill_2 FILLER_7_818 ();
 sg13g2_decap_8 FILLER_7_826 ();
 sg13g2_fill_2 FILLER_7_862 ();
 sg13g2_fill_1 FILLER_7_864 ();
 sg13g2_decap_8 FILLER_7_875 ();
 sg13g2_decap_8 FILLER_7_885 ();
 sg13g2_decap_8 FILLER_7_892 ();
 sg13g2_fill_1 FILLER_7_944 ();
 sg13g2_fill_1 FILLER_7_963 ();
 sg13g2_fill_1 FILLER_7_977 ();
 sg13g2_fill_2 FILLER_7_1018 ();
 sg13g2_decap_8 FILLER_7_1056 ();
 sg13g2_decap_8 FILLER_7_1063 ();
 sg13g2_decap_4 FILLER_7_1070 ();
 sg13g2_fill_2 FILLER_7_1074 ();
 sg13g2_fill_2 FILLER_7_1112 ();
 sg13g2_decap_8 FILLER_7_1140 ();
 sg13g2_decap_8 FILLER_7_1147 ();
 sg13g2_decap_8 FILLER_7_1154 ();
 sg13g2_decap_8 FILLER_7_1161 ();
 sg13g2_fill_2 FILLER_7_1168 ();
 sg13g2_decap_8 FILLER_7_1173 ();
 sg13g2_fill_1 FILLER_7_1190 ();
 sg13g2_fill_1 FILLER_7_1233 ();
 sg13g2_decap_8 FILLER_7_1257 ();
 sg13g2_fill_2 FILLER_7_1264 ();
 sg13g2_fill_1 FILLER_7_1266 ();
 sg13g2_decap_8 FILLER_7_1280 ();
 sg13g2_fill_1 FILLER_7_1287 ();
 sg13g2_decap_8 FILLER_7_1320 ();
 sg13g2_decap_8 FILLER_7_1327 ();
 sg13g2_decap_4 FILLER_7_1334 ();
 sg13g2_decap_8 FILLER_7_1348 ();
 sg13g2_decap_8 FILLER_7_1355 ();
 sg13g2_fill_2 FILLER_7_1362 ();
 sg13g2_decap_8 FILLER_7_1369 ();
 sg13g2_decap_8 FILLER_7_1376 ();
 sg13g2_fill_1 FILLER_7_1383 ();
 sg13g2_fill_1 FILLER_7_1390 ();
 sg13g2_fill_1 FILLER_7_1430 ();
 sg13g2_decap_4 FILLER_7_1441 ();
 sg13g2_fill_2 FILLER_7_1466 ();
 sg13g2_decap_4 FILLER_7_1500 ();
 sg13g2_decap_8 FILLER_7_1530 ();
 sg13g2_fill_1 FILLER_7_1537 ();
 sg13g2_fill_2 FILLER_7_1550 ();
 sg13g2_decap_8 FILLER_7_1578 ();
 sg13g2_fill_2 FILLER_7_1594 ();
 sg13g2_decap_8 FILLER_7_1602 ();
 sg13g2_decap_4 FILLER_7_1609 ();
 sg13g2_fill_1 FILLER_7_1613 ();
 sg13g2_decap_4 FILLER_7_1617 ();
 sg13g2_fill_2 FILLER_7_1621 ();
 sg13g2_fill_2 FILLER_7_1685 ();
 sg13g2_decap_8 FILLER_7_1749 ();
 sg13g2_fill_2 FILLER_7_1756 ();
 sg13g2_fill_1 FILLER_7_1791 ();
 sg13g2_fill_1 FILLER_7_1855 ();
 sg13g2_fill_1 FILLER_7_1901 ();
 sg13g2_fill_2 FILLER_7_1988 ();
 sg13g2_decap_4 FILLER_7_2029 ();
 sg13g2_fill_2 FILLER_7_2037 ();
 sg13g2_decap_4 FILLER_7_2048 ();
 sg13g2_fill_1 FILLER_7_2176 ();
 sg13g2_decap_4 FILLER_7_2419 ();
 sg13g2_fill_1 FILLER_7_2423 ();
 sg13g2_decap_8 FILLER_7_2497 ();
 sg13g2_decap_8 FILLER_7_2504 ();
 sg13g2_decap_8 FILLER_7_2511 ();
 sg13g2_decap_4 FILLER_7_2518 ();
 sg13g2_fill_1 FILLER_7_2522 ();
 sg13g2_fill_2 FILLER_7_2532 ();
 sg13g2_decap_4 FILLER_7_2573 ();
 sg13g2_fill_1 FILLER_7_2577 ();
 sg13g2_decap_8 FILLER_7_2586 ();
 sg13g2_decap_8 FILLER_7_2593 ();
 sg13g2_decap_8 FILLER_7_2600 ();
 sg13g2_decap_8 FILLER_7_2607 ();
 sg13g2_decap_8 FILLER_7_2614 ();
 sg13g2_decap_8 FILLER_7_2621 ();
 sg13g2_decap_8 FILLER_7_2628 ();
 sg13g2_decap_8 FILLER_7_2635 ();
 sg13g2_decap_8 FILLER_7_2642 ();
 sg13g2_decap_8 FILLER_7_2649 ();
 sg13g2_decap_8 FILLER_7_2656 ();
 sg13g2_decap_8 FILLER_7_2663 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_1 FILLER_8_7 ();
 sg13g2_fill_1 FILLER_8_16 ();
 sg13g2_fill_1 FILLER_8_21 ();
 sg13g2_fill_2 FILLER_8_48 ();
 sg13g2_decap_4 FILLER_8_84 ();
 sg13g2_fill_2 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_104 ();
 sg13g2_fill_2 FILLER_8_141 ();
 sg13g2_fill_1 FILLER_8_143 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_156 ();
 sg13g2_fill_1 FILLER_8_162 ();
 sg13g2_fill_2 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_176 ();
 sg13g2_fill_1 FILLER_8_181 ();
 sg13g2_fill_1 FILLER_8_187 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_4 FILLER_8_205 ();
 sg13g2_fill_1 FILLER_8_230 ();
 sg13g2_fill_1 FILLER_8_246 ();
 sg13g2_fill_2 FILLER_8_250 ();
 sg13g2_decap_4 FILLER_8_262 ();
 sg13g2_decap_4 FILLER_8_275 ();
 sg13g2_fill_1 FILLER_8_279 ();
 sg13g2_decap_4 FILLER_8_285 ();
 sg13g2_fill_1 FILLER_8_289 ();
 sg13g2_decap_4 FILLER_8_294 ();
 sg13g2_fill_2 FILLER_8_306 ();
 sg13g2_fill_2 FILLER_8_313 ();
 sg13g2_fill_1 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_339 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_fill_1 FILLER_8_360 ();
 sg13g2_fill_2 FILLER_8_365 ();
 sg13g2_fill_1 FILLER_8_375 ();
 sg13g2_fill_1 FILLER_8_380 ();
 sg13g2_fill_1 FILLER_8_386 ();
 sg13g2_fill_1 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_fill_1 FILLER_8_448 ();
 sg13g2_decap_4 FILLER_8_454 ();
 sg13g2_fill_2 FILLER_8_514 ();
 sg13g2_fill_1 FILLER_8_516 ();
 sg13g2_fill_1 FILLER_8_524 ();
 sg13g2_fill_1 FILLER_8_530 ();
 sg13g2_fill_1 FILLER_8_540 ();
 sg13g2_fill_1 FILLER_8_575 ();
 sg13g2_fill_2 FILLER_8_581 ();
 sg13g2_fill_1 FILLER_8_583 ();
 sg13g2_decap_4 FILLER_8_610 ();
 sg13g2_fill_1 FILLER_8_614 ();
 sg13g2_fill_1 FILLER_8_620 ();
 sg13g2_fill_2 FILLER_8_661 ();
 sg13g2_fill_2 FILLER_8_668 ();
 sg13g2_fill_2 FILLER_8_688 ();
 sg13g2_fill_2 FILLER_8_706 ();
 sg13g2_decap_4 FILLER_8_713 ();
 sg13g2_fill_2 FILLER_8_743 ();
 sg13g2_fill_2 FILLER_8_761 ();
 sg13g2_fill_2 FILLER_8_789 ();
 sg13g2_decap_8 FILLER_8_801 ();
 sg13g2_decap_4 FILLER_8_808 ();
 sg13g2_decap_4 FILLER_8_818 ();
 sg13g2_fill_2 FILLER_8_825 ();
 sg13g2_decap_8 FILLER_8_843 ();
 sg13g2_fill_2 FILLER_8_850 ();
 sg13g2_fill_2 FILLER_8_917 ();
 sg13g2_fill_2 FILLER_8_979 ();
 sg13g2_fill_1 FILLER_8_993 ();
 sg13g2_fill_2 FILLER_8_1007 ();
 sg13g2_fill_1 FILLER_8_1018 ();
 sg13g2_fill_2 FILLER_8_1028 ();
 sg13g2_decap_4 FILLER_8_1066 ();
 sg13g2_fill_2 FILLER_8_1114 ();
 sg13g2_fill_2 FILLER_8_1126 ();
 sg13g2_fill_1 FILLER_8_1128 ();
 sg13g2_fill_2 FILLER_8_1135 ();
 sg13g2_fill_1 FILLER_8_1137 ();
 sg13g2_fill_2 FILLER_8_1163 ();
 sg13g2_fill_1 FILLER_8_1191 ();
 sg13g2_fill_2 FILLER_8_1222 ();
 sg13g2_fill_2 FILLER_8_1260 ();
 sg13g2_decap_8 FILLER_8_1288 ();
 sg13g2_decap_4 FILLER_8_1295 ();
 sg13g2_decap_4 FILLER_8_1312 ();
 sg13g2_fill_2 FILLER_8_1316 ();
 sg13g2_fill_2 FILLER_8_1328 ();
 sg13g2_decap_8 FILLER_8_1356 ();
 sg13g2_fill_1 FILLER_8_1363 ();
 sg13g2_fill_2 FILLER_8_1377 ();
 sg13g2_fill_2 FILLER_8_1387 ();
 sg13g2_fill_2 FILLER_8_1453 ();
 sg13g2_fill_2 FILLER_8_1510 ();
 sg13g2_fill_1 FILLER_8_1512 ();
 sg13g2_decap_8 FILLER_8_1516 ();
 sg13g2_decap_4 FILLER_8_1523 ();
 sg13g2_decap_4 FILLER_8_1567 ();
 sg13g2_fill_1 FILLER_8_1571 ();
 sg13g2_fill_2 FILLER_8_1602 ();
 sg13g2_fill_1 FILLER_8_1617 ();
 sg13g2_fill_2 FILLER_8_1644 ();
 sg13g2_fill_1 FILLER_8_1672 ();
 sg13g2_fill_2 FILLER_8_1703 ();
 sg13g2_fill_1 FILLER_8_1718 ();
 sg13g2_decap_8 FILLER_8_1723 ();
 sg13g2_decap_4 FILLER_8_1730 ();
 sg13g2_fill_2 FILLER_8_1760 ();
 sg13g2_fill_1 FILLER_8_1762 ();
 sg13g2_fill_1 FILLER_8_1768 ();
 sg13g2_fill_2 FILLER_8_1773 ();
 sg13g2_fill_1 FILLER_8_1775 ();
 sg13g2_fill_2 FILLER_8_1780 ();
 sg13g2_fill_1 FILLER_8_1782 ();
 sg13g2_fill_1 FILLER_8_1829 ();
 sg13g2_fill_1 FILLER_8_1879 ();
 sg13g2_fill_1 FILLER_8_1915 ();
 sg13g2_fill_2 FILLER_8_1922 ();
 sg13g2_fill_1 FILLER_8_1930 ();
 sg13g2_fill_1 FILLER_8_1945 ();
 sg13g2_fill_1 FILLER_8_1975 ();
 sg13g2_fill_2 FILLER_8_2013 ();
 sg13g2_fill_1 FILLER_8_2015 ();
 sg13g2_fill_1 FILLER_8_2067 ();
 sg13g2_fill_2 FILLER_8_2078 ();
 sg13g2_fill_1 FILLER_8_2099 ();
 sg13g2_fill_1 FILLER_8_2126 ();
 sg13g2_fill_2 FILLER_8_2148 ();
 sg13g2_fill_1 FILLER_8_2182 ();
 sg13g2_fill_2 FILLER_8_2193 ();
 sg13g2_fill_2 FILLER_8_2238 ();
 sg13g2_fill_1 FILLER_8_2259 ();
 sg13g2_fill_2 FILLER_8_2301 ();
 sg13g2_fill_1 FILLER_8_2313 ();
 sg13g2_fill_1 FILLER_8_2351 ();
 sg13g2_fill_1 FILLER_8_2389 ();
 sg13g2_fill_2 FILLER_8_2400 ();
 sg13g2_fill_1 FILLER_8_2402 ();
 sg13g2_fill_2 FILLER_8_2407 ();
 sg13g2_fill_2 FILLER_8_2415 ();
 sg13g2_fill_2 FILLER_8_2423 ();
 sg13g2_fill_2 FILLER_8_2429 ();
 sg13g2_fill_2 FILLER_8_2460 ();
 sg13g2_fill_1 FILLER_8_2501 ();
 sg13g2_decap_4 FILLER_8_2546 ();
 sg13g2_fill_1 FILLER_8_2550 ();
 sg13g2_decap_4 FILLER_8_2559 ();
 sg13g2_decap_4 FILLER_8_2567 ();
 sg13g2_fill_2 FILLER_8_2571 ();
 sg13g2_decap_8 FILLER_8_2599 ();
 sg13g2_decap_8 FILLER_8_2606 ();
 sg13g2_decap_8 FILLER_8_2613 ();
 sg13g2_decap_8 FILLER_8_2620 ();
 sg13g2_decap_8 FILLER_8_2627 ();
 sg13g2_decap_8 FILLER_8_2634 ();
 sg13g2_decap_8 FILLER_8_2641 ();
 sg13g2_decap_8 FILLER_8_2648 ();
 sg13g2_decap_8 FILLER_8_2655 ();
 sg13g2_decap_8 FILLER_8_2662 ();
 sg13g2_fill_1 FILLER_8_2669 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_1 FILLER_9_28 ();
 sg13g2_fill_2 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_47 ();
 sg13g2_fill_2 FILLER_9_55 ();
 sg13g2_decap_8 FILLER_9_83 ();
 sg13g2_decap_8 FILLER_9_90 ();
 sg13g2_fill_1 FILLER_9_97 ();
 sg13g2_fill_2 FILLER_9_108 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_fill_1 FILLER_9_125 ();
 sg13g2_fill_2 FILLER_9_131 ();
 sg13g2_decap_4 FILLER_9_137 ();
 sg13g2_fill_1 FILLER_9_141 ();
 sg13g2_fill_1 FILLER_9_151 ();
 sg13g2_fill_2 FILLER_9_156 ();
 sg13g2_fill_2 FILLER_9_163 ();
 sg13g2_fill_2 FILLER_9_170 ();
 sg13g2_fill_1 FILLER_9_183 ();
 sg13g2_fill_2 FILLER_9_190 ();
 sg13g2_fill_1 FILLER_9_209 ();
 sg13g2_fill_2 FILLER_9_214 ();
 sg13g2_decap_4 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_234 ();
 sg13g2_fill_2 FILLER_9_258 ();
 sg13g2_fill_1 FILLER_9_260 ();
 sg13g2_fill_2 FILLER_9_268 ();
 sg13g2_fill_1 FILLER_9_270 ();
 sg13g2_fill_2 FILLER_9_281 ();
 sg13g2_fill_1 FILLER_9_283 ();
 sg13g2_fill_1 FILLER_9_290 ();
 sg13g2_fill_2 FILLER_9_299 ();
 sg13g2_fill_2 FILLER_9_318 ();
 sg13g2_decap_4 FILLER_9_325 ();
 sg13g2_fill_1 FILLER_9_329 ();
 sg13g2_decap_4 FILLER_9_334 ();
 sg13g2_decap_4 FILLER_9_365 ();
 sg13g2_fill_2 FILLER_9_369 ();
 sg13g2_fill_2 FILLER_9_381 ();
 sg13g2_fill_1 FILLER_9_383 ();
 sg13g2_fill_1 FILLER_9_394 ();
 sg13g2_fill_2 FILLER_9_403 ();
 sg13g2_fill_1 FILLER_9_405 ();
 sg13g2_decap_4 FILLER_9_419 ();
 sg13g2_decap_8 FILLER_9_432 ();
 sg13g2_decap_8 FILLER_9_439 ();
 sg13g2_decap_8 FILLER_9_446 ();
 sg13g2_fill_2 FILLER_9_458 ();
 sg13g2_decap_8 FILLER_9_523 ();
 sg13g2_decap_8 FILLER_9_530 ();
 sg13g2_decap_8 FILLER_9_537 ();
 sg13g2_fill_2 FILLER_9_544 ();
 sg13g2_fill_1 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_552 ();
 sg13g2_decap_8 FILLER_9_559 ();
 sg13g2_decap_4 FILLER_9_566 ();
 sg13g2_fill_1 FILLER_9_570 ();
 sg13g2_fill_2 FILLER_9_580 ();
 sg13g2_fill_1 FILLER_9_582 ();
 sg13g2_fill_1 FILLER_9_588 ();
 sg13g2_fill_1 FILLER_9_594 ();
 sg13g2_fill_2 FILLER_9_610 ();
 sg13g2_fill_2 FILLER_9_621 ();
 sg13g2_fill_2 FILLER_9_627 ();
 sg13g2_decap_8 FILLER_9_641 ();
 sg13g2_decap_4 FILLER_9_648 ();
 sg13g2_fill_2 FILLER_9_656 ();
 sg13g2_fill_2 FILLER_9_662 ();
 sg13g2_fill_1 FILLER_9_664 ();
 sg13g2_fill_1 FILLER_9_673 ();
 sg13g2_fill_2 FILLER_9_678 ();
 sg13g2_fill_1 FILLER_9_683 ();
 sg13g2_fill_1 FILLER_9_729 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_4 FILLER_9_812 ();
 sg13g2_fill_2 FILLER_9_828 ();
 sg13g2_fill_1 FILLER_9_830 ();
 sg13g2_decap_4 FILLER_9_843 ();
 sg13g2_fill_2 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_859 ();
 sg13g2_fill_2 FILLER_9_866 ();
 sg13g2_fill_2 FILLER_9_910 ();
 sg13g2_fill_2 FILLER_9_998 ();
 sg13g2_fill_2 FILLER_9_1027 ();
 sg13g2_fill_1 FILLER_9_1029 ();
 sg13g2_decap_8 FILLER_9_1047 ();
 sg13g2_fill_2 FILLER_9_1054 ();
 sg13g2_decap_4 FILLER_9_1072 ();
 sg13g2_fill_2 FILLER_9_1076 ();
 sg13g2_decap_8 FILLER_9_1083 ();
 sg13g2_fill_1 FILLER_9_1090 ();
 sg13g2_fill_2 FILLER_9_1101 ();
 sg13g2_fill_2 FILLER_9_1109 ();
 sg13g2_fill_1 FILLER_9_1111 ();
 sg13g2_decap_4 FILLER_9_1138 ();
 sg13g2_fill_2 FILLER_9_1142 ();
 sg13g2_fill_1 FILLER_9_1173 ();
 sg13g2_fill_2 FILLER_9_1187 ();
 sg13g2_decap_8 FILLER_9_1228 ();
 sg13g2_decap_8 FILLER_9_1235 ();
 sg13g2_decap_4 FILLER_9_1242 ();
 sg13g2_fill_1 FILLER_9_1246 ();
 sg13g2_fill_1 FILLER_9_1262 ();
 sg13g2_decap_8 FILLER_9_1299 ();
 sg13g2_decap_8 FILLER_9_1328 ();
 sg13g2_decap_4 FILLER_9_1335 ();
 sg13g2_decap_8 FILLER_9_1349 ();
 sg13g2_decap_8 FILLER_9_1356 ();
 sg13g2_fill_1 FILLER_9_1443 ();
 sg13g2_fill_1 FILLER_9_1472 ();
 sg13g2_decap_8 FILLER_9_1499 ();
 sg13g2_decap_8 FILLER_9_1506 ();
 sg13g2_decap_4 FILLER_9_1519 ();
 sg13g2_fill_1 FILLER_9_1526 ();
 sg13g2_fill_1 FILLER_9_1543 ();
 sg13g2_fill_1 FILLER_9_1589 ();
 sg13g2_fill_1 FILLER_9_1652 ();
 sg13g2_fill_1 FILLER_9_1671 ();
 sg13g2_fill_1 FILLER_9_1692 ();
 sg13g2_fill_1 FILLER_9_1719 ();
 sg13g2_decap_8 FILLER_9_1752 ();
 sg13g2_fill_1 FILLER_9_1759 ();
 sg13g2_fill_1 FILLER_9_1786 ();
 sg13g2_fill_2 FILLER_9_1794 ();
 sg13g2_decap_8 FILLER_9_1817 ();
 sg13g2_decap_8 FILLER_9_1824 ();
 sg13g2_fill_2 FILLER_9_1831 ();
 sg13g2_fill_1 FILLER_9_1847 ();
 sg13g2_fill_1 FILLER_9_1884 ();
 sg13g2_fill_2 FILLER_9_1895 ();
 sg13g2_fill_2 FILLER_9_1930 ();
 sg13g2_fill_2 FILLER_9_1985 ();
 sg13g2_fill_2 FILLER_9_2000 ();
 sg13g2_fill_1 FILLER_9_2015 ();
 sg13g2_fill_2 FILLER_9_2022 ();
 sg13g2_fill_1 FILLER_9_2033 ();
 sg13g2_fill_2 FILLER_9_2040 ();
 sg13g2_fill_1 FILLER_9_2051 ();
 sg13g2_fill_2 FILLER_9_2085 ();
 sg13g2_fill_2 FILLER_9_2109 ();
 sg13g2_fill_2 FILLER_9_2173 ();
 sg13g2_fill_1 FILLER_9_2201 ();
 sg13g2_fill_1 FILLER_9_2213 ();
 sg13g2_fill_1 FILLER_9_2226 ();
 sg13g2_fill_1 FILLER_9_2252 ();
 sg13g2_fill_2 FILLER_9_2292 ();
 sg13g2_fill_2 FILLER_9_2300 ();
 sg13g2_fill_1 FILLER_9_2311 ();
 sg13g2_decap_4 FILLER_9_2328 ();
 sg13g2_fill_1 FILLER_9_2332 ();
 sg13g2_fill_2 FILLER_9_2363 ();
 sg13g2_decap_8 FILLER_9_2385 ();
 sg13g2_decap_8 FILLER_9_2392 ();
 sg13g2_decap_8 FILLER_9_2399 ();
 sg13g2_fill_1 FILLER_9_2422 ();
 sg13g2_fill_2 FILLER_9_2427 ();
 sg13g2_fill_2 FILLER_9_2433 ();
 sg13g2_decap_8 FILLER_9_2494 ();
 sg13g2_fill_2 FILLER_9_2501 ();
 sg13g2_fill_1 FILLER_9_2503 ();
 sg13g2_fill_1 FILLER_9_2512 ();
 sg13g2_fill_1 FILLER_9_2539 ();
 sg13g2_fill_2 FILLER_9_2544 ();
 sg13g2_fill_1 FILLER_9_2554 ();
 sg13g2_decap_8 FILLER_9_2604 ();
 sg13g2_decap_8 FILLER_9_2611 ();
 sg13g2_decap_8 FILLER_9_2618 ();
 sg13g2_decap_8 FILLER_9_2625 ();
 sg13g2_decap_8 FILLER_9_2632 ();
 sg13g2_decap_8 FILLER_9_2639 ();
 sg13g2_decap_8 FILLER_9_2646 ();
 sg13g2_decap_8 FILLER_9_2653 ();
 sg13g2_decap_8 FILLER_9_2660 ();
 sg13g2_fill_2 FILLER_9_2667 ();
 sg13g2_fill_1 FILLER_9_2669 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_fill_1 FILLER_10_21 ();
 sg13g2_fill_1 FILLER_10_30 ();
 sg13g2_fill_1 FILLER_10_36 ();
 sg13g2_decap_4 FILLER_10_52 ();
 sg13g2_decap_4 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_73 ();
 sg13g2_fill_2 FILLER_10_80 ();
 sg13g2_decap_8 FILLER_10_86 ();
 sg13g2_decap_8 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_100 ();
 sg13g2_fill_1 FILLER_10_106 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_126 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_2 FILLER_10_189 ();
 sg13g2_fill_2 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_233 ();
 sg13g2_fill_1 FILLER_10_266 ();
 sg13g2_fill_1 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_2 FILLER_10_288 ();
 sg13g2_fill_1 FILLER_10_290 ();
 sg13g2_fill_2 FILLER_10_302 ();
 sg13g2_fill_2 FILLER_10_309 ();
 sg13g2_fill_2 FILLER_10_316 ();
 sg13g2_fill_1 FILLER_10_323 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_fill_2 FILLER_10_356 ();
 sg13g2_fill_2 FILLER_10_364 ();
 sg13g2_decap_4 FILLER_10_382 ();
 sg13g2_decap_4 FILLER_10_401 ();
 sg13g2_decap_8 FILLER_10_416 ();
 sg13g2_decap_8 FILLER_10_423 ();
 sg13g2_decap_8 FILLER_10_430 ();
 sg13g2_decap_4 FILLER_10_437 ();
 sg13g2_fill_2 FILLER_10_446 ();
 sg13g2_fill_1 FILLER_10_511 ();
 sg13g2_fill_2 FILLER_10_516 ();
 sg13g2_fill_2 FILLER_10_528 ();
 sg13g2_fill_1 FILLER_10_530 ();
 sg13g2_fill_2 FILLER_10_536 ();
 sg13g2_fill_1 FILLER_10_538 ();
 sg13g2_fill_1 FILLER_10_565 ();
 sg13g2_fill_1 FILLER_10_593 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_fill_2 FILLER_10_606 ();
 sg13g2_fill_2 FILLER_10_618 ();
 sg13g2_fill_2 FILLER_10_646 ();
 sg13g2_fill_2 FILLER_10_674 ();
 sg13g2_fill_1 FILLER_10_680 ();
 sg13g2_fill_1 FILLER_10_693 ();
 sg13g2_fill_2 FILLER_10_698 ();
 sg13g2_fill_2 FILLER_10_706 ();
 sg13g2_fill_2 FILLER_10_728 ();
 sg13g2_decap_4 FILLER_10_744 ();
 sg13g2_fill_1 FILLER_10_748 ();
 sg13g2_fill_2 FILLER_10_755 ();
 sg13g2_decap_4 FILLER_10_772 ();
 sg13g2_fill_2 FILLER_10_776 ();
 sg13g2_decap_8 FILLER_10_814 ();
 sg13g2_decap_8 FILLER_10_821 ();
 sg13g2_decap_4 FILLER_10_828 ();
 sg13g2_fill_1 FILLER_10_841 ();
 sg13g2_fill_1 FILLER_10_878 ();
 sg13g2_fill_2 FILLER_10_927 ();
 sg13g2_fill_2 FILLER_10_960 ();
 sg13g2_fill_1 FILLER_10_996 ();
 sg13g2_fill_1 FILLER_10_1032 ();
 sg13g2_decap_8 FILLER_10_1097 ();
 sg13g2_decap_8 FILLER_10_1112 ();
 sg13g2_fill_2 FILLER_10_1119 ();
 sg13g2_fill_1 FILLER_10_1126 ();
 sg13g2_fill_2 FILLER_10_1133 ();
 sg13g2_fill_1 FILLER_10_1140 ();
 sg13g2_fill_1 FILLER_10_1185 ();
 sg13g2_fill_1 FILLER_10_1198 ();
 sg13g2_decap_8 FILLER_10_1225 ();
 sg13g2_decap_8 FILLER_10_1232 ();
 sg13g2_decap_8 FILLER_10_1239 ();
 sg13g2_fill_2 FILLER_10_1246 ();
 sg13g2_decap_8 FILLER_10_1284 ();
 sg13g2_fill_1 FILLER_10_1291 ();
 sg13g2_decap_8 FILLER_10_1304 ();
 sg13g2_decap_8 FILLER_10_1311 ();
 sg13g2_decap_8 FILLER_10_1318 ();
 sg13g2_decap_8 FILLER_10_1325 ();
 sg13g2_decap_8 FILLER_10_1332 ();
 sg13g2_decap_8 FILLER_10_1339 ();
 sg13g2_decap_8 FILLER_10_1352 ();
 sg13g2_decap_4 FILLER_10_1359 ();
 sg13g2_fill_2 FILLER_10_1363 ();
 sg13g2_decap_8 FILLER_10_1369 ();
 sg13g2_decap_8 FILLER_10_1376 ();
 sg13g2_decap_8 FILLER_10_1383 ();
 sg13g2_decap_4 FILLER_10_1490 ();
 sg13g2_fill_1 FILLER_10_1494 ();
 sg13g2_fill_2 FILLER_10_1516 ();
 sg13g2_fill_1 FILLER_10_1526 ();
 sg13g2_fill_2 FILLER_10_1562 ();
 sg13g2_decap_8 FILLER_10_1631 ();
 sg13g2_decap_4 FILLER_10_1638 ();
 sg13g2_fill_1 FILLER_10_1642 ();
 sg13g2_decap_8 FILLER_10_1772 ();
 sg13g2_decap_8 FILLER_10_1779 ();
 sg13g2_fill_1 FILLER_10_1786 ();
 sg13g2_fill_2 FILLER_10_1796 ();
 sg13g2_decap_8 FILLER_10_1865 ();
 sg13g2_fill_1 FILLER_10_1891 ();
 sg13g2_fill_2 FILLER_10_1895 ();
 sg13g2_fill_2 FILLER_10_1942 ();
 sg13g2_fill_2 FILLER_10_1947 ();
 sg13g2_fill_1 FILLER_10_1978 ();
 sg13g2_decap_8 FILLER_10_1992 ();
 sg13g2_decap_4 FILLER_10_1999 ();
 sg13g2_fill_1 FILLER_10_2003 ();
 sg13g2_fill_1 FILLER_10_2024 ();
 sg13g2_fill_1 FILLER_10_2038 ();
 sg13g2_fill_2 FILLER_10_2058 ();
 sg13g2_fill_2 FILLER_10_2093 ();
 sg13g2_fill_1 FILLER_10_2134 ();
 sg13g2_fill_1 FILLER_10_2166 ();
 sg13g2_fill_1 FILLER_10_2176 ();
 sg13g2_fill_1 FILLER_10_2186 ();
 sg13g2_fill_1 FILLER_10_2229 ();
 sg13g2_fill_1 FILLER_10_2236 ();
 sg13g2_fill_1 FILLER_10_2272 ();
 sg13g2_fill_1 FILLER_10_2285 ();
 sg13g2_decap_8 FILLER_10_2289 ();
 sg13g2_fill_2 FILLER_10_2296 ();
 sg13g2_decap_8 FILLER_10_2332 ();
 sg13g2_fill_1 FILLER_10_2339 ();
 sg13g2_fill_2 FILLER_10_2344 ();
 sg13g2_fill_2 FILLER_10_2354 ();
 sg13g2_fill_1 FILLER_10_2390 ();
 sg13g2_fill_2 FILLER_10_2417 ();
 sg13g2_decap_4 FILLER_10_2445 ();
 sg13g2_decap_4 FILLER_10_2471 ();
 sg13g2_decap_4 FILLER_10_2479 ();
 sg13g2_fill_1 FILLER_10_2483 ();
 sg13g2_fill_2 FILLER_10_2492 ();
 sg13g2_fill_1 FILLER_10_2494 ();
 sg13g2_decap_4 FILLER_10_2500 ();
 sg13g2_fill_2 FILLER_10_2504 ();
 sg13g2_fill_1 FILLER_10_2511 ();
 sg13g2_fill_1 FILLER_10_2523 ();
 sg13g2_decap_8 FILLER_10_2532 ();
 sg13g2_fill_2 FILLER_10_2539 ();
 sg13g2_fill_1 FILLER_10_2552 ();
 sg13g2_fill_2 FILLER_10_2609 ();
 sg13g2_decap_8 FILLER_10_2637 ();
 sg13g2_decap_8 FILLER_10_2644 ();
 sg13g2_decap_8 FILLER_10_2651 ();
 sg13g2_decap_8 FILLER_10_2658 ();
 sg13g2_decap_4 FILLER_10_2665 ();
 sg13g2_fill_1 FILLER_10_2669 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_17 ();
 sg13g2_fill_1 FILLER_11_35 ();
 sg13g2_decap_4 FILLER_11_54 ();
 sg13g2_decap_4 FILLER_11_104 ();
 sg13g2_fill_2 FILLER_11_108 ();
 sg13g2_fill_2 FILLER_11_120 ();
 sg13g2_fill_1 FILLER_11_143 ();
 sg13g2_fill_1 FILLER_11_150 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_2 FILLER_11_182 ();
 sg13g2_fill_1 FILLER_11_184 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_198 ();
 sg13g2_fill_1 FILLER_11_214 ();
 sg13g2_decap_4 FILLER_11_220 ();
 sg13g2_fill_1 FILLER_11_229 ();
 sg13g2_fill_1 FILLER_11_246 ();
 sg13g2_fill_1 FILLER_11_252 ();
 sg13g2_fill_2 FILLER_11_268 ();
 sg13g2_fill_1 FILLER_11_277 ();
 sg13g2_fill_1 FILLER_11_283 ();
 sg13g2_fill_1 FILLER_11_289 ();
 sg13g2_decap_8 FILLER_11_311 ();
 sg13g2_fill_2 FILLER_11_323 ();
 sg13g2_decap_8 FILLER_11_330 ();
 sg13g2_fill_2 FILLER_11_337 ();
 sg13g2_decap_4 FILLER_11_343 ();
 sg13g2_fill_2 FILLER_11_347 ();
 sg13g2_fill_2 FILLER_11_395 ();
 sg13g2_fill_1 FILLER_11_402 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_decap_8 FILLER_11_435 ();
 sg13g2_decap_8 FILLER_11_442 ();
 sg13g2_decap_8 FILLER_11_449 ();
 sg13g2_fill_2 FILLER_11_456 ();
 sg13g2_fill_1 FILLER_11_458 ();
 sg13g2_fill_1 FILLER_11_477 ();
 sg13g2_fill_2 FILLER_11_481 ();
 sg13g2_fill_1 FILLER_11_492 ();
 sg13g2_fill_1 FILLER_11_505 ();
 sg13g2_fill_2 FILLER_11_518 ();
 sg13g2_fill_1 FILLER_11_520 ();
 sg13g2_decap_8 FILLER_11_526 ();
 sg13g2_decap_4 FILLER_11_533 ();
 sg13g2_fill_2 FILLER_11_537 ();
 sg13g2_fill_1 FILLER_11_565 ();
 sg13g2_fill_1 FILLER_11_570 ();
 sg13g2_fill_2 FILLER_11_575 ();
 sg13g2_decap_8 FILLER_11_601 ();
 sg13g2_decap_8 FILLER_11_622 ();
 sg13g2_decap_8 FILLER_11_629 ();
 sg13g2_decap_4 FILLER_11_636 ();
 sg13g2_fill_2 FILLER_11_640 ();
 sg13g2_fill_1 FILLER_11_652 ();
 sg13g2_fill_1 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_705 ();
 sg13g2_fill_2 FILLER_11_712 ();
 sg13g2_fill_1 FILLER_11_724 ();
 sg13g2_fill_1 FILLER_11_735 ();
 sg13g2_fill_1 FILLER_11_768 ();
 sg13g2_decap_8 FILLER_11_775 ();
 sg13g2_decap_8 FILLER_11_782 ();
 sg13g2_decap_4 FILLER_11_789 ();
 sg13g2_fill_1 FILLER_11_793 ();
 sg13g2_decap_4 FILLER_11_828 ();
 sg13g2_decap_8 FILLER_11_842 ();
 sg13g2_decap_4 FILLER_11_849 ();
 sg13g2_fill_2 FILLER_11_869 ();
 sg13g2_fill_1 FILLER_11_880 ();
 sg13g2_fill_1 FILLER_11_897 ();
 sg13g2_fill_2 FILLER_11_904 ();
 sg13g2_fill_2 FILLER_11_955 ();
 sg13g2_fill_2 FILLER_11_974 ();
 sg13g2_fill_2 FILLER_11_985 ();
 sg13g2_fill_2 FILLER_11_1032 ();
 sg13g2_fill_2 FILLER_11_1063 ();
 sg13g2_fill_1 FILLER_11_1080 ();
 sg13g2_fill_2 FILLER_11_1110 ();
 sg13g2_fill_1 FILLER_11_1153 ();
 sg13g2_fill_2 FILLER_11_1164 ();
 sg13g2_fill_2 FILLER_11_1172 ();
 sg13g2_fill_1 FILLER_11_1194 ();
 sg13g2_decap_8 FILLER_11_1224 ();
 sg13g2_decap_8 FILLER_11_1231 ();
 sg13g2_fill_1 FILLER_11_1238 ();
 sg13g2_fill_1 FILLER_11_1251 ();
 sg13g2_decap_8 FILLER_11_1260 ();
 sg13g2_fill_2 FILLER_11_1267 ();
 sg13g2_decap_8 FILLER_11_1277 ();
 sg13g2_fill_2 FILLER_11_1290 ();
 sg13g2_decap_4 FILLER_11_1336 ();
 sg13g2_fill_2 FILLER_11_1399 ();
 sg13g2_decap_8 FILLER_11_1427 ();
 sg13g2_fill_1 FILLER_11_1434 ();
 sg13g2_fill_1 FILLER_11_1459 ();
 sg13g2_fill_2 FILLER_11_1470 ();
 sg13g2_decap_4 FILLER_11_1544 ();
 sg13g2_fill_1 FILLER_11_1548 ();
 sg13g2_fill_1 FILLER_11_1561 ();
 sg13g2_decap_8 FILLER_11_1570 ();
 sg13g2_decap_8 FILLER_11_1577 ();
 sg13g2_decap_8 FILLER_11_1635 ();
 sg13g2_fill_1 FILLER_11_1642 ();
 sg13g2_fill_1 FILLER_11_1655 ();
 sg13g2_fill_1 FILLER_11_1682 ();
 sg13g2_fill_1 FILLER_11_1698 ();
 sg13g2_fill_1 FILLER_11_1725 ();
 sg13g2_fill_1 FILLER_11_1758 ();
 sg13g2_fill_2 FILLER_11_1764 ();
 sg13g2_fill_1 FILLER_11_1771 ();
 sg13g2_fill_1 FILLER_11_1798 ();
 sg13g2_fill_1 FILLER_11_1805 ();
 sg13g2_fill_2 FILLER_11_1825 ();
 sg13g2_fill_2 FILLER_11_1834 ();
 sg13g2_fill_2 FILLER_11_1860 ();
 sg13g2_fill_1 FILLER_11_1862 ();
 sg13g2_fill_2 FILLER_11_1924 ();
 sg13g2_fill_2 FILLER_11_1977 ();
 sg13g2_fill_1 FILLER_11_1979 ();
 sg13g2_fill_2 FILLER_11_2020 ();
 sg13g2_fill_2 FILLER_11_2030 ();
 sg13g2_fill_2 FILLER_11_2124 ();
 sg13g2_fill_1 FILLER_11_2156 ();
 sg13g2_fill_1 FILLER_11_2192 ();
 sg13g2_fill_1 FILLER_11_2207 ();
 sg13g2_fill_1 FILLER_11_2213 ();
 sg13g2_fill_1 FILLER_11_2233 ();
 sg13g2_fill_1 FILLER_11_2274 ();
 sg13g2_decap_8 FILLER_11_2297 ();
 sg13g2_decap_8 FILLER_11_2304 ();
 sg13g2_fill_2 FILLER_11_2311 ();
 sg13g2_decap_8 FILLER_11_2317 ();
 sg13g2_decap_8 FILLER_11_2324 ();
 sg13g2_decap_8 FILLER_11_2331 ();
 sg13g2_fill_2 FILLER_11_2338 ();
 sg13g2_decap_4 FILLER_11_2370 ();
 sg13g2_fill_2 FILLER_11_2378 ();
 sg13g2_fill_1 FILLER_11_2380 ();
 sg13g2_decap_4 FILLER_11_2415 ();
 sg13g2_fill_1 FILLER_11_2419 ();
 sg13g2_fill_1 FILLER_11_2435 ();
 sg13g2_decap_4 FILLER_11_2466 ();
 sg13g2_fill_1 FILLER_11_2470 ();
 sg13g2_fill_2 FILLER_11_2510 ();
 sg13g2_fill_2 FILLER_11_2533 ();
 sg13g2_fill_1 FILLER_11_2539 ();
 sg13g2_fill_2 FILLER_11_2570 ();
 sg13g2_decap_4 FILLER_11_2598 ();
 sg13g2_fill_1 FILLER_11_2602 ();
 sg13g2_decap_8 FILLER_11_2641 ();
 sg13g2_decap_8 FILLER_11_2648 ();
 sg13g2_decap_8 FILLER_11_2655 ();
 sg13g2_decap_8 FILLER_11_2662 ();
 sg13g2_fill_1 FILLER_11_2669 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_4 FILLER_12_7 ();
 sg13g2_fill_1 FILLER_12_11 ();
 sg13g2_fill_2 FILLER_12_54 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_4 FILLER_12_88 ();
 sg13g2_fill_1 FILLER_12_92 ();
 sg13g2_decap_4 FILLER_12_97 ();
 sg13g2_fill_2 FILLER_12_101 ();
 sg13g2_fill_1 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_150 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_165 ();
 sg13g2_fill_1 FILLER_12_197 ();
 sg13g2_fill_2 FILLER_12_202 ();
 sg13g2_fill_1 FILLER_12_209 ();
 sg13g2_fill_2 FILLER_12_221 ();
 sg13g2_fill_2 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_240 ();
 sg13g2_decap_8 FILLER_12_247 ();
 sg13g2_decap_4 FILLER_12_269 ();
 sg13g2_fill_1 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_316 ();
 sg13g2_decap_4 FILLER_12_323 ();
 sg13g2_fill_1 FILLER_12_361 ();
 sg13g2_decap_4 FILLER_12_371 ();
 sg13g2_fill_1 FILLER_12_385 ();
 sg13g2_fill_2 FILLER_12_390 ();
 sg13g2_fill_2 FILLER_12_397 ();
 sg13g2_fill_2 FILLER_12_404 ();
 sg13g2_decap_4 FILLER_12_419 ();
 sg13g2_fill_1 FILLER_12_456 ();
 sg13g2_fill_1 FILLER_12_483 ();
 sg13g2_fill_2 FILLER_12_496 ();
 sg13g2_fill_1 FILLER_12_503 ();
 sg13g2_fill_1 FILLER_12_517 ();
 sg13g2_decap_4 FILLER_12_522 ();
 sg13g2_decap_4 FILLER_12_535 ();
 sg13g2_fill_1 FILLER_12_539 ();
 sg13g2_fill_2 FILLER_12_547 ();
 sg13g2_fill_1 FILLER_12_549 ();
 sg13g2_fill_2 FILLER_12_558 ();
 sg13g2_fill_1 FILLER_12_560 ();
 sg13g2_decap_8 FILLER_12_567 ();
 sg13g2_fill_2 FILLER_12_574 ();
 sg13g2_fill_1 FILLER_12_576 ();
 sg13g2_fill_1 FILLER_12_590 ();
 sg13g2_fill_2 FILLER_12_637 ();
 sg13g2_fill_2 FILLER_12_648 ();
 sg13g2_decap_4 FILLER_12_655 ();
 sg13g2_fill_2 FILLER_12_659 ();
 sg13g2_fill_2 FILLER_12_671 ();
 sg13g2_fill_1 FILLER_12_673 ();
 sg13g2_decap_4 FILLER_12_787 ();
 sg13g2_decap_8 FILLER_12_794 ();
 sg13g2_fill_1 FILLER_12_801 ();
 sg13g2_fill_2 FILLER_12_828 ();
 sg13g2_fill_2 FILLER_12_840 ();
 sg13g2_fill_1 FILLER_12_929 ();
 sg13g2_fill_1 FILLER_12_956 ();
 sg13g2_fill_1 FILLER_12_965 ();
 sg13g2_fill_2 FILLER_12_1030 ();
 sg13g2_fill_2 FILLER_12_1057 ();
 sg13g2_fill_1 FILLER_12_1071 ();
 sg13g2_fill_2 FILLER_12_1079 ();
 sg13g2_fill_2 FILLER_12_1091 ();
 sg13g2_decap_8 FILLER_12_1119 ();
 sg13g2_decap_4 FILLER_12_1126 ();
 sg13g2_fill_1 FILLER_12_1130 ();
 sg13g2_decap_4 FILLER_12_1135 ();
 sg13g2_fill_2 FILLER_12_1139 ();
 sg13g2_decap_8 FILLER_12_1146 ();
 sg13g2_fill_2 FILLER_12_1153 ();
 sg13g2_fill_1 FILLER_12_1155 ();
 sg13g2_decap_8 FILLER_12_1182 ();
 sg13g2_decap_4 FILLER_12_1195 ();
 sg13g2_fill_2 FILLER_12_1199 ();
 sg13g2_decap_4 FILLER_12_1228 ();
 sg13g2_fill_2 FILLER_12_1232 ();
 sg13g2_fill_2 FILLER_12_1238 ();
 sg13g2_fill_1 FILLER_12_1240 ();
 sg13g2_decap_8 FILLER_12_1271 ();
 sg13g2_fill_2 FILLER_12_1304 ();
 sg13g2_fill_1 FILLER_12_1311 ();
 sg13g2_fill_2 FILLER_12_1357 ();
 sg13g2_fill_1 FILLER_12_1359 ();
 sg13g2_decap_4 FILLER_12_1363 ();
 sg13g2_fill_1 FILLER_12_1367 ();
 sg13g2_fill_1 FILLER_12_1371 ();
 sg13g2_fill_2 FILLER_12_1396 ();
 sg13g2_fill_1 FILLER_12_1413 ();
 sg13g2_fill_1 FILLER_12_1440 ();
 sg13g2_decap_4 FILLER_12_1517 ();
 sg13g2_fill_2 FILLER_12_1521 ();
 sg13g2_decap_8 FILLER_12_1526 ();
 sg13g2_decap_8 FILLER_12_1533 ();
 sg13g2_decap_4 FILLER_12_1540 ();
 sg13g2_fill_2 FILLER_12_1544 ();
 sg13g2_decap_8 FILLER_12_1585 ();
 sg13g2_fill_1 FILLER_12_1592 ();
 sg13g2_decap_8 FILLER_12_1611 ();
 sg13g2_fill_2 FILLER_12_1623 ();
 sg13g2_fill_1 FILLER_12_1661 ();
 sg13g2_fill_2 FILLER_12_1706 ();
 sg13g2_fill_2 FILLER_12_1730 ();
 sg13g2_fill_1 FILLER_12_1741 ();
 sg13g2_fill_2 FILLER_12_1759 ();
 sg13g2_fill_2 FILLER_12_1765 ();
 sg13g2_decap_8 FILLER_12_1774 ();
 sg13g2_decap_4 FILLER_12_1781 ();
 sg13g2_fill_2 FILLER_12_1785 ();
 sg13g2_decap_4 FILLER_12_1803 ();
 sg13g2_fill_2 FILLER_12_1807 ();
 sg13g2_fill_2 FILLER_12_1839 ();
 sg13g2_fill_1 FILLER_12_1850 ();
 sg13g2_fill_1 FILLER_12_1889 ();
 sg13g2_fill_1 FILLER_12_1898 ();
 sg13g2_fill_2 FILLER_12_1916 ();
 sg13g2_fill_1 FILLER_12_1947 ();
 sg13g2_fill_1 FILLER_12_1962 ();
 sg13g2_decap_4 FILLER_12_1977 ();
 sg13g2_decap_8 FILLER_12_1989 ();
 sg13g2_fill_1 FILLER_12_2019 ();
 sg13g2_fill_2 FILLER_12_2165 ();
 sg13g2_fill_2 FILLER_12_2197 ();
 sg13g2_fill_2 FILLER_12_2246 ();
 sg13g2_fill_1 FILLER_12_2285 ();
 sg13g2_decap_4 FILLER_12_2298 ();
 sg13g2_decap_8 FILLER_12_2332 ();
 sg13g2_decap_8 FILLER_12_2339 ();
 sg13g2_decap_8 FILLER_12_2346 ();
 sg13g2_decap_8 FILLER_12_2353 ();
 sg13g2_decap_8 FILLER_12_2360 ();
 sg13g2_decap_8 FILLER_12_2367 ();
 sg13g2_decap_8 FILLER_12_2374 ();
 sg13g2_decap_4 FILLER_12_2386 ();
 sg13g2_decap_8 FILLER_12_2404 ();
 sg13g2_decap_4 FILLER_12_2417 ();
 sg13g2_fill_1 FILLER_12_2425 ();
 sg13g2_fill_1 FILLER_12_2486 ();
 sg13g2_fill_1 FILLER_12_2491 ();
 sg13g2_decap_8 FILLER_12_2522 ();
 sg13g2_decap_8 FILLER_12_2529 ();
 sg13g2_decap_4 FILLER_12_2536 ();
 sg13g2_fill_2 FILLER_12_2548 ();
 sg13g2_decap_8 FILLER_12_2555 ();
 sg13g2_decap_4 FILLER_12_2562 ();
 sg13g2_fill_2 FILLER_12_2566 ();
 sg13g2_decap_8 FILLER_12_2572 ();
 sg13g2_decap_4 FILLER_12_2583 ();
 sg13g2_decap_8 FILLER_12_2590 ();
 sg13g2_fill_1 FILLER_12_2597 ();
 sg13g2_fill_2 FILLER_12_2625 ();
 sg13g2_fill_1 FILLER_12_2627 ();
 sg13g2_decap_8 FILLER_12_2654 ();
 sg13g2_decap_8 FILLER_12_2661 ();
 sg13g2_fill_2 FILLER_12_2668 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_4 FILLER_13_7 ();
 sg13g2_decap_4 FILLER_13_45 ();
 sg13g2_fill_1 FILLER_13_49 ();
 sg13g2_decap_4 FILLER_13_55 ();
 sg13g2_fill_1 FILLER_13_59 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_decap_8 FILLER_13_73 ();
 sg13g2_decap_8 FILLER_13_80 ();
 sg13g2_decap_8 FILLER_13_87 ();
 sg13g2_fill_2 FILLER_13_94 ();
 sg13g2_fill_1 FILLER_13_96 ();
 sg13g2_fill_1 FILLER_13_120 ();
 sg13g2_fill_1 FILLER_13_125 ();
 sg13g2_fill_2 FILLER_13_141 ();
 sg13g2_fill_1 FILLER_13_143 ();
 sg13g2_fill_1 FILLER_13_149 ();
 sg13g2_fill_1 FILLER_13_177 ();
 sg13g2_fill_1 FILLER_13_188 ();
 sg13g2_fill_2 FILLER_13_194 ();
 sg13g2_fill_1 FILLER_13_201 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_decap_4 FILLER_13_236 ();
 sg13g2_fill_2 FILLER_13_240 ();
 sg13g2_decap_8 FILLER_13_247 ();
 sg13g2_fill_1 FILLER_13_254 ();
 sg13g2_decap_4 FILLER_13_259 ();
 sg13g2_fill_1 FILLER_13_263 ();
 sg13g2_fill_2 FILLER_13_274 ();
 sg13g2_decap_8 FILLER_13_291 ();
 sg13g2_decap_4 FILLER_13_298 ();
 sg13g2_fill_2 FILLER_13_312 ();
 sg13g2_fill_2 FILLER_13_320 ();
 sg13g2_fill_1 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_332 ();
 sg13g2_decap_8 FILLER_13_339 ();
 sg13g2_decap_8 FILLER_13_346 ();
 sg13g2_fill_2 FILLER_13_353 ();
 sg13g2_fill_1 FILLER_13_355 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_fill_2 FILLER_13_411 ();
 sg13g2_decap_8 FILLER_13_417 ();
 sg13g2_fill_1 FILLER_13_424 ();
 sg13g2_decap_8 FILLER_13_433 ();
 sg13g2_decap_8 FILLER_13_440 ();
 sg13g2_decap_4 FILLER_13_447 ();
 sg13g2_fill_1 FILLER_13_455 ();
 sg13g2_decap_4 FILLER_13_469 ();
 sg13g2_fill_1 FILLER_13_481 ();
 sg13g2_fill_1 FILLER_13_500 ();
 sg13g2_fill_2 FILLER_13_506 ();
 sg13g2_decap_8 FILLER_13_512 ();
 sg13g2_decap_8 FILLER_13_519 ();
 sg13g2_decap_8 FILLER_13_526 ();
 sg13g2_decap_4 FILLER_13_533 ();
 sg13g2_decap_4 FILLER_13_577 ();
 sg13g2_decap_8 FILLER_13_585 ();
 sg13g2_decap_4 FILLER_13_592 ();
 sg13g2_fill_2 FILLER_13_596 ();
 sg13g2_decap_8 FILLER_13_603 ();
 sg13g2_decap_4 FILLER_13_610 ();
 sg13g2_fill_1 FILLER_13_614 ();
 sg13g2_fill_1 FILLER_13_620 ();
 sg13g2_fill_1 FILLER_13_637 ();
 sg13g2_decap_4 FILLER_13_666 ();
 sg13g2_fill_2 FILLER_13_670 ();
 sg13g2_fill_2 FILLER_13_676 ();
 sg13g2_fill_1 FILLER_13_678 ();
 sg13g2_fill_1 FILLER_13_694 ();
 sg13g2_fill_1 FILLER_13_703 ();
 sg13g2_fill_1 FILLER_13_740 ();
 sg13g2_decap_8 FILLER_13_753 ();
 sg13g2_decap_8 FILLER_13_760 ();
 sg13g2_decap_8 FILLER_13_767 ();
 sg13g2_decap_8 FILLER_13_774 ();
 sg13g2_fill_2 FILLER_13_799 ();
 sg13g2_fill_1 FILLER_13_801 ();
 sg13g2_decap_8 FILLER_13_815 ();
 sg13g2_decap_8 FILLER_13_822 ();
 sg13g2_decap_8 FILLER_13_829 ();
 sg13g2_fill_1 FILLER_13_836 ();
 sg13g2_fill_2 FILLER_13_841 ();
 sg13g2_fill_1 FILLER_13_843 ();
 sg13g2_fill_1 FILLER_13_870 ();
 sg13g2_fill_1 FILLER_13_874 ();
 sg13g2_fill_1 FILLER_13_909 ();
 sg13g2_fill_1 FILLER_13_928 ();
 sg13g2_fill_2 FILLER_13_948 ();
 sg13g2_fill_2 FILLER_13_976 ();
 sg13g2_fill_2 FILLER_13_1000 ();
 sg13g2_fill_2 FILLER_13_1023 ();
 sg13g2_decap_4 FILLER_13_1054 ();
 sg13g2_fill_1 FILLER_13_1058 ();
 sg13g2_fill_1 FILLER_13_1068 ();
 sg13g2_decap_4 FILLER_13_1109 ();
 sg13g2_fill_2 FILLER_13_1113 ();
 sg13g2_fill_2 FILLER_13_1121 ();
 sg13g2_fill_1 FILLER_13_1123 ();
 sg13g2_decap_8 FILLER_13_1144 ();
 sg13g2_decap_8 FILLER_13_1151 ();
 sg13g2_decap_4 FILLER_13_1158 ();
 sg13g2_decap_4 FILLER_13_1188 ();
 sg13g2_decap_4 FILLER_13_1218 ();
 sg13g2_fill_1 FILLER_13_1267 ();
 sg13g2_fill_1 FILLER_13_1302 ();
 sg13g2_decap_8 FILLER_13_1309 ();
 sg13g2_fill_2 FILLER_13_1363 ();
 sg13g2_fill_2 FILLER_13_1388 ();
 sg13g2_fill_2 FILLER_13_1408 ();
 sg13g2_fill_1 FILLER_13_1443 ();
 sg13g2_decap_8 FILLER_13_1482 ();
 sg13g2_decap_4 FILLER_13_1489 ();
 sg13g2_fill_1 FILLER_13_1505 ();
 sg13g2_decap_4 FILLER_13_1516 ();
 sg13g2_decap_4 FILLER_13_1546 ();
 sg13g2_fill_2 FILLER_13_1550 ();
 sg13g2_decap_8 FILLER_13_1558 ();
 sg13g2_decap_8 FILLER_13_1565 ();
 sg13g2_decap_8 FILLER_13_1572 ();
 sg13g2_decap_8 FILLER_13_1579 ();
 sg13g2_decap_8 FILLER_13_1586 ();
 sg13g2_fill_2 FILLER_13_1611 ();
 sg13g2_fill_1 FILLER_13_1613 ();
 sg13g2_decap_4 FILLER_13_1627 ();
 sg13g2_fill_1 FILLER_13_1631 ();
 sg13g2_fill_2 FILLER_13_1658 ();
 sg13g2_fill_2 FILLER_13_1666 ();
 sg13g2_fill_2 FILLER_13_1678 ();
 sg13g2_fill_1 FILLER_13_1712 ();
 sg13g2_fill_1 FILLER_13_1742 ();
 sg13g2_decap_8 FILLER_13_1783 ();
 sg13g2_decap_8 FILLER_13_1790 ();
 sg13g2_decap_8 FILLER_13_1797 ();
 sg13g2_decap_4 FILLER_13_1804 ();
 sg13g2_fill_2 FILLER_13_1808 ();
 sg13g2_fill_1 FILLER_13_1825 ();
 sg13g2_fill_2 FILLER_13_1874 ();
 sg13g2_fill_1 FILLER_13_1899 ();
 sg13g2_fill_2 FILLER_13_1908 ();
 sg13g2_fill_1 FILLER_13_1936 ();
 sg13g2_fill_2 FILLER_13_1969 ();
 sg13g2_fill_1 FILLER_13_1971 ();
 sg13g2_decap_4 FILLER_13_1986 ();
 sg13g2_fill_2 FILLER_13_2001 ();
 sg13g2_fill_1 FILLER_13_2003 ();
 sg13g2_fill_1 FILLER_13_2009 ();
 sg13g2_fill_1 FILLER_13_2035 ();
 sg13g2_fill_1 FILLER_13_2041 ();
 sg13g2_fill_2 FILLER_13_2045 ();
 sg13g2_fill_1 FILLER_13_2047 ();
 sg13g2_fill_1 FILLER_13_2072 ();
 sg13g2_fill_1 FILLER_13_2083 ();
 sg13g2_fill_2 FILLER_13_2117 ();
 sg13g2_fill_1 FILLER_13_2141 ();
 sg13g2_decap_4 FILLER_13_2188 ();
 sg13g2_fill_2 FILLER_13_2192 ();
 sg13g2_fill_1 FILLER_13_2236 ();
 sg13g2_fill_2 FILLER_13_2253 ();
 sg13g2_fill_2 FILLER_13_2272 ();
 sg13g2_decap_8 FILLER_13_2286 ();
 sg13g2_decap_8 FILLER_13_2293 ();
 sg13g2_fill_1 FILLER_13_2300 ();
 sg13g2_decap_8 FILLER_13_2331 ();
 sg13g2_decap_4 FILLER_13_2364 ();
 sg13g2_fill_2 FILLER_13_2398 ();
 sg13g2_fill_1 FILLER_13_2400 ();
 sg13g2_decap_4 FILLER_13_2412 ();
 sg13g2_fill_1 FILLER_13_2416 ();
 sg13g2_fill_1 FILLER_13_2461 ();
 sg13g2_fill_1 FILLER_13_2492 ();
 sg13g2_fill_2 FILLER_13_2501 ();
 sg13g2_decap_4 FILLER_13_2510 ();
 sg13g2_fill_2 FILLER_13_2514 ();
 sg13g2_decap_8 FILLER_13_2520 ();
 sg13g2_fill_1 FILLER_13_2527 ();
 sg13g2_decap_4 FILLER_13_2532 ();
 sg13g2_decap_4 FILLER_13_2571 ();
 sg13g2_fill_1 FILLER_13_2579 ();
 sg13g2_decap_8 FILLER_13_2653 ();
 sg13g2_decap_8 FILLER_13_2660 ();
 sg13g2_fill_2 FILLER_13_2667 ();
 sg13g2_fill_1 FILLER_13_2669 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_33 ();
 sg13g2_decap_8 FILLER_14_61 ();
 sg13g2_decap_8 FILLER_14_68 ();
 sg13g2_decap_8 FILLER_14_75 ();
 sg13g2_decap_8 FILLER_14_82 ();
 sg13g2_decap_4 FILLER_14_89 ();
 sg13g2_fill_1 FILLER_14_93 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_fill_1 FILLER_14_108 ();
 sg13g2_decap_4 FILLER_14_122 ();
 sg13g2_fill_2 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_136 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_fill_1 FILLER_14_172 ();
 sg13g2_fill_2 FILLER_14_190 ();
 sg13g2_fill_1 FILLER_14_192 ();
 sg13g2_fill_1 FILLER_14_204 ();
 sg13g2_fill_1 FILLER_14_218 ();
 sg13g2_fill_2 FILLER_14_223 ();
 sg13g2_fill_1 FILLER_14_234 ();
 sg13g2_fill_1 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_4 FILLER_14_292 ();
 sg13g2_fill_1 FILLER_14_296 ();
 sg13g2_fill_2 FILLER_14_305 ();
 sg13g2_fill_1 FILLER_14_307 ();
 sg13g2_decap_8 FILLER_14_317 ();
 sg13g2_decap_8 FILLER_14_324 ();
 sg13g2_decap_8 FILLER_14_331 ();
 sg13g2_decap_8 FILLER_14_338 ();
 sg13g2_decap_8 FILLER_14_345 ();
 sg13g2_decap_4 FILLER_14_352 ();
 sg13g2_decap_8 FILLER_14_391 ();
 sg13g2_decap_8 FILLER_14_398 ();
 sg13g2_decap_8 FILLER_14_405 ();
 sg13g2_decap_8 FILLER_14_412 ();
 sg13g2_fill_2 FILLER_14_419 ();
 sg13g2_fill_1 FILLER_14_426 ();
 sg13g2_fill_1 FILLER_14_453 ();
 sg13g2_fill_2 FILLER_14_457 ();
 sg13g2_decap_8 FILLER_14_475 ();
 sg13g2_decap_4 FILLER_14_482 ();
 sg13g2_fill_2 FILLER_14_486 ();
 sg13g2_fill_2 FILLER_14_516 ();
 sg13g2_fill_1 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_545 ();
 sg13g2_decap_8 FILLER_14_552 ();
 sg13g2_decap_8 FILLER_14_559 ();
 sg13g2_decap_8 FILLER_14_566 ();
 sg13g2_fill_1 FILLER_14_573 ();
 sg13g2_fill_2 FILLER_14_579 ();
 sg13g2_decap_4 FILLER_14_591 ();
 sg13g2_fill_2 FILLER_14_599 ();
 sg13g2_fill_1 FILLER_14_601 ();
 sg13g2_decap_8 FILLER_14_606 ();
 sg13g2_fill_2 FILLER_14_613 ();
 sg13g2_fill_1 FILLER_14_615 ();
 sg13g2_fill_1 FILLER_14_625 ();
 sg13g2_decap_4 FILLER_14_674 ();
 sg13g2_fill_1 FILLER_14_683 ();
 sg13g2_decap_4 FILLER_14_692 ();
 sg13g2_decap_8 FILLER_14_701 ();
 sg13g2_decap_4 FILLER_14_708 ();
 sg13g2_fill_1 FILLER_14_712 ();
 sg13g2_decap_4 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_745 ();
 sg13g2_decap_4 FILLER_14_752 ();
 sg13g2_fill_1 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_762 ();
 sg13g2_fill_1 FILLER_14_769 ();
 sg13g2_fill_2 FILLER_14_842 ();
 sg13g2_fill_1 FILLER_14_844 ();
 sg13g2_fill_1 FILLER_14_854 ();
 sg13g2_fill_2 FILLER_14_873 ();
 sg13g2_decap_4 FILLER_14_885 ();
 sg13g2_fill_2 FILLER_14_889 ();
 sg13g2_fill_1 FILLER_14_917 ();
 sg13g2_fill_1 FILLER_14_998 ();
 sg13g2_fill_2 FILLER_14_1016 ();
 sg13g2_fill_2 FILLER_14_1029 ();
 sg13g2_fill_2 FILLER_14_1063 ();
 sg13g2_fill_1 FILLER_14_1065 ();
 sg13g2_decap_8 FILLER_14_1076 ();
 sg13g2_fill_2 FILLER_14_1083 ();
 sg13g2_fill_1 FILLER_14_1085 ();
 sg13g2_fill_2 FILLER_14_1096 ();
 sg13g2_fill_1 FILLER_14_1098 ();
 sg13g2_fill_2 FILLER_14_1105 ();
 sg13g2_fill_1 FILLER_14_1133 ();
 sg13g2_decap_8 FILLER_14_1160 ();
 sg13g2_fill_1 FILLER_14_1167 ();
 sg13g2_fill_1 FILLER_14_1209 ();
 sg13g2_fill_2 FILLER_14_1258 ();
 sg13g2_fill_1 FILLER_14_1260 ();
 sg13g2_fill_2 FILLER_14_1284 ();
 sg13g2_fill_2 FILLER_14_1305 ();
 sg13g2_fill_2 FILLER_14_1343 ();
 sg13g2_fill_1 FILLER_14_1351 ();
 sg13g2_fill_2 FILLER_14_1378 ();
 sg13g2_fill_2 FILLER_14_1474 ();
 sg13g2_fill_1 FILLER_14_1476 ();
 sg13g2_decap_8 FILLER_14_1483 ();
 sg13g2_decap_4 FILLER_14_1490 ();
 sg13g2_decap_8 FILLER_14_1499 ();
 sg13g2_decap_8 FILLER_14_1506 ();
 sg13g2_decap_8 FILLER_14_1513 ();
 sg13g2_fill_1 FILLER_14_1520 ();
 sg13g2_fill_2 FILLER_14_1550 ();
 sg13g2_fill_2 FILLER_14_1555 ();
 sg13g2_decap_4 FILLER_14_1561 ();
 sg13g2_fill_2 FILLER_14_1565 ();
 sg13g2_fill_1 FILLER_14_1577 ();
 sg13g2_fill_2 FILLER_14_1604 ();
 sg13g2_decap_8 FILLER_14_1632 ();
 sg13g2_decap_8 FILLER_14_1639 ();
 sg13g2_decap_8 FILLER_14_1646 ();
 sg13g2_decap_4 FILLER_14_1653 ();
 sg13g2_fill_2 FILLER_14_1666 ();
 sg13g2_fill_2 FILLER_14_1808 ();
 sg13g2_fill_1 FILLER_14_1817 ();
 sg13g2_fill_1 FILLER_14_1828 ();
 sg13g2_decap_8 FILLER_14_1833 ();
 sg13g2_decap_8 FILLER_14_1840 ();
 sg13g2_fill_1 FILLER_14_1847 ();
 sg13g2_decap_4 FILLER_14_1856 ();
 sg13g2_fill_2 FILLER_14_1860 ();
 sg13g2_decap_8 FILLER_14_1876 ();
 sg13g2_fill_1 FILLER_14_1938 ();
 sg13g2_fill_1 FILLER_14_1963 ();
 sg13g2_decap_4 FILLER_14_1976 ();
 sg13g2_decap_4 FILLER_14_1990 ();
 sg13g2_fill_1 FILLER_14_2003 ();
 sg13g2_fill_1 FILLER_14_2009 ();
 sg13g2_fill_1 FILLER_14_2020 ();
 sg13g2_decap_4 FILLER_14_2025 ();
 sg13g2_fill_1 FILLER_14_2029 ();
 sg13g2_fill_2 FILLER_14_2044 ();
 sg13g2_fill_2 FILLER_14_2055 ();
 sg13g2_fill_1 FILLER_14_2057 ();
 sg13g2_fill_1 FILLER_14_2064 ();
 sg13g2_fill_2 FILLER_14_2077 ();
 sg13g2_fill_1 FILLER_14_2085 ();
 sg13g2_fill_1 FILLER_14_2100 ();
 sg13g2_fill_1 FILLER_14_2123 ();
 sg13g2_fill_2 FILLER_14_2180 ();
 sg13g2_fill_2 FILLER_14_2243 ();
 sg13g2_decap_8 FILLER_14_2271 ();
 sg13g2_decap_8 FILLER_14_2278 ();
 sg13g2_decap_8 FILLER_14_2285 ();
 sg13g2_decap_8 FILLER_14_2292 ();
 sg13g2_fill_2 FILLER_14_2299 ();
 sg13g2_fill_1 FILLER_14_2301 ();
 sg13g2_fill_1 FILLER_14_2308 ();
 sg13g2_fill_1 FILLER_14_2313 ();
 sg13g2_fill_1 FILLER_14_2318 ();
 sg13g2_fill_1 FILLER_14_2323 ();
 sg13g2_fill_2 FILLER_14_2385 ();
 sg13g2_fill_2 FILLER_14_2392 ();
 sg13g2_decap_8 FILLER_14_2407 ();
 sg13g2_decap_8 FILLER_14_2414 ();
 sg13g2_decap_4 FILLER_14_2421 ();
 sg13g2_fill_1 FILLER_14_2425 ();
 sg13g2_fill_2 FILLER_14_2430 ();
 sg13g2_decap_4 FILLER_14_2466 ();
 sg13g2_fill_1 FILLER_14_2490 ();
 sg13g2_decap_4 FILLER_14_2495 ();
 sg13g2_fill_1 FILLER_14_2512 ();
 sg13g2_fill_2 FILLER_14_2521 ();
 sg13g2_fill_1 FILLER_14_2523 ();
 sg13g2_fill_1 FILLER_14_2529 ();
 sg13g2_fill_1 FILLER_14_2535 ();
 sg13g2_fill_1 FILLER_14_2541 ();
 sg13g2_decap_8 FILLER_14_2568 ();
 sg13g2_decap_8 FILLER_14_2575 ();
 sg13g2_fill_2 FILLER_14_2582 ();
 sg13g2_fill_1 FILLER_14_2590 ();
 sg13g2_fill_2 FILLER_14_2597 ();
 sg13g2_fill_2 FILLER_14_2603 ();
 sg13g2_decap_8 FILLER_14_2609 ();
 sg13g2_fill_2 FILLER_14_2616 ();
 sg13g2_decap_8 FILLER_14_2640 ();
 sg13g2_decap_8 FILLER_14_2647 ();
 sg13g2_decap_8 FILLER_14_2654 ();
 sg13g2_decap_8 FILLER_14_2661 ();
 sg13g2_fill_2 FILLER_14_2668 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_fill_1 FILLER_15_7 ();
 sg13g2_fill_2 FILLER_15_33 ();
 sg13g2_fill_1 FILLER_15_35 ();
 sg13g2_decap_8 FILLER_15_43 ();
 sg13g2_fill_2 FILLER_15_50 ();
 sg13g2_decap_8 FILLER_15_56 ();
 sg13g2_decap_8 FILLER_15_63 ();
 sg13g2_decap_8 FILLER_15_70 ();
 sg13g2_decap_8 FILLER_15_77 ();
 sg13g2_decap_8 FILLER_15_84 ();
 sg13g2_decap_4 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_103 ();
 sg13g2_fill_2 FILLER_15_114 ();
 sg13g2_fill_1 FILLER_15_148 ();
 sg13g2_decap_4 FILLER_15_161 ();
 sg13g2_fill_2 FILLER_15_165 ();
 sg13g2_fill_2 FILLER_15_173 ();
 sg13g2_fill_1 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_203 ();
 sg13g2_fill_1 FILLER_15_205 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_decap_4 FILLER_15_289 ();
 sg13g2_fill_2 FILLER_15_293 ();
 sg13g2_fill_1 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_304 ();
 sg13g2_decap_4 FILLER_15_311 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_4 FILLER_15_355 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_4 FILLER_15_419 ();
 sg13g2_fill_1 FILLER_15_423 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_fill_2 FILLER_15_476 ();
 sg13g2_fill_1 FILLER_15_478 ();
 sg13g2_decap_8 FILLER_15_483 ();
 sg13g2_decap_8 FILLER_15_490 ();
 sg13g2_decap_4 FILLER_15_497 ();
 sg13g2_fill_1 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_505 ();
 sg13g2_fill_2 FILLER_15_512 ();
 sg13g2_fill_1 FILLER_15_514 ();
 sg13g2_decap_8 FILLER_15_525 ();
 sg13g2_decap_4 FILLER_15_566 ();
 sg13g2_fill_2 FILLER_15_570 ();
 sg13g2_fill_2 FILLER_15_577 ();
 sg13g2_fill_2 FILLER_15_620 ();
 sg13g2_fill_1 FILLER_15_627 ();
 sg13g2_fill_1 FILLER_15_640 ();
 sg13g2_fill_1 FILLER_15_648 ();
 sg13g2_fill_2 FILLER_15_670 ();
 sg13g2_fill_1 FILLER_15_677 ();
 sg13g2_decap_4 FILLER_15_696 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_fill_1 FILLER_15_795 ();
 sg13g2_fill_2 FILLER_15_822 ();
 sg13g2_fill_1 FILLER_15_824 ();
 sg13g2_fill_2 FILLER_15_867 ();
 sg13g2_fill_2 FILLER_15_879 ();
 sg13g2_fill_1 FILLER_15_891 ();
 sg13g2_fill_2 FILLER_15_916 ();
 sg13g2_fill_1 FILLER_15_931 ();
 sg13g2_decap_8 FILLER_15_935 ();
 sg13g2_fill_1 FILLER_15_985 ();
 sg13g2_fill_2 FILLER_15_1039 ();
 sg13g2_decap_4 FILLER_15_1096 ();
 sg13g2_fill_2 FILLER_15_1100 ();
 sg13g2_fill_2 FILLER_15_1112 ();
 sg13g2_fill_2 FILLER_15_1120 ();
 sg13g2_fill_2 FILLER_15_1130 ();
 sg13g2_fill_1 FILLER_15_1132 ();
 sg13g2_decap_8 FILLER_15_1169 ();
 sg13g2_fill_1 FILLER_15_1176 ();
 sg13g2_decap_4 FILLER_15_1252 ();
 sg13g2_fill_2 FILLER_15_1295 ();
 sg13g2_fill_1 FILLER_15_1329 ();
 sg13g2_fill_1 FILLER_15_1342 ();
 sg13g2_fill_2 FILLER_15_1359 ();
 sg13g2_fill_1 FILLER_15_1361 ();
 sg13g2_decap_8 FILLER_15_1455 ();
 sg13g2_fill_2 FILLER_15_1462 ();
 sg13g2_fill_1 FILLER_15_1464 ();
 sg13g2_decap_8 FILLER_15_1495 ();
 sg13g2_fill_2 FILLER_15_1502 ();
 sg13g2_fill_1 FILLER_15_1504 ();
 sg13g2_fill_2 FILLER_15_1545 ();
 sg13g2_decap_4 FILLER_15_1553 ();
 sg13g2_fill_2 FILLER_15_1557 ();
 sg13g2_decap_8 FILLER_15_1564 ();
 sg13g2_decap_4 FILLER_15_1584 ();
 sg13g2_fill_1 FILLER_15_1603 ();
 sg13g2_decap_4 FILLER_15_1625 ();
 sg13g2_fill_2 FILLER_15_1629 ();
 sg13g2_decap_8 FILLER_15_1639 ();
 sg13g2_fill_2 FILLER_15_1646 ();
 sg13g2_fill_1 FILLER_15_1665 ();
 sg13g2_fill_1 FILLER_15_1707 ();
 sg13g2_fill_1 FILLER_15_1765 ();
 sg13g2_decap_4 FILLER_15_1799 ();
 sg13g2_fill_2 FILLER_15_1803 ();
 sg13g2_decap_8 FILLER_15_1831 ();
 sg13g2_decap_4 FILLER_15_1838 ();
 sg13g2_fill_2 FILLER_15_1842 ();
 sg13g2_decap_4 FILLER_15_1849 ();
 sg13g2_fill_1 FILLER_15_1853 ();
 sg13g2_decap_8 FILLER_15_1864 ();
 sg13g2_decap_4 FILLER_15_1871 ();
 sg13g2_fill_2 FILLER_15_1887 ();
 sg13g2_fill_1 FILLER_15_1889 ();
 sg13g2_fill_1 FILLER_15_1900 ();
 sg13g2_fill_1 FILLER_15_1913 ();
 sg13g2_decap_8 FILLER_15_1927 ();
 sg13g2_decap_8 FILLER_15_1969 ();
 sg13g2_fill_2 FILLER_15_1976 ();
 sg13g2_fill_1 FILLER_15_1978 ();
 sg13g2_fill_1 FILLER_15_1983 ();
 sg13g2_fill_1 FILLER_15_1993 ();
 sg13g2_fill_1 FILLER_15_2002 ();
 sg13g2_fill_2 FILLER_15_2026 ();
 sg13g2_fill_1 FILLER_15_2028 ();
 sg13g2_decap_4 FILLER_15_2034 ();
 sg13g2_fill_1 FILLER_15_2038 ();
 sg13g2_decap_4 FILLER_15_2051 ();
 sg13g2_fill_2 FILLER_15_2055 ();
 sg13g2_decap_8 FILLER_15_2069 ();
 sg13g2_decap_4 FILLER_15_2076 ();
 sg13g2_fill_2 FILLER_15_2089 ();
 sg13g2_fill_1 FILLER_15_2091 ();
 sg13g2_decap_4 FILLER_15_2117 ();
 sg13g2_fill_2 FILLER_15_2152 ();
 sg13g2_fill_1 FILLER_15_2206 ();
 sg13g2_fill_1 FILLER_15_2222 ();
 sg13g2_fill_1 FILLER_15_2240 ();
 sg13g2_fill_2 FILLER_15_2251 ();
 sg13g2_decap_8 FILLER_15_2266 ();
 sg13g2_fill_2 FILLER_15_2283 ();
 sg13g2_fill_2 FILLER_15_2291 ();
 sg13g2_fill_1 FILLER_15_2293 ();
 sg13g2_fill_2 FILLER_15_2306 ();
 sg13g2_fill_1 FILLER_15_2308 ();
 sg13g2_fill_2 FILLER_15_2343 ();
 sg13g2_fill_1 FILLER_15_2345 ();
 sg13g2_fill_2 FILLER_15_2350 ();
 sg13g2_fill_2 FILLER_15_2356 ();
 sg13g2_fill_2 FILLER_15_2362 ();
 sg13g2_fill_2 FILLER_15_2376 ();
 sg13g2_fill_1 FILLER_15_2378 ();
 sg13g2_decap_4 FILLER_15_2388 ();
 sg13g2_decap_8 FILLER_15_2395 ();
 sg13g2_decap_8 FILLER_15_2402 ();
 sg13g2_fill_1 FILLER_15_2409 ();
 sg13g2_fill_2 FILLER_15_2415 ();
 sg13g2_fill_1 FILLER_15_2417 ();
 sg13g2_fill_1 FILLER_15_2430 ();
 sg13g2_decap_4 FILLER_15_2436 ();
 sg13g2_decap_8 FILLER_15_2444 ();
 sg13g2_decap_4 FILLER_15_2451 ();
 sg13g2_fill_2 FILLER_15_2468 ();
 sg13g2_fill_1 FILLER_15_2514 ();
 sg13g2_decap_8 FILLER_15_2559 ();
 sg13g2_fill_2 FILLER_15_2566 ();
 sg13g2_fill_1 FILLER_15_2576 ();
 sg13g2_decap_8 FILLER_15_2607 ();
 sg13g2_decap_8 FILLER_15_2614 ();
 sg13g2_decap_8 FILLER_15_2621 ();
 sg13g2_decap_8 FILLER_15_2628 ();
 sg13g2_decap_8 FILLER_15_2635 ();
 sg13g2_decap_8 FILLER_15_2642 ();
 sg13g2_decap_8 FILLER_15_2649 ();
 sg13g2_decap_8 FILLER_15_2656 ();
 sg13g2_decap_8 FILLER_15_2663 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_fill_2 FILLER_16_52 ();
 sg13g2_fill_1 FILLER_16_54 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_4 FILLER_16_91 ();
 sg13g2_fill_1 FILLER_16_100 ();
 sg13g2_fill_1 FILLER_16_146 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_162 ();
 sg13g2_fill_1 FILLER_16_181 ();
 sg13g2_fill_1 FILLER_16_188 ();
 sg13g2_fill_2 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_247 ();
 sg13g2_decap_4 FILLER_16_253 ();
 sg13g2_decap_4 FILLER_16_262 ();
 sg13g2_fill_1 FILLER_16_272 ();
 sg13g2_fill_1 FILLER_16_291 ();
 sg13g2_fill_1 FILLER_16_297 ();
 sg13g2_fill_2 FILLER_16_302 ();
 sg13g2_fill_1 FILLER_16_304 ();
 sg13g2_fill_1 FILLER_16_309 ();
 sg13g2_fill_2 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_326 ();
 sg13g2_decap_8 FILLER_16_333 ();
 sg13g2_decap_8 FILLER_16_340 ();
 sg13g2_decap_8 FILLER_16_347 ();
 sg13g2_decap_4 FILLER_16_354 ();
 sg13g2_decap_4 FILLER_16_363 ();
 sg13g2_fill_1 FILLER_16_367 ();
 sg13g2_fill_1 FILLER_16_381 ();
 sg13g2_fill_2 FILLER_16_395 ();
 sg13g2_fill_1 FILLER_16_397 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_4 FILLER_16_455 ();
 sg13g2_fill_2 FILLER_16_459 ();
 sg13g2_fill_1 FILLER_16_471 ();
 sg13g2_decap_8 FILLER_16_481 ();
 sg13g2_decap_8 FILLER_16_488 ();
 sg13g2_decap_8 FILLER_16_495 ();
 sg13g2_decap_8 FILLER_16_502 ();
 sg13g2_fill_1 FILLER_16_509 ();
 sg13g2_fill_1 FILLER_16_540 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_4 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_561 ();
 sg13g2_fill_2 FILLER_16_568 ();
 sg13g2_fill_1 FILLER_16_623 ();
 sg13g2_fill_1 FILLER_16_672 ();
 sg13g2_fill_1 FILLER_16_678 ();
 sg13g2_fill_1 FILLER_16_726 ();
 sg13g2_fill_1 FILLER_16_731 ();
 sg13g2_fill_2 FILLER_16_737 ();
 sg13g2_fill_1 FILLER_16_739 ();
 sg13g2_decap_8 FILLER_16_750 ();
 sg13g2_fill_2 FILLER_16_757 ();
 sg13g2_fill_2 FILLER_16_765 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_fill_1 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_816 ();
 sg13g2_decap_8 FILLER_16_823 ();
 sg13g2_decap_8 FILLER_16_830 ();
 sg13g2_decap_4 FILLER_16_837 ();
 sg13g2_fill_2 FILLER_16_841 ();
 sg13g2_decap_8 FILLER_16_852 ();
 sg13g2_fill_2 FILLER_16_859 ();
 sg13g2_fill_2 FILLER_16_864 ();
 sg13g2_decap_8 FILLER_16_901 ();
 sg13g2_fill_2 FILLER_16_908 ();
 sg13g2_fill_1 FILLER_16_910 ();
 sg13g2_decap_4 FILLER_16_926 ();
 sg13g2_fill_1 FILLER_16_930 ();
 sg13g2_fill_2 FILLER_16_944 ();
 sg13g2_fill_1 FILLER_16_946 ();
 sg13g2_fill_2 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_974 ();
 sg13g2_fill_2 FILLER_16_986 ();
 sg13g2_fill_1 FILLER_16_988 ();
 sg13g2_fill_1 FILLER_16_1015 ();
 sg13g2_fill_1 FILLER_16_1021 ();
 sg13g2_fill_2 FILLER_16_1081 ();
 sg13g2_fill_2 FILLER_16_1096 ();
 sg13g2_fill_1 FILLER_16_1098 ();
 sg13g2_decap_8 FILLER_16_1103 ();
 sg13g2_decap_4 FILLER_16_1110 ();
 sg13g2_fill_2 FILLER_16_1114 ();
 sg13g2_decap_4 FILLER_16_1121 ();
 sg13g2_fill_1 FILLER_16_1125 ();
 sg13g2_decap_8 FILLER_16_1136 ();
 sg13g2_decap_8 FILLER_16_1143 ();
 sg13g2_decap_4 FILLER_16_1150 ();
 sg13g2_decap_8 FILLER_16_1170 ();
 sg13g2_decap_8 FILLER_16_1177 ();
 sg13g2_fill_2 FILLER_16_1198 ();
 sg13g2_decap_8 FILLER_16_1203 ();
 sg13g2_fill_2 FILLER_16_1210 ();
 sg13g2_fill_1 FILLER_16_1212 ();
 sg13g2_decap_8 FILLER_16_1216 ();
 sg13g2_fill_1 FILLER_16_1223 ();
 sg13g2_fill_1 FILLER_16_1255 ();
 sg13g2_fill_2 FILLER_16_1318 ();
 sg13g2_decap_8 FILLER_16_1362 ();
 sg13g2_decap_8 FILLER_16_1395 ();
 sg13g2_fill_2 FILLER_16_1402 ();
 sg13g2_fill_1 FILLER_16_1404 ();
 sg13g2_decap_8 FILLER_16_1410 ();
 sg13g2_decap_8 FILLER_16_1422 ();
 sg13g2_fill_2 FILLER_16_1429 ();
 sg13g2_decap_8 FILLER_16_1447 ();
 sg13g2_decap_8 FILLER_16_1454 ();
 sg13g2_decap_8 FILLER_16_1461 ();
 sg13g2_fill_2 FILLER_16_1468 ();
 sg13g2_fill_1 FILLER_16_1470 ();
 sg13g2_decap_4 FILLER_16_1565 ();
 sg13g2_fill_2 FILLER_16_1569 ();
 sg13g2_decap_4 FILLER_16_1579 ();
 sg13g2_decap_8 FILLER_16_1599 ();
 sg13g2_decap_4 FILLER_16_1606 ();
 sg13g2_fill_1 FILLER_16_1610 ();
 sg13g2_decap_8 FILLER_16_1650 ();
 sg13g2_decap_4 FILLER_16_1657 ();
 sg13g2_fill_2 FILLER_16_1661 ();
 sg13g2_fill_2 FILLER_16_1673 ();
 sg13g2_fill_2 FILLER_16_1689 ();
 sg13g2_fill_1 FILLER_16_1712 ();
 sg13g2_fill_1 FILLER_16_1724 ();
 sg13g2_fill_1 FILLER_16_1734 ();
 sg13g2_fill_1 FILLER_16_1743 ();
 sg13g2_decap_4 FILLER_16_1814 ();
 sg13g2_fill_2 FILLER_16_1818 ();
 sg13g2_fill_1 FILLER_16_1826 ();
 sg13g2_decap_4 FILLER_16_1870 ();
 sg13g2_fill_1 FILLER_16_1874 ();
 sg13g2_fill_2 FILLER_16_1904 ();
 sg13g2_fill_1 FILLER_16_1906 ();
 sg13g2_fill_2 FILLER_16_1910 ();
 sg13g2_fill_1 FILLER_16_1912 ();
 sg13g2_decap_4 FILLER_16_1918 ();
 sg13g2_fill_1 FILLER_16_1922 ();
 sg13g2_fill_1 FILLER_16_1931 ();
 sg13g2_fill_1 FILLER_16_1940 ();
 sg13g2_fill_2 FILLER_16_2006 ();
 sg13g2_fill_1 FILLER_16_2027 ();
 sg13g2_fill_1 FILLER_16_2059 ();
 sg13g2_fill_2 FILLER_16_2076 ();
 sg13g2_fill_2 FILLER_16_2087 ();
 sg13g2_fill_1 FILLER_16_2097 ();
 sg13g2_fill_1 FILLER_16_2130 ();
 sg13g2_decap_8 FILLER_16_2154 ();
 sg13g2_fill_2 FILLER_16_2161 ();
 sg13g2_fill_2 FILLER_16_2168 ();
 sg13g2_fill_1 FILLER_16_2170 ();
 sg13g2_fill_2 FILLER_16_2178 ();
 sg13g2_decap_4 FILLER_16_2190 ();
 sg13g2_fill_2 FILLER_16_2206 ();
 sg13g2_fill_1 FILLER_16_2211 ();
 sg13g2_fill_1 FILLER_16_2252 ();
 sg13g2_fill_2 FILLER_16_2282 ();
 sg13g2_fill_1 FILLER_16_2284 ();
 sg13g2_fill_2 FILLER_16_2298 ();
 sg13g2_decap_8 FILLER_16_2314 ();
 sg13g2_decap_8 FILLER_16_2321 ();
 sg13g2_decap_8 FILLER_16_2328 ();
 sg13g2_decap_8 FILLER_16_2335 ();
 sg13g2_decap_8 FILLER_16_2342 ();
 sg13g2_fill_2 FILLER_16_2385 ();
 sg13g2_fill_2 FILLER_16_2413 ();
 sg13g2_fill_1 FILLER_16_2415 ();
 sg13g2_decap_8 FILLER_16_2442 ();
 sg13g2_fill_1 FILLER_16_2449 ();
 sg13g2_decap_8 FILLER_16_2489 ();
 sg13g2_fill_2 FILLER_16_2496 ();
 sg13g2_fill_1 FILLER_16_2498 ();
 sg13g2_decap_4 FILLER_16_2503 ();
 sg13g2_fill_2 FILLER_16_2507 ();
 sg13g2_decap_8 FILLER_16_2548 ();
 sg13g2_decap_4 FILLER_16_2612 ();
 sg13g2_fill_2 FILLER_16_2616 ();
 sg13g2_decap_8 FILLER_16_2622 ();
 sg13g2_decap_4 FILLER_16_2629 ();
 sg13g2_decap_8 FILLER_16_2663 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_2 FILLER_17_6 ();
 sg13g2_fill_1 FILLER_17_8 ();
 sg13g2_fill_1 FILLER_17_17 ();
 sg13g2_fill_2 FILLER_17_57 ();
 sg13g2_decap_4 FILLER_17_89 ();
 sg13g2_fill_2 FILLER_17_93 ();
 sg13g2_fill_2 FILLER_17_100 ();
 sg13g2_fill_1 FILLER_17_121 ();
 sg13g2_fill_2 FILLER_17_133 ();
 sg13g2_fill_1 FILLER_17_150 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_1 FILLER_17_168 ();
 sg13g2_fill_2 FILLER_17_184 ();
 sg13g2_fill_1 FILLER_17_191 ();
 sg13g2_fill_1 FILLER_17_197 ();
 sg13g2_fill_1 FILLER_17_203 ();
 sg13g2_fill_1 FILLER_17_210 ();
 sg13g2_decap_4 FILLER_17_247 ();
 sg13g2_fill_1 FILLER_17_251 ();
 sg13g2_fill_2 FILLER_17_278 ();
 sg13g2_fill_2 FILLER_17_303 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_decap_8 FILLER_17_324 ();
 sg13g2_decap_8 FILLER_17_331 ();
 sg13g2_fill_2 FILLER_17_338 ();
 sg13g2_decap_4 FILLER_17_366 ();
 sg13g2_fill_2 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_376 ();
 sg13g2_fill_1 FILLER_17_383 ();
 sg13g2_fill_2 FILLER_17_410 ();
 sg13g2_decap_4 FILLER_17_452 ();
 sg13g2_fill_1 FILLER_17_456 ();
 sg13g2_decap_8 FILLER_17_491 ();
 sg13g2_decap_8 FILLER_17_498 ();
 sg13g2_decap_8 FILLER_17_505 ();
 sg13g2_fill_2 FILLER_17_512 ();
 sg13g2_fill_1 FILLER_17_514 ();
 sg13g2_decap_4 FILLER_17_525 ();
 sg13g2_decap_8 FILLER_17_559 ();
 sg13g2_decap_8 FILLER_17_566 ();
 sg13g2_fill_2 FILLER_17_612 ();
 sg13g2_fill_1 FILLER_17_614 ();
 sg13g2_fill_1 FILLER_17_648 ();
 sg13g2_fill_2 FILLER_17_654 ();
 sg13g2_fill_1 FILLER_17_677 ();
 sg13g2_fill_2 FILLER_17_734 ();
 sg13g2_fill_1 FILLER_17_736 ();
 sg13g2_fill_1 FILLER_17_763 ();
 sg13g2_decap_4 FILLER_17_790 ();
 sg13g2_decap_8 FILLER_17_799 ();
 sg13g2_decap_8 FILLER_17_806 ();
 sg13g2_decap_4 FILLER_17_813 ();
 sg13g2_fill_2 FILLER_17_865 ();
 sg13g2_fill_1 FILLER_17_867 ();
 sg13g2_decap_4 FILLER_17_871 ();
 sg13g2_fill_1 FILLER_17_875 ();
 sg13g2_decap_8 FILLER_17_889 ();
 sg13g2_decap_8 FILLER_17_896 ();
 sg13g2_fill_2 FILLER_17_906 ();
 sg13g2_fill_1 FILLER_17_908 ();
 sg13g2_decap_4 FILLER_17_957 ();
 sg13g2_decap_8 FILLER_17_969 ();
 sg13g2_decap_4 FILLER_17_976 ();
 sg13g2_fill_2 FILLER_17_980 ();
 sg13g2_fill_1 FILLER_17_1014 ();
 sg13g2_fill_2 FILLER_17_1024 ();
 sg13g2_fill_1 FILLER_17_1035 ();
 sg13g2_fill_2 FILLER_17_1047 ();
 sg13g2_decap_8 FILLER_17_1064 ();
 sg13g2_fill_1 FILLER_17_1071 ();
 sg13g2_fill_1 FILLER_17_1083 ();
 sg13g2_fill_2 FILLER_17_1092 ();
 sg13g2_fill_2 FILLER_17_1097 ();
 sg13g2_fill_1 FILLER_17_1099 ();
 sg13g2_fill_2 FILLER_17_1126 ();
 sg13g2_fill_1 FILLER_17_1128 ();
 sg13g2_fill_2 FILLER_17_1135 ();
 sg13g2_fill_1 FILLER_17_1137 ();
 sg13g2_decap_8 FILLER_17_1151 ();
 sg13g2_decap_4 FILLER_17_1158 ();
 sg13g2_fill_1 FILLER_17_1162 ();
 sg13g2_decap_8 FILLER_17_1168 ();
 sg13g2_decap_8 FILLER_17_1175 ();
 sg13g2_decap_8 FILLER_17_1182 ();
 sg13g2_decap_8 FILLER_17_1189 ();
 sg13g2_fill_2 FILLER_17_1196 ();
 sg13g2_decap_4 FILLER_17_1224 ();
 sg13g2_decap_8 FILLER_17_1239 ();
 sg13g2_fill_1 FILLER_17_1246 ();
 sg13g2_decap_8 FILLER_17_1250 ();
 sg13g2_decap_4 FILLER_17_1257 ();
 sg13g2_fill_2 FILLER_17_1261 ();
 sg13g2_fill_1 FILLER_17_1285 ();
 sg13g2_fill_1 FILLER_17_1295 ();
 sg13g2_fill_2 FILLER_17_1301 ();
 sg13g2_fill_1 FILLER_17_1303 ();
 sg13g2_decap_8 FILLER_17_1308 ();
 sg13g2_decap_4 FILLER_17_1315 ();
 sg13g2_fill_1 FILLER_17_1319 ();
 sg13g2_fill_2 FILLER_17_1326 ();
 sg13g2_fill_1 FILLER_17_1328 ();
 sg13g2_decap_4 FILLER_17_1344 ();
 sg13g2_fill_2 FILLER_17_1348 ();
 sg13g2_decap_8 FILLER_17_1360 ();
 sg13g2_decap_8 FILLER_17_1367 ();
 sg13g2_decap_8 FILLER_17_1374 ();
 sg13g2_decap_4 FILLER_17_1381 ();
 sg13g2_fill_1 FILLER_17_1385 ();
 sg13g2_decap_8 FILLER_17_1389 ();
 sg13g2_decap_8 FILLER_17_1405 ();
 sg13g2_decap_8 FILLER_17_1412 ();
 sg13g2_decap_8 FILLER_17_1419 ();
 sg13g2_fill_2 FILLER_17_1426 ();
 sg13g2_decap_4 FILLER_17_1444 ();
 sg13g2_decap_8 FILLER_17_1454 ();
 sg13g2_fill_2 FILLER_17_1461 ();
 sg13g2_fill_1 FILLER_17_1463 ();
 sg13g2_fill_2 FILLER_17_1474 ();
 sg13g2_fill_2 FILLER_17_1486 ();
 sg13g2_fill_1 FILLER_17_1488 ();
 sg13g2_fill_2 FILLER_17_1495 ();
 sg13g2_fill_1 FILLER_17_1497 ();
 sg13g2_fill_1 FILLER_17_1514 ();
 sg13g2_fill_1 FILLER_17_1556 ();
 sg13g2_fill_2 FILLER_17_1583 ();
 sg13g2_fill_2 FILLER_17_1624 ();
 sg13g2_fill_2 FILLER_17_1629 ();
 sg13g2_fill_2 FILLER_17_1660 ();
 sg13g2_fill_1 FILLER_17_1662 ();
 sg13g2_fill_1 FILLER_17_1668 ();
 sg13g2_fill_1 FILLER_17_1738 ();
 sg13g2_decap_8 FILLER_17_1768 ();
 sg13g2_fill_2 FILLER_17_1775 ();
 sg13g2_decap_8 FILLER_17_1788 ();
 sg13g2_decap_4 FILLER_17_1795 ();
 sg13g2_fill_2 FILLER_17_1799 ();
 sg13g2_fill_2 FILLER_17_1804 ();
 sg13g2_fill_1 FILLER_17_1806 ();
 sg13g2_fill_2 FILLER_17_1815 ();
 sg13g2_fill_1 FILLER_17_1826 ();
 sg13g2_fill_1 FILLER_17_1860 ();
 sg13g2_fill_2 FILLER_17_1887 ();
 sg13g2_fill_2 FILLER_17_1897 ();
 sg13g2_decap_8 FILLER_17_1909 ();
 sg13g2_decap_8 FILLER_17_1916 ();
 sg13g2_decap_4 FILLER_17_1923 ();
 sg13g2_fill_2 FILLER_17_1931 ();
 sg13g2_decap_8 FILLER_17_1974 ();
 sg13g2_decap_4 FILLER_17_1985 ();
 sg13g2_fill_2 FILLER_17_1989 ();
 sg13g2_decap_4 FILLER_17_2001 ();
 sg13g2_fill_1 FILLER_17_2005 ();
 sg13g2_fill_2 FILLER_17_2014 ();
 sg13g2_fill_1 FILLER_17_2016 ();
 sg13g2_decap_8 FILLER_17_2020 ();
 sg13g2_decap_8 FILLER_17_2027 ();
 sg13g2_fill_1 FILLER_17_2034 ();
 sg13g2_fill_2 FILLER_17_2073 ();
 sg13g2_fill_1 FILLER_17_2075 ();
 sg13g2_decap_4 FILLER_17_2089 ();
 sg13g2_fill_1 FILLER_17_2106 ();
 sg13g2_decap_4 FILLER_17_2112 ();
 sg13g2_fill_2 FILLER_17_2116 ();
 sg13g2_decap_8 FILLER_17_2123 ();
 sg13g2_decap_4 FILLER_17_2130 ();
 sg13g2_decap_8 FILLER_17_2146 ();
 sg13g2_decap_8 FILLER_17_2153 ();
 sg13g2_decap_8 FILLER_17_2160 ();
 sg13g2_fill_1 FILLER_17_2167 ();
 sg13g2_decap_4 FILLER_17_2185 ();
 sg13g2_fill_1 FILLER_17_2189 ();
 sg13g2_decap_4 FILLER_17_2193 ();
 sg13g2_fill_2 FILLER_17_2233 ();
 sg13g2_fill_1 FILLER_17_2239 ();
 sg13g2_fill_2 FILLER_17_2263 ();
 sg13g2_fill_1 FILLER_17_2265 ();
 sg13g2_decap_4 FILLER_17_2292 ();
 sg13g2_fill_2 FILLER_17_2296 ();
 sg13g2_decap_8 FILLER_17_2304 ();
 sg13g2_decap_8 FILLER_17_2311 ();
 sg13g2_decap_8 FILLER_17_2318 ();
 sg13g2_decap_8 FILLER_17_2325 ();
 sg13g2_decap_4 FILLER_17_2332 ();
 sg13g2_fill_1 FILLER_17_2336 ();
 sg13g2_fill_1 FILLER_17_2375 ();
 sg13g2_fill_2 FILLER_17_2387 ();
 sg13g2_fill_2 FILLER_17_2415 ();
 sg13g2_fill_2 FILLER_17_2421 ();
 sg13g2_decap_8 FILLER_17_2453 ();
 sg13g2_decap_8 FILLER_17_2464 ();
 sg13g2_decap_8 FILLER_17_2471 ();
 sg13g2_decap_8 FILLER_17_2478 ();
 sg13g2_fill_2 FILLER_17_2485 ();
 sg13g2_fill_1 FILLER_17_2487 ();
 sg13g2_fill_2 FILLER_17_2523 ();
 sg13g2_fill_2 FILLER_17_2540 ();
 sg13g2_fill_1 FILLER_17_2558 ();
 sg13g2_decap_8 FILLER_17_2599 ();
 sg13g2_fill_1 FILLER_17_2606 ();
 sg13g2_decap_8 FILLER_17_2663 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_86 ();
 sg13g2_decap_8 FILLER_18_93 ();
 sg13g2_decap_8 FILLER_18_100 ();
 sg13g2_decap_8 FILLER_18_107 ();
 sg13g2_fill_2 FILLER_18_114 ();
 sg13g2_fill_1 FILLER_18_116 ();
 sg13g2_fill_2 FILLER_18_152 ();
 sg13g2_fill_1 FILLER_18_154 ();
 sg13g2_fill_2 FILLER_18_160 ();
 sg13g2_fill_1 FILLER_18_166 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_fill_1 FILLER_18_178 ();
 sg13g2_fill_2 FILLER_18_192 ();
 sg13g2_fill_1 FILLER_18_194 ();
 sg13g2_fill_1 FILLER_18_202 ();
 sg13g2_fill_2 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_277 ();
 sg13g2_fill_1 FILLER_18_289 ();
 sg13g2_fill_2 FILLER_18_295 ();
 sg13g2_decap_8 FILLER_18_302 ();
 sg13g2_decap_8 FILLER_18_309 ();
 sg13g2_decap_8 FILLER_18_316 ();
 sg13g2_decap_4 FILLER_18_323 ();
 sg13g2_fill_2 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_339 ();
 sg13g2_decap_8 FILLER_18_346 ();
 sg13g2_decap_8 FILLER_18_353 ();
 sg13g2_fill_2 FILLER_18_360 ();
 sg13g2_fill_1 FILLER_18_362 ();
 sg13g2_fill_2 FILLER_18_367 ();
 sg13g2_decap_8 FILLER_18_372 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_fill_2 FILLER_18_386 ();
 sg13g2_decap_8 FILLER_18_414 ();
 sg13g2_decap_8 FILLER_18_421 ();
 sg13g2_fill_1 FILLER_18_428 ();
 sg13g2_decap_4 FILLER_18_463 ();
 sg13g2_fill_1 FILLER_18_467 ();
 sg13g2_fill_2 FILLER_18_473 ();
 sg13g2_fill_1 FILLER_18_475 ();
 sg13g2_decap_4 FILLER_18_536 ();
 sg13g2_decap_8 FILLER_18_544 ();
 sg13g2_fill_1 FILLER_18_551 ();
 sg13g2_decap_4 FILLER_18_560 ();
 sg13g2_fill_2 FILLER_18_564 ();
 sg13g2_fill_1 FILLER_18_571 ();
 sg13g2_fill_1 FILLER_18_576 ();
 sg13g2_fill_1 FILLER_18_600 ();
 sg13g2_fill_2 FILLER_18_604 ();
 sg13g2_fill_1 FILLER_18_606 ();
 sg13g2_fill_1 FILLER_18_642 ();
 sg13g2_fill_1 FILLER_18_652 ();
 sg13g2_fill_1 FILLER_18_658 ();
 sg13g2_fill_1 FILLER_18_669 ();
 sg13g2_fill_2 FILLER_18_674 ();
 sg13g2_fill_1 FILLER_18_681 ();
 sg13g2_fill_2 FILLER_18_695 ();
 sg13g2_fill_2 FILLER_18_705 ();
 sg13g2_fill_2 FILLER_18_719 ();
 sg13g2_decap_4 FILLER_18_726 ();
 sg13g2_fill_1 FILLER_18_730 ();
 sg13g2_fill_2 FILLER_18_743 ();
 sg13g2_decap_4 FILLER_18_755 ();
 sg13g2_fill_2 FILLER_18_759 ();
 sg13g2_decap_8 FILLER_18_781 ();
 sg13g2_fill_2 FILLER_18_788 ();
 sg13g2_fill_1 FILLER_18_790 ();
 sg13g2_fill_2 FILLER_18_801 ();
 sg13g2_fill_1 FILLER_18_816 ();
 sg13g2_fill_2 FILLER_18_853 ();
 sg13g2_fill_2 FILLER_18_866 ();
 sg13g2_decap_8 FILLER_18_881 ();
 sg13g2_fill_2 FILLER_18_888 ();
 sg13g2_fill_1 FILLER_18_890 ();
 sg13g2_fill_2 FILLER_18_921 ();
 sg13g2_fill_2 FILLER_18_944 ();
 sg13g2_fill_1 FILLER_18_963 ();
 sg13g2_fill_2 FILLER_18_969 ();
 sg13g2_fill_2 FILLER_18_976 ();
 sg13g2_fill_1 FILLER_18_978 ();
 sg13g2_decap_8 FILLER_18_982 ();
 sg13g2_decap_8 FILLER_18_989 ();
 sg13g2_decap_8 FILLER_18_1005 ();
 sg13g2_fill_1 FILLER_18_1012 ();
 sg13g2_decap_4 FILLER_18_1017 ();
 sg13g2_fill_1 FILLER_18_1036 ();
 sg13g2_decap_8 FILLER_18_1046 ();
 sg13g2_decap_8 FILLER_18_1053 ();
 sg13g2_fill_1 FILLER_18_1060 ();
 sg13g2_fill_2 FILLER_18_1129 ();
 sg13g2_decap_8 FILLER_18_1192 ();
 sg13g2_fill_2 FILLER_18_1199 ();
 sg13g2_fill_1 FILLER_18_1201 ();
 sg13g2_decap_8 FILLER_18_1207 ();
 sg13g2_fill_2 FILLER_18_1214 ();
 sg13g2_fill_1 FILLER_18_1233 ();
 sg13g2_decap_8 FILLER_18_1242 ();
 sg13g2_decap_4 FILLER_18_1249 ();
 sg13g2_decap_8 FILLER_18_1258 ();
 sg13g2_decap_4 FILLER_18_1291 ();
 sg13g2_fill_1 FILLER_18_1300 ();
 sg13g2_decap_8 FILLER_18_1327 ();
 sg13g2_decap_8 FILLER_18_1334 ();
 sg13g2_fill_1 FILLER_18_1341 ();
 sg13g2_decap_4 FILLER_18_1368 ();
 sg13g2_fill_1 FILLER_18_1372 ();
 sg13g2_fill_2 FILLER_18_1402 ();
 sg13g2_fill_2 FILLER_18_1436 ();
 sg13g2_decap_4 FILLER_18_1493 ();
 sg13g2_fill_2 FILLER_18_1503 ();
 sg13g2_fill_2 FILLER_18_1547 ();
 sg13g2_fill_2 FILLER_18_1559 ();
 sg13g2_fill_1 FILLER_18_1561 ();
 sg13g2_fill_2 FILLER_18_1608 ();
 sg13g2_fill_1 FILLER_18_1676 ();
 sg13g2_fill_2 FILLER_18_1683 ();
 sg13g2_fill_1 FILLER_18_1691 ();
 sg13g2_fill_2 FILLER_18_1721 ();
 sg13g2_fill_1 FILLER_18_1806 ();
 sg13g2_fill_1 FILLER_18_1816 ();
 sg13g2_decap_8 FILLER_18_1830 ();
 sg13g2_fill_1 FILLER_18_1837 ();
 sg13g2_fill_1 FILLER_18_1853 ();
 sg13g2_fill_1 FILLER_18_1871 ();
 sg13g2_fill_2 FILLER_18_1904 ();
 sg13g2_decap_4 FILLER_18_1911 ();
 sg13g2_fill_2 FILLER_18_1915 ();
 sg13g2_fill_1 FILLER_18_1970 ();
 sg13g2_fill_2 FILLER_18_1981 ();
 sg13g2_decap_4 FILLER_18_1991 ();
 sg13g2_fill_1 FILLER_18_1995 ();
 sg13g2_decap_4 FILLER_18_2029 ();
 sg13g2_fill_2 FILLER_18_2033 ();
 sg13g2_decap_4 FILLER_18_2048 ();
 sg13g2_decap_8 FILLER_18_2066 ();
 sg13g2_decap_4 FILLER_18_2073 ();
 sg13g2_fill_2 FILLER_18_2108 ();
 sg13g2_fill_1 FILLER_18_2110 ();
 sg13g2_fill_1 FILLER_18_2142 ();
 sg13g2_decap_4 FILLER_18_2162 ();
 sg13g2_fill_1 FILLER_18_2166 ();
 sg13g2_fill_2 FILLER_18_2203 ();
 sg13g2_decap_4 FILLER_18_2249 ();
 sg13g2_decap_8 FILLER_18_2256 ();
 sg13g2_decap_8 FILLER_18_2263 ();
 sg13g2_decap_8 FILLER_18_2270 ();
 sg13g2_decap_4 FILLER_18_2277 ();
 sg13g2_fill_2 FILLER_18_2281 ();
 sg13g2_decap_4 FILLER_18_2292 ();
 sg13g2_fill_2 FILLER_18_2296 ();
 sg13g2_decap_4 FILLER_18_2407 ();
 sg13g2_decap_4 FILLER_18_2417 ();
 sg13g2_fill_2 FILLER_18_2421 ();
 sg13g2_decap_8 FILLER_18_2427 ();
 sg13g2_fill_1 FILLER_18_2434 ();
 sg13g2_decap_8 FILLER_18_2439 ();
 sg13g2_decap_8 FILLER_18_2446 ();
 sg13g2_decap_4 FILLER_18_2453 ();
 sg13g2_decap_4 FILLER_18_2492 ();
 sg13g2_fill_2 FILLER_18_2496 ();
 sg13g2_decap_8 FILLER_18_2560 ();
 sg13g2_fill_1 FILLER_18_2567 ();
 sg13g2_decap_4 FILLER_18_2572 ();
 sg13g2_fill_2 FILLER_18_2576 ();
 sg13g2_decap_4 FILLER_18_2586 ();
 sg13g2_fill_2 FILLER_18_2604 ();
 sg13g2_fill_2 FILLER_18_2642 ();
 sg13g2_fill_1 FILLER_18_2648 ();
 sg13g2_fill_2 FILLER_18_2653 ();
 sg13g2_decap_8 FILLER_18_2659 ();
 sg13g2_decap_4 FILLER_18_2666 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_4 FILLER_19_35 ();
 sg13g2_fill_1 FILLER_19_39 ();
 sg13g2_decap_8 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_50 ();
 sg13g2_fill_2 FILLER_19_59 ();
 sg13g2_fill_1 FILLER_19_61 ();
 sg13g2_fill_2 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_76 ();
 sg13g2_decap_8 FILLER_19_83 ();
 sg13g2_decap_8 FILLER_19_90 ();
 sg13g2_decap_8 FILLER_19_97 ();
 sg13g2_decap_8 FILLER_19_104 ();
 sg13g2_decap_8 FILLER_19_111 ();
 sg13g2_decap_8 FILLER_19_118 ();
 sg13g2_decap_4 FILLER_19_125 ();
 sg13g2_fill_2 FILLER_19_129 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_200 ();
 sg13g2_fill_2 FILLER_19_207 ();
 sg13g2_fill_1 FILLER_19_209 ();
 sg13g2_decap_4 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_297 ();
 sg13g2_decap_8 FILLER_19_304 ();
 sg13g2_decap_8 FILLER_19_311 ();
 sg13g2_fill_2 FILLER_19_318 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_390 ();
 sg13g2_decap_8 FILLER_19_397 ();
 sg13g2_fill_2 FILLER_19_404 ();
 sg13g2_fill_1 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_2 FILLER_19_429 ();
 sg13g2_fill_1 FILLER_19_431 ();
 sg13g2_decap_8 FILLER_19_452 ();
 sg13g2_decap_4 FILLER_19_459 ();
 sg13g2_decap_8 FILLER_19_489 ();
 sg13g2_decap_4 FILLER_19_496 ();
 sg13g2_fill_1 FILLER_19_500 ();
 sg13g2_fill_2 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_535 ();
 sg13g2_decap_8 FILLER_19_542 ();
 sg13g2_fill_2 FILLER_19_549 ();
 sg13g2_fill_1 FILLER_19_551 ();
 sg13g2_decap_8 FILLER_19_556 ();
 sg13g2_fill_2 FILLER_19_563 ();
 sg13g2_fill_2 FILLER_19_572 ();
 sg13g2_fill_1 FILLER_19_591 ();
 sg13g2_fill_1 FILLER_19_612 ();
 sg13g2_fill_2 FILLER_19_622 ();
 sg13g2_fill_1 FILLER_19_624 ();
 sg13g2_fill_1 FILLER_19_630 ();
 sg13g2_fill_1 FILLER_19_643 ();
 sg13g2_decap_8 FILLER_19_656 ();
 sg13g2_decap_4 FILLER_19_663 ();
 sg13g2_fill_1 FILLER_19_667 ();
 sg13g2_fill_1 FILLER_19_675 ();
 sg13g2_fill_1 FILLER_19_681 ();
 sg13g2_decap_4 FILLER_19_690 ();
 sg13g2_fill_1 FILLER_19_705 ();
 sg13g2_fill_1 FILLER_19_710 ();
 sg13g2_decap_8 FILLER_19_725 ();
 sg13g2_decap_4 FILLER_19_736 ();
 sg13g2_fill_2 FILLER_19_740 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_fill_2 FILLER_19_826 ();
 sg13g2_fill_1 FILLER_19_828 ();
 sg13g2_decap_8 FILLER_19_832 ();
 sg13g2_decap_4 FILLER_19_839 ();
 sg13g2_fill_2 FILLER_19_868 ();
 sg13g2_fill_1 FILLER_19_896 ();
 sg13g2_fill_1 FILLER_19_955 ();
 sg13g2_fill_1 FILLER_19_966 ();
 sg13g2_fill_1 FILLER_19_974 ();
 sg13g2_fill_1 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_999 ();
 sg13g2_decap_4 FILLER_19_1010 ();
 sg13g2_fill_1 FILLER_19_1014 ();
 sg13g2_decap_8 FILLER_19_1049 ();
 sg13g2_fill_1 FILLER_19_1060 ();
 sg13g2_decap_4 FILLER_19_1065 ();
 sg13g2_fill_1 FILLER_19_1069 ();
 sg13g2_fill_1 FILLER_19_1105 ();
 sg13g2_fill_2 FILLER_19_1116 ();
 sg13g2_fill_1 FILLER_19_1118 ();
 sg13g2_fill_2 FILLER_19_1127 ();
 sg13g2_fill_1 FILLER_19_1129 ();
 sg13g2_fill_2 FILLER_19_1156 ();
 sg13g2_fill_1 FILLER_19_1158 ();
 sg13g2_fill_1 FILLER_19_1163 ();
 sg13g2_fill_1 FILLER_19_1299 ();
 sg13g2_decap_8 FILLER_19_1331 ();
 sg13g2_decap_4 FILLER_19_1338 ();
 sg13g2_fill_1 FILLER_19_1342 ();
 sg13g2_decap_8 FILLER_19_1405 ();
 sg13g2_decap_4 FILLER_19_1412 ();
 sg13g2_fill_2 FILLER_19_1416 ();
 sg13g2_decap_4 FILLER_19_1487 ();
 sg13g2_decap_4 FILLER_19_1510 ();
 sg13g2_fill_1 FILLER_19_1514 ();
 sg13g2_fill_2 FILLER_19_1541 ();
 sg13g2_decap_4 FILLER_19_1554 ();
 sg13g2_fill_1 FILLER_19_1558 ();
 sg13g2_decap_8 FILLER_19_1575 ();
 sg13g2_fill_1 FILLER_19_1582 ();
 sg13g2_fill_2 FILLER_19_1664 ();
 sg13g2_fill_2 FILLER_19_1746 ();
 sg13g2_fill_2 FILLER_19_1769 ();
 sg13g2_fill_2 FILLER_19_1824 ();
 sg13g2_fill_1 FILLER_19_1826 ();
 sg13g2_fill_1 FILLER_19_1837 ();
 sg13g2_fill_2 FILLER_19_1842 ();
 sg13g2_decap_8 FILLER_19_1912 ();
 sg13g2_decap_4 FILLER_19_1919 ();
 sg13g2_fill_1 FILLER_19_1927 ();
 sg13g2_fill_1 FILLER_19_1953 ();
 sg13g2_fill_2 FILLER_19_1959 ();
 sg13g2_fill_1 FILLER_19_1965 ();
 sg13g2_fill_2 FILLER_19_1977 ();
 sg13g2_fill_1 FILLER_19_1979 ();
 sg13g2_decap_8 FILLER_19_1999 ();
 sg13g2_decap_4 FILLER_19_2006 ();
 sg13g2_fill_1 FILLER_19_2010 ();
 sg13g2_fill_2 FILLER_19_2026 ();
 sg13g2_decap_8 FILLER_19_2038 ();
 sg13g2_decap_8 FILLER_19_2045 ();
 sg13g2_decap_8 FILLER_19_2052 ();
 sg13g2_decap_4 FILLER_19_2059 ();
 sg13g2_fill_2 FILLER_19_2063 ();
 sg13g2_fill_1 FILLER_19_2183 ();
 sg13g2_decap_8 FILLER_19_2221 ();
 sg13g2_decap_8 FILLER_19_2234 ();
 sg13g2_fill_1 FILLER_19_2241 ();
 sg13g2_fill_2 FILLER_19_2289 ();
 sg13g2_fill_2 FILLER_19_2295 ();
 sg13g2_decap_8 FILLER_19_2307 ();
 sg13g2_decap_8 FILLER_19_2314 ();
 sg13g2_decap_4 FILLER_19_2321 ();
 sg13g2_fill_2 FILLER_19_2325 ();
 sg13g2_fill_2 FILLER_19_2331 ();
 sg13g2_fill_1 FILLER_19_2333 ();
 sg13g2_fill_2 FILLER_19_2342 ();
 sg13g2_fill_2 FILLER_19_2348 ();
 sg13g2_fill_1 FILLER_19_2350 ();
 sg13g2_fill_1 FILLER_19_2355 ();
 sg13g2_fill_2 FILLER_19_2360 ();
 sg13g2_fill_1 FILLER_19_2362 ();
 sg13g2_decap_8 FILLER_19_2367 ();
 sg13g2_decap_4 FILLER_19_2374 ();
 sg13g2_fill_1 FILLER_19_2378 ();
 sg13g2_decap_8 FILLER_19_2382 ();
 sg13g2_decap_8 FILLER_19_2389 ();
 sg13g2_fill_1 FILLER_19_2396 ();
 sg13g2_decap_8 FILLER_19_2427 ();
 sg13g2_decap_8 FILLER_19_2434 ();
 sg13g2_decap_8 FILLER_19_2441 ();
 sg13g2_decap_8 FILLER_19_2448 ();
 sg13g2_fill_2 FILLER_19_2455 ();
 sg13g2_decap_8 FILLER_19_2478 ();
 sg13g2_decap_8 FILLER_19_2485 ();
 sg13g2_decap_8 FILLER_19_2492 ();
 sg13g2_fill_2 FILLER_19_2556 ();
 sg13g2_fill_1 FILLER_19_2558 ();
 sg13g2_fill_1 FILLER_19_2598 ();
 sg13g2_decap_8 FILLER_19_2629 ();
 sg13g2_decap_8 FILLER_19_2636 ();
 sg13g2_decap_8 FILLER_19_2643 ();
 sg13g2_decap_8 FILLER_19_2650 ();
 sg13g2_decap_8 FILLER_19_2657 ();
 sg13g2_decap_4 FILLER_19_2664 ();
 sg13g2_fill_2 FILLER_19_2668 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_fill_1 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_19 ();
 sg13g2_fill_1 FILLER_20_26 ();
 sg13g2_decap_4 FILLER_20_31 ();
 sg13g2_fill_2 FILLER_20_39 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_48 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_4 FILLER_20_137 ();
 sg13g2_fill_1 FILLER_20_141 ();
 sg13g2_decap_4 FILLER_20_147 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_decap_8 FILLER_20_161 ();
 sg13g2_decap_8 FILLER_20_168 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_decap_4 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_decap_8 FILLER_20_196 ();
 sg13g2_decap_8 FILLER_20_203 ();
 sg13g2_decap_4 FILLER_20_210 ();
 sg13g2_fill_1 FILLER_20_214 ();
 sg13g2_fill_2 FILLER_20_219 ();
 sg13g2_fill_1 FILLER_20_221 ();
 sg13g2_decap_4 FILLER_20_230 ();
 sg13g2_fill_1 FILLER_20_234 ();
 sg13g2_decap_8 FILLER_20_240 ();
 sg13g2_decap_8 FILLER_20_247 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_268 ();
 sg13g2_decap_8 FILLER_20_275 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_decap_8 FILLER_20_296 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_332 ();
 sg13g2_fill_1 FILLER_20_360 ();
 sg13g2_fill_2 FILLER_20_416 ();
 sg13g2_fill_2 FILLER_20_428 ();
 sg13g2_decap_8 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_fill_2 FILLER_20_459 ();
 sg13g2_fill_1 FILLER_20_461 ();
 sg13g2_decap_4 FILLER_20_466 ();
 sg13g2_fill_2 FILLER_20_470 ();
 sg13g2_decap_8 FILLER_20_476 ();
 sg13g2_fill_2 FILLER_20_483 ();
 sg13g2_fill_2 FILLER_20_490 ();
 sg13g2_fill_1 FILLER_20_492 ();
 sg13g2_decap_8 FILLER_20_502 ();
 sg13g2_decap_8 FILLER_20_509 ();
 sg13g2_decap_8 FILLER_20_530 ();
 sg13g2_decap_8 FILLER_20_537 ();
 sg13g2_fill_2 FILLER_20_570 ();
 sg13g2_fill_1 FILLER_20_572 ();
 sg13g2_fill_2 FILLER_20_583 ();
 sg13g2_fill_1 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_591 ();
 sg13g2_decap_4 FILLER_20_598 ();
 sg13g2_fill_2 FILLER_20_602 ();
 sg13g2_fill_2 FILLER_20_608 ();
 sg13g2_fill_1 FILLER_20_610 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_4 FILLER_20_627 ();
 sg13g2_decap_4 FILLER_20_655 ();
 sg13g2_fill_1 FILLER_20_659 ();
 sg13g2_decap_8 FILLER_20_663 ();
 sg13g2_decap_8 FILLER_20_675 ();
 sg13g2_decap_8 FILLER_20_687 ();
 sg13g2_fill_2 FILLER_20_694 ();
 sg13g2_fill_1 FILLER_20_696 ();
 sg13g2_decap_8 FILLER_20_700 ();
 sg13g2_decap_8 FILLER_20_707 ();
 sg13g2_decap_4 FILLER_20_714 ();
 sg13g2_fill_1 FILLER_20_718 ();
 sg13g2_fill_1 FILLER_20_724 ();
 sg13g2_decap_8 FILLER_20_730 ();
 sg13g2_decap_8 FILLER_20_737 ();
 sg13g2_fill_2 FILLER_20_744 ();
 sg13g2_fill_1 FILLER_20_746 ();
 sg13g2_decap_4 FILLER_20_752 ();
 sg13g2_fill_1 FILLER_20_756 ();
 sg13g2_fill_1 FILLER_20_767 ();
 sg13g2_fill_2 FILLER_20_784 ();
 sg13g2_fill_2 FILLER_20_800 ();
 sg13g2_fill_1 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_839 ();
 sg13g2_fill_2 FILLER_20_846 ();
 sg13g2_fill_2 FILLER_20_872 ();
 sg13g2_decap_4 FILLER_20_946 ();
 sg13g2_fill_2 FILLER_20_950 ();
 sg13g2_fill_1 FILLER_20_960 ();
 sg13g2_decap_4 FILLER_20_966 ();
 sg13g2_fill_2 FILLER_20_999 ();
 sg13g2_fill_2 FILLER_20_1006 ();
 sg13g2_decap_4 FILLER_20_1012 ();
 sg13g2_fill_1 FILLER_20_1021 ();
 sg13g2_fill_1 FILLER_20_1026 ();
 sg13g2_decap_8 FILLER_20_1035 ();
 sg13g2_decap_8 FILLER_20_1051 ();
 sg13g2_fill_2 FILLER_20_1058 ();
 sg13g2_fill_1 FILLER_20_1060 ();
 sg13g2_fill_2 FILLER_20_1101 ();
 sg13g2_decap_8 FILLER_20_1132 ();
 sg13g2_fill_2 FILLER_20_1139 ();
 sg13g2_decap_8 FILLER_20_1144 ();
 sg13g2_decap_8 FILLER_20_1151 ();
 sg13g2_fill_2 FILLER_20_1158 ();
 sg13g2_fill_1 FILLER_20_1160 ();
 sg13g2_decap_8 FILLER_20_1200 ();
 sg13g2_fill_1 FILLER_20_1207 ();
 sg13g2_decap_4 FILLER_20_1212 ();
 sg13g2_decap_4 FILLER_20_1221 ();
 sg13g2_fill_2 FILLER_20_1251 ();
 sg13g2_fill_1 FILLER_20_1253 ();
 sg13g2_fill_2 FILLER_20_1272 ();
 sg13g2_fill_1 FILLER_20_1274 ();
 sg13g2_fill_1 FILLER_20_1286 ();
 sg13g2_decap_4 FILLER_20_1294 ();
 sg13g2_fill_1 FILLER_20_1298 ();
 sg13g2_decap_8 FILLER_20_1303 ();
 sg13g2_decap_8 FILLER_20_1336 ();
 sg13g2_decap_8 FILLER_20_1343 ();
 sg13g2_fill_1 FILLER_20_1350 ();
 sg13g2_fill_2 FILLER_20_1361 ();
 sg13g2_decap_8 FILLER_20_1408 ();
 sg13g2_decap_8 FILLER_20_1415 ();
 sg13g2_fill_2 FILLER_20_1422 ();
 sg13g2_decap_4 FILLER_20_1458 ();
 sg13g2_fill_1 FILLER_20_1462 ();
 sg13g2_fill_2 FILLER_20_1468 ();
 sg13g2_fill_1 FILLER_20_1470 ();
 sg13g2_fill_2 FILLER_20_1487 ();
 sg13g2_fill_1 FILLER_20_1495 ();
 sg13g2_decap_8 FILLER_20_1515 ();
 sg13g2_fill_2 FILLER_20_1522 ();
 sg13g2_fill_1 FILLER_20_1545 ();
 sg13g2_fill_2 FILLER_20_1554 ();
 sg13g2_fill_1 FILLER_20_1556 ();
 sg13g2_fill_2 FILLER_20_1582 ();
 sg13g2_decap_8 FILLER_20_1614 ();
 sg13g2_fill_1 FILLER_20_1621 ();
 sg13g2_fill_2 FILLER_20_1630 ();
 sg13g2_fill_2 FILLER_20_1648 ();
 sg13g2_fill_1 FILLER_20_1658 ();
 sg13g2_fill_1 FILLER_20_1694 ();
 sg13g2_fill_1 FILLER_20_1720 ();
 sg13g2_fill_1 FILLER_20_1732 ();
 sg13g2_fill_2 FILLER_20_1803 ();
 sg13g2_decap_8 FILLER_20_1809 ();
 sg13g2_fill_1 FILLER_20_1816 ();
 sg13g2_fill_2 FILLER_20_1826 ();
 sg13g2_decap_8 FILLER_20_1834 ();
 sg13g2_decap_4 FILLER_20_1841 ();
 sg13g2_fill_1 FILLER_20_1845 ();
 sg13g2_fill_2 FILLER_20_1862 ();
 sg13g2_decap_8 FILLER_20_1900 ();
 sg13g2_decap_8 FILLER_20_1907 ();
 sg13g2_fill_2 FILLER_20_1914 ();
 sg13g2_fill_1 FILLER_20_1942 ();
 sg13g2_decap_8 FILLER_20_1972 ();
 sg13g2_decap_8 FILLER_20_1979 ();
 sg13g2_decap_8 FILLER_20_1986 ();
 sg13g2_decap_8 FILLER_20_1993 ();
 sg13g2_decap_8 FILLER_20_2000 ();
 sg13g2_fill_2 FILLER_20_2012 ();
 sg13g2_fill_1 FILLER_20_2022 ();
 sg13g2_decap_8 FILLER_20_2028 ();
 sg13g2_fill_1 FILLER_20_2035 ();
 sg13g2_fill_1 FILLER_20_2040 ();
 sg13g2_fill_2 FILLER_20_2045 ();
 sg13g2_fill_2 FILLER_20_2051 ();
 sg13g2_decap_8 FILLER_20_2058 ();
 sg13g2_decap_8 FILLER_20_2065 ();
 sg13g2_decap_8 FILLER_20_2072 ();
 sg13g2_decap_4 FILLER_20_2079 ();
 sg13g2_fill_2 FILLER_20_2175 ();
 sg13g2_fill_2 FILLER_20_2193 ();
 sg13g2_fill_2 FILLER_20_2285 ();
 sg13g2_fill_1 FILLER_20_2287 ();
 sg13g2_fill_2 FILLER_20_2296 ();
 sg13g2_fill_2 FILLER_20_2303 ();
 sg13g2_fill_1 FILLER_20_2305 ();
 sg13g2_fill_1 FILLER_20_2348 ();
 sg13g2_fill_2 FILLER_20_2375 ();
 sg13g2_fill_1 FILLER_20_2377 ();
 sg13g2_decap_8 FILLER_20_2382 ();
 sg13g2_decap_8 FILLER_20_2389 ();
 sg13g2_decap_8 FILLER_20_2435 ();
 sg13g2_fill_2 FILLER_20_2442 ();
 sg13g2_fill_1 FILLER_20_2444 ();
 sg13g2_fill_2 FILLER_20_2546 ();
 sg13g2_decap_4 FILLER_20_2552 ();
 sg13g2_fill_1 FILLER_20_2556 ();
 sg13g2_decap_4 FILLER_20_2562 ();
 sg13g2_fill_1 FILLER_20_2566 ();
 sg13g2_fill_2 FILLER_20_2571 ();
 sg13g2_fill_1 FILLER_20_2599 ();
 sg13g2_fill_2 FILLER_20_2614 ();
 sg13g2_fill_1 FILLER_20_2616 ();
 sg13g2_fill_2 FILLER_20_2621 ();
 sg13g2_fill_1 FILLER_20_2623 ();
 sg13g2_decap_8 FILLER_20_2628 ();
 sg13g2_decap_8 FILLER_20_2635 ();
 sg13g2_decap_8 FILLER_20_2642 ();
 sg13g2_decap_8 FILLER_20_2649 ();
 sg13g2_decap_8 FILLER_20_2656 ();
 sg13g2_decap_8 FILLER_20_2663 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_47 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_decap_8 FILLER_21_95 ();
 sg13g2_decap_8 FILLER_21_102 ();
 sg13g2_decap_8 FILLER_21_109 ();
 sg13g2_decap_8 FILLER_21_116 ();
 sg13g2_decap_8 FILLER_21_123 ();
 sg13g2_decap_8 FILLER_21_130 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_decap_8 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_8 FILLER_21_158 ();
 sg13g2_decap_8 FILLER_21_165 ();
 sg13g2_decap_8 FILLER_21_172 ();
 sg13g2_decap_8 FILLER_21_179 ();
 sg13g2_decap_8 FILLER_21_186 ();
 sg13g2_decap_8 FILLER_21_193 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_decap_8 FILLER_21_207 ();
 sg13g2_decap_8 FILLER_21_214 ();
 sg13g2_decap_8 FILLER_21_221 ();
 sg13g2_decap_8 FILLER_21_228 ();
 sg13g2_decap_8 FILLER_21_235 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_fill_1 FILLER_21_294 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_342 ();
 sg13g2_decap_8 FILLER_21_349 ();
 sg13g2_fill_2 FILLER_21_356 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_4 FILLER_21_415 ();
 sg13g2_fill_1 FILLER_21_440 ();
 sg13g2_fill_2 FILLER_21_446 ();
 sg13g2_fill_1 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_458 ();
 sg13g2_decap_8 FILLER_21_465 ();
 sg13g2_fill_2 FILLER_21_472 ();
 sg13g2_fill_1 FILLER_21_474 ();
 sg13g2_decap_8 FILLER_21_479 ();
 sg13g2_decap_8 FILLER_21_486 ();
 sg13g2_decap_8 FILLER_21_493 ();
 sg13g2_fill_1 FILLER_21_500 ();
 sg13g2_decap_8 FILLER_21_530 ();
 sg13g2_fill_2 FILLER_21_537 ();
 sg13g2_fill_1 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_545 ();
 sg13g2_decap_8 FILLER_21_556 ();
 sg13g2_fill_1 FILLER_21_563 ();
 sg13g2_fill_1 FILLER_21_569 ();
 sg13g2_decap_4 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_583 ();
 sg13g2_fill_1 FILLER_21_590 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_613 ();
 sg13g2_decap_8 FILLER_21_620 ();
 sg13g2_decap_8 FILLER_21_627 ();
 sg13g2_decap_8 FILLER_21_634 ();
 sg13g2_fill_2 FILLER_21_641 ();
 sg13g2_fill_1 FILLER_21_643 ();
 sg13g2_decap_8 FILLER_21_655 ();
 sg13g2_fill_2 FILLER_21_662 ();
 sg13g2_fill_1 FILLER_21_670 ();
 sg13g2_fill_1 FILLER_21_676 ();
 sg13g2_decap_4 FILLER_21_694 ();
 sg13g2_fill_1 FILLER_21_704 ();
 sg13g2_decap_8 FILLER_21_711 ();
 sg13g2_decap_8 FILLER_21_718 ();
 sg13g2_decap_8 FILLER_21_725 ();
 sg13g2_decap_8 FILLER_21_732 ();
 sg13g2_decap_4 FILLER_21_739 ();
 sg13g2_fill_2 FILLER_21_743 ();
 sg13g2_fill_2 FILLER_21_760 ();
 sg13g2_fill_2 FILLER_21_771 ();
 sg13g2_decap_8 FILLER_21_789 ();
 sg13g2_decap_8 FILLER_21_796 ();
 sg13g2_decap_4 FILLER_21_803 ();
 sg13g2_decap_8 FILLER_21_820 ();
 sg13g2_fill_1 FILLER_21_827 ();
 sg13g2_fill_1 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_4 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_884 ();
 sg13g2_fill_2 FILLER_21_891 ();
 sg13g2_fill_1 FILLER_21_893 ();
 sg13g2_fill_2 FILLER_21_921 ();
 sg13g2_fill_1 FILLER_21_933 ();
 sg13g2_decap_4 FILLER_21_938 ();
 sg13g2_decap_8 FILLER_21_946 ();
 sg13g2_decap_8 FILLER_21_953 ();
 sg13g2_decap_8 FILLER_21_960 ();
 sg13g2_fill_1 FILLER_21_980 ();
 sg13g2_fill_1 FILLER_21_984 ();
 sg13g2_fill_2 FILLER_21_990 ();
 sg13g2_fill_1 FILLER_21_992 ();
 sg13g2_decap_8 FILLER_21_998 ();
 sg13g2_decap_8 FILLER_21_1005 ();
 sg13g2_fill_2 FILLER_21_1021 ();
 sg13g2_fill_1 FILLER_21_1023 ();
 sg13g2_fill_1 FILLER_21_1033 ();
 sg13g2_decap_4 FILLER_21_1038 ();
 sg13g2_fill_2 FILLER_21_1112 ();
 sg13g2_fill_1 FILLER_21_1122 ();
 sg13g2_fill_2 FILLER_21_1127 ();
 sg13g2_decap_8 FILLER_21_1134 ();
 sg13g2_fill_2 FILLER_21_1150 ();
 sg13g2_fill_1 FILLER_21_1152 ();
 sg13g2_decap_8 FILLER_21_1159 ();
 sg13g2_decap_8 FILLER_21_1166 ();
 sg13g2_decap_8 FILLER_21_1173 ();
 sg13g2_decap_8 FILLER_21_1189 ();
 sg13g2_decap_8 FILLER_21_1196 ();
 sg13g2_decap_8 FILLER_21_1203 ();
 sg13g2_decap_4 FILLER_21_1215 ();
 sg13g2_fill_2 FILLER_21_1219 ();
 sg13g2_decap_8 FILLER_21_1225 ();
 sg13g2_decap_8 FILLER_21_1232 ();
 sg13g2_decap_8 FILLER_21_1239 ();
 sg13g2_decap_4 FILLER_21_1246 ();
 sg13g2_fill_1 FILLER_21_1250 ();
 sg13g2_decap_4 FILLER_21_1260 ();
 sg13g2_fill_1 FILLER_21_1264 ();
 sg13g2_decap_4 FILLER_21_1273 ();
 sg13g2_fill_1 FILLER_21_1277 ();
 sg13g2_decap_8 FILLER_21_1295 ();
 sg13g2_decap_8 FILLER_21_1302 ();
 sg13g2_decap_8 FILLER_21_1309 ();
 sg13g2_decap_8 FILLER_21_1356 ();
 sg13g2_decap_8 FILLER_21_1363 ();
 sg13g2_decap_8 FILLER_21_1370 ();
 sg13g2_decap_8 FILLER_21_1377 ();
 sg13g2_decap_4 FILLER_21_1384 ();
 sg13g2_fill_1 FILLER_21_1388 ();
 sg13g2_decap_8 FILLER_21_1398 ();
 sg13g2_decap_8 FILLER_21_1405 ();
 sg13g2_decap_8 FILLER_21_1412 ();
 sg13g2_fill_2 FILLER_21_1419 ();
 sg13g2_decap_8 FILLER_21_1463 ();
 sg13g2_decap_8 FILLER_21_1470 ();
 sg13g2_decap_8 FILLER_21_1477 ();
 sg13g2_fill_2 FILLER_21_1484 ();
 sg13g2_fill_2 FILLER_21_1496 ();
 sg13g2_fill_1 FILLER_21_1498 ();
 sg13g2_decap_4 FILLER_21_1519 ();
 sg13g2_fill_1 FILLER_21_1523 ();
 sg13g2_decap_8 FILLER_21_1560 ();
 sg13g2_decap_8 FILLER_21_1567 ();
 sg13g2_fill_2 FILLER_21_1574 ();
 sg13g2_fill_1 FILLER_21_1576 ();
 sg13g2_decap_8 FILLER_21_1583 ();
 sg13g2_decap_8 FILLER_21_1590 ();
 sg13g2_decap_8 FILLER_21_1597 ();
 sg13g2_decap_8 FILLER_21_1604 ();
 sg13g2_decap_4 FILLER_21_1611 ();
 sg13g2_fill_1 FILLER_21_1634 ();
 sg13g2_fill_1 FILLER_21_1638 ();
 sg13g2_fill_1 FILLER_21_1712 ();
 sg13g2_fill_1 FILLER_21_1761 ();
 sg13g2_decap_8 FILLER_21_1782 ();
 sg13g2_decap_8 FILLER_21_1789 ();
 sg13g2_decap_8 FILLER_21_1796 ();
 sg13g2_decap_8 FILLER_21_1803 ();
 sg13g2_decap_8 FILLER_21_1810 ();
 sg13g2_decap_8 FILLER_21_1817 ();
 sg13g2_decap_8 FILLER_21_1824 ();
 sg13g2_fill_2 FILLER_21_1831 ();
 sg13g2_fill_1 FILLER_21_1833 ();
 sg13g2_fill_2 FILLER_21_1893 ();
 sg13g2_fill_1 FILLER_21_1911 ();
 sg13g2_decap_8 FILLER_21_1916 ();
 sg13g2_decap_8 FILLER_21_1923 ();
 sg13g2_fill_1 FILLER_21_1930 ();
 sg13g2_fill_2 FILLER_21_1940 ();
 sg13g2_fill_1 FILLER_21_1946 ();
 sg13g2_decap_8 FILLER_21_1956 ();
 sg13g2_decap_8 FILLER_21_1967 ();
 sg13g2_decap_4 FILLER_21_1974 ();
 sg13g2_fill_1 FILLER_21_1978 ();
 sg13g2_decap_4 FILLER_21_1985 ();
 sg13g2_fill_2 FILLER_21_2091 ();
 sg13g2_fill_1 FILLER_21_2119 ();
 sg13g2_fill_1 FILLER_21_2156 ();
 sg13g2_fill_1 FILLER_21_2200 ();
 sg13g2_fill_1 FILLER_21_2227 ();
 sg13g2_fill_2 FILLER_21_2266 ();
 sg13g2_fill_1 FILLER_21_2268 ();
 sg13g2_fill_2 FILLER_21_2277 ();
 sg13g2_decap_4 FILLER_21_2310 ();
 sg13g2_fill_2 FILLER_21_2314 ();
 sg13g2_decap_8 FILLER_21_2320 ();
 sg13g2_decap_8 FILLER_21_2327 ();
 sg13g2_fill_1 FILLER_21_2334 ();
 sg13g2_fill_2 FILLER_21_2350 ();
 sg13g2_fill_1 FILLER_21_2352 ();
 sg13g2_fill_1 FILLER_21_2409 ();
 sg13g2_fill_1 FILLER_21_2414 ();
 sg13g2_fill_2 FILLER_21_2484 ();
 sg13g2_decap_8 FILLER_21_2490 ();
 sg13g2_decap_8 FILLER_21_2497 ();
 sg13g2_decap_4 FILLER_21_2504 ();
 sg13g2_fill_1 FILLER_21_2508 ();
 sg13g2_fill_2 FILLER_21_2513 ();
 sg13g2_fill_1 FILLER_21_2515 ();
 sg13g2_decap_8 FILLER_21_2520 ();
 sg13g2_decap_8 FILLER_21_2527 ();
 sg13g2_decap_8 FILLER_21_2534 ();
 sg13g2_decap_8 FILLER_21_2541 ();
 sg13g2_fill_1 FILLER_21_2558 ();
 sg13g2_decap_8 FILLER_21_2593 ();
 sg13g2_decap_8 FILLER_21_2600 ();
 sg13g2_decap_8 FILLER_21_2607 ();
 sg13g2_decap_8 FILLER_21_2614 ();
 sg13g2_decap_8 FILLER_21_2621 ();
 sg13g2_decap_4 FILLER_21_2628 ();
 sg13g2_fill_2 FILLER_21_2632 ();
 sg13g2_fill_2 FILLER_21_2668 ();
 sg13g2_fill_2 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_48 ();
 sg13g2_fill_1 FILLER_22_50 ();
 sg13g2_fill_2 FILLER_22_62 ();
 sg13g2_fill_1 FILLER_22_64 ();
 sg13g2_decap_4 FILLER_22_69 ();
 sg13g2_fill_1 FILLER_22_73 ();
 sg13g2_fill_2 FILLER_22_82 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_4 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_113 ();
 sg13g2_fill_1 FILLER_22_148 ();
 sg13g2_decap_8 FILLER_22_159 ();
 sg13g2_decap_8 FILLER_22_166 ();
 sg13g2_decap_8 FILLER_22_173 ();
 sg13g2_decap_8 FILLER_22_180 ();
 sg13g2_decap_8 FILLER_22_187 ();
 sg13g2_decap_8 FILLER_22_194 ();
 sg13g2_decap_8 FILLER_22_201 ();
 sg13g2_decap_4 FILLER_22_208 ();
 sg13g2_fill_1 FILLER_22_212 ();
 sg13g2_fill_2 FILLER_22_216 ();
 sg13g2_fill_2 FILLER_22_230 ();
 sg13g2_decap_8 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_262 ();
 sg13g2_decap_8 FILLER_22_269 ();
 sg13g2_decap_8 FILLER_22_276 ();
 sg13g2_fill_2 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_285 ();
 sg13g2_fill_1 FILLER_22_312 ();
 sg13g2_decap_4 FILLER_22_318 ();
 sg13g2_fill_2 FILLER_22_322 ();
 sg13g2_decap_8 FILLER_22_350 ();
 sg13g2_fill_2 FILLER_22_357 ();
 sg13g2_fill_1 FILLER_22_359 ();
 sg13g2_fill_1 FILLER_22_384 ();
 sg13g2_fill_2 FILLER_22_390 ();
 sg13g2_fill_1 FILLER_22_392 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_4 FILLER_22_417 ();
 sg13g2_fill_2 FILLER_22_421 ();
 sg13g2_fill_1 FILLER_22_428 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_4 FILLER_22_445 ();
 sg13g2_fill_1 FILLER_22_449 ();
 sg13g2_decap_8 FILLER_22_455 ();
 sg13g2_decap_8 FILLER_22_462 ();
 sg13g2_decap_8 FILLER_22_469 ();
 sg13g2_decap_8 FILLER_22_476 ();
 sg13g2_decap_4 FILLER_22_513 ();
 sg13g2_fill_1 FILLER_22_517 ();
 sg13g2_decap_8 FILLER_22_544 ();
 sg13g2_decap_8 FILLER_22_551 ();
 sg13g2_fill_1 FILLER_22_558 ();
 sg13g2_decap_8 FILLER_22_563 ();
 sg13g2_fill_2 FILLER_22_582 ();
 sg13g2_fill_1 FILLER_22_584 ();
 sg13g2_decap_8 FILLER_22_611 ();
 sg13g2_decap_4 FILLER_22_652 ();
 sg13g2_fill_2 FILLER_22_665 ();
 sg13g2_fill_1 FILLER_22_670 ();
 sg13g2_fill_1 FILLER_22_676 ();
 sg13g2_fill_1 FILLER_22_681 ();
 sg13g2_fill_1 FILLER_22_704 ();
 sg13g2_fill_1 FILLER_22_791 ();
 sg13g2_fill_2 FILLER_22_841 ();
 sg13g2_fill_1 FILLER_22_843 ();
 sg13g2_fill_2 FILLER_22_858 ();
 sg13g2_fill_2 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_896 ();
 sg13g2_fill_2 FILLER_22_903 ();
 sg13g2_fill_1 FILLER_22_934 ();
 sg13g2_fill_1 FILLER_22_961 ();
 sg13g2_decap_4 FILLER_22_967 ();
 sg13g2_fill_1 FILLER_22_971 ();
 sg13g2_fill_2 FILLER_22_986 ();
 sg13g2_decap_4 FILLER_22_993 ();
 sg13g2_fill_2 FILLER_22_1010 ();
 sg13g2_fill_1 FILLER_22_1023 ();
 sg13g2_fill_2 FILLER_22_1033 ();
 sg13g2_fill_1 FILLER_22_1035 ();
 sg13g2_fill_1 FILLER_22_1041 ();
 sg13g2_decap_8 FILLER_22_1047 ();
 sg13g2_fill_2 FILLER_22_1054 ();
 sg13g2_fill_2 FILLER_22_1061 ();
 sg13g2_fill_1 FILLER_22_1063 ();
 sg13g2_fill_1 FILLER_22_1083 ();
 sg13g2_fill_1 FILLER_22_1090 ();
 sg13g2_fill_1 FILLER_22_1094 ();
 sg13g2_decap_4 FILLER_22_1099 ();
 sg13g2_fill_2 FILLER_22_1103 ();
 sg13g2_decap_8 FILLER_22_1114 ();
 sg13g2_decap_8 FILLER_22_1121 ();
 sg13g2_decap_8 FILLER_22_1128 ();
 sg13g2_decap_8 FILLER_22_1171 ();
 sg13g2_decap_8 FILLER_22_1184 ();
 sg13g2_decap_8 FILLER_22_1191 ();
 sg13g2_fill_1 FILLER_22_1198 ();
 sg13g2_decap_4 FILLER_22_1202 ();
 sg13g2_decap_4 FILLER_22_1232 ();
 sg13g2_fill_1 FILLER_22_1236 ();
 sg13g2_decap_4 FILLER_22_1241 ();
 sg13g2_fill_2 FILLER_22_1245 ();
 sg13g2_fill_1 FILLER_22_1278 ();
 sg13g2_decap_4 FILLER_22_1283 ();
 sg13g2_fill_2 FILLER_22_1295 ();
 sg13g2_decap_8 FILLER_22_1306 ();
 sg13g2_decap_4 FILLER_22_1313 ();
 sg13g2_decap_8 FILLER_22_1325 ();
 sg13g2_decap_4 FILLER_22_1332 ();
 sg13g2_fill_2 FILLER_22_1348 ();
 sg13g2_fill_1 FILLER_22_1350 ();
 sg13g2_decap_8 FILLER_22_1355 ();
 sg13g2_fill_1 FILLER_22_1362 ();
 sg13g2_decap_8 FILLER_22_1394 ();
 sg13g2_decap_8 FILLER_22_1401 ();
 sg13g2_decap_4 FILLER_22_1408 ();
 sg13g2_fill_2 FILLER_22_1412 ();
 sg13g2_decap_4 FILLER_22_1433 ();
 sg13g2_fill_1 FILLER_22_1437 ();
 sg13g2_fill_2 FILLER_22_1526 ();
 sg13g2_fill_2 FILLER_22_1590 ();
 sg13g2_fill_1 FILLER_22_1592 ();
 sg13g2_fill_2 FILLER_22_1598 ();
 sg13g2_fill_1 FILLER_22_1600 ();
 sg13g2_fill_2 FILLER_22_1605 ();
 sg13g2_decap_4 FILLER_22_1612 ();
 sg13g2_fill_2 FILLER_22_1616 ();
 sg13g2_fill_1 FILLER_22_1695 ();
 sg13g2_fill_1 FILLER_22_1718 ();
 sg13g2_fill_2 FILLER_22_1771 ();
 sg13g2_decap_8 FILLER_22_1799 ();
 sg13g2_decap_8 FILLER_22_1806 ();
 sg13g2_decap_4 FILLER_22_1813 ();
 sg13g2_fill_2 FILLER_22_1817 ();
 sg13g2_fill_1 FILLER_22_1823 ();
 sg13g2_fill_2 FILLER_22_1841 ();
 sg13g2_fill_2 FILLER_22_1855 ();
 sg13g2_fill_2 FILLER_22_1863 ();
 sg13g2_fill_1 FILLER_22_1966 ();
 sg13g2_decap_4 FILLER_22_2003 ();
 sg13g2_fill_2 FILLER_22_2025 ();
 sg13g2_fill_2 FILLER_22_2044 ();
 sg13g2_fill_2 FILLER_22_2072 ();
 sg13g2_fill_1 FILLER_22_2074 ();
 sg13g2_decap_8 FILLER_22_2085 ();
 sg13g2_fill_2 FILLER_22_2101 ();
 sg13g2_fill_2 FILLER_22_2109 ();
 sg13g2_fill_1 FILLER_22_2126 ();
 sg13g2_decap_4 FILLER_22_2152 ();
 sg13g2_decap_8 FILLER_22_2159 ();
 sg13g2_decap_4 FILLER_22_2166 ();
 sg13g2_decap_8 FILLER_22_2176 ();
 sg13g2_fill_2 FILLER_22_2183 ();
 sg13g2_fill_1 FILLER_22_2193 ();
 sg13g2_decap_8 FILLER_22_2204 ();
 sg13g2_decap_8 FILLER_22_2211 ();
 sg13g2_decap_4 FILLER_22_2224 ();
 sg13g2_fill_2 FILLER_22_2228 ();
 sg13g2_fill_2 FILLER_22_2236 ();
 sg13g2_fill_1 FILLER_22_2245 ();
 sg13g2_decap_8 FILLER_22_2260 ();
 sg13g2_decap_8 FILLER_22_2267 ();
 sg13g2_decap_4 FILLER_22_2274 ();
 sg13g2_fill_1 FILLER_22_2278 ();
 sg13g2_fill_2 FILLER_22_2300 ();
 sg13g2_fill_2 FILLER_22_2306 ();
 sg13g2_fill_2 FILLER_22_2334 ();
 sg13g2_fill_1 FILLER_22_2336 ();
 sg13g2_fill_2 FILLER_22_2363 ();
 sg13g2_fill_1 FILLER_22_2365 ();
 sg13g2_fill_2 FILLER_22_2372 ();
 sg13g2_decap_8 FILLER_22_2404 ();
 sg13g2_decap_8 FILLER_22_2411 ();
 sg13g2_decap_8 FILLER_22_2418 ();
 sg13g2_decap_8 FILLER_22_2425 ();
 sg13g2_decap_4 FILLER_22_2432 ();
 sg13g2_fill_1 FILLER_22_2436 ();
 sg13g2_fill_2 FILLER_22_2476 ();
 sg13g2_decap_4 FILLER_22_2508 ();
 sg13g2_fill_1 FILLER_22_2512 ();
 sg13g2_decap_8 FILLER_22_2519 ();
 sg13g2_decap_8 FILLER_22_2526 ();
 sg13g2_decap_4 FILLER_22_2533 ();
 sg13g2_fill_2 FILLER_22_2537 ();
 sg13g2_decap_8 FILLER_22_2543 ();
 sg13g2_decap_4 FILLER_22_2550 ();
 sg13g2_fill_2 FILLER_22_2554 ();
 sg13g2_decap_8 FILLER_22_2561 ();
 sg13g2_fill_2 FILLER_22_2568 ();
 sg13g2_decap_4 FILLER_22_2574 ();
 sg13g2_fill_1 FILLER_22_2578 ();
 sg13g2_fill_2 FILLER_22_2583 ();
 sg13g2_fill_1 FILLER_22_2585 ();
 sg13g2_decap_8 FILLER_22_2599 ();
 sg13g2_decap_8 FILLER_22_2606 ();
 sg13g2_decap_8 FILLER_22_2613 ();
 sg13g2_fill_2 FILLER_22_2620 ();
 sg13g2_fill_1 FILLER_22_2622 ();
 sg13g2_decap_4 FILLER_22_2665 ();
 sg13g2_fill_1 FILLER_22_2669 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_fill_1 FILLER_23_32 ();
 sg13g2_fill_1 FILLER_23_39 ();
 sg13g2_decap_4 FILLER_23_58 ();
 sg13g2_fill_2 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_85 ();
 sg13g2_decap_8 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_99 ();
 sg13g2_fill_2 FILLER_23_152 ();
 sg13g2_fill_1 FILLER_23_154 ();
 sg13g2_fill_2 FILLER_23_185 ();
 sg13g2_fill_1 FILLER_23_187 ();
 sg13g2_fill_1 FILLER_23_192 ();
 sg13g2_decap_8 FILLER_23_197 ();
 sg13g2_fill_2 FILLER_23_204 ();
 sg13g2_fill_1 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_268 ();
 sg13g2_decap_8 FILLER_23_275 ();
 sg13g2_decap_8 FILLER_23_282 ();
 sg13g2_decap_4 FILLER_23_289 ();
 sg13g2_fill_2 FILLER_23_293 ();
 sg13g2_fill_1 FILLER_23_316 ();
 sg13g2_decap_8 FILLER_23_327 ();
 sg13g2_decap_8 FILLER_23_334 ();
 sg13g2_decap_4 FILLER_23_341 ();
 sg13g2_fill_2 FILLER_23_376 ();
 sg13g2_decap_8 FILLER_23_393 ();
 sg13g2_fill_2 FILLER_23_400 ();
 sg13g2_fill_1 FILLER_23_402 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_1 FILLER_23_409 ();
 sg13g2_decap_4 FILLER_23_414 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_4 FILLER_23_483 ();
 sg13g2_fill_2 FILLER_23_487 ();
 sg13g2_decap_4 FILLER_23_530 ();
 sg13g2_fill_1 FILLER_23_538 ();
 sg13g2_fill_1 FILLER_23_543 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_4 FILLER_23_574 ();
 sg13g2_fill_2 FILLER_23_578 ();
 sg13g2_decap_8 FILLER_23_590 ();
 sg13g2_decap_8 FILLER_23_597 ();
 sg13g2_fill_1 FILLER_23_604 ();
 sg13g2_decap_4 FILLER_23_641 ();
 sg13g2_fill_2 FILLER_23_649 ();
 sg13g2_fill_1 FILLER_23_651 ();
 sg13g2_fill_1 FILLER_23_695 ();
 sg13g2_fill_1 FILLER_23_755 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_decap_8 FILLER_23_882 ();
 sg13g2_fill_1 FILLER_23_889 ();
 sg13g2_fill_1 FILLER_23_896 ();
 sg13g2_fill_2 FILLER_23_936 ();
 sg13g2_fill_1 FILLER_23_938 ();
 sg13g2_fill_2 FILLER_23_944 ();
 sg13g2_decap_4 FILLER_23_981 ();
 sg13g2_fill_2 FILLER_23_985 ();
 sg13g2_fill_2 FILLER_23_997 ();
 sg13g2_fill_2 FILLER_23_1003 ();
 sg13g2_fill_1 FILLER_23_1005 ();
 sg13g2_fill_2 FILLER_23_1036 ();
 sg13g2_fill_1 FILLER_23_1038 ();
 sg13g2_fill_1 FILLER_23_1047 ();
 sg13g2_fill_2 FILLER_23_1061 ();
 sg13g2_fill_1 FILLER_23_1063 ();
 sg13g2_decap_4 FILLER_23_1069 ();
 sg13g2_decap_4 FILLER_23_1078 ();
 sg13g2_decap_4 FILLER_23_1087 ();
 sg13g2_fill_1 FILLER_23_1122 ();
 sg13g2_decap_8 FILLER_23_1149 ();
 sg13g2_fill_1 FILLER_23_1156 ();
 sg13g2_fill_1 FILLER_23_1187 ();
 sg13g2_fill_2 FILLER_23_1194 ();
 sg13g2_fill_1 FILLER_23_1209 ();
 sg13g2_decap_8 FILLER_23_1233 ();
 sg13g2_decap_8 FILLER_23_1240 ();
 sg13g2_decap_8 FILLER_23_1247 ();
 sg13g2_decap_8 FILLER_23_1254 ();
 sg13g2_decap_8 FILLER_23_1261 ();
 sg13g2_decap_8 FILLER_23_1268 ();
 sg13g2_decap_8 FILLER_23_1280 ();
 sg13g2_fill_1 FILLER_23_1287 ();
 sg13g2_fill_2 FILLER_23_1319 ();
 sg13g2_decap_8 FILLER_23_1353 ();
 sg13g2_decap_8 FILLER_23_1360 ();
 sg13g2_decap_8 FILLER_23_1367 ();
 sg13g2_decap_8 FILLER_23_1374 ();
 sg13g2_fill_2 FILLER_23_1381 ();
 sg13g2_fill_1 FILLER_23_1387 ();
 sg13g2_fill_1 FILLER_23_1394 ();
 sg13g2_fill_1 FILLER_23_1399 ();
 sg13g2_fill_1 FILLER_23_1405 ();
 sg13g2_fill_2 FILLER_23_1467 ();
 sg13g2_decap_8 FILLER_23_1495 ();
 sg13g2_fill_1 FILLER_23_1542 ();
 sg13g2_fill_1 FILLER_23_1560 ();
 sg13g2_fill_1 FILLER_23_1580 ();
 sg13g2_fill_1 FILLER_23_1653 ();
 sg13g2_fill_1 FILLER_23_1663 ();
 sg13g2_fill_1 FILLER_23_1737 ();
 sg13g2_fill_2 FILLER_23_1755 ();
 sg13g2_decap_8 FILLER_23_1778 ();
 sg13g2_decap_8 FILLER_23_1785 ();
 sg13g2_fill_1 FILLER_23_1792 ();
 sg13g2_decap_8 FILLER_23_1797 ();
 sg13g2_decap_4 FILLER_23_1804 ();
 sg13g2_fill_2 FILLER_23_1854 ();
 sg13g2_fill_1 FILLER_23_1856 ();
 sg13g2_fill_1 FILLER_23_1863 ();
 sg13g2_decap_8 FILLER_23_1869 ();
 sg13g2_decap_8 FILLER_23_1876 ();
 sg13g2_decap_4 FILLER_23_1883 ();
 sg13g2_fill_2 FILLER_23_1887 ();
 sg13g2_fill_1 FILLER_23_1894 ();
 sg13g2_fill_1 FILLER_23_1903 ();
 sg13g2_fill_1 FILLER_23_1910 ();
 sg13g2_fill_1 FILLER_23_1917 ();
 sg13g2_fill_1 FILLER_23_1931 ();
 sg13g2_fill_2 FILLER_23_1935 ();
 sg13g2_fill_2 FILLER_23_1946 ();
 sg13g2_fill_1 FILLER_23_1948 ();
 sg13g2_fill_1 FILLER_23_2029 ();
 sg13g2_decap_4 FILLER_23_2048 ();
 sg13g2_decap_4 FILLER_23_2057 ();
 sg13g2_fill_2 FILLER_23_2061 ();
 sg13g2_decap_4 FILLER_23_2067 ();
 sg13g2_decap_4 FILLER_23_2076 ();
 sg13g2_fill_2 FILLER_23_2080 ();
 sg13g2_fill_2 FILLER_23_2098 ();
 sg13g2_fill_2 FILLER_23_2118 ();
 sg13g2_fill_1 FILLER_23_2128 ();
 sg13g2_decap_8 FILLER_23_2166 ();
 sg13g2_decap_8 FILLER_23_2173 ();
 sg13g2_fill_1 FILLER_23_2180 ();
 sg13g2_fill_2 FILLER_23_2186 ();
 sg13g2_fill_1 FILLER_23_2188 ();
 sg13g2_decap_8 FILLER_23_2211 ();
 sg13g2_fill_2 FILLER_23_2266 ();
 sg13g2_fill_1 FILLER_23_2268 ();
 sg13g2_decap_8 FILLER_23_2324 ();
 sg13g2_fill_1 FILLER_23_2331 ();
 sg13g2_decap_8 FILLER_23_2336 ();
 sg13g2_fill_1 FILLER_23_2343 ();
 sg13g2_decap_4 FILLER_23_2348 ();
 sg13g2_decap_8 FILLER_23_2356 ();
 sg13g2_fill_1 FILLER_23_2363 ();
 sg13g2_decap_8 FILLER_23_2368 ();
 sg13g2_decap_8 FILLER_23_2375 ();
 sg13g2_decap_4 FILLER_23_2393 ();
 sg13g2_fill_1 FILLER_23_2401 ();
 sg13g2_fill_2 FILLER_23_2428 ();
 sg13g2_fill_1 FILLER_23_2435 ();
 sg13g2_decap_4 FILLER_23_2449 ();
 sg13g2_fill_1 FILLER_23_2453 ();
 sg13g2_fill_2 FILLER_23_2459 ();
 sg13g2_decap_8 FILLER_23_2465 ();
 sg13g2_decap_4 FILLER_23_2472 ();
 sg13g2_fill_1 FILLER_23_2476 ();
 sg13g2_decap_8 FILLER_23_2602 ();
 sg13g2_decap_8 FILLER_23_2609 ();
 sg13g2_fill_2 FILLER_23_2616 ();
 sg13g2_fill_1 FILLER_23_2618 ();
 sg13g2_fill_1 FILLER_23_2634 ();
 sg13g2_fill_1 FILLER_23_2669 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_1 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_27 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_1 FILLER_24_43 ();
 sg13g2_fill_1 FILLER_24_53 ();
 sg13g2_fill_1 FILLER_24_60 ();
 sg13g2_decap_4 FILLER_24_99 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_1 FILLER_24_142 ();
 sg13g2_decap_4 FILLER_24_169 ();
 sg13g2_fill_1 FILLER_24_177 ();
 sg13g2_fill_2 FILLER_24_196 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_1 FILLER_24_238 ();
 sg13g2_fill_2 FILLER_24_273 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_fill_2 FILLER_24_305 ();
 sg13g2_fill_1 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_317 ();
 sg13g2_decap_4 FILLER_24_324 ();
 sg13g2_fill_2 FILLER_24_328 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_4 FILLER_24_340 ();
 sg13g2_fill_2 FILLER_24_344 ();
 sg13g2_decap_4 FILLER_24_392 ();
 sg13g2_fill_2 FILLER_24_396 ();
 sg13g2_fill_1 FILLER_24_440 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_fill_1 FILLER_24_487 ();
 sg13g2_fill_2 FILLER_24_505 ();
 sg13g2_fill_1 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_531 ();
 sg13g2_decap_8 FILLER_24_538 ();
 sg13g2_fill_2 FILLER_24_545 ();
 sg13g2_decap_4 FILLER_24_587 ();
 sg13g2_fill_1 FILLER_24_595 ();
 sg13g2_fill_2 FILLER_24_601 ();
 sg13g2_fill_1 FILLER_24_613 ();
 sg13g2_fill_1 FILLER_24_619 ();
 sg13g2_decap_4 FILLER_24_630 ();
 sg13g2_fill_1 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_647 ();
 sg13g2_decap_8 FILLER_24_654 ();
 sg13g2_fill_2 FILLER_24_661 ();
 sg13g2_fill_1 FILLER_24_663 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_751 ();
 sg13g2_decap_8 FILLER_24_758 ();
 sg13g2_decap_8 FILLER_24_765 ();
 sg13g2_decap_4 FILLER_24_772 ();
 sg13g2_fill_1 FILLER_24_776 ();
 sg13g2_decap_8 FILLER_24_787 ();
 sg13g2_decap_4 FILLER_24_794 ();
 sg13g2_fill_1 FILLER_24_798 ();
 sg13g2_fill_1 FILLER_24_866 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_fill_2 FILLER_24_907 ();
 sg13g2_fill_1 FILLER_24_909 ();
 sg13g2_fill_2 FILLER_24_927 ();
 sg13g2_decap_4 FILLER_24_963 ();
 sg13g2_fill_2 FILLER_24_967 ();
 sg13g2_decap_4 FILLER_24_973 ();
 sg13g2_fill_1 FILLER_24_1016 ();
 sg13g2_decap_4 FILLER_24_1029 ();
 sg13g2_fill_1 FILLER_24_1033 ();
 sg13g2_fill_1 FILLER_24_1044 ();
 sg13g2_fill_1 FILLER_24_1050 ();
 sg13g2_fill_2 FILLER_24_1056 ();
 sg13g2_fill_1 FILLER_24_1064 ();
 sg13g2_decap_4 FILLER_24_1087 ();
 sg13g2_fill_2 FILLER_24_1091 ();
 sg13g2_decap_4 FILLER_24_1098 ();
 sg13g2_decap_8 FILLER_24_1106 ();
 sg13g2_decap_8 FILLER_24_1118 ();
 sg13g2_decap_8 FILLER_24_1125 ();
 sg13g2_decap_8 FILLER_24_1132 ();
 sg13g2_decap_8 FILLER_24_1139 ();
 sg13g2_decap_8 FILLER_24_1146 ();
 sg13g2_decap_4 FILLER_24_1153 ();
 sg13g2_fill_1 FILLER_24_1157 ();
 sg13g2_decap_8 FILLER_24_1163 ();
 sg13g2_fill_1 FILLER_24_1170 ();
 sg13g2_fill_2 FILLER_24_1197 ();
 sg13g2_decap_4 FILLER_24_1252 ();
 sg13g2_decap_8 FILLER_24_1260 ();
 sg13g2_fill_1 FILLER_24_1267 ();
 sg13g2_fill_2 FILLER_24_1312 ();
 sg13g2_fill_2 FILLER_24_1320 ();
 sg13g2_fill_1 FILLER_24_1322 ();
 sg13g2_decap_8 FILLER_24_1354 ();
 sg13g2_fill_2 FILLER_24_1361 ();
 sg13g2_fill_1 FILLER_24_1363 ();
 sg13g2_fill_2 FILLER_24_1399 ();
 sg13g2_fill_1 FILLER_24_1401 ();
 sg13g2_fill_1 FILLER_24_1408 ();
 sg13g2_decap_8 FILLER_24_1413 ();
 sg13g2_fill_2 FILLER_24_1420 ();
 sg13g2_fill_1 FILLER_24_1422 ();
 sg13g2_fill_1 FILLER_24_1458 ();
 sg13g2_fill_2 FILLER_24_1501 ();
 sg13g2_decap_4 FILLER_24_1529 ();
 sg13g2_fill_2 FILLER_24_1533 ();
 sg13g2_decap_8 FILLER_24_1544 ();
 sg13g2_fill_1 FILLER_24_1570 ();
 sg13g2_decap_4 FILLER_24_1618 ();
 sg13g2_fill_1 FILLER_24_1631 ();
 sg13g2_fill_1 FILLER_24_1695 ();
 sg13g2_fill_1 FILLER_24_1751 ();
 sg13g2_fill_2 FILLER_24_1898 ();
 sg13g2_fill_1 FILLER_24_1900 ();
 sg13g2_decap_8 FILLER_24_1906 ();
 sg13g2_fill_2 FILLER_24_1913 ();
 sg13g2_fill_1 FILLER_24_1946 ();
 sg13g2_decap_8 FILLER_24_1960 ();
 sg13g2_decap_8 FILLER_24_1967 ();
 sg13g2_decap_8 FILLER_24_1974 ();
 sg13g2_decap_4 FILLER_24_1981 ();
 sg13g2_fill_1 FILLER_24_1985 ();
 sg13g2_fill_1 FILLER_24_1991 ();
 sg13g2_decap_4 FILLER_24_2024 ();
 sg13g2_fill_1 FILLER_24_2028 ();
 sg13g2_decap_8 FILLER_24_2033 ();
 sg13g2_decap_4 FILLER_24_2040 ();
 sg13g2_fill_2 FILLER_24_2044 ();
 sg13g2_fill_1 FILLER_24_2052 ();
 sg13g2_fill_2 FILLER_24_2063 ();
 sg13g2_fill_1 FILLER_24_2065 ();
 sg13g2_fill_2 FILLER_24_2103 ();
 sg13g2_fill_1 FILLER_24_2105 ();
 sg13g2_fill_1 FILLER_24_2114 ();
 sg13g2_fill_2 FILLER_24_2153 ();
 sg13g2_fill_1 FILLER_24_2155 ();
 sg13g2_decap_8 FILLER_24_2182 ();
 sg13g2_decap_8 FILLER_24_2189 ();
 sg13g2_fill_2 FILLER_24_2196 ();
 sg13g2_fill_1 FILLER_24_2198 ();
 sg13g2_fill_2 FILLER_24_2229 ();
 sg13g2_fill_1 FILLER_24_2279 ();
 sg13g2_decap_4 FILLER_24_2294 ();
 sg13g2_fill_2 FILLER_24_2303 ();
 sg13g2_decap_8 FILLER_24_2313 ();
 sg13g2_decap_8 FILLER_24_2320 ();
 sg13g2_decap_8 FILLER_24_2327 ();
 sg13g2_decap_8 FILLER_24_2334 ();
 sg13g2_decap_8 FILLER_24_2341 ();
 sg13g2_fill_2 FILLER_24_2348 ();
 sg13g2_fill_1 FILLER_24_2350 ();
 sg13g2_fill_2 FILLER_24_2384 ();
 sg13g2_decap_8 FILLER_24_2432 ();
 sg13g2_decap_8 FILLER_24_2439 ();
 sg13g2_decap_8 FILLER_24_2446 ();
 sg13g2_decap_8 FILLER_24_2453 ();
 sg13g2_fill_2 FILLER_24_2460 ();
 sg13g2_fill_1 FILLER_24_2462 ();
 sg13g2_fill_1 FILLER_24_2493 ();
 sg13g2_fill_2 FILLER_24_2509 ();
 sg13g2_fill_1 FILLER_24_2540 ();
 sg13g2_decap_4 FILLER_24_2567 ();
 sg13g2_decap_8 FILLER_24_2604 ();
 sg13g2_fill_2 FILLER_24_2611 ();
 sg13g2_decap_8 FILLER_24_2657 ();
 sg13g2_decap_4 FILLER_24_2664 ();
 sg13g2_fill_2 FILLER_24_2668 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_fill_2 FILLER_25_39 ();
 sg13g2_fill_2 FILLER_25_45 ();
 sg13g2_fill_1 FILLER_25_47 ();
 sg13g2_decap_8 FILLER_25_90 ();
 sg13g2_decap_8 FILLER_25_97 ();
 sg13g2_decap_8 FILLER_25_104 ();
 sg13g2_decap_8 FILLER_25_111 ();
 sg13g2_fill_1 FILLER_25_130 ();
 sg13g2_fill_1 FILLER_25_137 ();
 sg13g2_fill_1 FILLER_25_142 ();
 sg13g2_fill_1 FILLER_25_148 ();
 sg13g2_fill_1 FILLER_25_184 ();
 sg13g2_fill_2 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_220 ();
 sg13g2_fill_2 FILLER_25_252 ();
 sg13g2_decap_4 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_295 ();
 sg13g2_fill_1 FILLER_25_323 ();
 sg13g2_fill_1 FILLER_25_334 ();
 sg13g2_fill_2 FILLER_25_396 ();
 sg13g2_fill_1 FILLER_25_398 ();
 sg13g2_fill_2 FILLER_25_404 ();
 sg13g2_fill_2 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_25_421 ();
 sg13g2_decap_4 FILLER_25_431 ();
 sg13g2_fill_1 FILLER_25_435 ();
 sg13g2_decap_8 FILLER_25_444 ();
 sg13g2_decap_8 FILLER_25_451 ();
 sg13g2_decap_4 FILLER_25_458 ();
 sg13g2_decap_4 FILLER_25_480 ();
 sg13g2_fill_2 FILLER_25_484 ();
 sg13g2_fill_1 FILLER_25_495 ();
 sg13g2_fill_1 FILLER_25_499 ();
 sg13g2_fill_1 FILLER_25_508 ();
 sg13g2_fill_2 FILLER_25_529 ();
 sg13g2_decap_8 FILLER_25_541 ();
 sg13g2_fill_2 FILLER_25_548 ();
 sg13g2_fill_1 FILLER_25_550 ();
 sg13g2_decap_8 FILLER_25_582 ();
 sg13g2_fill_2 FILLER_25_589 ();
 sg13g2_fill_1 FILLER_25_591 ();
 sg13g2_decap_4 FILLER_25_597 ();
 sg13g2_fill_1 FILLER_25_606 ();
 sg13g2_fill_2 FILLER_25_616 ();
 sg13g2_fill_2 FILLER_25_623 ();
 sg13g2_fill_1 FILLER_25_625 ();
 sg13g2_decap_8 FILLER_25_634 ();
 sg13g2_decap_4 FILLER_25_641 ();
 sg13g2_fill_2 FILLER_25_650 ();
 sg13g2_fill_2 FILLER_25_668 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_4 FILLER_25_747 ();
 sg13g2_fill_1 FILLER_25_751 ();
 sg13g2_decap_8 FILLER_25_778 ();
 sg13g2_decap_8 FILLER_25_785 ();
 sg13g2_decap_8 FILLER_25_792 ();
 sg13g2_decap_4 FILLER_25_799 ();
 sg13g2_decap_8 FILLER_25_807 ();
 sg13g2_fill_2 FILLER_25_814 ();
 sg13g2_decap_4 FILLER_25_886 ();
 sg13g2_fill_1 FILLER_25_890 ();
 sg13g2_decap_8 FILLER_25_895 ();
 sg13g2_fill_2 FILLER_25_902 ();
 sg13g2_decap_8 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_4 FILLER_25_973 ();
 sg13g2_fill_1 FILLER_25_977 ();
 sg13g2_decap_8 FILLER_25_982 ();
 sg13g2_decap_8 FILLER_25_989 ();
 sg13g2_decap_8 FILLER_25_996 ();
 sg13g2_fill_2 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1028 ();
 sg13g2_decap_4 FILLER_25_1040 ();
 sg13g2_fill_1 FILLER_25_1048 ();
 sg13g2_decap_4 FILLER_25_1088 ();
 sg13g2_fill_1 FILLER_25_1092 ();
 sg13g2_fill_2 FILLER_25_1096 ();
 sg13g2_fill_1 FILLER_25_1098 ();
 sg13g2_decap_8 FILLER_25_1124 ();
 sg13g2_decap_8 FILLER_25_1131 ();
 sg13g2_decap_8 FILLER_25_1138 ();
 sg13g2_decap_4 FILLER_25_1145 ();
 sg13g2_fill_2 FILLER_25_1149 ();
 sg13g2_fill_2 FILLER_25_1155 ();
 sg13g2_fill_1 FILLER_25_1157 ();
 sg13g2_fill_2 FILLER_25_1164 ();
 sg13g2_fill_2 FILLER_25_1171 ();
 sg13g2_fill_1 FILLER_25_1173 ();
 sg13g2_fill_1 FILLER_25_1178 ();
 sg13g2_fill_1 FILLER_25_1183 ();
 sg13g2_fill_2 FILLER_25_1204 ();
 sg13g2_fill_1 FILLER_25_1217 ();
 sg13g2_fill_1 FILLER_25_1224 ();
 sg13g2_fill_2 FILLER_25_1231 ();
 sg13g2_decap_4 FILLER_25_1259 ();
 sg13g2_fill_2 FILLER_25_1263 ();
 sg13g2_decap_8 FILLER_25_1297 ();
 sg13g2_decap_8 FILLER_25_1313 ();
 sg13g2_decap_8 FILLER_25_1320 ();
 sg13g2_decap_4 FILLER_25_1327 ();
 sg13g2_fill_1 FILLER_25_1336 ();
 sg13g2_decap_8 FILLER_25_1341 ();
 sg13g2_fill_1 FILLER_25_1348 ();
 sg13g2_decap_4 FILLER_25_1353 ();
 sg13g2_fill_1 FILLER_25_1357 ();
 sg13g2_fill_1 FILLER_25_1362 ();
 sg13g2_decap_4 FILLER_25_1368 ();
 sg13g2_fill_1 FILLER_25_1372 ();
 sg13g2_decap_8 FILLER_25_1379 ();
 sg13g2_decap_4 FILLER_25_1390 ();
 sg13g2_fill_1 FILLER_25_1394 ();
 sg13g2_decap_8 FILLER_25_1421 ();
 sg13g2_decap_8 FILLER_25_1428 ();
 sg13g2_decap_8 FILLER_25_1451 ();
 sg13g2_decap_8 FILLER_25_1458 ();
 sg13g2_decap_8 FILLER_25_1465 ();
 sg13g2_decap_8 FILLER_25_1472 ();
 sg13g2_decap_8 FILLER_25_1479 ();
 sg13g2_decap_4 FILLER_25_1486 ();
 sg13g2_fill_2 FILLER_25_1515 ();
 sg13g2_fill_1 FILLER_25_1517 ();
 sg13g2_decap_8 FILLER_25_1521 ();
 sg13g2_fill_1 FILLER_25_1528 ();
 sg13g2_decap_8 FILLER_25_1539 ();
 sg13g2_decap_8 FILLER_25_1546 ();
 sg13g2_decap_8 FILLER_25_1553 ();
 sg13g2_decap_8 FILLER_25_1560 ();
 sg13g2_fill_1 FILLER_25_1567 ();
 sg13g2_decap_8 FILLER_25_1577 ();
 sg13g2_fill_1 FILLER_25_1584 ();
 sg13g2_fill_1 FILLER_25_1634 ();
 sg13g2_fill_2 FILLER_25_1653 ();
 sg13g2_fill_2 FILLER_25_1687 ();
 sg13g2_fill_1 FILLER_25_1741 ();
 sg13g2_fill_1 FILLER_25_1747 ();
 sg13g2_fill_1 FILLER_25_1777 ();
 sg13g2_fill_2 FILLER_25_1823 ();
 sg13g2_decap_8 FILLER_25_1829 ();
 sg13g2_fill_1 FILLER_25_1836 ();
 sg13g2_fill_2 FILLER_25_1843 ();
 sg13g2_decap_8 FILLER_25_1850 ();
 sg13g2_fill_2 FILLER_25_1857 ();
 sg13g2_fill_1 FILLER_25_1859 ();
 sg13g2_fill_2 FILLER_25_1870 ();
 sg13g2_fill_2 FILLER_25_1883 ();
 sg13g2_fill_2 FILLER_25_1943 ();
 sg13g2_decap_8 FILLER_25_1959 ();
 sg13g2_decap_8 FILLER_25_1966 ();
 sg13g2_fill_2 FILLER_25_1973 ();
 sg13g2_decap_8 FILLER_25_2018 ();
 sg13g2_decap_8 FILLER_25_2025 ();
 sg13g2_decap_4 FILLER_25_2032 ();
 sg13g2_fill_1 FILLER_25_2036 ();
 sg13g2_fill_1 FILLER_25_2100 ();
 sg13g2_fill_2 FILLER_25_2112 ();
 sg13g2_fill_2 FILLER_25_2138 ();
 sg13g2_fill_1 FILLER_25_2140 ();
 sg13g2_fill_2 FILLER_25_2156 ();
 sg13g2_fill_1 FILLER_25_2158 ();
 sg13g2_fill_2 FILLER_25_2185 ();
 sg13g2_fill_1 FILLER_25_2187 ();
 sg13g2_decap_8 FILLER_25_2214 ();
 sg13g2_fill_1 FILLER_25_2233 ();
 sg13g2_fill_2 FILLER_25_2240 ();
 sg13g2_fill_2 FILLER_25_2296 ();
 sg13g2_decap_8 FILLER_25_2314 ();
 sg13g2_decap_8 FILLER_25_2321 ();
 sg13g2_decap_4 FILLER_25_2328 ();
 sg13g2_decap_8 FILLER_25_2340 ();
 sg13g2_decap_8 FILLER_25_2347 ();
 sg13g2_fill_2 FILLER_25_2354 ();
 sg13g2_fill_1 FILLER_25_2356 ();
 sg13g2_decap_4 FILLER_25_2365 ();
 sg13g2_fill_1 FILLER_25_2369 ();
 sg13g2_fill_2 FILLER_25_2382 ();
 sg13g2_decap_8 FILLER_25_2424 ();
 sg13g2_fill_1 FILLER_25_2431 ();
 sg13g2_decap_8 FILLER_25_2458 ();
 sg13g2_decap_4 FILLER_25_2465 ();
 sg13g2_fill_2 FILLER_25_2492 ();
 sg13g2_decap_4 FILLER_25_2562 ();
 sg13g2_fill_1 FILLER_25_2566 ();
 sg13g2_decap_4 FILLER_25_2577 ();
 sg13g2_fill_1 FILLER_25_2581 ();
 sg13g2_fill_1 FILLER_25_2615 ();
 sg13g2_fill_1 FILLER_25_2638 ();
 sg13g2_fill_2 FILLER_25_2658 ();
 sg13g2_fill_1 FILLER_25_2660 ();
 sg13g2_decap_4 FILLER_25_2665 ();
 sg13g2_fill_1 FILLER_25_2669 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_4 FILLER_26_14 ();
 sg13g2_fill_1 FILLER_26_18 ();
 sg13g2_fill_2 FILLER_26_45 ();
 sg13g2_fill_1 FILLER_26_47 ();
 sg13g2_fill_2 FILLER_26_69 ();
 sg13g2_decap_8 FILLER_26_87 ();
 sg13g2_decap_8 FILLER_26_94 ();
 sg13g2_decap_4 FILLER_26_101 ();
 sg13g2_decap_8 FILLER_26_109 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_125 ();
 sg13g2_fill_1 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_4 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_192 ();
 sg13g2_fill_2 FILLER_26_213 ();
 sg13g2_fill_1 FILLER_26_232 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_2 FILLER_26_301 ();
 sg13g2_fill_1 FILLER_26_329 ();
 sg13g2_decap_4 FILLER_26_355 ();
 sg13g2_fill_2 FILLER_26_359 ();
 sg13g2_fill_2 FILLER_26_382 ();
 sg13g2_fill_1 FILLER_26_384 ();
 sg13g2_decap_4 FILLER_26_428 ();
 sg13g2_fill_2 FILLER_26_432 ();
 sg13g2_decap_8 FILLER_26_439 ();
 sg13g2_fill_1 FILLER_26_446 ();
 sg13g2_decap_4 FILLER_26_452 ();
 sg13g2_fill_2 FILLER_26_456 ();
 sg13g2_fill_2 FILLER_26_484 ();
 sg13g2_fill_1 FILLER_26_525 ();
 sg13g2_fill_1 FILLER_26_535 ();
 sg13g2_decap_8 FILLER_26_541 ();
 sg13g2_decap_8 FILLER_26_561 ();
 sg13g2_decap_4 FILLER_26_568 ();
 sg13g2_decap_8 FILLER_26_582 ();
 sg13g2_decap_4 FILLER_26_589 ();
 sg13g2_fill_2 FILLER_26_597 ();
 sg13g2_fill_1 FILLER_26_599 ();
 sg13g2_fill_2 FILLER_26_650 ();
 sg13g2_decap_4 FILLER_26_674 ();
 sg13g2_fill_1 FILLER_26_678 ();
 sg13g2_fill_1 FILLER_26_709 ();
 sg13g2_decap_8 FILLER_26_722 ();
 sg13g2_decap_8 FILLER_26_729 ();
 sg13g2_decap_8 FILLER_26_736 ();
 sg13g2_decap_8 FILLER_26_743 ();
 sg13g2_decap_4 FILLER_26_750 ();
 sg13g2_decap_4 FILLER_26_759 ();
 sg13g2_fill_1 FILLER_26_763 ();
 sg13g2_decap_4 FILLER_26_768 ();
 sg13g2_fill_2 FILLER_26_772 ();
 sg13g2_fill_1 FILLER_26_818 ();
 sg13g2_fill_1 FILLER_26_824 ();
 sg13g2_fill_2 FILLER_26_829 ();
 sg13g2_fill_1 FILLER_26_870 ();
 sg13g2_decap_8 FILLER_26_891 ();
 sg13g2_decap_8 FILLER_26_898 ();
 sg13g2_fill_1 FILLER_26_905 ();
 sg13g2_decap_8 FILLER_26_915 ();
 sg13g2_decap_8 FILLER_26_922 ();
 sg13g2_fill_1 FILLER_26_929 ();
 sg13g2_decap_4 FILLER_26_943 ();
 sg13g2_fill_2 FILLER_26_947 ();
 sg13g2_fill_2 FILLER_26_961 ();
 sg13g2_fill_2 FILLER_26_989 ();
 sg13g2_fill_1 FILLER_26_1021 ();
 sg13g2_decap_8 FILLER_26_1031 ();
 sg13g2_decap_4 FILLER_26_1078 ();
 sg13g2_fill_2 FILLER_26_1082 ();
 sg13g2_decap_4 FILLER_26_1120 ();
 sg13g2_decap_8 FILLER_26_1181 ();
 sg13g2_fill_2 FILLER_26_1188 ();
 sg13g2_fill_1 FILLER_26_1190 ();
 sg13g2_decap_4 FILLER_26_1230 ();
 sg13g2_fill_2 FILLER_26_1234 ();
 sg13g2_decap_8 FILLER_26_1241 ();
 sg13g2_fill_1 FILLER_26_1258 ();
 sg13g2_fill_1 FILLER_26_1267 ();
 sg13g2_decap_4 FILLER_26_1276 ();
 sg13g2_fill_1 FILLER_26_1293 ();
 sg13g2_decap_4 FILLER_26_1320 ();
 sg13g2_fill_1 FILLER_26_1324 ();
 sg13g2_decap_8 FILLER_26_1374 ();
 sg13g2_fill_2 FILLER_26_1386 ();
 sg13g2_fill_1 FILLER_26_1388 ();
 sg13g2_fill_2 FILLER_26_1411 ();
 sg13g2_decap_8 FILLER_26_1464 ();
 sg13g2_decap_4 FILLER_26_1471 ();
 sg13g2_fill_2 FILLER_26_1475 ();
 sg13g2_fill_1 FILLER_26_1489 ();
 sg13g2_fill_2 FILLER_26_1496 ();
 sg13g2_fill_1 FILLER_26_1498 ();
 sg13g2_fill_2 FILLER_26_1530 ();
 sg13g2_fill_1 FILLER_26_1532 ();
 sg13g2_fill_2 FILLER_26_1543 ();
 sg13g2_fill_1 FILLER_26_1545 ();
 sg13g2_fill_2 FILLER_26_1560 ();
 sg13g2_fill_1 FILLER_26_1562 ();
 sg13g2_decap_8 FILLER_26_1571 ();
 sg13g2_decap_8 FILLER_26_1578 ();
 sg13g2_decap_8 FILLER_26_1585 ();
 sg13g2_decap_4 FILLER_26_1592 ();
 sg13g2_fill_1 FILLER_26_1596 ();
 sg13g2_fill_2 FILLER_26_1601 ();
 sg13g2_fill_2 FILLER_26_1609 ();
 sg13g2_fill_2 FILLER_26_1642 ();
 sg13g2_fill_2 FILLER_26_1660 ();
 sg13g2_fill_1 FILLER_26_1692 ();
 sg13g2_fill_1 FILLER_26_1711 ();
 sg13g2_fill_2 FILLER_26_1731 ();
 sg13g2_fill_1 FILLER_26_1754 ();
 sg13g2_decap_8 FILLER_26_1781 ();
 sg13g2_fill_2 FILLER_26_1788 ();
 sg13g2_fill_2 FILLER_26_1800 ();
 sg13g2_fill_1 FILLER_26_1802 ();
 sg13g2_decap_8 FILLER_26_1808 ();
 sg13g2_decap_4 FILLER_26_1815 ();
 sg13g2_fill_2 FILLER_26_1819 ();
 sg13g2_fill_2 FILLER_26_1830 ();
 sg13g2_decap_4 FILLER_26_1842 ();
 sg13g2_decap_8 FILLER_26_1855 ();
 sg13g2_decap_8 FILLER_26_1862 ();
 sg13g2_fill_2 FILLER_26_1889 ();
 sg13g2_fill_1 FILLER_26_1891 ();
 sg13g2_fill_2 FILLER_26_1906 ();
 sg13g2_fill_1 FILLER_26_1908 ();
 sg13g2_fill_2 FILLER_26_1943 ();
 sg13g2_fill_1 FILLER_26_1945 ();
 sg13g2_decap_8 FILLER_26_1959 ();
 sg13g2_decap_8 FILLER_26_1966 ();
 sg13g2_fill_2 FILLER_26_1973 ();
 sg13g2_decap_8 FILLER_26_2001 ();
 sg13g2_decap_8 FILLER_26_2008 ();
 sg13g2_decap_4 FILLER_26_2015 ();
 sg13g2_decap_4 FILLER_26_2027 ();
 sg13g2_fill_1 FILLER_26_2057 ();
 sg13g2_fill_1 FILLER_26_2094 ();
 sg13g2_fill_2 FILLER_26_2116 ();
 sg13g2_fill_1 FILLER_26_2118 ();
 sg13g2_fill_1 FILLER_26_2125 ();
 sg13g2_decap_4 FILLER_26_2132 ();
 sg13g2_fill_2 FILLER_26_2136 ();
 sg13g2_decap_8 FILLER_26_2143 ();
 sg13g2_fill_1 FILLER_26_2150 ();
 sg13g2_fill_2 FILLER_26_2177 ();
 sg13g2_decap_8 FILLER_26_2188 ();
 sg13g2_decap_4 FILLER_26_2195 ();
 sg13g2_decap_8 FILLER_26_2208 ();
 sg13g2_decap_4 FILLER_26_2215 ();
 sg13g2_fill_2 FILLER_26_2219 ();
 sg13g2_fill_2 FILLER_26_2247 ();
 sg13g2_fill_2 FILLER_26_2281 ();
 sg13g2_fill_2 FILLER_26_2361 ();
 sg13g2_fill_1 FILLER_26_2377 ();
 sg13g2_fill_1 FILLER_26_2383 ();
 sg13g2_fill_2 FILLER_26_2408 ();
 sg13g2_decap_8 FILLER_26_2415 ();
 sg13g2_fill_2 FILLER_26_2422 ();
 sg13g2_decap_4 FILLER_26_2454 ();
 sg13g2_decap_8 FILLER_26_2462 ();
 sg13g2_decap_8 FILLER_26_2469 ();
 sg13g2_fill_2 FILLER_26_2476 ();
 sg13g2_fill_1 FILLER_26_2478 ();
 sg13g2_fill_1 FILLER_26_2497 ();
 sg13g2_fill_1 FILLER_26_2528 ();
 sg13g2_decap_8 FILLER_26_2543 ();
 sg13g2_decap_4 FILLER_26_2550 ();
 sg13g2_fill_2 FILLER_26_2554 ();
 sg13g2_fill_2 FILLER_26_2595 ();
 sg13g2_fill_2 FILLER_26_2668 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_fill_2 FILLER_27_14 ();
 sg13g2_fill_2 FILLER_27_54 ();
 sg13g2_fill_1 FILLER_27_56 ();
 sg13g2_fill_2 FILLER_27_96 ();
 sg13g2_decap_8 FILLER_27_133 ();
 sg13g2_decap_8 FILLER_27_140 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_8 FILLER_27_154 ();
 sg13g2_decap_8 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_168 ();
 sg13g2_fill_1 FILLER_27_173 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_193 ();
 sg13g2_fill_2 FILLER_27_235 ();
 sg13g2_fill_1 FILLER_27_246 ();
 sg13g2_fill_1 FILLER_27_335 ();
 sg13g2_decap_4 FILLER_27_374 ();
 sg13g2_decap_8 FILLER_27_381 ();
 sg13g2_decap_8 FILLER_27_388 ();
 sg13g2_decap_8 FILLER_27_395 ();
 sg13g2_fill_2 FILLER_27_414 ();
 sg13g2_fill_2 FILLER_27_420 ();
 sg13g2_decap_8 FILLER_27_429 ();
 sg13g2_fill_1 FILLER_27_436 ();
 sg13g2_decap_8 FILLER_27_442 ();
 sg13g2_fill_2 FILLER_27_453 ();
 sg13g2_fill_1 FILLER_27_455 ();
 sg13g2_fill_1 FILLER_27_461 ();
 sg13g2_decap_4 FILLER_27_465 ();
 sg13g2_fill_1 FILLER_27_491 ();
 sg13g2_fill_2 FILLER_27_505 ();
 sg13g2_fill_1 FILLER_27_507 ();
 sg13g2_fill_1 FILLER_27_523 ();
 sg13g2_fill_1 FILLER_27_540 ();
 sg13g2_fill_1 FILLER_27_546 ();
 sg13g2_fill_2 FILLER_27_587 ();
 sg13g2_decap_4 FILLER_27_620 ();
 sg13g2_fill_1 FILLER_27_624 ();
 sg13g2_fill_1 FILLER_27_638 ();
 sg13g2_fill_1 FILLER_27_658 ();
 sg13g2_fill_1 FILLER_27_662 ();
 sg13g2_fill_2 FILLER_27_666 ();
 sg13g2_fill_2 FILLER_27_671 ();
 sg13g2_fill_2 FILLER_27_687 ();
 sg13g2_fill_1 FILLER_27_689 ();
 sg13g2_decap_8 FILLER_27_731 ();
 sg13g2_decap_8 FILLER_27_738 ();
 sg13g2_decap_4 FILLER_27_745 ();
 sg13g2_fill_2 FILLER_27_749 ();
 sg13g2_fill_2 FILLER_27_777 ();
 sg13g2_fill_1 FILLER_27_814 ();
 sg13g2_fill_2 FILLER_27_819 ();
 sg13g2_fill_1 FILLER_27_830 ();
 sg13g2_fill_2 FILLER_27_857 ();
 sg13g2_fill_2 FILLER_27_903 ();
 sg13g2_decap_8 FILLER_27_909 ();
 sg13g2_fill_2 FILLER_27_916 ();
 sg13g2_decap_4 FILLER_27_975 ();
 sg13g2_fill_1 FILLER_27_979 ();
 sg13g2_decap_8 FILLER_27_989 ();
 sg13g2_decap_4 FILLER_27_996 ();
 sg13g2_fill_1 FILLER_27_1008 ();
 sg13g2_decap_8 FILLER_27_1025 ();
 sg13g2_decap_8 FILLER_27_1032 ();
 sg13g2_decap_8 FILLER_27_1039 ();
 sg13g2_decap_4 FILLER_27_1050 ();
 sg13g2_fill_2 FILLER_27_1061 ();
 sg13g2_decap_8 FILLER_27_1066 ();
 sg13g2_decap_8 FILLER_27_1073 ();
 sg13g2_fill_1 FILLER_27_1080 ();
 sg13g2_fill_1 FILLER_27_1122 ();
 sg13g2_fill_1 FILLER_27_1128 ();
 sg13g2_fill_1 FILLER_27_1155 ();
 sg13g2_fill_1 FILLER_27_1162 ();
 sg13g2_fill_2 FILLER_27_1169 ();
 sg13g2_fill_2 FILLER_27_1175 ();
 sg13g2_decap_8 FILLER_27_1183 ();
 sg13g2_fill_1 FILLER_27_1190 ();
 sg13g2_decap_4 FILLER_27_1196 ();
 sg13g2_decap_4 FILLER_27_1204 ();
 sg13g2_fill_2 FILLER_27_1208 ();
 sg13g2_fill_2 FILLER_27_1236 ();
 sg13g2_decap_4 FILLER_27_1264 ();
 sg13g2_fill_1 FILLER_27_1287 ();
 sg13g2_decap_4 FILLER_27_1303 ();
 sg13g2_fill_2 FILLER_27_1307 ();
 sg13g2_decap_8 FILLER_27_1335 ();
 sg13g2_decap_8 FILLER_27_1342 ();
 sg13g2_decap_8 FILLER_27_1384 ();
 sg13g2_decap_8 FILLER_27_1391 ();
 sg13g2_decap_4 FILLER_27_1398 ();
 sg13g2_fill_2 FILLER_27_1402 ();
 sg13g2_decap_8 FILLER_27_1407 ();
 sg13g2_decap_8 FILLER_27_1414 ();
 sg13g2_fill_2 FILLER_27_1421 ();
 sg13g2_fill_1 FILLER_27_1436 ();
 sg13g2_fill_2 FILLER_27_1449 ();
 sg13g2_fill_1 FILLER_27_1527 ();
 sg13g2_fill_1 FILLER_27_1557 ();
 sg13g2_fill_2 FILLER_27_1584 ();
 sg13g2_fill_1 FILLER_27_1586 ();
 sg13g2_decap_8 FILLER_27_1590 ();
 sg13g2_fill_2 FILLER_27_1597 ();
 sg13g2_fill_1 FILLER_27_1599 ();
 sg13g2_decap_4 FILLER_27_1609 ();
 sg13g2_fill_1 FILLER_27_1613 ();
 sg13g2_fill_2 FILLER_27_1641 ();
 sg13g2_fill_1 FILLER_27_1695 ();
 sg13g2_fill_2 FILLER_27_1716 ();
 sg13g2_decap_4 FILLER_27_1748 ();
 sg13g2_fill_2 FILLER_27_1752 ();
 sg13g2_decap_4 FILLER_27_1795 ();
 sg13g2_decap_4 FILLER_27_1804 ();
 sg13g2_fill_1 FILLER_27_1812 ();
 sg13g2_decap_8 FILLER_27_1835 ();
 sg13g2_decap_8 FILLER_27_1842 ();
 sg13g2_decap_8 FILLER_27_1849 ();
 sg13g2_decap_4 FILLER_27_1856 ();
 sg13g2_decap_8 FILLER_27_1895 ();
 sg13g2_decap_8 FILLER_27_1902 ();
 sg13g2_decap_8 FILLER_27_1909 ();
 sg13g2_fill_2 FILLER_27_1916 ();
 sg13g2_fill_1 FILLER_27_1918 ();
 sg13g2_decap_8 FILLER_27_1925 ();
 sg13g2_fill_2 FILLER_27_1932 ();
 sg13g2_fill_1 FILLER_27_1934 ();
 sg13g2_decap_4 FILLER_27_1948 ();
 sg13g2_fill_2 FILLER_27_1995 ();
 sg13g2_fill_2 FILLER_27_2011 ();
 sg13g2_fill_1 FILLER_27_2039 ();
 sg13g2_fill_1 FILLER_27_2072 ();
 sg13g2_fill_2 FILLER_27_2118 ();
 sg13g2_fill_1 FILLER_27_2120 ();
 sg13g2_decap_8 FILLER_27_2160 ();
 sg13g2_decap_4 FILLER_27_2167 ();
 sg13g2_decap_8 FILLER_27_2176 ();
 sg13g2_decap_8 FILLER_27_2183 ();
 sg13g2_decap_8 FILLER_27_2190 ();
 sg13g2_decap_8 FILLER_27_2197 ();
 sg13g2_decap_8 FILLER_27_2204 ();
 sg13g2_fill_1 FILLER_27_2211 ();
 sg13g2_decap_8 FILLER_27_2284 ();
 sg13g2_decap_8 FILLER_27_2291 ();
 sg13g2_decap_8 FILLER_27_2298 ();
 sg13g2_decap_4 FILLER_27_2305 ();
 sg13g2_fill_1 FILLER_27_2334 ();
 sg13g2_fill_1 FILLER_27_2399 ();
 sg13g2_fill_2 FILLER_27_2404 ();
 sg13g2_fill_1 FILLER_27_2406 ();
 sg13g2_fill_2 FILLER_27_2416 ();
 sg13g2_decap_4 FILLER_27_2424 ();
 sg13g2_decap_4 FILLER_27_2432 ();
 sg13g2_fill_1 FILLER_27_2440 ();
 sg13g2_fill_2 FILLER_27_2449 ();
 sg13g2_decap_8 FILLER_27_2481 ();
 sg13g2_fill_2 FILLER_27_2493 ();
 sg13g2_fill_1 FILLER_27_2525 ();
 sg13g2_decap_8 FILLER_27_2541 ();
 sg13g2_fill_2 FILLER_27_2548 ();
 sg13g2_fill_1 FILLER_27_2550 ();
 sg13g2_fill_1 FILLER_27_2555 ();
 sg13g2_fill_1 FILLER_27_2616 ();
 sg13g2_fill_1 FILLER_27_2622 ();
 sg13g2_fill_2 FILLER_27_2635 ();
 sg13g2_fill_1 FILLER_27_2647 ();
 sg13g2_decap_8 FILLER_27_2653 ();
 sg13g2_decap_8 FILLER_27_2660 ();
 sg13g2_fill_2 FILLER_27_2667 ();
 sg13g2_fill_1 FILLER_27_2669 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_4 FILLER_28_21 ();
 sg13g2_fill_2 FILLER_28_25 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_80 ();
 sg13g2_decap_8 FILLER_28_87 ();
 sg13g2_decap_8 FILLER_28_94 ();
 sg13g2_decap_8 FILLER_28_101 ();
 sg13g2_decap_8 FILLER_28_108 ();
 sg13g2_decap_8 FILLER_28_115 ();
 sg13g2_decap_8 FILLER_28_122 ();
 sg13g2_decap_8 FILLER_28_129 ();
 sg13g2_decap_8 FILLER_28_136 ();
 sg13g2_fill_2 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_149 ();
 sg13g2_decap_8 FILLER_28_156 ();
 sg13g2_fill_2 FILLER_28_163 ();
 sg13g2_fill_1 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_260 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_2 FILLER_28_275 ();
 sg13g2_fill_1 FILLER_28_295 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_4 FILLER_28_308 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_decap_8 FILLER_28_318 ();
 sg13g2_decap_4 FILLER_28_325 ();
 sg13g2_fill_1 FILLER_28_329 ();
 sg13g2_decap_4 FILLER_28_342 ();
 sg13g2_fill_2 FILLER_28_346 ();
 sg13g2_decap_8 FILLER_28_351 ();
 sg13g2_decap_8 FILLER_28_358 ();
 sg13g2_decap_8 FILLER_28_365 ();
 sg13g2_decap_8 FILLER_28_372 ();
 sg13g2_decap_8 FILLER_28_384 ();
 sg13g2_fill_2 FILLER_28_396 ();
 sg13g2_fill_1 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_28_421 ();
 sg13g2_decap_4 FILLER_28_429 ();
 sg13g2_fill_2 FILLER_28_433 ();
 sg13g2_fill_1 FILLER_28_465 ();
 sg13g2_fill_1 FILLER_28_495 ();
 sg13g2_fill_1 FILLER_28_501 ();
 sg13g2_fill_1 FILLER_28_510 ();
 sg13g2_fill_2 FILLER_28_548 ();
 sg13g2_fill_1 FILLER_28_550 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_fill_1 FILLER_28_567 ();
 sg13g2_fill_1 FILLER_28_572 ();
 sg13g2_fill_2 FILLER_28_578 ();
 sg13g2_fill_1 FILLER_28_580 ();
 sg13g2_decap_8 FILLER_28_596 ();
 sg13g2_decap_4 FILLER_28_603 ();
 sg13g2_fill_2 FILLER_28_607 ();
 sg13g2_fill_2 FILLER_28_628 ();
 sg13g2_fill_1 FILLER_28_647 ();
 sg13g2_fill_2 FILLER_28_656 ();
 sg13g2_fill_2 FILLER_28_664 ();
 sg13g2_decap_8 FILLER_28_682 ();
 sg13g2_fill_1 FILLER_28_689 ();
 sg13g2_fill_2 FILLER_28_695 ();
 sg13g2_fill_1 FILLER_28_725 ();
 sg13g2_decap_4 FILLER_28_731 ();
 sg13g2_decap_8 FILLER_28_740 ();
 sg13g2_fill_2 FILLER_28_747 ();
 sg13g2_decap_8 FILLER_28_762 ();
 sg13g2_fill_2 FILLER_28_769 ();
 sg13g2_fill_1 FILLER_28_771 ();
 sg13g2_decap_4 FILLER_28_806 ();
 sg13g2_decap_4 FILLER_28_829 ();
 sg13g2_fill_2 FILLER_28_833 ();
 sg13g2_fill_2 FILLER_28_862 ();
 sg13g2_decap_8 FILLER_28_909 ();
 sg13g2_decap_8 FILLER_28_916 ();
 sg13g2_decap_4 FILLER_28_923 ();
 sg13g2_fill_1 FILLER_28_927 ();
 sg13g2_fill_2 FILLER_28_949 ();
 sg13g2_decap_4 FILLER_28_991 ();
 sg13g2_fill_2 FILLER_28_995 ();
 sg13g2_fill_2 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1045 ();
 sg13g2_fill_2 FILLER_28_1052 ();
 sg13g2_fill_1 FILLER_28_1054 ();
 sg13g2_fill_1 FILLER_28_1090 ();
 sg13g2_fill_2 FILLER_28_1122 ();
 sg13g2_fill_1 FILLER_28_1124 ();
 sg13g2_fill_2 FILLER_28_1129 ();
 sg13g2_fill_1 FILLER_28_1131 ();
 sg13g2_fill_1 FILLER_28_1137 ();
 sg13g2_fill_1 FILLER_28_1142 ();
 sg13g2_fill_1 FILLER_28_1169 ();
 sg13g2_decap_8 FILLER_28_1196 ();
 sg13g2_decap_8 FILLER_28_1203 ();
 sg13g2_decap_8 FILLER_28_1210 ();
 sg13g2_decap_8 FILLER_28_1217 ();
 sg13g2_fill_1 FILLER_28_1224 ();
 sg13g2_fill_1 FILLER_28_1230 ();
 sg13g2_fill_1 FILLER_28_1240 ();
 sg13g2_fill_1 FILLER_28_1273 ();
 sg13g2_fill_1 FILLER_28_1326 ();
 sg13g2_fill_1 FILLER_28_1332 ();
 sg13g2_decap_8 FILLER_28_1337 ();
 sg13g2_fill_2 FILLER_28_1344 ();
 sg13g2_fill_1 FILLER_28_1346 ();
 sg13g2_fill_2 FILLER_28_1352 ();
 sg13g2_decap_8 FILLER_28_1389 ();
 sg13g2_decap_8 FILLER_28_1396 ();
 sg13g2_fill_1 FILLER_28_1403 ();
 sg13g2_decap_8 FILLER_28_1472 ();
 sg13g2_decap_8 FILLER_28_1479 ();
 sg13g2_decap_4 FILLER_28_1486 ();
 sg13g2_fill_1 FILLER_28_1499 ();
 sg13g2_fill_2 FILLER_28_1503 ();
 sg13g2_decap_8 FILLER_28_1531 ();
 sg13g2_decap_8 FILLER_28_1538 ();
 sg13g2_fill_2 FILLER_28_1545 ();
 sg13g2_fill_1 FILLER_28_1547 ();
 sg13g2_fill_1 FILLER_28_1562 ();
 sg13g2_decap_8 FILLER_28_1567 ();
 sg13g2_decap_4 FILLER_28_1574 ();
 sg13g2_fill_1 FILLER_28_1578 ();
 sg13g2_fill_1 FILLER_28_1583 ();
 sg13g2_fill_2 FILLER_28_1603 ();
 sg13g2_fill_2 FILLER_28_1617 ();
 sg13g2_fill_2 FILLER_28_1626 ();
 sg13g2_fill_2 FILLER_28_1698 ();
 sg13g2_fill_1 FILLER_28_1726 ();
 sg13g2_decap_8 FILLER_28_1763 ();
 sg13g2_decap_8 FILLER_28_1770 ();
 sg13g2_decap_4 FILLER_28_1777 ();
 sg13g2_fill_2 FILLER_28_1781 ();
 sg13g2_fill_1 FILLER_28_1819 ();
 sg13g2_fill_1 FILLER_28_1886 ();
 sg13g2_decap_8 FILLER_28_1892 ();
 sg13g2_fill_2 FILLER_28_1899 ();
 sg13g2_fill_1 FILLER_28_1901 ();
 sg13g2_fill_2 FILLER_28_1917 ();
 sg13g2_fill_1 FILLER_28_1967 ();
 sg13g2_fill_2 FILLER_28_1978 ();
 sg13g2_decap_8 FILLER_28_2001 ();
 sg13g2_decap_4 FILLER_28_2022 ();
 sg13g2_fill_1 FILLER_28_2026 ();
 sg13g2_fill_1 FILLER_28_2036 ();
 sg13g2_fill_2 FILLER_28_2057 ();
 sg13g2_decap_4 FILLER_28_2067 ();
 sg13g2_fill_2 FILLER_28_2071 ();
 sg13g2_decap_8 FILLER_28_2081 ();
 sg13g2_fill_1 FILLER_28_2088 ();
 sg13g2_fill_2 FILLER_28_2107 ();
 sg13g2_decap_8 FILLER_28_2114 ();
 sg13g2_decap_4 FILLER_28_2121 ();
 sg13g2_fill_2 FILLER_28_2125 ();
 sg13g2_decap_8 FILLER_28_2180 ();
 sg13g2_fill_2 FILLER_28_2187 ();
 sg13g2_fill_1 FILLER_28_2189 ();
 sg13g2_decap_4 FILLER_28_2199 ();
 sg13g2_fill_1 FILLER_28_2217 ();
 sg13g2_fill_1 FILLER_28_2251 ();
 sg13g2_fill_2 FILLER_28_2261 ();
 sg13g2_decap_8 FILLER_28_2289 ();
 sg13g2_decap_8 FILLER_28_2296 ();
 sg13g2_decap_8 FILLER_28_2333 ();
 sg13g2_fill_2 FILLER_28_2340 ();
 sg13g2_fill_1 FILLER_28_2342 ();
 sg13g2_fill_2 FILLER_28_2347 ();
 sg13g2_fill_2 FILLER_28_2375 ();
 sg13g2_fill_1 FILLER_28_2377 ();
 sg13g2_fill_1 FILLER_28_2382 ();
 sg13g2_fill_1 FILLER_28_2387 ();
 sg13g2_fill_1 FILLER_28_2392 ();
 sg13g2_fill_1 FILLER_28_2413 ();
 sg13g2_fill_1 FILLER_28_2445 ();
 sg13g2_fill_2 FILLER_28_2476 ();
 sg13g2_fill_1 FILLER_28_2478 ();
 sg13g2_fill_1 FILLER_28_2489 ();
 sg13g2_fill_1 FILLER_28_2516 ();
 sg13g2_fill_2 FILLER_28_2521 ();
 sg13g2_fill_1 FILLER_28_2523 ();
 sg13g2_decap_4 FILLER_28_2533 ();
 sg13g2_fill_2 FILLER_28_2537 ();
 sg13g2_fill_1 FILLER_28_2587 ();
 sg13g2_fill_2 FILLER_28_2596 ();
 sg13g2_fill_2 FILLER_28_2667 ();
 sg13g2_fill_1 FILLER_28_2669 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_fill_1 FILLER_29_49 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_decap_8 FILLER_29_70 ();
 sg13g2_decap_8 FILLER_29_77 ();
 sg13g2_decap_8 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_91 ();
 sg13g2_decap_8 FILLER_29_98 ();
 sg13g2_decap_8 FILLER_29_105 ();
 sg13g2_decap_8 FILLER_29_112 ();
 sg13g2_decap_8 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_126 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_fill_1 FILLER_29_164 ();
 sg13g2_fill_2 FILLER_29_197 ();
 sg13g2_fill_1 FILLER_29_246 ();
 sg13g2_fill_1 FILLER_29_255 ();
 sg13g2_decap_8 FILLER_29_308 ();
 sg13g2_decap_8 FILLER_29_315 ();
 sg13g2_decap_8 FILLER_29_348 ();
 sg13g2_decap_8 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_29_435 ();
 sg13g2_decap_8 FILLER_29_442 ();
 sg13g2_decap_8 FILLER_29_449 ();
 sg13g2_decap_8 FILLER_29_456 ();
 sg13g2_decap_4 FILLER_29_463 ();
 sg13g2_fill_1 FILLER_29_467 ();
 sg13g2_fill_2 FILLER_29_498 ();
 sg13g2_fill_2 FILLER_29_505 ();
 sg13g2_fill_2 FILLER_29_528 ();
 sg13g2_fill_1 FILLER_29_530 ();
 sg13g2_decap_4 FILLER_29_536 ();
 sg13g2_fill_1 FILLER_29_540 ();
 sg13g2_fill_2 FILLER_29_579 ();
 sg13g2_decap_4 FILLER_29_586 ();
 sg13g2_fill_2 FILLER_29_602 ();
 sg13g2_fill_1 FILLER_29_604 ();
 sg13g2_fill_2 FILLER_29_615 ();
 sg13g2_fill_1 FILLER_29_656 ();
 sg13g2_fill_1 FILLER_29_666 ();
 sg13g2_decap_4 FILLER_29_681 ();
 sg13g2_fill_1 FILLER_29_685 ();
 sg13g2_decap_8 FILLER_29_696 ();
 sg13g2_fill_1 FILLER_29_703 ();
 sg13g2_fill_2 FILLER_29_716 ();
 sg13g2_fill_1 FILLER_29_718 ();
 sg13g2_fill_1 FILLER_29_724 ();
 sg13g2_decap_8 FILLER_29_729 ();
 sg13g2_decap_4 FILLER_29_736 ();
 sg13g2_fill_2 FILLER_29_740 ();
 sg13g2_fill_1 FILLER_29_773 ();
 sg13g2_fill_1 FILLER_29_818 ();
 sg13g2_fill_2 FILLER_29_832 ();
 sg13g2_fill_1 FILLER_29_842 ();
 sg13g2_fill_2 FILLER_29_851 ();
 sg13g2_fill_1 FILLER_29_886 ();
 sg13g2_decap_4 FILLER_29_897 ();
 sg13g2_fill_2 FILLER_29_907 ();
 sg13g2_fill_1 FILLER_29_909 ();
 sg13g2_fill_2 FILLER_29_915 ();
 sg13g2_fill_2 FILLER_29_943 ();
 sg13g2_fill_2 FILLER_29_989 ();
 sg13g2_fill_1 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_997 ();
 sg13g2_fill_2 FILLER_29_1004 ();
 sg13g2_decap_8 FILLER_29_1024 ();
 sg13g2_decap_8 FILLER_29_1031 ();
 sg13g2_decap_8 FILLER_29_1038 ();
 sg13g2_decap_4 FILLER_29_1045 ();
 sg13g2_fill_2 FILLER_29_1058 ();
 sg13g2_fill_1 FILLER_29_1094 ();
 sg13g2_fill_2 FILLER_29_1106 ();
 sg13g2_fill_1 FILLER_29_1108 ();
 sg13g2_decap_4 FILLER_29_1140 ();
 sg13g2_fill_2 FILLER_29_1144 ();
 sg13g2_fill_1 FILLER_29_1169 ();
 sg13g2_decap_4 FILLER_29_1184 ();
 sg13g2_fill_1 FILLER_29_1196 ();
 sg13g2_fill_2 FILLER_29_1202 ();
 sg13g2_decap_8 FILLER_29_1230 ();
 sg13g2_decap_8 FILLER_29_1237 ();
 sg13g2_fill_1 FILLER_29_1244 ();
 sg13g2_fill_2 FILLER_29_1255 ();
 sg13g2_fill_2 FILLER_29_1304 ();
 sg13g2_fill_1 FILLER_29_1311 ();
 sg13g2_fill_1 FILLER_29_1316 ();
 sg13g2_fill_2 FILLER_29_1323 ();
 sg13g2_fill_1 FILLER_29_1325 ();
 sg13g2_fill_2 FILLER_29_1331 ();
 sg13g2_decap_8 FILLER_29_1337 ();
 sg13g2_decap_8 FILLER_29_1344 ();
 sg13g2_fill_2 FILLER_29_1351 ();
 sg13g2_fill_1 FILLER_29_1353 ();
 sg13g2_decap_4 FILLER_29_1359 ();
 sg13g2_fill_1 FILLER_29_1363 ();
 sg13g2_fill_1 FILLER_29_1370 ();
 sg13g2_fill_1 FILLER_29_1379 ();
 sg13g2_decap_8 FILLER_29_1423 ();
 sg13g2_fill_2 FILLER_29_1430 ();
 sg13g2_fill_1 FILLER_29_1432 ();
 sg13g2_decap_8 FILLER_29_1448 ();
 sg13g2_fill_2 FILLER_29_1455 ();
 sg13g2_fill_1 FILLER_29_1457 ();
 sg13g2_fill_1 FILLER_29_1489 ();
 sg13g2_decap_8 FILLER_29_1535 ();
 sg13g2_decap_4 FILLER_29_1542 ();
 sg13g2_fill_1 FILLER_29_1546 ();
 sg13g2_decap_8 FILLER_29_1553 ();
 sg13g2_fill_2 FILLER_29_1560 ();
 sg13g2_fill_2 FILLER_29_1588 ();
 sg13g2_fill_2 FILLER_29_1607 ();
 sg13g2_fill_1 FILLER_29_1725 ();
 sg13g2_decap_8 FILLER_29_1731 ();
 sg13g2_fill_1 FILLER_29_1738 ();
 sg13g2_decap_4 FILLER_29_1743 ();
 sg13g2_fill_1 FILLER_29_1747 ();
 sg13g2_decap_8 FILLER_29_1752 ();
 sg13g2_decap_8 FILLER_29_1759 ();
 sg13g2_decap_8 FILLER_29_1766 ();
 sg13g2_decap_8 FILLER_29_1773 ();
 sg13g2_fill_2 FILLER_29_1780 ();
 sg13g2_decap_8 FILLER_29_1812 ();
 sg13g2_fill_2 FILLER_29_1862 ();
 sg13g2_fill_1 FILLER_29_1864 ();
 sg13g2_fill_2 FILLER_29_1887 ();
 sg13g2_decap_4 FILLER_29_1925 ();
 sg13g2_fill_2 FILLER_29_1929 ();
 sg13g2_fill_1 FILLER_29_1944 ();
 sg13g2_decap_4 FILLER_29_1972 ();
 sg13g2_fill_2 FILLER_29_1976 ();
 sg13g2_fill_2 FILLER_29_2004 ();
 sg13g2_fill_1 FILLER_29_2016 ();
 sg13g2_fill_2 FILLER_29_2022 ();
 sg13g2_decap_4 FILLER_29_2064 ();
 sg13g2_decap_4 FILLER_29_2072 ();
 sg13g2_fill_2 FILLER_29_2079 ();
 sg13g2_fill_2 FILLER_29_2086 ();
 sg13g2_fill_1 FILLER_29_2088 ();
 sg13g2_decap_4 FILLER_29_2133 ();
 sg13g2_fill_1 FILLER_29_2150 ();
 sg13g2_decap_8 FILLER_29_2157 ();
 sg13g2_decap_8 FILLER_29_2164 ();
 sg13g2_fill_2 FILLER_29_2171 ();
 sg13g2_fill_1 FILLER_29_2173 ();
 sg13g2_fill_2 FILLER_29_2225 ();
 sg13g2_fill_2 FILLER_29_2230 ();
 sg13g2_fill_2 FILLER_29_2285 ();
 sg13g2_fill_2 FILLER_29_2293 ();
 sg13g2_fill_1 FILLER_29_2295 ();
 sg13g2_decap_8 FILLER_29_2326 ();
 sg13g2_decap_4 FILLER_29_2333 ();
 sg13g2_fill_2 FILLER_29_2337 ();
 sg13g2_decap_8 FILLER_29_2343 ();
 sg13g2_decap_4 FILLER_29_2354 ();
 sg13g2_decap_8 FILLER_29_2362 ();
 sg13g2_decap_8 FILLER_29_2369 ();
 sg13g2_decap_8 FILLER_29_2376 ();
 sg13g2_fill_1 FILLER_29_2383 ();
 sg13g2_decap_4 FILLER_29_2388 ();
 sg13g2_fill_1 FILLER_29_2392 ();
 sg13g2_decap_8 FILLER_29_2398 ();
 sg13g2_decap_4 FILLER_29_2405 ();
 sg13g2_fill_1 FILLER_29_2409 ();
 sg13g2_fill_2 FILLER_29_2436 ();
 sg13g2_fill_2 FILLER_29_2459 ();
 sg13g2_fill_1 FILLER_29_2461 ();
 sg13g2_fill_2 FILLER_29_2510 ();
 sg13g2_decap_8 FILLER_29_2517 ();
 sg13g2_fill_2 FILLER_29_2524 ();
 sg13g2_fill_1 FILLER_29_2526 ();
 sg13g2_fill_1 FILLER_29_2535 ();
 sg13g2_fill_2 FILLER_29_2575 ();
 sg13g2_fill_2 FILLER_29_2599 ();
 sg13g2_fill_2 FILLER_29_2619 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_fill_2 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_53 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_decap_8 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_107 ();
 sg13g2_fill_2 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_116 ();
 sg13g2_fill_1 FILLER_30_158 ();
 sg13g2_fill_2 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_303 ();
 sg13g2_decap_8 FILLER_30_317 ();
 sg13g2_decap_4 FILLER_30_324 ();
 sg13g2_decap_8 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_339 ();
 sg13g2_decap_8 FILLER_30_346 ();
 sg13g2_decap_4 FILLER_30_353 ();
 sg13g2_fill_1 FILLER_30_357 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_decap_4 FILLER_30_376 ();
 sg13g2_fill_1 FILLER_30_380 ();
 sg13g2_decap_4 FILLER_30_389 ();
 sg13g2_fill_1 FILLER_30_393 ();
 sg13g2_fill_2 FILLER_30_397 ();
 sg13g2_fill_1 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_447 ();
 sg13g2_decap_8 FILLER_30_454 ();
 sg13g2_fill_2 FILLER_30_461 ();
 sg13g2_fill_1 FILLER_30_463 ();
 sg13g2_fill_1 FILLER_30_472 ();
 sg13g2_fill_2 FILLER_30_480 ();
 sg13g2_fill_2 FILLER_30_485 ();
 sg13g2_fill_2 FILLER_30_492 ();
 sg13g2_fill_2 FILLER_30_498 ();
 sg13g2_fill_1 FILLER_30_500 ();
 sg13g2_fill_1 FILLER_30_505 ();
 sg13g2_decap_8 FILLER_30_510 ();
 sg13g2_decap_8 FILLER_30_517 ();
 sg13g2_decap_4 FILLER_30_524 ();
 sg13g2_fill_1 FILLER_30_528 ();
 sg13g2_decap_8 FILLER_30_542 ();
 sg13g2_decap_8 FILLER_30_549 ();
 sg13g2_decap_4 FILLER_30_566 ();
 sg13g2_fill_2 FILLER_30_575 ();
 sg13g2_decap_4 FILLER_30_601 ();
 sg13g2_fill_1 FILLER_30_627 ();
 sg13g2_fill_1 FILLER_30_646 ();
 sg13g2_decap_8 FILLER_30_678 ();
 sg13g2_decap_4 FILLER_30_685 ();
 sg13g2_fill_1 FILLER_30_689 ();
 sg13g2_fill_1 FILLER_30_698 ();
 sg13g2_fill_2 FILLER_30_708 ();
 sg13g2_fill_1 FILLER_30_710 ();
 sg13g2_fill_2 FILLER_30_733 ();
 sg13g2_decap_4 FILLER_30_745 ();
 sg13g2_fill_1 FILLER_30_749 ();
 sg13g2_fill_2 FILLER_30_818 ();
 sg13g2_fill_1 FILLER_30_820 ();
 sg13g2_fill_1 FILLER_30_847 ();
 sg13g2_fill_2 FILLER_30_855 ();
 sg13g2_fill_1 FILLER_30_862 ();
 sg13g2_fill_2 FILLER_30_867 ();
 sg13g2_fill_2 FILLER_30_877 ();
 sg13g2_fill_1 FILLER_30_879 ();
 sg13g2_fill_2 FILLER_30_901 ();
 sg13g2_fill_1 FILLER_30_903 ();
 sg13g2_fill_1 FILLER_30_913 ();
 sg13g2_decap_8 FILLER_30_919 ();
 sg13g2_fill_1 FILLER_30_936 ();
 sg13g2_fill_2 FILLER_30_941 ();
 sg13g2_fill_1 FILLER_30_951 ();
 sg13g2_decap_4 FILLER_30_963 ();
 sg13g2_fill_2 FILLER_30_972 ();
 sg13g2_fill_1 FILLER_30_974 ();
 sg13g2_decap_8 FILLER_30_979 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_fill_2 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1027 ();
 sg13g2_fill_2 FILLER_30_1034 ();
 sg13g2_decap_4 FILLER_30_1040 ();
 sg13g2_fill_1 FILLER_30_1044 ();
 sg13g2_fill_1 FILLER_30_1056 ();
 sg13g2_fill_2 FILLER_30_1061 ();
 sg13g2_fill_1 FILLER_30_1068 ();
 sg13g2_fill_2 FILLER_30_1095 ();
 sg13g2_fill_2 FILLER_30_1102 ();
 sg13g2_decap_8 FILLER_30_1118 ();
 sg13g2_decap_8 FILLER_30_1125 ();
 sg13g2_fill_1 FILLER_30_1136 ();
 sg13g2_fill_2 FILLER_30_1152 ();
 sg13g2_fill_2 FILLER_30_1159 ();
 sg13g2_fill_2 FILLER_30_1166 ();
 sg13g2_decap_4 FILLER_30_1173 ();
 sg13g2_fill_2 FILLER_30_1177 ();
 sg13g2_decap_4 FILLER_30_1190 ();
 sg13g2_fill_2 FILLER_30_1214 ();
 sg13g2_fill_1 FILLER_30_1216 ();
 sg13g2_fill_1 FILLER_30_1222 ();
 sg13g2_fill_1 FILLER_30_1232 ();
 sg13g2_decap_8 FILLER_30_1259 ();
 sg13g2_fill_2 FILLER_30_1266 ();
 sg13g2_fill_1 FILLER_30_1268 ();
 sg13g2_fill_1 FILLER_30_1277 ();
 sg13g2_fill_1 FILLER_30_1308 ();
 sg13g2_fill_1 FILLER_30_1320 ();
 sg13g2_decap_8 FILLER_30_1351 ();
 sg13g2_decap_8 FILLER_30_1358 ();
 sg13g2_decap_8 FILLER_30_1365 ();
 sg13g2_fill_2 FILLER_30_1372 ();
 sg13g2_fill_1 FILLER_30_1374 ();
 sg13g2_decap_4 FILLER_30_1379 ();
 sg13g2_fill_2 FILLER_30_1383 ();
 sg13g2_decap_8 FILLER_30_1389 ();
 sg13g2_decap_8 FILLER_30_1396 ();
 sg13g2_decap_8 FILLER_30_1403 ();
 sg13g2_fill_2 FILLER_30_1410 ();
 sg13g2_fill_1 FILLER_30_1412 ();
 sg13g2_fill_2 FILLER_30_1419 ();
 sg13g2_decap_8 FILLER_30_1430 ();
 sg13g2_decap_8 FILLER_30_1437 ();
 sg13g2_decap_8 FILLER_30_1444 ();
 sg13g2_decap_8 FILLER_30_1451 ();
 sg13g2_fill_1 FILLER_30_1478 ();
 sg13g2_fill_1 FILLER_30_1490 ();
 sg13g2_fill_1 FILLER_30_1540 ();
 sg13g2_fill_2 FILLER_30_1546 ();
 sg13g2_fill_2 FILLER_30_1554 ();
 sg13g2_fill_1 FILLER_30_1556 ();
 sg13g2_decap_4 FILLER_30_1567 ();
 sg13g2_fill_2 FILLER_30_1571 ();
 sg13g2_decap_4 FILLER_30_1582 ();
 sg13g2_fill_1 FILLER_30_1586 ();
 sg13g2_fill_2 FILLER_30_1625 ();
 sg13g2_decap_8 FILLER_30_1636 ();
 sg13g2_decap_8 FILLER_30_1643 ();
 sg13g2_fill_2 FILLER_30_1650 ();
 sg13g2_fill_1 FILLER_30_1661 ();
 sg13g2_fill_1 FILLER_30_1672 ();
 sg13g2_decap_4 FILLER_30_1735 ();
 sg13g2_fill_2 FILLER_30_1747 ();
 sg13g2_decap_8 FILLER_30_1783 ();
 sg13g2_decap_4 FILLER_30_1790 ();
 sg13g2_fill_1 FILLER_30_1794 ();
 sg13g2_decap_8 FILLER_30_1798 ();
 sg13g2_decap_8 FILLER_30_1805 ();
 sg13g2_fill_2 FILLER_30_1812 ();
 sg13g2_fill_1 FILLER_30_1819 ();
 sg13g2_fill_2 FILLER_30_1830 ();
 sg13g2_decap_4 FILLER_30_1842 ();
 sg13g2_decap_8 FILLER_30_1904 ();
 sg13g2_decap_8 FILLER_30_1911 ();
 sg13g2_decap_4 FILLER_30_1918 ();
 sg13g2_fill_2 FILLER_30_1922 ();
 sg13g2_decap_4 FILLER_30_1958 ();
 sg13g2_fill_1 FILLER_30_1962 ();
 sg13g2_fill_2 FILLER_30_1973 ();
 sg13g2_fill_1 FILLER_30_1975 ();
 sg13g2_decap_4 FILLER_30_1981 ();
 sg13g2_fill_1 FILLER_30_1985 ();
 sg13g2_decap_4 FILLER_30_1990 ();
 sg13g2_decap_8 FILLER_30_1999 ();
 sg13g2_fill_2 FILLER_30_2006 ();
 sg13g2_fill_1 FILLER_30_2008 ();
 sg13g2_decap_8 FILLER_30_2019 ();
 sg13g2_decap_4 FILLER_30_2026 ();
 sg13g2_fill_2 FILLER_30_2030 ();
 sg13g2_fill_2 FILLER_30_2041 ();
 sg13g2_decap_8 FILLER_30_2046 ();
 sg13g2_decap_4 FILLER_30_2053 ();
 sg13g2_decap_8 FILLER_30_2065 ();
 sg13g2_decap_4 FILLER_30_2072 ();
 sg13g2_fill_1 FILLER_30_2076 ();
 sg13g2_decap_8 FILLER_30_2083 ();
 sg13g2_decap_8 FILLER_30_2090 ();
 sg13g2_fill_2 FILLER_30_2097 ();
 sg13g2_fill_1 FILLER_30_2099 ();
 sg13g2_fill_2 FILLER_30_2135 ();
 sg13g2_fill_1 FILLER_30_2137 ();
 sg13g2_decap_8 FILLER_30_2143 ();
 sg13g2_decap_8 FILLER_30_2150 ();
 sg13g2_decap_8 FILLER_30_2157 ();
 sg13g2_decap_8 FILLER_30_2164 ();
 sg13g2_decap_4 FILLER_30_2171 ();
 sg13g2_decap_8 FILLER_30_2216 ();
 sg13g2_decap_4 FILLER_30_2223 ();
 sg13g2_fill_2 FILLER_30_2241 ();
 sg13g2_decap_8 FILLER_30_2297 ();
 sg13g2_decap_8 FILLER_30_2304 ();
 sg13g2_decap_8 FILLER_30_2311 ();
 sg13g2_decap_8 FILLER_30_2318 ();
 sg13g2_decap_8 FILLER_30_2325 ();
 sg13g2_fill_2 FILLER_30_2340 ();
 sg13g2_fill_1 FILLER_30_2342 ();
 sg13g2_fill_2 FILLER_30_2369 ();
 sg13g2_fill_2 FILLER_30_2384 ();
 sg13g2_fill_1 FILLER_30_2386 ();
 sg13g2_fill_1 FILLER_30_2400 ();
 sg13g2_decap_8 FILLER_30_2420 ();
 sg13g2_fill_2 FILLER_30_2427 ();
 sg13g2_fill_1 FILLER_30_2429 ();
 sg13g2_decap_4 FILLER_30_2434 ();
 sg13g2_fill_1 FILLER_30_2438 ();
 sg13g2_decap_8 FILLER_30_2444 ();
 sg13g2_decap_8 FILLER_30_2451 ();
 sg13g2_decap_4 FILLER_30_2466 ();
 sg13g2_fill_2 FILLER_30_2470 ();
 sg13g2_decap_4 FILLER_30_2476 ();
 sg13g2_fill_2 FILLER_30_2484 ();
 sg13g2_fill_1 FILLER_30_2486 ();
 sg13g2_fill_2 FILLER_30_2518 ();
 sg13g2_fill_2 FILLER_30_2590 ();
 sg13g2_fill_2 FILLER_30_2622 ();
 sg13g2_decap_8 FILLER_30_2663 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_2 FILLER_31_11 ();
 sg13g2_fill_2 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_55 ();
 sg13g2_decap_8 FILLER_31_62 ();
 sg13g2_decap_8 FILLER_31_69 ();
 sg13g2_decap_4 FILLER_31_76 ();
 sg13g2_fill_1 FILLER_31_80 ();
 sg13g2_fill_1 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_1 FILLER_31_141 ();
 sg13g2_fill_2 FILLER_31_163 ();
 sg13g2_fill_1 FILLER_31_165 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_decap_8 FILLER_31_177 ();
 sg13g2_decap_8 FILLER_31_184 ();
 sg13g2_fill_2 FILLER_31_191 ();
 sg13g2_fill_2 FILLER_31_196 ();
 sg13g2_fill_1 FILLER_31_228 ();
 sg13g2_fill_1 FILLER_31_274 ();
 sg13g2_fill_1 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_311 ();
 sg13g2_decap_8 FILLER_31_318 ();
 sg13g2_decap_8 FILLER_31_325 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_1 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_380 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_4 FILLER_31_401 ();
 sg13g2_fill_2 FILLER_31_405 ();
 sg13g2_decap_8 FILLER_31_424 ();
 sg13g2_decap_8 FILLER_31_431 ();
 sg13g2_decap_8 FILLER_31_438 ();
 sg13g2_fill_2 FILLER_31_445 ();
 sg13g2_fill_1 FILLER_31_447 ();
 sg13g2_decap_8 FILLER_31_453 ();
 sg13g2_decap_8 FILLER_31_460 ();
 sg13g2_decap_8 FILLER_31_467 ();
 sg13g2_decap_8 FILLER_31_474 ();
 sg13g2_fill_1 FILLER_31_481 ();
 sg13g2_decap_8 FILLER_31_491 ();
 sg13g2_decap_4 FILLER_31_498 ();
 sg13g2_decap_8 FILLER_31_507 ();
 sg13g2_fill_2 FILLER_31_514 ();
 sg13g2_fill_1 FILLER_31_516 ();
 sg13g2_fill_2 FILLER_31_521 ();
 sg13g2_decap_8 FILLER_31_528 ();
 sg13g2_decap_4 FILLER_31_535 ();
 sg13g2_fill_2 FILLER_31_539 ();
 sg13g2_fill_2 FILLER_31_544 ();
 sg13g2_fill_1 FILLER_31_546 ();
 sg13g2_fill_1 FILLER_31_552 ();
 sg13g2_decap_4 FILLER_31_567 ();
 sg13g2_fill_1 FILLER_31_571 ();
 sg13g2_fill_2 FILLER_31_626 ();
 sg13g2_fill_1 FILLER_31_641 ();
 sg13g2_fill_1 FILLER_31_709 ();
 sg13g2_fill_2 FILLER_31_736 ();
 sg13g2_fill_1 FILLER_31_738 ();
 sg13g2_decap_8 FILLER_31_744 ();
 sg13g2_decap_8 FILLER_31_751 ();
 sg13g2_fill_2 FILLER_31_758 ();
 sg13g2_fill_2 FILLER_31_781 ();
 sg13g2_fill_1 FILLER_31_783 ();
 sg13g2_decap_4 FILLER_31_824 ();
 sg13g2_fill_1 FILLER_31_841 ();
 sg13g2_decap_4 FILLER_31_866 ();
 sg13g2_fill_1 FILLER_31_886 ();
 sg13g2_fill_2 FILLER_31_919 ();
 sg13g2_decap_8 FILLER_31_950 ();
 sg13g2_decap_4 FILLER_31_983 ();
 sg13g2_fill_2 FILLER_31_987 ();
 sg13g2_fill_2 FILLER_31_997 ();
 sg13g2_fill_2 FILLER_31_1012 ();
 sg13g2_fill_1 FILLER_31_1014 ();
 sg13g2_fill_2 FILLER_31_1019 ();
 sg13g2_fill_1 FILLER_31_1021 ();
 sg13g2_decap_4 FILLER_31_1034 ();
 sg13g2_fill_2 FILLER_31_1038 ();
 sg13g2_fill_1 FILLER_31_1044 ();
 sg13g2_fill_1 FILLER_31_1092 ();
 sg13g2_fill_2 FILLER_31_1119 ();
 sg13g2_fill_2 FILLER_31_1126 ();
 sg13g2_fill_1 FILLER_31_1128 ();
 sg13g2_decap_4 FILLER_31_1135 ();
 sg13g2_decap_4 FILLER_31_1144 ();
 sg13g2_fill_2 FILLER_31_1193 ();
 sg13g2_decap_4 FILLER_31_1221 ();
 sg13g2_decap_4 FILLER_31_1230 ();
 sg13g2_fill_1 FILLER_31_1239 ();
 sg13g2_fill_2 FILLER_31_1283 ();
 sg13g2_fill_1 FILLER_31_1285 ();
 sg13g2_decap_8 FILLER_31_1295 ();
 sg13g2_decap_8 FILLER_31_1302 ();
 sg13g2_decap_8 FILLER_31_1309 ();
 sg13g2_decap_8 FILLER_31_1320 ();
 sg13g2_decap_8 FILLER_31_1327 ();
 sg13g2_decap_4 FILLER_31_1334 ();
 sg13g2_fill_2 FILLER_31_1369 ();
 sg13g2_fill_1 FILLER_31_1371 ();
 sg13g2_fill_2 FILLER_31_1381 ();
 sg13g2_fill_1 FILLER_31_1383 ();
 sg13g2_fill_2 FILLER_31_1398 ();
 sg13g2_fill_1 FILLER_31_1400 ();
 sg13g2_fill_1 FILLER_31_1406 ();
 sg13g2_decap_8 FILLER_31_1433 ();
 sg13g2_fill_1 FILLER_31_1440 ();
 sg13g2_decap_8 FILLER_31_1446 ();
 sg13g2_decap_4 FILLER_31_1453 ();
 sg13g2_fill_2 FILLER_31_1457 ();
 sg13g2_decap_4 FILLER_31_1468 ();
 sg13g2_decap_8 FILLER_31_1503 ();
 sg13g2_decap_8 FILLER_31_1510 ();
 sg13g2_fill_1 FILLER_31_1517 ();
 sg13g2_fill_2 FILLER_31_1524 ();
 sg13g2_fill_1 FILLER_31_1526 ();
 sg13g2_decap_8 FILLER_31_1540 ();
 sg13g2_decap_8 FILLER_31_1547 ();
 sg13g2_decap_8 FILLER_31_1554 ();
 sg13g2_decap_8 FILLER_31_1561 ();
 sg13g2_decap_8 FILLER_31_1568 ();
 sg13g2_fill_2 FILLER_31_1575 ();
 sg13g2_fill_1 FILLER_31_1577 ();
 sg13g2_decap_8 FILLER_31_1591 ();
 sg13g2_decap_4 FILLER_31_1602 ();
 sg13g2_fill_1 FILLER_31_1606 ();
 sg13g2_fill_2 FILLER_31_1615 ();
 sg13g2_decap_8 FILLER_31_1643 ();
 sg13g2_decap_4 FILLER_31_1650 ();
 sg13g2_fill_2 FILLER_31_1654 ();
 sg13g2_fill_1 FILLER_31_1679 ();
 sg13g2_fill_1 FILLER_31_1683 ();
 sg13g2_fill_2 FILLER_31_1689 ();
 sg13g2_decap_4 FILLER_31_1723 ();
 sg13g2_fill_1 FILLER_31_1727 ();
 sg13g2_decap_4 FILLER_31_1785 ();
 sg13g2_fill_2 FILLER_31_1800 ();
 sg13g2_decap_8 FILLER_31_1806 ();
 sg13g2_decap_8 FILLER_31_1813 ();
 sg13g2_decap_8 FILLER_31_1820 ();
 sg13g2_decap_8 FILLER_31_1827 ();
 sg13g2_decap_8 FILLER_31_1834 ();
 sg13g2_decap_8 FILLER_31_1841 ();
 sg13g2_decap_8 FILLER_31_1848 ();
 sg13g2_decap_4 FILLER_31_1855 ();
 sg13g2_fill_2 FILLER_31_1859 ();
 sg13g2_decap_8 FILLER_31_1865 ();
 sg13g2_decap_8 FILLER_31_1872 ();
 sg13g2_decap_4 FILLER_31_1879 ();
 sg13g2_fill_1 FILLER_31_1883 ();
 sg13g2_decap_8 FILLER_31_1925 ();
 sg13g2_fill_2 FILLER_31_1932 ();
 sg13g2_decap_8 FILLER_31_1940 ();
 sg13g2_fill_2 FILLER_31_1947 ();
 sg13g2_fill_1 FILLER_31_1949 ();
 sg13g2_fill_1 FILLER_31_1990 ();
 sg13g2_decap_8 FILLER_31_1999 ();
 sg13g2_fill_2 FILLER_31_2006 ();
 sg13g2_fill_1 FILLER_31_2008 ();
 sg13g2_fill_2 FILLER_31_2014 ();
 sg13g2_fill_2 FILLER_31_2049 ();
 sg13g2_decap_8 FILLER_31_2103 ();
 sg13g2_decap_8 FILLER_31_2110 ();
 sg13g2_decap_4 FILLER_31_2117 ();
 sg13g2_fill_2 FILLER_31_2121 ();
 sg13g2_fill_1 FILLER_31_2133 ();
 sg13g2_decap_4 FILLER_31_2142 ();
 sg13g2_fill_2 FILLER_31_2172 ();
 sg13g2_decap_4 FILLER_31_2180 ();
 sg13g2_decap_8 FILLER_31_2200 ();
 sg13g2_fill_2 FILLER_31_2219 ();
 sg13g2_fill_2 FILLER_31_2230 ();
 sg13g2_decap_4 FILLER_31_2236 ();
 sg13g2_fill_1 FILLER_31_2240 ();
 sg13g2_fill_2 FILLER_31_2276 ();
 sg13g2_fill_1 FILLER_31_2278 ();
 sg13g2_fill_1 FILLER_31_2287 ();
 sg13g2_decap_8 FILLER_31_2294 ();
 sg13g2_fill_2 FILLER_31_2301 ();
 sg13g2_decap_4 FILLER_31_2359 ();
 sg13g2_fill_2 FILLER_31_2363 ();
 sg13g2_fill_2 FILLER_31_2371 ();
 sg13g2_fill_1 FILLER_31_2373 ();
 sg13g2_fill_1 FILLER_31_2400 ();
 sg13g2_fill_2 FILLER_31_2406 ();
 sg13g2_fill_1 FILLER_31_2408 ();
 sg13g2_decap_8 FILLER_31_2415 ();
 sg13g2_decap_8 FILLER_31_2422 ();
 sg13g2_decap_8 FILLER_31_2429 ();
 sg13g2_decap_8 FILLER_31_2436 ();
 sg13g2_decap_8 FILLER_31_2443 ();
 sg13g2_fill_1 FILLER_31_2450 ();
 sg13g2_fill_2 FILLER_31_2485 ();
 sg13g2_fill_1 FILLER_31_2500 ();
 sg13g2_decap_8 FILLER_31_2505 ();
 sg13g2_decap_8 FILLER_31_2512 ();
 sg13g2_decap_8 FILLER_31_2519 ();
 sg13g2_decap_4 FILLER_31_2526 ();
 sg13g2_fill_1 FILLER_31_2530 ();
 sg13g2_decap_8 FILLER_31_2539 ();
 sg13g2_decap_8 FILLER_31_2546 ();
 sg13g2_decap_8 FILLER_31_2553 ();
 sg13g2_decap_8 FILLER_31_2560 ();
 sg13g2_decap_4 FILLER_31_2567 ();
 sg13g2_fill_1 FILLER_31_2575 ();
 sg13g2_decap_4 FILLER_31_2580 ();
 sg13g2_fill_2 FILLER_31_2584 ();
 sg13g2_fill_1 FILLER_31_2631 ();
 sg13g2_fill_2 FILLER_31_2639 ();
 sg13g2_fill_1 FILLER_31_2641 ();
 sg13g2_decap_4 FILLER_31_2645 ();
 sg13g2_decap_8 FILLER_31_2653 ();
 sg13g2_decap_8 FILLER_31_2660 ();
 sg13g2_fill_2 FILLER_31_2667 ();
 sg13g2_fill_1 FILLER_31_2669 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_7 ();
 sg13g2_fill_1 FILLER_32_9 ();
 sg13g2_fill_1 FILLER_32_44 ();
 sg13g2_fill_2 FILLER_32_58 ();
 sg13g2_fill_1 FILLER_32_110 ();
 sg13g2_decap_4 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_1 FILLER_32_153 ();
 sg13g2_decap_8 FILLER_32_159 ();
 sg13g2_decap_8 FILLER_32_166 ();
 sg13g2_decap_8 FILLER_32_173 ();
 sg13g2_decap_4 FILLER_32_180 ();
 sg13g2_fill_1 FILLER_32_184 ();
 sg13g2_decap_8 FILLER_32_189 ();
 sg13g2_decap_4 FILLER_32_196 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_fill_1 FILLER_32_236 ();
 sg13g2_fill_1 FILLER_32_288 ();
 sg13g2_fill_2 FILLER_32_295 ();
 sg13g2_decap_8 FILLER_32_323 ();
 sg13g2_decap_8 FILLER_32_330 ();
 sg13g2_decap_8 FILLER_32_337 ();
 sg13g2_decap_8 FILLER_32_344 ();
 sg13g2_decap_4 FILLER_32_351 ();
 sg13g2_fill_1 FILLER_32_358 ();
 sg13g2_fill_2 FILLER_32_369 ();
 sg13g2_decap_4 FILLER_32_376 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_4 FILLER_32_396 ();
 sg13g2_fill_2 FILLER_32_400 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_413 ();
 sg13g2_fill_2 FILLER_32_442 ();
 sg13g2_fill_1 FILLER_32_444 ();
 sg13g2_fill_2 FILLER_32_450 ();
 sg13g2_fill_1 FILLER_32_452 ();
 sg13g2_fill_2 FILLER_32_463 ();
 sg13g2_fill_1 FILLER_32_465 ();
 sg13g2_fill_1 FILLER_32_478 ();
 sg13g2_decap_4 FILLER_32_484 ();
 sg13g2_fill_1 FILLER_32_502 ();
 sg13g2_fill_1 FILLER_32_508 ();
 sg13g2_fill_2 FILLER_32_528 ();
 sg13g2_decap_8 FILLER_32_548 ();
 sg13g2_decap_8 FILLER_32_555 ();
 sg13g2_decap_8 FILLER_32_562 ();
 sg13g2_fill_1 FILLER_32_574 ();
 sg13g2_fill_1 FILLER_32_586 ();
 sg13g2_fill_1 FILLER_32_592 ();
 sg13g2_fill_1 FILLER_32_597 ();
 sg13g2_fill_1 FILLER_32_603 ();
 sg13g2_fill_1 FILLER_32_609 ();
 sg13g2_fill_1 FILLER_32_615 ();
 sg13g2_fill_1 FILLER_32_620 ();
 sg13g2_fill_1 FILLER_32_629 ();
 sg13g2_fill_2 FILLER_32_634 ();
 sg13g2_fill_2 FILLER_32_640 ();
 sg13g2_fill_1 FILLER_32_653 ();
 sg13g2_fill_2 FILLER_32_657 ();
 sg13g2_fill_1 FILLER_32_667 ();
 sg13g2_fill_1 FILLER_32_735 ();
 sg13g2_decap_8 FILLER_32_745 ();
 sg13g2_decap_8 FILLER_32_752 ();
 sg13g2_decap_8 FILLER_32_759 ();
 sg13g2_decap_4 FILLER_32_766 ();
 sg13g2_decap_4 FILLER_32_781 ();
 sg13g2_fill_2 FILLER_32_794 ();
 sg13g2_fill_2 FILLER_32_801 ();
 sg13g2_fill_1 FILLER_32_803 ();
 sg13g2_fill_1 FILLER_32_809 ();
 sg13g2_decap_4 FILLER_32_816 ();
 sg13g2_fill_1 FILLER_32_820 ();
 sg13g2_decap_8 FILLER_32_861 ();
 sg13g2_fill_2 FILLER_32_868 ();
 sg13g2_fill_1 FILLER_32_875 ();
 sg13g2_fill_2 FILLER_32_915 ();
 sg13g2_fill_1 FILLER_32_917 ();
 sg13g2_fill_2 FILLER_32_926 ();
 sg13g2_fill_1 FILLER_32_931 ();
 sg13g2_decap_4 FILLER_32_942 ();
 sg13g2_decap_8 FILLER_32_950 ();
 sg13g2_fill_1 FILLER_32_957 ();
 sg13g2_decap_4 FILLER_32_968 ();
 sg13g2_fill_2 FILLER_32_1036 ();
 sg13g2_fill_1 FILLER_32_1038 ();
 sg13g2_decap_4 FILLER_32_1048 ();
 sg13g2_fill_2 FILLER_32_1052 ();
 sg13g2_decap_4 FILLER_32_1060 ();
 sg13g2_fill_1 FILLER_32_1068 ();
 sg13g2_decap_8 FILLER_32_1090 ();
 sg13g2_decap_8 FILLER_32_1097 ();
 sg13g2_decap_4 FILLER_32_1104 ();
 sg13g2_fill_1 FILLER_32_1108 ();
 sg13g2_fill_2 FILLER_32_1139 ();
 sg13g2_fill_1 FILLER_32_1141 ();
 sg13g2_decap_8 FILLER_32_1147 ();
 sg13g2_decap_8 FILLER_32_1157 ();
 sg13g2_decap_8 FILLER_32_1164 ();
 sg13g2_fill_2 FILLER_32_1171 ();
 sg13g2_fill_1 FILLER_32_1173 ();
 sg13g2_fill_1 FILLER_32_1214 ();
 sg13g2_fill_2 FILLER_32_1219 ();
 sg13g2_fill_1 FILLER_32_1221 ();
 sg13g2_decap_8 FILLER_32_1226 ();
 sg13g2_decap_8 FILLER_32_1233 ();
 sg13g2_decap_4 FILLER_32_1240 ();
 sg13g2_fill_2 FILLER_32_1244 ();
 sg13g2_decap_8 FILLER_32_1256 ();
 sg13g2_fill_2 FILLER_32_1263 ();
 sg13g2_fill_1 FILLER_32_1265 ();
 sg13g2_decap_8 FILLER_32_1338 ();
 sg13g2_decap_4 FILLER_32_1345 ();
 sg13g2_decap_4 FILLER_32_1355 ();
 sg13g2_fill_1 FILLER_32_1429 ();
 sg13g2_fill_2 FILLER_32_1456 ();
 sg13g2_decap_8 FILLER_32_1494 ();
 sg13g2_decap_8 FILLER_32_1501 ();
 sg13g2_fill_1 FILLER_32_1544 ();
 sg13g2_decap_8 FILLER_32_1548 ();
 sg13g2_decap_8 FILLER_32_1555 ();
 sg13g2_decap_8 FILLER_32_1562 ();
 sg13g2_decap_8 FILLER_32_1569 ();
 sg13g2_fill_2 FILLER_32_1576 ();
 sg13g2_fill_1 FILLER_32_1578 ();
 sg13g2_fill_2 FILLER_32_1589 ();
 sg13g2_fill_1 FILLER_32_1591 ();
 sg13g2_decap_4 FILLER_32_1595 ();
 sg13g2_fill_1 FILLER_32_1599 ();
 sg13g2_decap_8 FILLER_32_1603 ();
 sg13g2_fill_2 FILLER_32_1610 ();
 sg13g2_fill_2 FILLER_32_1635 ();
 sg13g2_fill_2 FILLER_32_1718 ();
 sg13g2_decap_8 FILLER_32_1733 ();
 sg13g2_decap_8 FILLER_32_1740 ();
 sg13g2_fill_2 FILLER_32_1747 ();
 sg13g2_decap_8 FILLER_32_1759 ();
 sg13g2_decap_8 FILLER_32_1766 ();
 sg13g2_decap_4 FILLER_32_1773 ();
 sg13g2_decap_8 FILLER_32_1808 ();
 sg13g2_decap_8 FILLER_32_1815 ();
 sg13g2_fill_1 FILLER_32_1822 ();
 sg13g2_decap_4 FILLER_32_1837 ();
 sg13g2_fill_1 FILLER_32_1841 ();
 sg13g2_fill_2 FILLER_32_1846 ();
 sg13g2_fill_1 FILLER_32_1848 ();
 sg13g2_decap_8 FILLER_32_1861 ();
 sg13g2_decap_8 FILLER_32_1868 ();
 sg13g2_decap_4 FILLER_32_1920 ();
 sg13g2_fill_1 FILLER_32_1924 ();
 sg13g2_decap_8 FILLER_32_1951 ();
 sg13g2_decap_8 FILLER_32_1958 ();
 sg13g2_fill_2 FILLER_32_2001 ();
 sg13g2_decap_8 FILLER_32_2009 ();
 sg13g2_fill_1 FILLER_32_2022 ();
 sg13g2_fill_1 FILLER_32_2028 ();
 sg13g2_decap_8 FILLER_32_2035 ();
 sg13g2_fill_1 FILLER_32_2042 ();
 sg13g2_decap_8 FILLER_32_2049 ();
 sg13g2_decap_4 FILLER_32_2064 ();
 sg13g2_fill_2 FILLER_32_2068 ();
 sg13g2_decap_8 FILLER_32_2074 ();
 sg13g2_decap_8 FILLER_32_2081 ();
 sg13g2_decap_8 FILLER_32_2091 ();
 sg13g2_decap_4 FILLER_32_2098 ();
 sg13g2_fill_2 FILLER_32_2111 ();
 sg13g2_fill_1 FILLER_32_2121 ();
 sg13g2_decap_8 FILLER_32_2148 ();
 sg13g2_decap_4 FILLER_32_2181 ();
 sg13g2_fill_1 FILLER_32_2185 ();
 sg13g2_fill_2 FILLER_32_2191 ();
 sg13g2_fill_1 FILLER_32_2193 ();
 sg13g2_decap_8 FILLER_32_2200 ();
 sg13g2_fill_2 FILLER_32_2207 ();
 sg13g2_fill_1 FILLER_32_2209 ();
 sg13g2_fill_2 FILLER_32_2237 ();
 sg13g2_fill_1 FILLER_32_2239 ();
 sg13g2_fill_2 FILLER_32_2259 ();
 sg13g2_fill_1 FILLER_32_2261 ();
 sg13g2_decap_4 FILLER_32_2267 ();
 sg13g2_fill_1 FILLER_32_2271 ();
 sg13g2_decap_8 FILLER_32_2286 ();
 sg13g2_decap_8 FILLER_32_2293 ();
 sg13g2_decap_4 FILLER_32_2314 ();
 sg13g2_fill_1 FILLER_32_2322 ();
 sg13g2_fill_1 FILLER_32_2327 ();
 sg13g2_fill_2 FILLER_32_2354 ();
 sg13g2_fill_1 FILLER_32_2356 ();
 sg13g2_fill_1 FILLER_32_2361 ();
 sg13g2_fill_1 FILLER_32_2423 ();
 sg13g2_decap_8 FILLER_32_2432 ();
 sg13g2_fill_2 FILLER_32_2449 ();
 sg13g2_fill_1 FILLER_32_2451 ();
 sg13g2_fill_1 FILLER_32_2504 ();
 sg13g2_fill_2 FILLER_32_2517 ();
 sg13g2_fill_1 FILLER_32_2519 ();
 sg13g2_decap_8 FILLER_32_2533 ();
 sg13g2_decap_8 FILLER_32_2540 ();
 sg13g2_decap_8 FILLER_32_2547 ();
 sg13g2_decap_8 FILLER_32_2554 ();
 sg13g2_decap_4 FILLER_32_2561 ();
 sg13g2_fill_1 FILLER_32_2599 ();
 sg13g2_decap_8 FILLER_32_2629 ();
 sg13g2_decap_8 FILLER_32_2636 ();
 sg13g2_decap_8 FILLER_32_2643 ();
 sg13g2_decap_8 FILLER_32_2650 ();
 sg13g2_decap_8 FILLER_32_2657 ();
 sg13g2_decap_4 FILLER_32_2664 ();
 sg13g2_fill_2 FILLER_32_2668 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_18 ();
 sg13g2_decap_4 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_29 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_fill_1 FILLER_33_53 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_fill_2 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_fill_1 FILLER_33_91 ();
 sg13g2_decap_4 FILLER_33_116 ();
 sg13g2_fill_1 FILLER_33_120 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_decap_8 FILLER_33_157 ();
 sg13g2_decap_8 FILLER_33_164 ();
 sg13g2_decap_8 FILLER_33_171 ();
 sg13g2_decap_8 FILLER_33_186 ();
 sg13g2_decap_8 FILLER_33_193 ();
 sg13g2_decap_8 FILLER_33_200 ();
 sg13g2_fill_1 FILLER_33_207 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_fill_1 FILLER_33_218 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_2 FILLER_33_295 ();
 sg13g2_fill_2 FILLER_33_305 ();
 sg13g2_fill_1 FILLER_33_307 ();
 sg13g2_fill_2 FILLER_33_321 ();
 sg13g2_fill_1 FILLER_33_323 ();
 sg13g2_decap_4 FILLER_33_333 ();
 sg13g2_fill_2 FILLER_33_337 ();
 sg13g2_decap_8 FILLER_33_347 ();
 sg13g2_decap_4 FILLER_33_354 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_387 ();
 sg13g2_fill_1 FILLER_33_391 ();
 sg13g2_decap_4 FILLER_33_400 ();
 sg13g2_fill_1 FILLER_33_419 ();
 sg13g2_fill_1 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_447 ();
 sg13g2_decap_8 FILLER_33_454 ();
 sg13g2_decap_8 FILLER_33_466 ();
 sg13g2_fill_2 FILLER_33_473 ();
 sg13g2_fill_1 FILLER_33_475 ();
 sg13g2_decap_4 FILLER_33_480 ();
 sg13g2_fill_2 FILLER_33_484 ();
 sg13g2_fill_2 FILLER_33_491 ();
 sg13g2_fill_1 FILLER_33_497 ();
 sg13g2_fill_2 FILLER_33_502 ();
 sg13g2_decap_8 FILLER_33_530 ();
 sg13g2_decap_8 FILLER_33_537 ();
 sg13g2_decap_8 FILLER_33_544 ();
 sg13g2_decap_8 FILLER_33_551 ();
 sg13g2_fill_1 FILLER_33_580 ();
 sg13g2_fill_1 FILLER_33_593 ();
 sg13g2_fill_2 FILLER_33_599 ();
 sg13g2_fill_1 FILLER_33_601 ();
 sg13g2_fill_1 FILLER_33_606 ();
 sg13g2_fill_2 FILLER_33_635 ();
 sg13g2_fill_1 FILLER_33_646 ();
 sg13g2_fill_1 FILLER_33_672 ();
 sg13g2_fill_1 FILLER_33_692 ();
 sg13g2_fill_2 FILLER_33_705 ();
 sg13g2_fill_1 FILLER_33_707 ();
 sg13g2_fill_2 FILLER_33_717 ();
 sg13g2_fill_1 FILLER_33_719 ();
 sg13g2_fill_2 FILLER_33_737 ();
 sg13g2_fill_1 FILLER_33_739 ();
 sg13g2_decap_8 FILLER_33_745 ();
 sg13g2_decap_8 FILLER_33_752 ();
 sg13g2_decap_8 FILLER_33_759 ();
 sg13g2_decap_8 FILLER_33_766 ();
 sg13g2_decap_8 FILLER_33_776 ();
 sg13g2_fill_2 FILLER_33_783 ();
 sg13g2_fill_1 FILLER_33_790 ();
 sg13g2_fill_2 FILLER_33_811 ();
 sg13g2_fill_1 FILLER_33_853 ();
 sg13g2_fill_2 FILLER_33_884 ();
 sg13g2_fill_1 FILLER_33_886 ();
 sg13g2_fill_1 FILLER_33_936 ();
 sg13g2_decap_8 FILLER_33_981 ();
 sg13g2_decap_4 FILLER_33_988 ();
 sg13g2_fill_2 FILLER_33_1003 ();
 sg13g2_decap_8 FILLER_33_1019 ();
 sg13g2_decap_8 FILLER_33_1026 ();
 sg13g2_decap_8 FILLER_33_1033 ();
 sg13g2_fill_2 FILLER_33_1048 ();
 sg13g2_fill_1 FILLER_33_1050 ();
 sg13g2_fill_2 FILLER_33_1062 ();
 sg13g2_fill_1 FILLER_33_1068 ();
 sg13g2_decap_8 FILLER_33_1084 ();
 sg13g2_decap_8 FILLER_33_1091 ();
 sg13g2_fill_2 FILLER_33_1098 ();
 sg13g2_fill_1 FILLER_33_1100 ();
 sg13g2_decap_4 FILLER_33_1142 ();
 sg13g2_fill_2 FILLER_33_1171 ();
 sg13g2_decap_8 FILLER_33_1209 ();
 sg13g2_decap_8 FILLER_33_1216 ();
 sg13g2_decap_8 FILLER_33_1223 ();
 sg13g2_fill_2 FILLER_33_1230 ();
 sg13g2_fill_1 FILLER_33_1246 ();
 sg13g2_decap_4 FILLER_33_1277 ();
 sg13g2_fill_1 FILLER_33_1281 ();
 sg13g2_decap_8 FILLER_33_1324 ();
 sg13g2_fill_1 FILLER_33_1336 ();
 sg13g2_decap_8 FILLER_33_1393 ();
 sg13g2_decap_8 FILLER_33_1400 ();
 sg13g2_decap_8 FILLER_33_1407 ();
 sg13g2_decap_8 FILLER_33_1420 ();
 sg13g2_fill_1 FILLER_33_1427 ();
 sg13g2_fill_2 FILLER_33_1438 ();
 sg13g2_fill_1 FILLER_33_1440 ();
 sg13g2_fill_2 FILLER_33_1467 ();
 sg13g2_decap_4 FILLER_33_1474 ();
 sg13g2_fill_2 FILLER_33_1504 ();
 sg13g2_decap_4 FILLER_33_1516 ();
 sg13g2_decap_8 FILLER_33_1526 ();
 sg13g2_decap_8 FILLER_33_1533 ();
 sg13g2_fill_1 FILLER_33_1544 ();
 sg13g2_fill_2 FILLER_33_1550 ();
 sg13g2_fill_1 FILLER_33_1552 ();
 sg13g2_decap_4 FILLER_33_1558 ();
 sg13g2_fill_1 FILLER_33_1566 ();
 sg13g2_fill_2 FILLER_33_1572 ();
 sg13g2_fill_1 FILLER_33_1574 ();
 sg13g2_fill_2 FILLER_33_1597 ();
 sg13g2_fill_1 FILLER_33_1599 ();
 sg13g2_decap_8 FILLER_33_1604 ();
 sg13g2_decap_4 FILLER_33_1611 ();
 sg13g2_fill_2 FILLER_33_1615 ();
 sg13g2_fill_1 FILLER_33_1622 ();
 sg13g2_fill_2 FILLER_33_1649 ();
 sg13g2_fill_1 FILLER_33_1651 ();
 sg13g2_decap_8 FILLER_33_1656 ();
 sg13g2_decap_4 FILLER_33_1663 ();
 sg13g2_fill_1 FILLER_33_1667 ();
 sg13g2_decap_8 FILLER_33_1681 ();
 sg13g2_decap_4 FILLER_33_1688 ();
 sg13g2_fill_1 FILLER_33_1692 ();
 sg13g2_decap_8 FILLER_33_1700 ();
 sg13g2_decap_4 FILLER_33_1707 ();
 sg13g2_fill_2 FILLER_33_1711 ();
 sg13g2_decap_8 FILLER_33_1764 ();
 sg13g2_fill_1 FILLER_33_1771 ();
 sg13g2_decap_8 FILLER_33_1806 ();
 sg13g2_fill_2 FILLER_33_1813 ();
 sg13g2_fill_1 FILLER_33_1815 ();
 sg13g2_fill_1 FILLER_33_1824 ();
 sg13g2_fill_1 FILLER_33_1833 ();
 sg13g2_fill_1 FILLER_33_1860 ();
 sg13g2_fill_2 FILLER_33_1865 ();
 sg13g2_fill_2 FILLER_33_1884 ();
 sg13g2_fill_1 FILLER_33_1886 ();
 sg13g2_fill_2 FILLER_33_1892 ();
 sg13g2_fill_2 FILLER_33_1898 ();
 sg13g2_fill_2 FILLER_33_1904 ();
 sg13g2_fill_1 FILLER_33_1906 ();
 sg13g2_decap_8 FILLER_33_1938 ();
 sg13g2_decap_8 FILLER_33_1945 ();
 sg13g2_fill_2 FILLER_33_1952 ();
 sg13g2_fill_1 FILLER_33_1982 ();
 sg13g2_fill_2 FILLER_33_2020 ();
 sg13g2_fill_2 FILLER_33_2032 ();
 sg13g2_fill_1 FILLER_33_2034 ();
 sg13g2_fill_2 FILLER_33_2059 ();
 sg13g2_fill_2 FILLER_33_2066 ();
 sg13g2_fill_1 FILLER_33_2073 ();
 sg13g2_fill_2 FILLER_33_2107 ();
 sg13g2_fill_1 FILLER_33_2109 ();
 sg13g2_fill_2 FILLER_33_2139 ();
 sg13g2_decap_8 FILLER_33_2163 ();
 sg13g2_decap_8 FILLER_33_2170 ();
 sg13g2_decap_8 FILLER_33_2177 ();
 sg13g2_decap_8 FILLER_33_2184 ();
 sg13g2_decap_8 FILLER_33_2191 ();
 sg13g2_decap_4 FILLER_33_2198 ();
 sg13g2_decap_8 FILLER_33_2207 ();
 sg13g2_decap_4 FILLER_33_2214 ();
 sg13g2_fill_2 FILLER_33_2244 ();
 sg13g2_fill_1 FILLER_33_2246 ();
 sg13g2_fill_2 FILLER_33_2253 ();
 sg13g2_decap_4 FILLER_33_2296 ();
 sg13g2_decap_8 FILLER_33_2359 ();
 sg13g2_fill_2 FILLER_33_2366 ();
 sg13g2_decap_8 FILLER_33_2372 ();
 sg13g2_fill_1 FILLER_33_2379 ();
 sg13g2_decap_8 FILLER_33_2388 ();
 sg13g2_fill_2 FILLER_33_2395 ();
 sg13g2_fill_1 FILLER_33_2431 ();
 sg13g2_decap_8 FILLER_33_2436 ();
 sg13g2_decap_4 FILLER_33_2443 ();
 sg13g2_fill_2 FILLER_33_2447 ();
 sg13g2_decap_4 FILLER_33_2453 ();
 sg13g2_fill_2 FILLER_33_2465 ();
 sg13g2_fill_1 FILLER_33_2467 ();
 sg13g2_fill_2 FILLER_33_2479 ();
 sg13g2_fill_2 FILLER_33_2528 ();
 sg13g2_fill_2 FILLER_33_2561 ();
 sg13g2_decap_8 FILLER_33_2567 ();
 sg13g2_decap_8 FILLER_33_2574 ();
 sg13g2_decap_8 FILLER_33_2581 ();
 sg13g2_decap_4 FILLER_33_2588 ();
 sg13g2_fill_1 FILLER_33_2592 ();
 sg13g2_decap_8 FILLER_33_2618 ();
 sg13g2_decap_8 FILLER_33_2625 ();
 sg13g2_decap_8 FILLER_33_2632 ();
 sg13g2_decap_8 FILLER_33_2639 ();
 sg13g2_decap_8 FILLER_33_2646 ();
 sg13g2_decap_8 FILLER_33_2653 ();
 sg13g2_decap_8 FILLER_33_2660 ();
 sg13g2_fill_2 FILLER_33_2667 ();
 sg13g2_fill_1 FILLER_33_2669 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_4 FILLER_34_7 ();
 sg13g2_fill_1 FILLER_34_11 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_decap_4 FILLER_34_94 ();
 sg13g2_fill_1 FILLER_34_98 ();
 sg13g2_decap_4 FILLER_34_125 ();
 sg13g2_fill_1 FILLER_34_129 ();
 sg13g2_decap_8 FILLER_34_152 ();
 sg13g2_decap_8 FILLER_34_159 ();
 sg13g2_decap_8 FILLER_34_166 ();
 sg13g2_decap_4 FILLER_34_199 ();
 sg13g2_fill_2 FILLER_34_233 ();
 sg13g2_fill_1 FILLER_34_241 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_4 FILLER_34_298 ();
 sg13g2_fill_2 FILLER_34_302 ();
 sg13g2_decap_8 FILLER_34_308 ();
 sg13g2_decap_8 FILLER_34_315 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_fill_2 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_4 FILLER_34_357 ();
 sg13g2_fill_2 FILLER_34_361 ();
 sg13g2_fill_2 FILLER_34_376 ();
 sg13g2_decap_4 FILLER_34_413 ();
 sg13g2_fill_2 FILLER_34_417 ();
 sg13g2_fill_2 FILLER_34_433 ();
 sg13g2_fill_1 FILLER_34_440 ();
 sg13g2_decap_8 FILLER_34_447 ();
 sg13g2_fill_2 FILLER_34_463 ();
 sg13g2_decap_8 FILLER_34_470 ();
 sg13g2_decap_8 FILLER_34_477 ();
 sg13g2_decap_8 FILLER_34_484 ();
 sg13g2_decap_8 FILLER_34_491 ();
 sg13g2_fill_1 FILLER_34_518 ();
 sg13g2_fill_2 FILLER_34_525 ();
 sg13g2_fill_2 FILLER_34_538 ();
 sg13g2_fill_1 FILLER_34_540 ();
 sg13g2_fill_2 FILLER_34_575 ();
 sg13g2_fill_1 FILLER_34_577 ();
 sg13g2_fill_1 FILLER_34_586 ();
 sg13g2_fill_1 FILLER_34_592 ();
 sg13g2_decap_4 FILLER_34_608 ();
 sg13g2_fill_1 FILLER_34_612 ();
 sg13g2_fill_2 FILLER_34_617 ();
 sg13g2_fill_2 FILLER_34_652 ();
 sg13g2_fill_2 FILLER_34_675 ();
 sg13g2_decap_8 FILLER_34_692 ();
 sg13g2_decap_8 FILLER_34_699 ();
 sg13g2_fill_2 FILLER_34_706 ();
 sg13g2_fill_2 FILLER_34_712 ();
 sg13g2_decap_8 FILLER_34_741 ();
 sg13g2_decap_8 FILLER_34_748 ();
 sg13g2_decap_8 FILLER_34_755 ();
 sg13g2_decap_8 FILLER_34_762 ();
 sg13g2_decap_4 FILLER_34_769 ();
 sg13g2_fill_2 FILLER_34_806 ();
 sg13g2_fill_2 FILLER_34_826 ();
 sg13g2_fill_2 FILLER_34_832 ();
 sg13g2_fill_2 FILLER_34_843 ();
 sg13g2_decap_8 FILLER_34_849 ();
 sg13g2_decap_8 FILLER_34_856 ();
 sg13g2_decap_4 FILLER_34_863 ();
 sg13g2_fill_2 FILLER_34_871 ();
 sg13g2_fill_1 FILLER_34_873 ();
 sg13g2_fill_1 FILLER_34_900 ();
 sg13g2_fill_2 FILLER_34_931 ();
 sg13g2_fill_1 FILLER_34_933 ();
 sg13g2_fill_1 FILLER_34_939 ();
 sg13g2_fill_1 FILLER_34_944 ();
 sg13g2_fill_1 FILLER_34_971 ();
 sg13g2_decap_8 FILLER_34_977 ();
 sg13g2_decap_8 FILLER_34_984 ();
 sg13g2_decap_4 FILLER_34_991 ();
 sg13g2_decap_4 FILLER_34_999 ();
 sg13g2_decap_4 FILLER_34_1012 ();
 sg13g2_decap_8 FILLER_34_1025 ();
 sg13g2_decap_8 FILLER_34_1032 ();
 sg13g2_decap_8 FILLER_34_1039 ();
 sg13g2_decap_8 FILLER_34_1046 ();
 sg13g2_fill_1 FILLER_34_1053 ();
 sg13g2_fill_2 FILLER_34_1057 ();
 sg13g2_fill_2 FILLER_34_1064 ();
 sg13g2_decap_8 FILLER_34_1070 ();
 sg13g2_decap_8 FILLER_34_1077 ();
 sg13g2_decap_8 FILLER_34_1084 ();
 sg13g2_decap_8 FILLER_34_1091 ();
 sg13g2_fill_2 FILLER_34_1118 ();
 sg13g2_decap_8 FILLER_34_1156 ();
 sg13g2_fill_1 FILLER_34_1163 ();
 sg13g2_fill_1 FILLER_34_1167 ();
 sg13g2_fill_2 FILLER_34_1182 ();
 sg13g2_fill_1 FILLER_34_1184 ();
 sg13g2_decap_4 FILLER_34_1194 ();
 sg13g2_fill_2 FILLER_34_1198 ();
 sg13g2_fill_2 FILLER_34_1205 ();
 sg13g2_decap_8 FILLER_34_1211 ();
 sg13g2_fill_1 FILLER_34_1218 ();
 sg13g2_decap_4 FILLER_34_1224 ();
 sg13g2_decap_8 FILLER_34_1270 ();
 sg13g2_decap_8 FILLER_34_1277 ();
 sg13g2_fill_2 FILLER_34_1284 ();
 sg13g2_fill_1 FILLER_34_1286 ();
 sg13g2_decap_4 FILLER_34_1292 ();
 sg13g2_fill_2 FILLER_34_1309 ();
 sg13g2_fill_2 FILLER_34_1316 ();
 sg13g2_fill_1 FILLER_34_1318 ();
 sg13g2_decap_4 FILLER_34_1323 ();
 sg13g2_fill_2 FILLER_34_1327 ();
 sg13g2_decap_8 FILLER_34_1337 ();
 sg13g2_fill_1 FILLER_34_1344 ();
 sg13g2_decap_8 FILLER_34_1348 ();
 sg13g2_fill_2 FILLER_34_1355 ();
 sg13g2_decap_8 FILLER_34_1383 ();
 sg13g2_decap_8 FILLER_34_1390 ();
 sg13g2_decap_4 FILLER_34_1397 ();
 sg13g2_fill_2 FILLER_34_1427 ();
 sg13g2_decap_4 FILLER_34_1439 ();
 sg13g2_fill_2 FILLER_34_1505 ();
 sg13g2_fill_1 FILLER_34_1507 ();
 sg13g2_decap_8 FILLER_34_1534 ();
 sg13g2_decap_8 FILLER_34_1541 ();
 sg13g2_decap_4 FILLER_34_1548 ();
 sg13g2_fill_1 FILLER_34_1552 ();
 sg13g2_fill_1 FILLER_34_1576 ();
 sg13g2_fill_1 FILLER_34_1592 ();
 sg13g2_decap_8 FILLER_34_1612 ();
 sg13g2_decap_4 FILLER_34_1619 ();
 sg13g2_fill_1 FILLER_34_1659 ();
 sg13g2_fill_1 FILLER_34_1666 ();
 sg13g2_decap_8 FILLER_34_1671 ();
 sg13g2_fill_2 FILLER_34_1678 ();
 sg13g2_fill_1 FILLER_34_1680 ();
 sg13g2_fill_2 FILLER_34_1685 ();
 sg13g2_fill_1 FILLER_34_1687 ();
 sg13g2_decap_8 FILLER_34_1723 ();
 sg13g2_decap_8 FILLER_34_1730 ();
 sg13g2_decap_8 FILLER_34_1737 ();
 sg13g2_decap_8 FILLER_34_1744 ();
 sg13g2_decap_8 FILLER_34_1751 ();
 sg13g2_decap_8 FILLER_34_1758 ();
 sg13g2_decap_8 FILLER_34_1765 ();
 sg13g2_fill_1 FILLER_34_1772 ();
 sg13g2_fill_1 FILLER_34_1778 ();
 sg13g2_decap_4 FILLER_34_1784 ();
 sg13g2_fill_2 FILLER_34_1788 ();
 sg13g2_decap_8 FILLER_34_1794 ();
 sg13g2_decap_8 FILLER_34_1801 ();
 sg13g2_fill_2 FILLER_34_1808 ();
 sg13g2_fill_1 FILLER_34_1810 ();
 sg13g2_fill_1 FILLER_34_1815 ();
 sg13g2_fill_2 FILLER_34_1828 ();
 sg13g2_fill_2 FILLER_34_1833 ();
 sg13g2_fill_1 FILLER_34_1835 ();
 sg13g2_fill_1 FILLER_34_1845 ();
 sg13g2_decap_8 FILLER_34_1850 ();
 sg13g2_fill_2 FILLER_34_1857 ();
 sg13g2_fill_1 FILLER_34_1859 ();
 sg13g2_decap_4 FILLER_34_1895 ();
 sg13g2_fill_1 FILLER_34_1899 ();
 sg13g2_fill_2 FILLER_34_1905 ();
 sg13g2_fill_1 FILLER_34_1907 ();
 sg13g2_fill_1 FILLER_34_1912 ();
 sg13g2_fill_2 FILLER_34_1921 ();
 sg13g2_fill_1 FILLER_34_1923 ();
 sg13g2_fill_1 FILLER_34_1950 ();
 sg13g2_fill_1 FILLER_34_1955 ();
 sg13g2_fill_2 FILLER_34_1992 ();
 sg13g2_decap_8 FILLER_34_2002 ();
 sg13g2_decap_8 FILLER_34_2009 ();
 sg13g2_fill_2 FILLER_34_2016 ();
 sg13g2_fill_1 FILLER_34_2023 ();
 sg13g2_fill_1 FILLER_34_2043 ();
 sg13g2_fill_2 FILLER_34_2048 ();
 sg13g2_fill_1 FILLER_34_2055 ();
 sg13g2_decap_8 FILLER_34_2082 ();
 sg13g2_fill_2 FILLER_34_2089 ();
 sg13g2_fill_1 FILLER_34_2091 ();
 sg13g2_decap_4 FILLER_34_2096 ();
 sg13g2_fill_2 FILLER_34_2105 ();
 sg13g2_decap_4 FILLER_34_2124 ();
 sg13g2_fill_2 FILLER_34_2131 ();
 sg13g2_fill_1 FILLER_34_2133 ();
 sg13g2_fill_1 FILLER_34_2164 ();
 sg13g2_fill_2 FILLER_34_2196 ();
 sg13g2_fill_1 FILLER_34_2198 ();
 sg13g2_decap_8 FILLER_34_2229 ();
 sg13g2_decap_8 FILLER_34_2302 ();
 sg13g2_decap_8 FILLER_34_2309 ();
 sg13g2_fill_1 FILLER_34_2316 ();
 sg13g2_decap_8 FILLER_34_2351 ();
 sg13g2_decap_8 FILLER_34_2358 ();
 sg13g2_fill_2 FILLER_34_2365 ();
 sg13g2_decap_8 FILLER_34_2376 ();
 sg13g2_decap_8 FILLER_34_2383 ();
 sg13g2_decap_8 FILLER_34_2390 ();
 sg13g2_decap_8 FILLER_34_2397 ();
 sg13g2_fill_1 FILLER_34_2404 ();
 sg13g2_decap_8 FILLER_34_2409 ();
 sg13g2_fill_2 FILLER_34_2416 ();
 sg13g2_decap_4 FILLER_34_2422 ();
 sg13g2_fill_2 FILLER_34_2426 ();
 sg13g2_fill_2 FILLER_34_2458 ();
 sg13g2_fill_1 FILLER_34_2460 ();
 sg13g2_fill_2 FILLER_34_2498 ();
 sg13g2_decap_8 FILLER_34_2504 ();
 sg13g2_decap_8 FILLER_34_2511 ();
 sg13g2_fill_2 FILLER_34_2518 ();
 sg13g2_fill_1 FILLER_34_2526 ();
 sg13g2_decap_4 FILLER_34_2560 ();
 sg13g2_fill_2 FILLER_34_2564 ();
 sg13g2_decap_8 FILLER_34_2592 ();
 sg13g2_fill_1 FILLER_34_2599 ();
 sg13g2_decap_8 FILLER_34_2629 ();
 sg13g2_decap_8 FILLER_34_2636 ();
 sg13g2_decap_8 FILLER_34_2643 ();
 sg13g2_decap_8 FILLER_34_2650 ();
 sg13g2_decap_8 FILLER_34_2657 ();
 sg13g2_decap_4 FILLER_34_2664 ();
 sg13g2_fill_2 FILLER_34_2668 ();
 sg13g2_decap_4 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_4 ();
 sg13g2_decap_4 FILLER_35_43 ();
 sg13g2_decap_8 FILLER_35_89 ();
 sg13g2_fill_2 FILLER_35_96 ();
 sg13g2_decap_8 FILLER_35_128 ();
 sg13g2_fill_1 FILLER_35_135 ();
 sg13g2_fill_2 FILLER_35_144 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_decap_4 FILLER_35_200 ();
 sg13g2_fill_2 FILLER_35_233 ();
 sg13g2_fill_1 FILLER_35_235 ();
 sg13g2_fill_1 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_4 FILLER_35_294 ();
 sg13g2_fill_1 FILLER_35_298 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_fill_2 FILLER_35_309 ();
 sg13g2_fill_1 FILLER_35_311 ();
 sg13g2_fill_2 FILLER_35_366 ();
 sg13g2_fill_1 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_412 ();
 sg13g2_decap_8 FILLER_35_419 ();
 sg13g2_fill_1 FILLER_35_426 ();
 sg13g2_decap_4 FILLER_35_431 ();
 sg13g2_fill_2 FILLER_35_435 ();
 sg13g2_decap_8 FILLER_35_440 ();
 sg13g2_decap_8 FILLER_35_447 ();
 sg13g2_decap_8 FILLER_35_487 ();
 sg13g2_decap_8 FILLER_35_494 ();
 sg13g2_fill_1 FILLER_35_501 ();
 sg13g2_decap_4 FILLER_35_516 ();
 sg13g2_fill_1 FILLER_35_538 ();
 sg13g2_decap_8 FILLER_35_544 ();
 sg13g2_decap_8 FILLER_35_551 ();
 sg13g2_decap_8 FILLER_35_558 ();
 sg13g2_decap_8 FILLER_35_565 ();
 sg13g2_decap_8 FILLER_35_572 ();
 sg13g2_fill_1 FILLER_35_579 ();
 sg13g2_fill_2 FILLER_35_598 ();
 sg13g2_fill_1 FILLER_35_620 ();
 sg13g2_fill_1 FILLER_35_631 ();
 sg13g2_decap_4 FILLER_35_651 ();
 sg13g2_fill_2 FILLER_35_655 ();
 sg13g2_fill_1 FILLER_35_661 ();
 sg13g2_decap_4 FILLER_35_688 ();
 sg13g2_fill_2 FILLER_35_692 ();
 sg13g2_decap_8 FILLER_35_697 ();
 sg13g2_decap_4 FILLER_35_704 ();
 sg13g2_fill_2 FILLER_35_708 ();
 sg13g2_fill_2 FILLER_35_714 ();
 sg13g2_fill_1 FILLER_35_716 ();
 sg13g2_fill_2 FILLER_35_725 ();
 sg13g2_decap_4 FILLER_35_750 ();
 sg13g2_fill_1 FILLER_35_754 ();
 sg13g2_fill_2 FILLER_35_781 ();
 sg13g2_fill_1 FILLER_35_811 ();
 sg13g2_fill_1 FILLER_35_846 ();
 sg13g2_decap_8 FILLER_35_856 ();
 sg13g2_fill_2 FILLER_35_863 ();
 sg13g2_decap_8 FILLER_35_869 ();
 sg13g2_fill_1 FILLER_35_876 ();
 sg13g2_fill_1 FILLER_35_934 ();
 sg13g2_fill_1 FILLER_35_982 ();
 sg13g2_fill_2 FILLER_35_987 ();
 sg13g2_fill_1 FILLER_35_997 ();
 sg13g2_fill_2 FILLER_35_1011 ();
 sg13g2_fill_2 FILLER_35_1017 ();
 sg13g2_fill_2 FILLER_35_1045 ();
 sg13g2_decap_4 FILLER_35_1073 ();
 sg13g2_fill_2 FILLER_35_1100 ();
 sg13g2_fill_1 FILLER_35_1102 ();
 sg13g2_fill_2 FILLER_35_1120 ();
 sg13g2_fill_1 FILLER_35_1134 ();
 sg13g2_fill_2 FILLER_35_1161 ();
 sg13g2_fill_1 FILLER_35_1163 ();
 sg13g2_decap_8 FILLER_35_1170 ();
 sg13g2_fill_1 FILLER_35_1242 ();
 sg13g2_fill_1 FILLER_35_1250 ();
 sg13g2_decap_8 FILLER_35_1265 ();
 sg13g2_decap_8 FILLER_35_1272 ();
 sg13g2_fill_1 FILLER_35_1279 ();
 sg13g2_decap_8 FILLER_35_1312 ();
 sg13g2_decap_8 FILLER_35_1319 ();
 sg13g2_decap_8 FILLER_35_1326 ();
 sg13g2_decap_8 FILLER_35_1333 ();
 sg13g2_decap_4 FILLER_35_1340 ();
 sg13g2_fill_1 FILLER_35_1344 ();
 sg13g2_decap_4 FILLER_35_1368 ();
 sg13g2_fill_2 FILLER_35_1372 ();
 sg13g2_fill_1 FILLER_35_1383 ();
 sg13g2_fill_1 FILLER_35_1394 ();
 sg13g2_decap_4 FILLER_35_1421 ();
 sg13g2_decap_8 FILLER_35_1443 ();
 sg13g2_fill_1 FILLER_35_1450 ();
 sg13g2_decap_8 FILLER_35_1457 ();
 sg13g2_decap_4 FILLER_35_1464 ();
 sg13g2_fill_1 FILLER_35_1468 ();
 sg13g2_fill_2 FILLER_35_1486 ();
 sg13g2_fill_2 FILLER_35_1494 ();
 sg13g2_fill_1 FILLER_35_1496 ();
 sg13g2_decap_8 FILLER_35_1518 ();
 sg13g2_decap_8 FILLER_35_1525 ();
 sg13g2_decap_4 FILLER_35_1532 ();
 sg13g2_fill_2 FILLER_35_1536 ();
 sg13g2_fill_2 FILLER_35_1561 ();
 sg13g2_fill_2 FILLER_35_1571 ();
 sg13g2_fill_1 FILLER_35_1578 ();
 sg13g2_fill_1 FILLER_35_1602 ();
 sg13g2_fill_1 FILLER_35_1608 ();
 sg13g2_fill_2 FILLER_35_1614 ();
 sg13g2_fill_1 FILLER_35_1629 ();
 sg13g2_fill_2 FILLER_35_1663 ();
 sg13g2_decap_8 FILLER_35_1732 ();
 sg13g2_fill_1 FILLER_35_1739 ();
 sg13g2_fill_2 FILLER_35_1776 ();
 sg13g2_decap_8 FILLER_35_1787 ();
 sg13g2_decap_8 FILLER_35_1794 ();
 sg13g2_decap_8 FILLER_35_1801 ();
 sg13g2_decap_4 FILLER_35_1808 ();
 sg13g2_decap_8 FILLER_35_1817 ();
 sg13g2_decap_4 FILLER_35_1824 ();
 sg13g2_fill_2 FILLER_35_1828 ();
 sg13g2_decap_4 FILLER_35_1834 ();
 sg13g2_fill_1 FILLER_35_1838 ();
 sg13g2_decap_8 FILLER_35_1852 ();
 sg13g2_decap_8 FILLER_35_1859 ();
 sg13g2_decap_8 FILLER_35_1866 ();
 sg13g2_decap_4 FILLER_35_1873 ();
 sg13g2_fill_2 FILLER_35_1877 ();
 sg13g2_decap_8 FILLER_35_1883 ();
 sg13g2_decap_4 FILLER_35_1890 ();
 sg13g2_fill_2 FILLER_35_1902 ();
 sg13g2_decap_8 FILLER_35_1936 ();
 sg13g2_decap_8 FILLER_35_1943 ();
 sg13g2_decap_8 FILLER_35_1950 ();
 sg13g2_decap_8 FILLER_35_1957 ();
 sg13g2_decap_8 FILLER_35_1964 ();
 sg13g2_decap_8 FILLER_35_1971 ();
 sg13g2_fill_1 FILLER_35_1983 ();
 sg13g2_decap_8 FILLER_35_1988 ();
 sg13g2_decap_8 FILLER_35_1995 ();
 sg13g2_fill_1 FILLER_35_2002 ();
 sg13g2_decap_8 FILLER_35_2060 ();
 sg13g2_decap_4 FILLER_35_2067 ();
 sg13g2_fill_1 FILLER_35_2071 ();
 sg13g2_decap_8 FILLER_35_2076 ();
 sg13g2_fill_1 FILLER_35_2083 ();
 sg13g2_fill_2 FILLER_35_2113 ();
 sg13g2_fill_1 FILLER_35_2115 ();
 sg13g2_decap_8 FILLER_35_2121 ();
 sg13g2_fill_2 FILLER_35_2128 ();
 sg13g2_fill_1 FILLER_35_2130 ();
 sg13g2_fill_1 FILLER_35_2137 ();
 sg13g2_decap_8 FILLER_35_2143 ();
 sg13g2_decap_8 FILLER_35_2150 ();
 sg13g2_fill_1 FILLER_35_2157 ();
 sg13g2_decap_4 FILLER_35_2169 ();
 sg13g2_decap_8 FILLER_35_2177 ();
 sg13g2_fill_2 FILLER_35_2184 ();
 sg13g2_decap_8 FILLER_35_2196 ();
 sg13g2_fill_2 FILLER_35_2203 ();
 sg13g2_fill_1 FILLER_35_2205 ();
 sg13g2_fill_2 FILLER_35_2215 ();
 sg13g2_decap_8 FILLER_35_2222 ();
 sg13g2_fill_2 FILLER_35_2229 ();
 sg13g2_fill_1 FILLER_35_2231 ();
 sg13g2_fill_2 FILLER_35_2242 ();
 sg13g2_fill_1 FILLER_35_2244 ();
 sg13g2_fill_2 FILLER_35_2255 ();
 sg13g2_fill_1 FILLER_35_2257 ();
 sg13g2_decap_8 FILLER_35_2268 ();
 sg13g2_fill_2 FILLER_35_2275 ();
 sg13g2_decap_8 FILLER_35_2309 ();
 sg13g2_decap_4 FILLER_35_2316 ();
 sg13g2_fill_1 FILLER_35_2320 ();
 sg13g2_decap_8 FILLER_35_2351 ();
 sg13g2_decap_4 FILLER_35_2358 ();
 sg13g2_fill_2 FILLER_35_2362 ();
 sg13g2_decap_4 FILLER_35_2377 ();
 sg13g2_fill_2 FILLER_35_2381 ();
 sg13g2_decap_4 FILLER_35_2392 ();
 sg13g2_fill_1 FILLER_35_2396 ();
 sg13g2_fill_1 FILLER_35_2402 ();
 sg13g2_decap_8 FILLER_35_2447 ();
 sg13g2_decap_8 FILLER_35_2454 ();
 sg13g2_fill_1 FILLER_35_2494 ();
 sg13g2_fill_1 FILLER_35_2537 ();
 sg13g2_decap_4 FILLER_35_2546 ();
 sg13g2_fill_1 FILLER_35_2550 ();
 sg13g2_fill_2 FILLER_35_2581 ();
 sg13g2_fill_1 FILLER_35_2583 ();
 sg13g2_decap_8 FILLER_35_2614 ();
 sg13g2_decap_8 FILLER_35_2621 ();
 sg13g2_fill_2 FILLER_35_2628 ();
 sg13g2_fill_1 FILLER_35_2669 ();
 sg13g2_decap_4 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_4 ();
 sg13g2_decap_8 FILLER_36_36 ();
 sg13g2_decap_8 FILLER_36_43 ();
 sg13g2_decap_4 FILLER_36_50 ();
 sg13g2_decap_8 FILLER_36_62 ();
 sg13g2_decap_8 FILLER_36_69 ();
 sg13g2_decap_4 FILLER_36_76 ();
 sg13g2_fill_2 FILLER_36_80 ();
 sg13g2_decap_8 FILLER_36_86 ();
 sg13g2_decap_8 FILLER_36_93 ();
 sg13g2_decap_8 FILLER_36_100 ();
 sg13g2_decap_8 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_114 ();
 sg13g2_fill_2 FILLER_36_150 ();
 sg13g2_fill_2 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_171 ();
 sg13g2_decap_4 FILLER_36_184 ();
 sg13g2_fill_1 FILLER_36_188 ();
 sg13g2_fill_2 FILLER_36_192 ();
 sg13g2_fill_1 FILLER_36_194 ();
 sg13g2_fill_1 FILLER_36_204 ();
 sg13g2_fill_1 FILLER_36_260 ();
 sg13g2_fill_1 FILLER_36_267 ();
 sg13g2_decap_8 FILLER_36_275 ();
 sg13g2_decap_8 FILLER_36_282 ();
 sg13g2_decap_4 FILLER_36_289 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_decap_4 FILLER_36_358 ();
 sg13g2_fill_2 FILLER_36_429 ();
 sg13g2_fill_1 FILLER_36_431 ();
 sg13g2_fill_2 FILLER_36_458 ();
 sg13g2_fill_1 FILLER_36_479 ();
 sg13g2_decap_8 FILLER_36_484 ();
 sg13g2_decap_4 FILLER_36_491 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_fill_2 FILLER_36_511 ();
 sg13g2_fill_1 FILLER_36_513 ();
 sg13g2_decap_8 FILLER_36_519 ();
 sg13g2_fill_2 FILLER_36_526 ();
 sg13g2_fill_2 FILLER_36_532 ();
 sg13g2_fill_1 FILLER_36_534 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_fill_1 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_565 ();
 sg13g2_decap_8 FILLER_36_572 ();
 sg13g2_decap_8 FILLER_36_584 ();
 sg13g2_fill_1 FILLER_36_591 ();
 sg13g2_fill_2 FILLER_36_602 ();
 sg13g2_fill_1 FILLER_36_622 ();
 sg13g2_fill_1 FILLER_36_628 ();
 sg13g2_fill_2 FILLER_36_646 ();
 sg13g2_fill_1 FILLER_36_648 ();
 sg13g2_decap_8 FILLER_36_654 ();
 sg13g2_decap_8 FILLER_36_661 ();
 sg13g2_decap_4 FILLER_36_668 ();
 sg13g2_decap_4 FILLER_36_675 ();
 sg13g2_fill_2 FILLER_36_679 ();
 sg13g2_fill_1 FILLER_36_695 ();
 sg13g2_fill_2 FILLER_36_700 ();
 sg13g2_fill_2 FILLER_36_710 ();
 sg13g2_fill_2 FILLER_36_722 ();
 sg13g2_fill_2 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_752 ();
 sg13g2_decap_8 FILLER_36_759 ();
 sg13g2_decap_4 FILLER_36_766 ();
 sg13g2_fill_2 FILLER_36_770 ();
 sg13g2_fill_1 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_821 ();
 sg13g2_fill_1 FILLER_36_828 ();
 sg13g2_decap_4 FILLER_36_839 ();
 sg13g2_fill_1 FILLER_36_843 ();
 sg13g2_fill_1 FILLER_36_849 ();
 sg13g2_decap_8 FILLER_36_860 ();
 sg13g2_decap_8 FILLER_36_867 ();
 sg13g2_decap_8 FILLER_36_879 ();
 sg13g2_decap_8 FILLER_36_886 ();
 sg13g2_fill_1 FILLER_36_893 ();
 sg13g2_fill_1 FILLER_36_906 ();
 sg13g2_fill_1 FILLER_36_913 ();
 sg13g2_fill_1 FILLER_36_958 ();
 sg13g2_decap_4 FILLER_36_963 ();
 sg13g2_fill_1 FILLER_36_967 ();
 sg13g2_fill_2 FILLER_36_973 ();
 sg13g2_fill_1 FILLER_36_975 ();
 sg13g2_fill_2 FILLER_36_982 ();
 sg13g2_fill_1 FILLER_36_1045 ();
 sg13g2_fill_2 FILLER_36_1098 ();
 sg13g2_fill_1 FILLER_36_1109 ();
 sg13g2_fill_1 FILLER_36_1153 ();
 sg13g2_decap_8 FILLER_36_1158 ();
 sg13g2_fill_1 FILLER_36_1165 ();
 sg13g2_decap_8 FILLER_36_1170 ();
 sg13g2_decap_8 FILLER_36_1177 ();
 sg13g2_decap_8 FILLER_36_1184 ();
 sg13g2_fill_2 FILLER_36_1191 ();
 sg13g2_fill_2 FILLER_36_1202 ();
 sg13g2_fill_1 FILLER_36_1204 ();
 sg13g2_fill_2 FILLER_36_1213 ();
 sg13g2_fill_1 FILLER_36_1241 ();
 sg13g2_fill_1 FILLER_36_1246 ();
 sg13g2_decap_4 FILLER_36_1261 ();
 sg13g2_fill_1 FILLER_36_1265 ();
 sg13g2_fill_2 FILLER_36_1275 ();
 sg13g2_fill_1 FILLER_36_1277 ();
 sg13g2_decap_8 FILLER_36_1309 ();
 sg13g2_decap_8 FILLER_36_1316 ();
 sg13g2_fill_1 FILLER_36_1323 ();
 sg13g2_decap_4 FILLER_36_1330 ();
 sg13g2_fill_1 FILLER_36_1334 ();
 sg13g2_decap_4 FILLER_36_1388 ();
 sg13g2_fill_1 FILLER_36_1392 ();
 sg13g2_decap_4 FILLER_36_1419 ();
 sg13g2_decap_8 FILLER_36_1438 ();
 sg13g2_decap_4 FILLER_36_1445 ();
 sg13g2_fill_2 FILLER_36_1449 ();
 sg13g2_decap_8 FILLER_36_1487 ();
 sg13g2_fill_2 FILLER_36_1494 ();
 sg13g2_fill_1 FILLER_36_1496 ();
 sg13g2_decap_8 FILLER_36_1523 ();
 sg13g2_fill_1 FILLER_36_1530 ();
 sg13g2_fill_1 FILLER_36_1536 ();
 sg13g2_decap_8 FILLER_36_1547 ();
 sg13g2_fill_2 FILLER_36_1554 ();
 sg13g2_fill_2 FILLER_36_1560 ();
 sg13g2_fill_2 FILLER_36_1568 ();
 sg13g2_fill_1 FILLER_36_1570 ();
 sg13g2_fill_2 FILLER_36_1582 ();
 sg13g2_fill_1 FILLER_36_1590 ();
 sg13g2_fill_2 FILLER_36_1600 ();
 sg13g2_fill_2 FILLER_36_1607 ();
 sg13g2_fill_2 FILLER_36_1614 ();
 sg13g2_fill_2 FILLER_36_1620 ();
 sg13g2_fill_1 FILLER_36_1622 ();
 sg13g2_decap_4 FILLER_36_1637 ();
 sg13g2_fill_2 FILLER_36_1650 ();
 sg13g2_fill_1 FILLER_36_1652 ();
 sg13g2_decap_8 FILLER_36_1659 ();
 sg13g2_decap_8 FILLER_36_1666 ();
 sg13g2_fill_2 FILLER_36_1673 ();
 sg13g2_fill_1 FILLER_36_1675 ();
 sg13g2_decap_8 FILLER_36_1680 ();
 sg13g2_decap_4 FILLER_36_1687 ();
 sg13g2_fill_2 FILLER_36_1718 ();
 sg13g2_fill_2 FILLER_36_1746 ();
 sg13g2_fill_2 FILLER_36_1751 ();
 sg13g2_decap_4 FILLER_36_1786 ();
 sg13g2_decap_4 FILLER_36_1794 ();
 sg13g2_fill_1 FILLER_36_1798 ();
 sg13g2_decap_4 FILLER_36_1805 ();
 sg13g2_fill_2 FILLER_36_1809 ();
 sg13g2_decap_8 FILLER_36_1816 ();
 sg13g2_decap_4 FILLER_36_1823 ();
 sg13g2_decap_8 FILLER_36_1857 ();
 sg13g2_decap_8 FILLER_36_1864 ();
 sg13g2_fill_2 FILLER_36_1871 ();
 sg13g2_fill_1 FILLER_36_1873 ();
 sg13g2_decap_8 FILLER_36_1883 ();
 sg13g2_decap_8 FILLER_36_1890 ();
 sg13g2_fill_1 FILLER_36_1897 ();
 sg13g2_decap_8 FILLER_36_1942 ();
 sg13g2_fill_1 FILLER_36_1949 ();
 sg13g2_fill_1 FILLER_36_1955 ();
 sg13g2_decap_4 FILLER_36_2001 ();
 sg13g2_decap_8 FILLER_36_2070 ();
 sg13g2_decap_8 FILLER_36_2077 ();
 sg13g2_fill_2 FILLER_36_2084 ();
 sg13g2_fill_1 FILLER_36_2086 ();
 sg13g2_decap_8 FILLER_36_2100 ();
 sg13g2_fill_1 FILLER_36_2107 ();
 sg13g2_decap_4 FILLER_36_2117 ();
 sg13g2_fill_2 FILLER_36_2121 ();
 sg13g2_decap_4 FILLER_36_2131 ();
 sg13g2_fill_1 FILLER_36_2135 ();
 sg13g2_fill_2 FILLER_36_2141 ();
 sg13g2_fill_1 FILLER_36_2199 ();
 sg13g2_decap_4 FILLER_36_2204 ();
 sg13g2_fill_2 FILLER_36_2208 ();
 sg13g2_decap_4 FILLER_36_2214 ();
 sg13g2_fill_2 FILLER_36_2244 ();
 sg13g2_decap_8 FILLER_36_2254 ();
 sg13g2_decap_8 FILLER_36_2274 ();
 sg13g2_decap_8 FILLER_36_2281 ();
 sg13g2_fill_1 FILLER_36_2288 ();
 sg13g2_decap_8 FILLER_36_2295 ();
 sg13g2_decap_4 FILLER_36_2302 ();
 sg13g2_fill_1 FILLER_36_2306 ();
 sg13g2_fill_1 FILLER_36_2341 ();
 sg13g2_decap_4 FILLER_36_2346 ();
 sg13g2_fill_1 FILLER_36_2350 ();
 sg13g2_decap_8 FILLER_36_2361 ();
 sg13g2_decap_4 FILLER_36_2368 ();
 sg13g2_fill_1 FILLER_36_2372 ();
 sg13g2_decap_4 FILLER_36_2386 ();
 sg13g2_fill_1 FILLER_36_2416 ();
 sg13g2_fill_2 FILLER_36_2434 ();
 sg13g2_fill_2 FILLER_36_2462 ();
 sg13g2_decap_8 FILLER_36_2472 ();
 sg13g2_decap_4 FILLER_36_2543 ();
 sg13g2_fill_1 FILLER_36_2547 ();
 sg13g2_fill_2 FILLER_36_2554 ();
 sg13g2_fill_1 FILLER_36_2556 ();
 sg13g2_fill_2 FILLER_36_2563 ();
 sg13g2_fill_2 FILLER_36_2569 ();
 sg13g2_fill_1 FILLER_36_2571 ();
 sg13g2_fill_2 FILLER_36_2589 ();
 sg13g2_decap_8 FILLER_36_2617 ();
 sg13g2_decap_4 FILLER_36_2624 ();
 sg13g2_decap_8 FILLER_36_2662 ();
 sg13g2_fill_1 FILLER_36_2669 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_4 FILLER_37_14 ();
 sg13g2_fill_2 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_41 ();
 sg13g2_decap_4 FILLER_37_48 ();
 sg13g2_fill_1 FILLER_37_52 ();
 sg13g2_decap_8 FILLER_37_66 ();
 sg13g2_decap_8 FILLER_37_73 ();
 sg13g2_decap_8 FILLER_37_80 ();
 sg13g2_decap_8 FILLER_37_87 ();
 sg13g2_decap_8 FILLER_37_94 ();
 sg13g2_decap_8 FILLER_37_101 ();
 sg13g2_decap_8 FILLER_37_108 ();
 sg13g2_decap_8 FILLER_37_115 ();
 sg13g2_decap_8 FILLER_37_122 ();
 sg13g2_decap_8 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_136 ();
 sg13g2_fill_2 FILLER_37_145 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_4 FILLER_37_200 ();
 sg13g2_fill_1 FILLER_37_243 ();
 sg13g2_fill_1 FILLER_37_248 ();
 sg13g2_fill_2 FILLER_37_253 ();
 sg13g2_fill_1 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_305 ();
 sg13g2_fill_2 FILLER_37_314 ();
 sg13g2_decap_4 FILLER_37_329 ();
 sg13g2_fill_2 FILLER_37_377 ();
 sg13g2_fill_1 FILLER_37_403 ();
 sg13g2_fill_1 FILLER_37_409 ();
 sg13g2_fill_1 FILLER_37_414 ();
 sg13g2_fill_2 FILLER_37_420 ();
 sg13g2_decap_8 FILLER_37_449 ();
 sg13g2_decap_4 FILLER_37_456 ();
 sg13g2_fill_1 FILLER_37_460 ();
 sg13g2_decap_8 FILLER_37_487 ();
 sg13g2_decap_8 FILLER_37_494 ();
 sg13g2_fill_1 FILLER_37_528 ();
 sg13g2_decap_8 FILLER_37_538 ();
 sg13g2_decap_4 FILLER_37_545 ();
 sg13g2_fill_2 FILLER_37_549 ();
 sg13g2_fill_2 FILLER_37_561 ();
 sg13g2_fill_1 FILLER_37_577 ();
 sg13g2_fill_2 FILLER_37_582 ();
 sg13g2_decap_4 FILLER_37_593 ();
 sg13g2_decap_4 FILLER_37_612 ();
 sg13g2_fill_2 FILLER_37_616 ();
 sg13g2_fill_2 FILLER_37_622 ();
 sg13g2_fill_1 FILLER_37_631 ();
 sg13g2_decap_4 FILLER_37_635 ();
 sg13g2_fill_1 FILLER_37_649 ();
 sg13g2_fill_1 FILLER_37_659 ();
 sg13g2_fill_1 FILLER_37_668 ();
 sg13g2_fill_2 FILLER_37_712 ();
 sg13g2_fill_2 FILLER_37_730 ();
 sg13g2_fill_2 FILLER_37_737 ();
 sg13g2_fill_2 FILLER_37_745 ();
 sg13g2_fill_1 FILLER_37_776 ();
 sg13g2_fill_1 FILLER_37_782 ();
 sg13g2_decap_4 FILLER_37_788 ();
 sg13g2_fill_1 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_829 ();
 sg13g2_decap_8 FILLER_37_867 ();
 sg13g2_decap_4 FILLER_37_874 ();
 sg13g2_fill_2 FILLER_37_878 ();
 sg13g2_decap_4 FILLER_37_889 ();
 sg13g2_decap_8 FILLER_37_919 ();
 sg13g2_decap_8 FILLER_37_926 ();
 sg13g2_decap_4 FILLER_37_933 ();
 sg13g2_fill_2 FILLER_37_937 ();
 sg13g2_fill_2 FILLER_37_951 ();
 sg13g2_decap_8 FILLER_37_959 ();
 sg13g2_decap_8 FILLER_37_966 ();
 sg13g2_fill_2 FILLER_37_973 ();
 sg13g2_fill_1 FILLER_37_975 ();
 sg13g2_fill_2 FILLER_37_984 ();
 sg13g2_fill_2 FILLER_37_1026 ();
 sg13g2_fill_2 FILLER_37_1033 ();
 sg13g2_fill_1 FILLER_37_1035 ();
 sg13g2_decap_4 FILLER_37_1049 ();
 sg13g2_fill_1 FILLER_37_1053 ();
 sg13g2_decap_8 FILLER_37_1063 ();
 sg13g2_fill_1 FILLER_37_1070 ();
 sg13g2_fill_2 FILLER_37_1076 ();
 sg13g2_decap_8 FILLER_37_1114 ();
 sg13g2_fill_1 FILLER_37_1121 ();
 sg13g2_fill_2 FILLER_37_1130 ();
 sg13g2_fill_1 FILLER_37_1141 ();
 sg13g2_decap_8 FILLER_37_1155 ();
 sg13g2_decap_8 FILLER_37_1162 ();
 sg13g2_decap_4 FILLER_37_1169 ();
 sg13g2_fill_1 FILLER_37_1173 ();
 sg13g2_decap_8 FILLER_37_1178 ();
 sg13g2_decap_4 FILLER_37_1185 ();
 sg13g2_decap_4 FILLER_37_1193 ();
 sg13g2_fill_2 FILLER_37_1197 ();
 sg13g2_decap_8 FILLER_37_1218 ();
 sg13g2_decap_8 FILLER_37_1225 ();
 sg13g2_fill_1 FILLER_37_1297 ();
 sg13g2_fill_2 FILLER_37_1302 ();
 sg13g2_fill_1 FILLER_37_1304 ();
 sg13g2_decap_8 FILLER_37_1339 ();
 sg13g2_decap_8 FILLER_37_1346 ();
 sg13g2_decap_8 FILLER_37_1353 ();
 sg13g2_decap_4 FILLER_37_1360 ();
 sg13g2_fill_1 FILLER_37_1364 ();
 sg13g2_decap_4 FILLER_37_1416 ();
 sg13g2_fill_1 FILLER_37_1420 ();
 sg13g2_decap_4 FILLER_37_1447 ();
 sg13g2_decap_4 FILLER_37_1468 ();
 sg13g2_fill_1 FILLER_37_1472 ();
 sg13g2_decap_8 FILLER_37_1479 ();
 sg13g2_decap_8 FILLER_37_1486 ();
 sg13g2_decap_8 FILLER_37_1493 ();
 sg13g2_decap_8 FILLER_37_1500 ();
 sg13g2_decap_8 FILLER_37_1507 ();
 sg13g2_decap_8 FILLER_37_1514 ();
 sg13g2_fill_2 FILLER_37_1521 ();
 sg13g2_decap_4 FILLER_37_1529 ();
 sg13g2_fill_1 FILLER_37_1562 ();
 sg13g2_fill_2 FILLER_37_1568 ();
 sg13g2_fill_1 FILLER_37_1576 ();
 sg13g2_fill_1 FILLER_37_1599 ();
 sg13g2_fill_1 FILLER_37_1618 ();
 sg13g2_fill_2 FILLER_37_1636 ();
 sg13g2_fill_1 FILLER_37_1638 ();
 sg13g2_decap_8 FILLER_37_1652 ();
 sg13g2_fill_2 FILLER_37_1659 ();
 sg13g2_fill_1 FILLER_37_1661 ();
 sg13g2_decap_8 FILLER_37_1667 ();
 sg13g2_decap_8 FILLER_37_1674 ();
 sg13g2_fill_2 FILLER_37_1740 ();
 sg13g2_fill_2 FILLER_37_1769 ();
 sg13g2_fill_1 FILLER_37_1771 ();
 sg13g2_fill_2 FILLER_37_1776 ();
 sg13g2_decap_8 FILLER_37_1782 ();
 sg13g2_decap_8 FILLER_37_1789 ();
 sg13g2_fill_2 FILLER_37_1800 ();
 sg13g2_fill_1 FILLER_37_1802 ();
 sg13g2_fill_1 FILLER_37_1808 ();
 sg13g2_fill_2 FILLER_37_1814 ();
 sg13g2_decap_4 FILLER_37_1820 ();
 sg13g2_decap_8 FILLER_37_1834 ();
 sg13g2_decap_4 FILLER_37_1841 ();
 sg13g2_decap_8 FILLER_37_1849 ();
 sg13g2_decap_4 FILLER_37_1856 ();
 sg13g2_fill_2 FILLER_37_1860 ();
 sg13g2_decap_8 FILLER_37_1893 ();
 sg13g2_fill_2 FILLER_37_1900 ();
 sg13g2_fill_1 FILLER_37_1902 ();
 sg13g2_fill_1 FILLER_37_1934 ();
 sg13g2_decap_8 FILLER_37_1965 ();
 sg13g2_decap_8 FILLER_37_1972 ();
 sg13g2_decap_8 FILLER_37_1979 ();
 sg13g2_decap_8 FILLER_37_1990 ();
 sg13g2_decap_8 FILLER_37_1997 ();
 sg13g2_decap_4 FILLER_37_2004 ();
 sg13g2_fill_2 FILLER_37_2008 ();
 sg13g2_decap_8 FILLER_37_2069 ();
 sg13g2_fill_2 FILLER_37_2076 ();
 sg13g2_fill_1 FILLER_37_2078 ();
 sg13g2_fill_1 FILLER_37_2106 ();
 sg13g2_decap_8 FILLER_37_2124 ();
 sg13g2_fill_2 FILLER_37_2131 ();
 sg13g2_fill_2 FILLER_37_2141 ();
 sg13g2_decap_8 FILLER_37_2148 ();
 sg13g2_fill_1 FILLER_37_2155 ();
 sg13g2_decap_8 FILLER_37_2160 ();
 sg13g2_fill_1 FILLER_37_2172 ();
 sg13g2_fill_2 FILLER_37_2187 ();
 sg13g2_fill_1 FILLER_37_2189 ();
 sg13g2_decap_8 FILLER_37_2204 ();
 sg13g2_decap_8 FILLER_37_2211 ();
 sg13g2_fill_2 FILLER_37_2243 ();
 sg13g2_decap_8 FILLER_37_2254 ();
 sg13g2_decap_4 FILLER_37_2261 ();
 sg13g2_fill_2 FILLER_37_2265 ();
 sg13g2_fill_2 FILLER_37_2271 ();
 sg13g2_decap_8 FILLER_37_2290 ();
 sg13g2_fill_2 FILLER_37_2297 ();
 sg13g2_decap_8 FILLER_37_2313 ();
 sg13g2_fill_2 FILLER_37_2320 ();
 sg13g2_decap_8 FILLER_37_2328 ();
 sg13g2_decap_4 FILLER_37_2335 ();
 sg13g2_decap_8 FILLER_37_2375 ();
 sg13g2_decap_4 FILLER_37_2382 ();
 sg13g2_fill_1 FILLER_37_2386 ();
 sg13g2_fill_2 FILLER_37_2392 ();
 sg13g2_fill_1 FILLER_37_2394 ();
 sg13g2_decap_4 FILLER_37_2405 ();
 sg13g2_fill_2 FILLER_37_2409 ();
 sg13g2_decap_4 FILLER_37_2415 ();
 sg13g2_fill_1 FILLER_37_2419 ();
 sg13g2_fill_1 FILLER_37_2438 ();
 sg13g2_fill_2 FILLER_37_2471 ();
 sg13g2_fill_1 FILLER_37_2473 ();
 sg13g2_decap_8 FILLER_37_2482 ();
 sg13g2_fill_2 FILLER_37_2489 ();
 sg13g2_fill_1 FILLER_37_2494 ();
 sg13g2_decap_4 FILLER_37_2499 ();
 sg13g2_fill_2 FILLER_37_2507 ();
 sg13g2_decap_8 FILLER_37_2522 ();
 sg13g2_decap_8 FILLER_37_2529 ();
 sg13g2_decap_8 FILLER_37_2540 ();
 sg13g2_decap_8 FILLER_37_2560 ();
 sg13g2_decap_8 FILLER_37_2567 ();
 sg13g2_decap_8 FILLER_37_2574 ();
 sg13g2_fill_1 FILLER_37_2581 ();
 sg13g2_decap_8 FILLER_37_2602 ();
 sg13g2_fill_1 FILLER_37_2609 ();
 sg13g2_decap_8 FILLER_37_2638 ();
 sg13g2_decap_4 FILLER_37_2645 ();
 sg13g2_fill_2 FILLER_37_2649 ();
 sg13g2_decap_4 FILLER_37_2664 ();
 sg13g2_fill_2 FILLER_37_2668 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_fill_2 FILLER_38_28 ();
 sg13g2_fill_1 FILLER_38_30 ();
 sg13g2_decap_8 FILLER_38_34 ();
 sg13g2_decap_4 FILLER_38_41 ();
 sg13g2_fill_2 FILLER_38_45 ();
 sg13g2_decap_8 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_95 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_fill_2 FILLER_38_129 ();
 sg13g2_fill_1 FILLER_38_131 ();
 sg13g2_fill_1 FILLER_38_140 ();
 sg13g2_decap_4 FILLER_38_189 ();
 sg13g2_fill_2 FILLER_38_193 ();
 sg13g2_decap_8 FILLER_38_243 ();
 sg13g2_decap_8 FILLER_38_250 ();
 sg13g2_decap_4 FILLER_38_257 ();
 sg13g2_fill_1 FILLER_38_284 ();
 sg13g2_decap_4 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_330 ();
 sg13g2_decap_8 FILLER_38_354 ();
 sg13g2_decap_8 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_381 ();
 sg13g2_decap_4 FILLER_38_390 ();
 sg13g2_fill_2 FILLER_38_394 ();
 sg13g2_fill_2 FILLER_38_401 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_1 FILLER_38_442 ();
 sg13g2_fill_2 FILLER_38_448 ();
 sg13g2_fill_1 FILLER_38_450 ();
 sg13g2_fill_2 FILLER_38_456 ();
 sg13g2_decap_8 FILLER_38_479 ();
 sg13g2_decap_4 FILLER_38_486 ();
 sg13g2_decap_8 FILLER_38_496 ();
 sg13g2_fill_1 FILLER_38_503 ();
 sg13g2_decap_4 FILLER_38_508 ();
 sg13g2_decap_4 FILLER_38_520 ();
 sg13g2_fill_2 FILLER_38_524 ();
 sg13g2_decap_8 FILLER_38_531 ();
 sg13g2_decap_8 FILLER_38_538 ();
 sg13g2_decap_8 FILLER_38_545 ();
 sg13g2_decap_8 FILLER_38_552 ();
 sg13g2_fill_1 FILLER_38_583 ();
 sg13g2_fill_1 FILLER_38_595 ();
 sg13g2_fill_1 FILLER_38_606 ();
 sg13g2_fill_1 FILLER_38_612 ();
 sg13g2_decap_4 FILLER_38_642 ();
 sg13g2_fill_1 FILLER_38_649 ();
 sg13g2_fill_2 FILLER_38_653 ();
 sg13g2_fill_1 FILLER_38_664 ();
 sg13g2_fill_2 FILLER_38_673 ();
 sg13g2_fill_1 FILLER_38_695 ();
 sg13g2_fill_2 FILLER_38_750 ();
 sg13g2_fill_1 FILLER_38_757 ();
 sg13g2_fill_1 FILLER_38_763 ();
 sg13g2_fill_2 FILLER_38_772 ();
 sg13g2_fill_2 FILLER_38_778 ();
 sg13g2_decap_8 FILLER_38_827 ();
 sg13g2_fill_1 FILLER_38_860 ();
 sg13g2_fill_1 FILLER_38_865 ();
 sg13g2_decap_8 FILLER_38_892 ();
 sg13g2_decap_4 FILLER_38_899 ();
 sg13g2_decap_8 FILLER_38_912 ();
 sg13g2_decap_8 FILLER_38_919 ();
 sg13g2_decap_8 FILLER_38_926 ();
 sg13g2_decap_8 FILLER_38_933 ();
 sg13g2_fill_2 FILLER_38_940 ();
 sg13g2_fill_1 FILLER_38_942 ();
 sg13g2_decap_8 FILLER_38_951 ();
 sg13g2_decap_8 FILLER_38_984 ();
 sg13g2_decap_8 FILLER_38_996 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_fill_2 FILLER_38_1015 ();
 sg13g2_fill_1 FILLER_38_1036 ();
 sg13g2_fill_2 FILLER_38_1051 ();
 sg13g2_fill_2 FILLER_38_1057 ();
 sg13g2_decap_8 FILLER_38_1068 ();
 sg13g2_decap_4 FILLER_38_1075 ();
 sg13g2_fill_2 FILLER_38_1087 ();
 sg13g2_fill_1 FILLER_38_1089 ();
 sg13g2_fill_1 FILLER_38_1099 ();
 sg13g2_decap_8 FILLER_38_1114 ();
 sg13g2_fill_1 FILLER_38_1169 ();
 sg13g2_decap_4 FILLER_38_1201 ();
 sg13g2_fill_1 FILLER_38_1205 ();
 sg13g2_fill_2 FILLER_38_1211 ();
 sg13g2_decap_4 FILLER_38_1218 ();
 sg13g2_decap_8 FILLER_38_1230 ();
 sg13g2_decap_8 FILLER_38_1237 ();
 sg13g2_decap_8 FILLER_38_1247 ();
 sg13g2_fill_1 FILLER_38_1254 ();
 sg13g2_decap_4 FILLER_38_1258 ();
 sg13g2_fill_1 FILLER_38_1262 ();
 sg13g2_fill_2 FILLER_38_1298 ();
 sg13g2_fill_1 FILLER_38_1300 ();
 sg13g2_fill_1 FILLER_38_1310 ();
 sg13g2_fill_2 FILLER_38_1402 ();
 sg13g2_decap_8 FILLER_38_1417 ();
 sg13g2_decap_8 FILLER_38_1424 ();
 sg13g2_decap_8 FILLER_38_1431 ();
 sg13g2_decap_8 FILLER_38_1438 ();
 sg13g2_decap_4 FILLER_38_1445 ();
 sg13g2_fill_2 FILLER_38_1449 ();
 sg13g2_fill_1 FILLER_38_1460 ();
 sg13g2_decap_8 FILLER_38_1474 ();
 sg13g2_decap_8 FILLER_38_1481 ();
 sg13g2_decap_8 FILLER_38_1488 ();
 sg13g2_decap_8 FILLER_38_1495 ();
 sg13g2_decap_8 FILLER_38_1502 ();
 sg13g2_decap_8 FILLER_38_1515 ();
 sg13g2_fill_1 FILLER_38_1527 ();
 sg13g2_fill_2 FILLER_38_1533 ();
 sg13g2_fill_1 FILLER_38_1547 ();
 sg13g2_fill_1 FILLER_38_1553 ();
 sg13g2_fill_2 FILLER_38_1560 ();
 sg13g2_fill_2 FILLER_38_1568 ();
 sg13g2_fill_1 FILLER_38_1570 ();
 sg13g2_fill_2 FILLER_38_1576 ();
 sg13g2_fill_1 FILLER_38_1578 ();
 sg13g2_fill_2 FILLER_38_1589 ();
 sg13g2_fill_1 FILLER_38_1591 ();
 sg13g2_fill_1 FILLER_38_1597 ();
 sg13g2_fill_2 FILLER_38_1605 ();
 sg13g2_fill_1 FILLER_38_1607 ();
 sg13g2_decap_4 FILLER_38_1621 ();
 sg13g2_fill_2 FILLER_38_1666 ();
 sg13g2_decap_4 FILLER_38_1673 ();
 sg13g2_fill_2 FILLER_38_1697 ();
 sg13g2_fill_2 FILLER_38_1747 ();
 sg13g2_decap_8 FILLER_38_1779 ();
 sg13g2_fill_2 FILLER_38_1786 ();
 sg13g2_fill_2 FILLER_38_1792 ();
 sg13g2_decap_8 FILLER_38_1840 ();
 sg13g2_decap_8 FILLER_38_1847 ();
 sg13g2_decap_8 FILLER_38_1854 ();
 sg13g2_decap_4 FILLER_38_1861 ();
 sg13g2_fill_2 FILLER_38_1865 ();
 sg13g2_fill_1 FILLER_38_1897 ();
 sg13g2_decap_4 FILLER_38_1917 ();
 sg13g2_fill_2 FILLER_38_1927 ();
 sg13g2_decap_8 FILLER_38_1968 ();
 sg13g2_decap_8 FILLER_38_1975 ();
 sg13g2_decap_8 FILLER_38_1991 ();
 sg13g2_decap_8 FILLER_38_1998 ();
 sg13g2_decap_4 FILLER_38_2005 ();
 sg13g2_fill_1 FILLER_38_2009 ();
 sg13g2_fill_2 FILLER_38_2014 ();
 sg13g2_fill_1 FILLER_38_2016 ();
 sg13g2_fill_2 FILLER_38_2025 ();
 sg13g2_decap_8 FILLER_38_2065 ();
 sg13g2_decap_8 FILLER_38_2072 ();
 sg13g2_decap_4 FILLER_38_2079 ();
 sg13g2_fill_1 FILLER_38_2089 ();
 sg13g2_fill_2 FILLER_38_2126 ();
 sg13g2_fill_1 FILLER_38_2128 ();
 sg13g2_decap_4 FILLER_38_2138 ();
 sg13g2_fill_2 FILLER_38_2142 ();
 sg13g2_decap_8 FILLER_38_2182 ();
 sg13g2_decap_4 FILLER_38_2189 ();
 sg13g2_fill_1 FILLER_38_2193 ();
 sg13g2_fill_2 FILLER_38_2202 ();
 sg13g2_fill_1 FILLER_38_2212 ();
 sg13g2_fill_2 FILLER_38_2227 ();
 sg13g2_fill_1 FILLER_38_2238 ();
 sg13g2_decap_8 FILLER_38_2244 ();
 sg13g2_decap_4 FILLER_38_2251 ();
 sg13g2_decap_4 FILLER_38_2261 ();
 sg13g2_fill_2 FILLER_38_2265 ();
 sg13g2_decap_8 FILLER_38_2276 ();
 sg13g2_fill_2 FILLER_38_2283 ();
 sg13g2_decap_8 FILLER_38_2315 ();
 sg13g2_fill_1 FILLER_38_2322 ();
 sg13g2_decap_8 FILLER_38_2328 ();
 sg13g2_decap_4 FILLER_38_2335 ();
 sg13g2_fill_2 FILLER_38_2339 ();
 sg13g2_fill_2 FILLER_38_2345 ();
 sg13g2_fill_1 FILLER_38_2347 ();
 sg13g2_fill_2 FILLER_38_2352 ();
 sg13g2_fill_1 FILLER_38_2354 ();
 sg13g2_fill_1 FILLER_38_2371 ();
 sg13g2_fill_1 FILLER_38_2376 ();
 sg13g2_fill_1 FILLER_38_2387 ();
 sg13g2_fill_1 FILLER_38_2392 ();
 sg13g2_decap_8 FILLER_38_2398 ();
 sg13g2_decap_4 FILLER_38_2410 ();
 sg13g2_decap_8 FILLER_38_2418 ();
 sg13g2_decap_8 FILLER_38_2425 ();
 sg13g2_decap_4 FILLER_38_2432 ();
 sg13g2_fill_1 FILLER_38_2436 ();
 sg13g2_fill_2 FILLER_38_2447 ();
 sg13g2_decap_8 FILLER_38_2483 ();
 sg13g2_fill_1 FILLER_38_2490 ();
 sg13g2_decap_4 FILLER_38_2494 ();
 sg13g2_fill_1 FILLER_38_2498 ();
 sg13g2_fill_2 FILLER_38_2512 ();
 sg13g2_fill_1 FILLER_38_2514 ();
 sg13g2_decap_4 FILLER_38_2546 ();
 sg13g2_fill_1 FILLER_38_2550 ();
 sg13g2_decap_8 FILLER_38_2560 ();
 sg13g2_decap_8 FILLER_38_2567 ();
 sg13g2_fill_2 FILLER_38_2632 ();
 sg13g2_decap_8 FILLER_38_2655 ();
 sg13g2_decap_8 FILLER_38_2662 ();
 sg13g2_fill_1 FILLER_38_2669 ();
 sg13g2_decap_4 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_98 ();
 sg13g2_decap_8 FILLER_39_105 ();
 sg13g2_decap_8 FILLER_39_112 ();
 sg13g2_decap_8 FILLER_39_119 ();
 sg13g2_fill_2 FILLER_39_126 ();
 sg13g2_fill_1 FILLER_39_128 ();
 sg13g2_fill_2 FILLER_39_142 ();
 sg13g2_fill_2 FILLER_39_173 ();
 sg13g2_fill_1 FILLER_39_178 ();
 sg13g2_decap_8 FILLER_39_191 ();
 sg13g2_decap_8 FILLER_39_198 ();
 sg13g2_decap_4 FILLER_39_205 ();
 sg13g2_fill_1 FILLER_39_212 ();
 sg13g2_decap_8 FILLER_39_229 ();
 sg13g2_decap_4 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_240 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_decap_4 FILLER_39_252 ();
 sg13g2_fill_1 FILLER_39_256 ();
 sg13g2_decap_8 FILLER_39_283 ();
 sg13g2_decap_4 FILLER_39_290 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_decap_4 FILLER_39_329 ();
 sg13g2_fill_1 FILLER_39_333 ();
 sg13g2_fill_1 FILLER_39_342 ();
 sg13g2_decap_8 FILLER_39_359 ();
 sg13g2_decap_4 FILLER_39_366 ();
 sg13g2_fill_2 FILLER_39_374 ();
 sg13g2_fill_1 FILLER_39_376 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_4 FILLER_39_396 ();
 sg13g2_fill_1 FILLER_39_400 ();
 sg13g2_decap_4 FILLER_39_419 ();
 sg13g2_fill_2 FILLER_39_423 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_39_482 ();
 sg13g2_decap_4 FILLER_39_489 ();
 sg13g2_fill_1 FILLER_39_493 ();
 sg13g2_fill_2 FILLER_39_498 ();
 sg13g2_fill_1 FILLER_39_500 ();
 sg13g2_decap_8 FILLER_39_504 ();
 sg13g2_fill_1 FILLER_39_511 ();
 sg13g2_fill_2 FILLER_39_530 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_4 FILLER_39_550 ();
 sg13g2_fill_2 FILLER_39_554 ();
 sg13g2_fill_2 FILLER_39_579 ();
 sg13g2_fill_1 FILLER_39_586 ();
 sg13g2_decap_4 FILLER_39_597 ();
 sg13g2_fill_2 FILLER_39_611 ();
 sg13g2_fill_1 FILLER_39_613 ();
 sg13g2_fill_1 FILLER_39_624 ();
 sg13g2_fill_1 FILLER_39_629 ();
 sg13g2_decap_4 FILLER_39_637 ();
 sg13g2_decap_8 FILLER_39_659 ();
 sg13g2_fill_1 FILLER_39_666 ();
 sg13g2_fill_2 FILLER_39_697 ();
 sg13g2_fill_1 FILLER_39_720 ();
 sg13g2_fill_1 FILLER_39_726 ();
 sg13g2_fill_1 FILLER_39_734 ();
 sg13g2_fill_2 FILLER_39_743 ();
 sg13g2_fill_2 FILLER_39_752 ();
 sg13g2_decap_8 FILLER_39_767 ();
 sg13g2_decap_8 FILLER_39_782 ();
 sg13g2_decap_8 FILLER_39_789 ();
 sg13g2_fill_1 FILLER_39_796 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_4 FILLER_39_809 ();
 sg13g2_fill_1 FILLER_39_813 ();
 sg13g2_decap_8 FILLER_39_819 ();
 sg13g2_decap_4 FILLER_39_826 ();
 sg13g2_decap_8 FILLER_39_897 ();
 sg13g2_decap_8 FILLER_39_904 ();
 sg13g2_decap_8 FILLER_39_911 ();
 sg13g2_fill_2 FILLER_39_918 ();
 sg13g2_fill_1 FILLER_39_920 ();
 sg13g2_decap_4 FILLER_39_926 ();
 sg13g2_fill_1 FILLER_39_930 ();
 sg13g2_fill_2 FILLER_39_966 ();
 sg13g2_fill_1 FILLER_39_972 ();
 sg13g2_fill_2 FILLER_39_985 ();
 sg13g2_fill_1 FILLER_39_996 ();
 sg13g2_fill_1 FILLER_39_1036 ();
 sg13g2_fill_2 FILLER_39_1045 ();
 sg13g2_fill_1 FILLER_39_1073 ();
 sg13g2_fill_2 FILLER_39_1082 ();
 sg13g2_fill_1 FILLER_39_1084 ();
 sg13g2_decap_8 FILLER_39_1090 ();
 sg13g2_fill_2 FILLER_39_1097 ();
 sg13g2_fill_2 FILLER_39_1109 ();
 sg13g2_decap_4 FILLER_39_1124 ();
 sg13g2_fill_2 FILLER_39_1128 ();
 sg13g2_decap_8 FILLER_39_1172 ();
 sg13g2_fill_2 FILLER_39_1179 ();
 sg13g2_decap_4 FILLER_39_1185 ();
 sg13g2_fill_1 FILLER_39_1189 ();
 sg13g2_decap_8 FILLER_39_1196 ();
 sg13g2_decap_8 FILLER_39_1211 ();
 sg13g2_fill_1 FILLER_39_1227 ();
 sg13g2_decap_4 FILLER_39_1234 ();
 sg13g2_fill_2 FILLER_39_1249 ();
 sg13g2_fill_1 FILLER_39_1259 ();
 sg13g2_decap_4 FILLER_39_1265 ();
 sg13g2_decap_8 FILLER_39_1279 ();
 sg13g2_fill_2 FILLER_39_1295 ();
 sg13g2_fill_2 FILLER_39_1308 ();
 sg13g2_fill_1 FILLER_39_1310 ();
 sg13g2_fill_1 FILLER_39_1337 ();
 sg13g2_decap_4 FILLER_39_1374 ();
 sg13g2_fill_2 FILLER_39_1378 ();
 sg13g2_fill_1 FILLER_39_1419 ();
 sg13g2_fill_2 FILLER_39_1470 ();
 sg13g2_decap_8 FILLER_39_1485 ();
 sg13g2_decap_4 FILLER_39_1492 ();
 sg13g2_fill_2 FILLER_39_1501 ();
 sg13g2_decap_4 FILLER_39_1525 ();
 sg13g2_fill_1 FILLER_39_1529 ();
 sg13g2_fill_2 FILLER_39_1552 ();
 sg13g2_fill_1 FILLER_39_1554 ();
 sg13g2_fill_2 FILLER_39_1579 ();
 sg13g2_decap_4 FILLER_39_1591 ();
 sg13g2_fill_1 FILLER_39_1595 ();
 sg13g2_decap_8 FILLER_39_1601 ();
 sg13g2_fill_2 FILLER_39_1608 ();
 sg13g2_fill_1 FILLER_39_1610 ();
 sg13g2_decap_8 FILLER_39_1619 ();
 sg13g2_decap_4 FILLER_39_1626 ();
 sg13g2_decap_8 FILLER_39_1643 ();
 sg13g2_decap_8 FILLER_39_1650 ();
 sg13g2_fill_1 FILLER_39_1657 ();
 sg13g2_fill_2 FILLER_39_1665 ();
 sg13g2_fill_2 FILLER_39_1730 ();
 sg13g2_decap_4 FILLER_39_1745 ();
 sg13g2_fill_2 FILLER_39_1749 ();
 sg13g2_decap_8 FILLER_39_1763 ();
 sg13g2_decap_4 FILLER_39_1770 ();
 sg13g2_decap_8 FILLER_39_1778 ();
 sg13g2_fill_2 FILLER_39_1785 ();
 sg13g2_fill_2 FILLER_39_1835 ();
 sg13g2_fill_1 FILLER_39_1837 ();
 sg13g2_fill_2 FILLER_39_1842 ();
 sg13g2_fill_2 FILLER_39_1848 ();
 sg13g2_fill_1 FILLER_39_1850 ();
 sg13g2_fill_1 FILLER_39_1890 ();
 sg13g2_fill_2 FILLER_39_1895 ();
 sg13g2_fill_2 FILLER_39_1911 ();
 sg13g2_fill_1 FILLER_39_1913 ();
 sg13g2_fill_1 FILLER_39_1926 ();
 sg13g2_fill_1 FILLER_39_1945 ();
 sg13g2_fill_1 FILLER_39_1954 ();
 sg13g2_fill_2 FILLER_39_2007 ();
 sg13g2_decap_8 FILLER_39_2014 ();
 sg13g2_fill_2 FILLER_39_2039 ();
 sg13g2_fill_2 FILLER_39_2080 ();
 sg13g2_fill_1 FILLER_39_2082 ();
 sg13g2_fill_1 FILLER_39_2094 ();
 sg13g2_fill_2 FILLER_39_2099 ();
 sg13g2_fill_2 FILLER_39_2106 ();
 sg13g2_fill_1 FILLER_39_2118 ();
 sg13g2_fill_1 FILLER_39_2128 ();
 sg13g2_fill_1 FILLER_39_2133 ();
 sg13g2_fill_1 FILLER_39_2178 ();
 sg13g2_decap_4 FILLER_39_2189 ();
 sg13g2_fill_1 FILLER_39_2193 ();
 sg13g2_fill_1 FILLER_39_2199 ();
 sg13g2_fill_2 FILLER_39_2230 ();
 sg13g2_fill_1 FILLER_39_2232 ();
 sg13g2_decap_4 FILLER_39_2242 ();
 sg13g2_decap_8 FILLER_39_2331 ();
 sg13g2_decap_4 FILLER_39_2338 ();
 sg13g2_fill_2 FILLER_39_2342 ();
 sg13g2_decap_8 FILLER_39_2367 ();
 sg13g2_decap_8 FILLER_39_2374 ();
 sg13g2_fill_1 FILLER_39_2381 ();
 sg13g2_fill_1 FILLER_39_2387 ();
 sg13g2_fill_2 FILLER_39_2394 ();
 sg13g2_fill_1 FILLER_39_2396 ();
 sg13g2_decap_8 FILLER_39_2401 ();
 sg13g2_decap_4 FILLER_39_2408 ();
 sg13g2_fill_2 FILLER_39_2412 ();
 sg13g2_decap_4 FILLER_39_2418 ();
 sg13g2_fill_1 FILLER_39_2422 ();
 sg13g2_decap_8 FILLER_39_2428 ();
 sg13g2_fill_2 FILLER_39_2435 ();
 sg13g2_fill_1 FILLER_39_2437 ();
 sg13g2_decap_8 FILLER_39_2445 ();
 sg13g2_decap_4 FILLER_39_2452 ();
 sg13g2_fill_2 FILLER_39_2456 ();
 sg13g2_decap_8 FILLER_39_2488 ();
 sg13g2_decap_4 FILLER_39_2495 ();
 sg13g2_fill_1 FILLER_39_2538 ();
 sg13g2_fill_1 FILLER_39_2557 ();
 sg13g2_decap_4 FILLER_39_2638 ();
 sg13g2_fill_2 FILLER_39_2668 ();
 sg13g2_decap_4 FILLER_40_0 ();
 sg13g2_fill_1 FILLER_40_4 ();
 sg13g2_fill_1 FILLER_40_41 ();
 sg13g2_fill_2 FILLER_40_73 ();
 sg13g2_fill_2 FILLER_40_90 ();
 sg13g2_decap_8 FILLER_40_118 ();
 sg13g2_decap_8 FILLER_40_125 ();
 sg13g2_decap_8 FILLER_40_132 ();
 sg13g2_fill_2 FILLER_40_139 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_fill_1 FILLER_40_203 ();
 sg13g2_fill_2 FILLER_40_230 ();
 sg13g2_decap_4 FILLER_40_272 ();
 sg13g2_fill_2 FILLER_40_276 ();
 sg13g2_decap_4 FILLER_40_281 ();
 sg13g2_fill_2 FILLER_40_285 ();
 sg13g2_fill_1 FILLER_40_292 ();
 sg13g2_decap_4 FILLER_40_298 ();
 sg13g2_fill_2 FILLER_40_306 ();
 sg13g2_decap_8 FILLER_40_318 ();
 sg13g2_decap_8 FILLER_40_325 ();
 sg13g2_decap_8 FILLER_40_332 ();
 sg13g2_decap_8 FILLER_40_339 ();
 sg13g2_decap_8 FILLER_40_346 ();
 sg13g2_decap_8 FILLER_40_353 ();
 sg13g2_decap_4 FILLER_40_360 ();
 sg13g2_fill_1 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_374 ();
 sg13g2_fill_2 FILLER_40_381 ();
 sg13g2_decap_4 FILLER_40_388 ();
 sg13g2_decap_8 FILLER_40_405 ();
 sg13g2_decap_8 FILLER_40_412 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_2 FILLER_40_438 ();
 sg13g2_fill_1 FILLER_40_445 ();
 sg13g2_fill_1 FILLER_40_450 ();
 sg13g2_fill_1 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_471 ();
 sg13g2_fill_1 FILLER_40_478 ();
 sg13g2_decap_4 FILLER_40_488 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_fill_1 FILLER_40_563 ();
 sg13g2_fill_2 FILLER_40_568 ();
 sg13g2_decap_4 FILLER_40_577 ();
 sg13g2_fill_1 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_586 ();
 sg13g2_decap_8 FILLER_40_593 ();
 sg13g2_decap_8 FILLER_40_600 ();
 sg13g2_decap_4 FILLER_40_607 ();
 sg13g2_fill_1 FILLER_40_611 ();
 sg13g2_decap_4 FILLER_40_622 ();
 sg13g2_fill_2 FILLER_40_626 ();
 sg13g2_fill_1 FILLER_40_649 ();
 sg13g2_decap_8 FILLER_40_653 ();
 sg13g2_decap_8 FILLER_40_660 ();
 sg13g2_decap_8 FILLER_40_667 ();
 sg13g2_decap_8 FILLER_40_674 ();
 sg13g2_fill_1 FILLER_40_714 ();
 sg13g2_fill_2 FILLER_40_723 ();
 sg13g2_fill_1 FILLER_40_738 ();
 sg13g2_fill_2 FILLER_40_744 ();
 sg13g2_fill_2 FILLER_40_757 ();
 sg13g2_fill_2 FILLER_40_785 ();
 sg13g2_decap_4 FILLER_40_791 ();
 sg13g2_fill_2 FILLER_40_821 ();
 sg13g2_fill_1 FILLER_40_862 ();
 sg13g2_fill_2 FILLER_40_869 ();
 sg13g2_fill_1 FILLER_40_880 ();
 sg13g2_decap_4 FILLER_40_912 ();
 sg13g2_fill_1 FILLER_40_916 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_fill_1 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_1000 ();
 sg13g2_decap_8 FILLER_40_1007 ();
 sg13g2_decap_4 FILLER_40_1014 ();
 sg13g2_fill_1 FILLER_40_1018 ();
 sg13g2_decap_8 FILLER_40_1040 ();
 sg13g2_decap_8 FILLER_40_1047 ();
 sg13g2_decap_8 FILLER_40_1060 ();
 sg13g2_decap_8 FILLER_40_1067 ();
 sg13g2_fill_2 FILLER_40_1087 ();
 sg13g2_fill_1 FILLER_40_1089 ();
 sg13g2_fill_1 FILLER_40_1121 ();
 sg13g2_decap_4 FILLER_40_1127 ();
 sg13g2_fill_1 FILLER_40_1131 ();
 sg13g2_fill_1 FILLER_40_1136 ();
 sg13g2_fill_1 FILLER_40_1141 ();
 sg13g2_fill_2 FILLER_40_1152 ();
 sg13g2_fill_1 FILLER_40_1189 ();
 sg13g2_fill_2 FILLER_40_1236 ();
 sg13g2_fill_1 FILLER_40_1238 ();
 sg13g2_decap_8 FILLER_40_1245 ();
 sg13g2_decap_4 FILLER_40_1252 ();
 sg13g2_fill_1 FILLER_40_1256 ();
 sg13g2_fill_2 FILLER_40_1261 ();
 sg13g2_decap_8 FILLER_40_1289 ();
 sg13g2_decap_8 FILLER_40_1350 ();
 sg13g2_decap_4 FILLER_40_1357 ();
 sg13g2_fill_2 FILLER_40_1361 ();
 sg13g2_decap_8 FILLER_40_1367 ();
 sg13g2_decap_4 FILLER_40_1374 ();
 sg13g2_fill_2 FILLER_40_1378 ();
 sg13g2_decap_8 FILLER_40_1420 ();
 sg13g2_decap_4 FILLER_40_1427 ();
 sg13g2_fill_2 FILLER_40_1431 ();
 sg13g2_fill_2 FILLER_40_1443 ();
 sg13g2_fill_1 FILLER_40_1445 ();
 sg13g2_fill_1 FILLER_40_1450 ();
 sg13g2_fill_1 FILLER_40_1505 ();
 sg13g2_decap_8 FILLER_40_1513 ();
 sg13g2_fill_1 FILLER_40_1520 ();
 sg13g2_fill_1 FILLER_40_1536 ();
 sg13g2_fill_2 FILLER_40_1542 ();
 sg13g2_fill_2 FILLER_40_1563 ();
 sg13g2_decap_4 FILLER_40_1574 ();
 sg13g2_fill_2 FILLER_40_1578 ();
 sg13g2_decap_8 FILLER_40_1595 ();
 sg13g2_decap_8 FILLER_40_1602 ();
 sg13g2_fill_2 FILLER_40_1609 ();
 sg13g2_decap_8 FILLER_40_1619 ();
 sg13g2_decap_8 FILLER_40_1626 ();
 sg13g2_decap_8 FILLER_40_1633 ();
 sg13g2_decap_4 FILLER_40_1640 ();
 sg13g2_decap_8 FILLER_40_1649 ();
 sg13g2_decap_4 FILLER_40_1656 ();
 sg13g2_decap_8 FILLER_40_1673 ();
 sg13g2_fill_2 FILLER_40_1685 ();
 sg13g2_fill_1 FILLER_40_1687 ();
 sg13g2_fill_2 FILLER_40_1702 ();
 sg13g2_fill_1 FILLER_40_1713 ();
 sg13g2_fill_1 FILLER_40_1718 ();
 sg13g2_fill_1 FILLER_40_1728 ();
 sg13g2_decap_8 FILLER_40_1734 ();
 sg13g2_decap_8 FILLER_40_1741 ();
 sg13g2_decap_8 FILLER_40_1748 ();
 sg13g2_decap_8 FILLER_40_1755 ();
 sg13g2_decap_4 FILLER_40_1762 ();
 sg13g2_fill_1 FILLER_40_1766 ();
 sg13g2_decap_8 FILLER_40_1772 ();
 sg13g2_decap_8 FILLER_40_1779 ();
 sg13g2_decap_8 FILLER_40_1786 ();
 sg13g2_decap_4 FILLER_40_1793 ();
 sg13g2_fill_1 FILLER_40_1797 ();
 sg13g2_fill_2 FILLER_40_1807 ();
 sg13g2_fill_2 FILLER_40_1814 ();
 sg13g2_fill_1 FILLER_40_1816 ();
 sg13g2_decap_4 FILLER_40_1822 ();
 sg13g2_fill_1 FILLER_40_1862 ();
 sg13g2_decap_8 FILLER_40_1872 ();
 sg13g2_decap_4 FILLER_40_1879 ();
 sg13g2_fill_1 FILLER_40_1883 ();
 sg13g2_decap_8 FILLER_40_1894 ();
 sg13g2_decap_8 FILLER_40_1939 ();
 sg13g2_fill_2 FILLER_40_1946 ();
 sg13g2_fill_1 FILLER_40_1948 ();
 sg13g2_decap_4 FILLER_40_1966 ();
 sg13g2_fill_2 FILLER_40_1970 ();
 sg13g2_decap_4 FILLER_40_1981 ();
 sg13g2_fill_2 FILLER_40_1985 ();
 sg13g2_decap_4 FILLER_40_1991 ();
 sg13g2_fill_2 FILLER_40_1995 ();
 sg13g2_decap_8 FILLER_40_2003 ();
 sg13g2_decap_8 FILLER_40_2010 ();
 sg13g2_decap_8 FILLER_40_2017 ();
 sg13g2_fill_2 FILLER_40_2024 ();
 sg13g2_fill_1 FILLER_40_2026 ();
 sg13g2_fill_1 FILLER_40_2031 ();
 sg13g2_fill_1 FILLER_40_2043 ();
 sg13g2_decap_8 FILLER_40_2063 ();
 sg13g2_decap_8 FILLER_40_2070 ();
 sg13g2_fill_2 FILLER_40_2077 ();
 sg13g2_decap_4 FILLER_40_2088 ();
 sg13g2_fill_1 FILLER_40_2092 ();
 sg13g2_decap_4 FILLER_40_2098 ();
 sg13g2_fill_2 FILLER_40_2107 ();
 sg13g2_fill_1 FILLER_40_2109 ();
 sg13g2_decap_4 FILLER_40_2116 ();
 sg13g2_fill_2 FILLER_40_2124 ();
 sg13g2_decap_4 FILLER_40_2134 ();
 sg13g2_decap_4 FILLER_40_2188 ();
 sg13g2_fill_2 FILLER_40_2192 ();
 sg13g2_decap_8 FILLER_40_2204 ();
 sg13g2_fill_2 FILLER_40_2223 ();
 sg13g2_decap_4 FILLER_40_2228 ();
 sg13g2_decap_4 FILLER_40_2237 ();
 sg13g2_fill_1 FILLER_40_2241 ();
 sg13g2_decap_8 FILLER_40_2251 ();
 sg13g2_decap_8 FILLER_40_2258 ();
 sg13g2_decap_8 FILLER_40_2265 ();
 sg13g2_decap_8 FILLER_40_2272 ();
 sg13g2_decap_8 FILLER_40_2279 ();
 sg13g2_decap_4 FILLER_40_2286 ();
 sg13g2_decap_4 FILLER_40_2296 ();
 sg13g2_fill_2 FILLER_40_2300 ();
 sg13g2_fill_1 FILLER_40_2306 ();
 sg13g2_fill_1 FILLER_40_2333 ();
 sg13g2_decap_8 FILLER_40_2338 ();
 sg13g2_decap_8 FILLER_40_2345 ();
 sg13g2_decap_8 FILLER_40_2352 ();
 sg13g2_decap_8 FILLER_40_2359 ();
 sg13g2_decap_4 FILLER_40_2374 ();
 sg13g2_fill_1 FILLER_40_2378 ();
 sg13g2_fill_1 FILLER_40_2388 ();
 sg13g2_decap_4 FILLER_40_2394 ();
 sg13g2_fill_1 FILLER_40_2398 ();
 sg13g2_decap_4 FILLER_40_2403 ();
 sg13g2_fill_2 FILLER_40_2407 ();
 sg13g2_fill_2 FILLER_40_2413 ();
 sg13g2_fill_1 FILLER_40_2415 ();
 sg13g2_decap_8 FILLER_40_2420 ();
 sg13g2_decap_8 FILLER_40_2427 ();
 sg13g2_fill_1 FILLER_40_2434 ();
 sg13g2_fill_2 FILLER_40_2441 ();
 sg13g2_fill_2 FILLER_40_2447 ();
 sg13g2_fill_2 FILLER_40_2462 ();
 sg13g2_fill_1 FILLER_40_2464 ();
 sg13g2_fill_2 FILLER_40_2474 ();
 sg13g2_fill_1 FILLER_40_2476 ();
 sg13g2_decap_8 FILLER_40_2481 ();
 sg13g2_decap_4 FILLER_40_2488 ();
 sg13g2_fill_2 FILLER_40_2492 ();
 sg13g2_fill_2 FILLER_40_2501 ();
 sg13g2_decap_8 FILLER_40_2599 ();
 sg13g2_fill_1 FILLER_40_2606 ();
 sg13g2_decap_8 FILLER_40_2659 ();
 sg13g2_decap_4 FILLER_40_2666 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_4 FILLER_41_7 ();
 sg13g2_decap_4 FILLER_41_37 ();
 sg13g2_fill_1 FILLER_41_41 ();
 sg13g2_fill_1 FILLER_41_52 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_4 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_82 ();
 sg13g2_decap_4 FILLER_41_89 ();
 sg13g2_fill_1 FILLER_41_93 ();
 sg13g2_decap_8 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_111 ();
 sg13g2_decap_8 FILLER_41_122 ();
 sg13g2_decap_8 FILLER_41_129 ();
 sg13g2_decap_8 FILLER_41_136 ();
 sg13g2_decap_4 FILLER_41_143 ();
 sg13g2_decap_8 FILLER_41_157 ();
 sg13g2_decap_8 FILLER_41_164 ();
 sg13g2_decap_8 FILLER_41_171 ();
 sg13g2_decap_8 FILLER_41_184 ();
 sg13g2_decap_8 FILLER_41_191 ();
 sg13g2_decap_4 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_212 ();
 sg13g2_fill_1 FILLER_41_214 ();
 sg13g2_fill_1 FILLER_41_248 ();
 sg13g2_decap_8 FILLER_41_272 ();
 sg13g2_fill_2 FILLER_41_279 ();
 sg13g2_fill_1 FILLER_41_294 ();
 sg13g2_fill_2 FILLER_41_321 ();
 sg13g2_decap_8 FILLER_41_328 ();
 sg13g2_decap_4 FILLER_41_335 ();
 sg13g2_decap_4 FILLER_41_374 ();
 sg13g2_fill_1 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_fill_1 FILLER_41_420 ();
 sg13g2_decap_4 FILLER_41_426 ();
 sg13g2_fill_2 FILLER_41_437 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_fill_1 FILLER_41_455 ();
 sg13g2_fill_1 FILLER_41_460 ();
 sg13g2_fill_2 FILLER_41_467 ();
 sg13g2_fill_1 FILLER_41_469 ();
 sg13g2_fill_2 FILLER_41_502 ();
 sg13g2_decap_8 FILLER_41_537 ();
 sg13g2_decap_8 FILLER_41_544 ();
 sg13g2_decap_8 FILLER_41_577 ();
 sg13g2_fill_2 FILLER_41_584 ();
 sg13g2_decap_8 FILLER_41_592 ();
 sg13g2_decap_8 FILLER_41_599 ();
 sg13g2_decap_4 FILLER_41_606 ();
 sg13g2_fill_2 FILLER_41_614 ();
 sg13g2_fill_2 FILLER_41_625 ();
 sg13g2_fill_1 FILLER_41_627 ();
 sg13g2_decap_8 FILLER_41_648 ();
 sg13g2_fill_2 FILLER_41_655 ();
 sg13g2_decap_4 FILLER_41_668 ();
 sg13g2_fill_1 FILLER_41_672 ();
 sg13g2_fill_2 FILLER_41_684 ();
 sg13g2_fill_2 FILLER_41_702 ();
 sg13g2_fill_1 FILLER_41_726 ();
 sg13g2_fill_2 FILLER_41_734 ();
 sg13g2_fill_1 FILLER_41_743 ();
 sg13g2_fill_1 FILLER_41_767 ();
 sg13g2_fill_2 FILLER_41_773 ();
 sg13g2_fill_1 FILLER_41_775 ();
 sg13g2_fill_2 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_824 ();
 sg13g2_decap_8 FILLER_41_831 ();
 sg13g2_decap_4 FILLER_41_838 ();
 sg13g2_fill_2 FILLER_41_842 ();
 sg13g2_decap_8 FILLER_41_853 ();
 sg13g2_fill_2 FILLER_41_860 ();
 sg13g2_decap_4 FILLER_41_868 ();
 sg13g2_fill_1 FILLER_41_872 ();
 sg13g2_fill_2 FILLER_41_883 ();
 sg13g2_fill_1 FILLER_41_885 ();
 sg13g2_fill_1 FILLER_41_923 ();
 sg13g2_fill_2 FILLER_41_959 ();
 sg13g2_fill_1 FILLER_41_961 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_989 ();
 sg13g2_decap_8 FILLER_41_996 ();
 sg13g2_decap_8 FILLER_41_1003 ();
 sg13g2_decap_8 FILLER_41_1010 ();
 sg13g2_decap_4 FILLER_41_1017 ();
 sg13g2_fill_2 FILLER_41_1021 ();
 sg13g2_fill_1 FILLER_41_1065 ();
 sg13g2_fill_2 FILLER_41_1071 ();
 sg13g2_fill_2 FILLER_41_1083 ();
 sg13g2_fill_1 FILLER_41_1085 ();
 sg13g2_decap_8 FILLER_41_1104 ();
 sg13g2_decap_8 FILLER_41_1111 ();
 sg13g2_decap_4 FILLER_41_1118 ();
 sg13g2_fill_1 FILLER_41_1122 ();
 sg13g2_decap_4 FILLER_41_1158 ();
 sg13g2_fill_2 FILLER_41_1165 ();
 sg13g2_fill_2 FILLER_41_1205 ();
 sg13g2_fill_1 FILLER_41_1213 ();
 sg13g2_fill_1 FILLER_41_1218 ();
 sg13g2_fill_2 FILLER_41_1228 ();
 sg13g2_fill_1 FILLER_41_1230 ();
 sg13g2_fill_2 FILLER_41_1237 ();
 sg13g2_fill_1 FILLER_41_1239 ();
 sg13g2_fill_2 FILLER_41_1258 ();
 sg13g2_fill_1 FILLER_41_1260 ();
 sg13g2_fill_2 FILLER_41_1292 ();
 sg13g2_fill_1 FILLER_41_1294 ();
 sg13g2_fill_2 FILLER_41_1304 ();
 sg13g2_fill_2 FILLER_41_1341 ();
 sg13g2_fill_2 FILLER_41_1369 ();
 sg13g2_decap_8 FILLER_41_1383 ();
 sg13g2_decap_8 FILLER_41_1390 ();
 sg13g2_fill_2 FILLER_41_1397 ();
 sg13g2_fill_2 FILLER_41_1411 ();
 sg13g2_decap_8 FILLER_41_1420 ();
 sg13g2_decap_8 FILLER_41_1427 ();
 sg13g2_decap_8 FILLER_41_1434 ();
 sg13g2_fill_2 FILLER_41_1441 ();
 sg13g2_fill_1 FILLER_41_1443 ();
 sg13g2_decap_4 FILLER_41_1449 ();
 sg13g2_fill_1 FILLER_41_1453 ();
 sg13g2_decap_8 FILLER_41_1457 ();
 sg13g2_fill_1 FILLER_41_1464 ();
 sg13g2_decap_4 FILLER_41_1473 ();
 sg13g2_fill_1 FILLER_41_1477 ();
 sg13g2_decap_8 FILLER_41_1482 ();
 sg13g2_decap_8 FILLER_41_1519 ();
 sg13g2_decap_8 FILLER_41_1526 ();
 sg13g2_fill_2 FILLER_41_1533 ();
 sg13g2_fill_1 FILLER_41_1535 ();
 sg13g2_fill_2 FILLER_41_1542 ();
 sg13g2_fill_1 FILLER_41_1549 ();
 sg13g2_decap_8 FILLER_41_1554 ();
 sg13g2_fill_1 FILLER_41_1561 ();
 sg13g2_decap_8 FILLER_41_1572 ();
 sg13g2_decap_4 FILLER_41_1579 ();
 sg13g2_fill_1 FILLER_41_1583 ();
 sg13g2_decap_8 FILLER_41_1619 ();
 sg13g2_decap_4 FILLER_41_1626 ();
 sg13g2_fill_1 FILLER_41_1630 ();
 sg13g2_decap_4 FILLER_41_1639 ();
 sg13g2_fill_1 FILLER_41_1643 ();
 sg13g2_decap_8 FILLER_41_1670 ();
 sg13g2_fill_1 FILLER_41_1677 ();
 sg13g2_decap_4 FILLER_41_1687 ();
 sg13g2_fill_2 FILLER_41_1691 ();
 sg13g2_fill_2 FILLER_41_1708 ();
 sg13g2_decap_4 FILLER_41_1740 ();
 sg13g2_fill_1 FILLER_41_1744 ();
 sg13g2_decap_4 FILLER_41_1750 ();
 sg13g2_fill_2 FILLER_41_1758 ();
 sg13g2_decap_8 FILLER_41_1764 ();
 sg13g2_decap_8 FILLER_41_1771 ();
 sg13g2_decap_8 FILLER_41_1778 ();
 sg13g2_decap_8 FILLER_41_1785 ();
 sg13g2_decap_8 FILLER_41_1792 ();
 sg13g2_decap_8 FILLER_41_1799 ();
 sg13g2_fill_1 FILLER_41_1806 ();
 sg13g2_fill_2 FILLER_41_1849 ();
 sg13g2_decap_4 FILLER_41_1859 ();
 sg13g2_fill_2 FILLER_41_1867 ();
 sg13g2_decap_4 FILLER_41_1877 ();
 sg13g2_fill_1 FILLER_41_1881 ();
 sg13g2_fill_1 FILLER_41_1901 ();
 sg13g2_fill_2 FILLER_41_1907 ();
 sg13g2_decap_4 FILLER_41_1913 ();
 sg13g2_decap_8 FILLER_41_1923 ();
 sg13g2_fill_2 FILLER_41_1930 ();
 sg13g2_fill_2 FILLER_41_1958 ();
 sg13g2_fill_1 FILLER_41_1960 ();
 sg13g2_decap_8 FILLER_41_1992 ();
 sg13g2_fill_2 FILLER_41_1999 ();
 sg13g2_fill_1 FILLER_41_2001 ();
 sg13g2_decap_4 FILLER_41_2007 ();
 sg13g2_fill_2 FILLER_41_2011 ();
 sg13g2_fill_2 FILLER_41_2025 ();
 sg13g2_fill_1 FILLER_41_2030 ();
 sg13g2_decap_8 FILLER_41_2067 ();
 sg13g2_decap_8 FILLER_41_2074 ();
 sg13g2_fill_2 FILLER_41_2081 ();
 sg13g2_fill_1 FILLER_41_2083 ();
 sg13g2_fill_2 FILLER_41_2087 ();
 sg13g2_decap_8 FILLER_41_2107 ();
 sg13g2_decap_8 FILLER_41_2114 ();
 sg13g2_decap_8 FILLER_41_2121 ();
 sg13g2_decap_8 FILLER_41_2132 ();
 sg13g2_fill_2 FILLER_41_2145 ();
 sg13g2_fill_1 FILLER_41_2147 ();
 sg13g2_fill_1 FILLER_41_2184 ();
 sg13g2_fill_1 FILLER_41_2195 ();
 sg13g2_fill_2 FILLER_41_2235 ();
 sg13g2_fill_1 FILLER_41_2237 ();
 sg13g2_decap_8 FILLER_41_2278 ();
 sg13g2_decap_8 FILLER_41_2285 ();
 sg13g2_decap_4 FILLER_41_2297 ();
 sg13g2_decap_8 FILLER_41_2321 ();
 sg13g2_fill_2 FILLER_41_2328 ();
 sg13g2_fill_1 FILLER_41_2330 ();
 sg13g2_decap_8 FILLER_41_2363 ();
 sg13g2_decap_4 FILLER_41_2370 ();
 sg13g2_fill_1 FILLER_41_2374 ();
 sg13g2_fill_2 FILLER_41_2381 ();
 sg13g2_fill_2 FILLER_41_2399 ();
 sg13g2_fill_1 FILLER_41_2401 ();
 sg13g2_fill_2 FILLER_41_2428 ();
 sg13g2_decap_8 FILLER_41_2464 ();
 sg13g2_decap_8 FILLER_41_2471 ();
 sg13g2_decap_8 FILLER_41_2478 ();
 sg13g2_fill_2 FILLER_41_2485 ();
 sg13g2_fill_1 FILLER_41_2487 ();
 sg13g2_decap_8 FILLER_41_2493 ();
 sg13g2_fill_2 FILLER_41_2500 ();
 sg13g2_decap_8 FILLER_41_2540 ();
 sg13g2_fill_1 FILLER_41_2551 ();
 sg13g2_fill_2 FILLER_41_2556 ();
 sg13g2_decap_8 FILLER_41_2584 ();
 sg13g2_decap_8 FILLER_41_2591 ();
 sg13g2_decap_8 FILLER_41_2598 ();
 sg13g2_decap_8 FILLER_41_2605 ();
 sg13g2_decap_8 FILLER_41_2612 ();
 sg13g2_fill_2 FILLER_41_2619 ();
 sg13g2_decap_8 FILLER_41_2643 ();
 sg13g2_decap_8 FILLER_41_2650 ();
 sg13g2_decap_8 FILLER_41_2657 ();
 sg13g2_decap_4 FILLER_41_2664 ();
 sg13g2_fill_2 FILLER_41_2668 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_52 ();
 sg13g2_decap_8 FILLER_42_59 ();
 sg13g2_decap_8 FILLER_42_66 ();
 sg13g2_decap_8 FILLER_42_73 ();
 sg13g2_decap_8 FILLER_42_80 ();
 sg13g2_decap_8 FILLER_42_87 ();
 sg13g2_decap_8 FILLER_42_94 ();
 sg13g2_decap_8 FILLER_42_101 ();
 sg13g2_fill_1 FILLER_42_108 ();
 sg13g2_decap_8 FILLER_42_135 ();
 sg13g2_decap_4 FILLER_42_142 ();
 sg13g2_fill_2 FILLER_42_146 ();
 sg13g2_fill_2 FILLER_42_187 ();
 sg13g2_fill_1 FILLER_42_225 ();
 sg13g2_fill_1 FILLER_42_234 ();
 sg13g2_fill_2 FILLER_42_242 ();
 sg13g2_fill_1 FILLER_42_244 ();
 sg13g2_fill_1 FILLER_42_284 ();
 sg13g2_fill_1 FILLER_42_308 ();
 sg13g2_decap_8 FILLER_42_322 ();
 sg13g2_decap_8 FILLER_42_329 ();
 sg13g2_decap_8 FILLER_42_336 ();
 sg13g2_decap_4 FILLER_42_343 ();
 sg13g2_decap_8 FILLER_42_350 ();
 sg13g2_decap_8 FILLER_42_357 ();
 sg13g2_decap_4 FILLER_42_364 ();
 sg13g2_fill_1 FILLER_42_373 ();
 sg13g2_decap_4 FILLER_42_408 ();
 sg13g2_fill_1 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_fill_1 FILLER_42_424 ();
 sg13g2_fill_1 FILLER_42_430 ();
 sg13g2_fill_2 FILLER_42_440 ();
 sg13g2_fill_1 FILLER_42_442 ();
 sg13g2_fill_1 FILLER_42_469 ();
 sg13g2_decap_4 FILLER_42_545 ();
 sg13g2_fill_1 FILLER_42_549 ();
 sg13g2_decap_8 FILLER_42_565 ();
 sg13g2_decap_8 FILLER_42_572 ();
 sg13g2_decap_8 FILLER_42_579 ();
 sg13g2_fill_2 FILLER_42_586 ();
 sg13g2_fill_1 FILLER_42_588 ();
 sg13g2_decap_4 FILLER_42_609 ();
 sg13g2_fill_1 FILLER_42_613 ();
 sg13g2_decap_4 FILLER_42_618 ();
 sg13g2_fill_1 FILLER_42_636 ();
 sg13g2_fill_1 FILLER_42_640 ();
 sg13g2_decap_8 FILLER_42_646 ();
 sg13g2_decap_8 FILLER_42_653 ();
 sg13g2_decap_8 FILLER_42_660 ();
 sg13g2_fill_2 FILLER_42_667 ();
 sg13g2_decap_4 FILLER_42_674 ();
 sg13g2_fill_1 FILLER_42_683 ();
 sg13g2_fill_1 FILLER_42_735 ();
 sg13g2_decap_4 FILLER_42_739 ();
 sg13g2_fill_1 FILLER_42_743 ();
 sg13g2_fill_1 FILLER_42_747 ();
 sg13g2_decap_4 FILLER_42_782 ();
 sg13g2_fill_1 FILLER_42_786 ();
 sg13g2_fill_2 FILLER_42_792 ();
 sg13g2_decap_8 FILLER_42_798 ();
 sg13g2_decap_8 FILLER_42_805 ();
 sg13g2_decap_8 FILLER_42_812 ();
 sg13g2_decap_4 FILLER_42_819 ();
 sg13g2_fill_1 FILLER_42_828 ();
 sg13g2_fill_2 FILLER_42_833 ();
 sg13g2_fill_1 FILLER_42_835 ();
 sg13g2_decap_4 FILLER_42_840 ();
 sg13g2_fill_2 FILLER_42_844 ();
 sg13g2_decap_4 FILLER_42_855 ();
 sg13g2_fill_2 FILLER_42_859 ();
 sg13g2_decap_8 FILLER_42_864 ();
 sg13g2_decap_4 FILLER_42_871 ();
 sg13g2_fill_2 FILLER_42_875 ();
 sg13g2_decap_8 FILLER_42_917 ();
 sg13g2_decap_8 FILLER_42_934 ();
 sg13g2_fill_2 FILLER_42_941 ();
 sg13g2_fill_1 FILLER_42_943 ();
 sg13g2_decap_8 FILLER_42_948 ();
 sg13g2_fill_2 FILLER_42_955 ();
 sg13g2_decap_4 FILLER_42_962 ();
 sg13g2_decap_8 FILLER_42_995 ();
 sg13g2_fill_2 FILLER_42_1002 ();
 sg13g2_decap_8 FILLER_42_1056 ();
 sg13g2_fill_1 FILLER_42_1093 ();
 sg13g2_decap_8 FILLER_42_1107 ();
 sg13g2_fill_1 FILLER_42_1114 ();
 sg13g2_fill_2 FILLER_42_1124 ();
 sg13g2_fill_2 FILLER_42_1129 ();
 sg13g2_fill_2 FILLER_42_1157 ();
 sg13g2_fill_2 FILLER_42_1183 ();
 sg13g2_fill_2 FILLER_42_1211 ();
 sg13g2_fill_2 FILLER_42_1254 ();
 sg13g2_fill_1 FILLER_42_1256 ();
 sg13g2_decap_8 FILLER_42_1262 ();
 sg13g2_fill_2 FILLER_42_1269 ();
 sg13g2_decap_8 FILLER_42_1307 ();
 sg13g2_decap_8 FILLER_42_1330 ();
 sg13g2_decap_8 FILLER_42_1337 ();
 sg13g2_decap_4 FILLER_42_1344 ();
 sg13g2_decap_4 FILLER_42_1353 ();
 sg13g2_decap_4 FILLER_42_1361 ();
 sg13g2_fill_2 FILLER_42_1365 ();
 sg13g2_decap_8 FILLER_42_1379 ();
 sg13g2_decap_4 FILLER_42_1391 ();
 sg13g2_decap_8 FILLER_42_1399 ();
 sg13g2_fill_2 FILLER_42_1406 ();
 sg13g2_decap_8 FILLER_42_1470 ();
 sg13g2_decap_8 FILLER_42_1477 ();
 sg13g2_decap_8 FILLER_42_1484 ();
 sg13g2_decap_4 FILLER_42_1491 ();
 sg13g2_fill_1 FILLER_42_1495 ();
 sg13g2_decap_8 FILLER_42_1505 ();
 sg13g2_decap_8 FILLER_42_1512 ();
 sg13g2_decap_8 FILLER_42_1519 ();
 sg13g2_fill_1 FILLER_42_1526 ();
 sg13g2_decap_4 FILLER_42_1531 ();
 sg13g2_fill_2 FILLER_42_1535 ();
 sg13g2_decap_8 FILLER_42_1552 ();
 sg13g2_decap_8 FILLER_42_1559 ();
 sg13g2_fill_1 FILLER_42_1566 ();
 sg13g2_decap_8 FILLER_42_1576 ();
 sg13g2_fill_1 FILLER_42_1583 ();
 sg13g2_fill_2 FILLER_42_1628 ();
 sg13g2_fill_2 FILLER_42_1635 ();
 sg13g2_fill_1 FILLER_42_1637 ();
 sg13g2_decap_8 FILLER_42_1643 ();
 sg13g2_decap_4 FILLER_42_1650 ();
 sg13g2_fill_1 FILLER_42_1654 ();
 sg13g2_decap_8 FILLER_42_1662 ();
 sg13g2_decap_4 FILLER_42_1669 ();
 sg13g2_fill_1 FILLER_42_1673 ();
 sg13g2_fill_2 FILLER_42_1679 ();
 sg13g2_fill_1 FILLER_42_1681 ();
 sg13g2_decap_8 FILLER_42_1739 ();
 sg13g2_fill_1 FILLER_42_1746 ();
 sg13g2_fill_2 FILLER_42_1785 ();
 sg13g2_fill_1 FILLER_42_1794 ();
 sg13g2_decap_8 FILLER_42_1798 ();
 sg13g2_decap_4 FILLER_42_1805 ();
 sg13g2_fill_1 FILLER_42_1809 ();
 sg13g2_fill_1 FILLER_42_1815 ();
 sg13g2_decap_4 FILLER_42_1830 ();
 sg13g2_fill_1 FILLER_42_1834 ();
 sg13g2_decap_4 FILLER_42_1839 ();
 sg13g2_decap_4 FILLER_42_1846 ();
 sg13g2_fill_2 FILLER_42_1850 ();
 sg13g2_decap_8 FILLER_42_1858 ();
 sg13g2_fill_1 FILLER_42_1865 ();
 sg13g2_fill_1 FILLER_42_1900 ();
 sg13g2_fill_1 FILLER_42_1932 ();
 sg13g2_decap_8 FILLER_42_1977 ();
 sg13g2_decap_8 FILLER_42_1984 ();
 sg13g2_fill_2 FILLER_42_1991 ();
 sg13g2_fill_1 FILLER_42_1993 ();
 sg13g2_decap_8 FILLER_42_1998 ();
 sg13g2_fill_1 FILLER_42_2005 ();
 sg13g2_decap_8 FILLER_42_2045 ();
 sg13g2_fill_2 FILLER_42_2052 ();
 sg13g2_fill_2 FILLER_42_2057 ();
 sg13g2_decap_4 FILLER_42_2074 ();
 sg13g2_fill_2 FILLER_42_2078 ();
 sg13g2_decap_4 FILLER_42_2115 ();
 sg13g2_fill_1 FILLER_42_2119 ();
 sg13g2_decap_8 FILLER_42_2138 ();
 sg13g2_decap_8 FILLER_42_2145 ();
 sg13g2_decap_4 FILLER_42_2152 ();
 sg13g2_fill_2 FILLER_42_2156 ();
 sg13g2_fill_2 FILLER_42_2162 ();
 sg13g2_decap_8 FILLER_42_2170 ();
 sg13g2_decap_8 FILLER_42_2177 ();
 sg13g2_decap_8 FILLER_42_2223 ();
 sg13g2_fill_1 FILLER_42_2230 ();
 sg13g2_fill_1 FILLER_42_2249 ();
 sg13g2_fill_1 FILLER_42_2269 ();
 sg13g2_decap_8 FILLER_42_2286 ();
 sg13g2_decap_8 FILLER_42_2293 ();
 sg13g2_decap_8 FILLER_42_2300 ();
 sg13g2_fill_2 FILLER_42_2307 ();
 sg13g2_decap_8 FILLER_42_2313 ();
 sg13g2_decap_8 FILLER_42_2320 ();
 sg13g2_decap_8 FILLER_42_2327 ();
 sg13g2_decap_8 FILLER_42_2334 ();
 sg13g2_fill_2 FILLER_42_2341 ();
 sg13g2_decap_8 FILLER_42_2373 ();
 sg13g2_fill_1 FILLER_42_2392 ();
 sg13g2_decap_8 FILLER_42_2397 ();
 sg13g2_decap_8 FILLER_42_2468 ();
 sg13g2_fill_1 FILLER_42_2475 ();
 sg13g2_decap_8 FILLER_42_2502 ();
 sg13g2_decap_4 FILLER_42_2513 ();
 sg13g2_fill_2 FILLER_42_2517 ();
 sg13g2_decap_8 FILLER_42_2527 ();
 sg13g2_decap_8 FILLER_42_2534 ();
 sg13g2_decap_8 FILLER_42_2541 ();
 sg13g2_decap_8 FILLER_42_2548 ();
 sg13g2_decap_4 FILLER_42_2555 ();
 sg13g2_fill_1 FILLER_42_2559 ();
 sg13g2_fill_1 FILLER_42_2568 ();
 sg13g2_decap_8 FILLER_42_2577 ();
 sg13g2_decap_8 FILLER_42_2584 ();
 sg13g2_decap_8 FILLER_42_2591 ();
 sg13g2_decap_8 FILLER_42_2598 ();
 sg13g2_decap_8 FILLER_42_2605 ();
 sg13g2_decap_8 FILLER_42_2612 ();
 sg13g2_decap_8 FILLER_42_2619 ();
 sg13g2_fill_1 FILLER_42_2626 ();
 sg13g2_decap_8 FILLER_42_2643 ();
 sg13g2_decap_8 FILLER_42_2650 ();
 sg13g2_decap_8 FILLER_42_2657 ();
 sg13g2_decap_4 FILLER_42_2664 ();
 sg13g2_fill_2 FILLER_42_2668 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_fill_1 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_39 ();
 sg13g2_decap_8 FILLER_43_46 ();
 sg13g2_decap_8 FILLER_43_53 ();
 sg13g2_decap_8 FILLER_43_101 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_decap_8 FILLER_43_115 ();
 sg13g2_decap_8 FILLER_43_122 ();
 sg13g2_fill_2 FILLER_43_129 ();
 sg13g2_fill_1 FILLER_43_131 ();
 sg13g2_decap_8 FILLER_43_158 ();
 sg13g2_fill_2 FILLER_43_165 ();
 sg13g2_fill_1 FILLER_43_203 ();
 sg13g2_fill_2 FILLER_43_207 ();
 sg13g2_decap_8 FILLER_43_212 ();
 sg13g2_decap_4 FILLER_43_219 ();
 sg13g2_fill_2 FILLER_43_223 ();
 sg13g2_decap_4 FILLER_43_233 ();
 sg13g2_fill_1 FILLER_43_237 ();
 sg13g2_fill_1 FILLER_43_249 ();
 sg13g2_fill_1 FILLER_43_263 ();
 sg13g2_decap_4 FILLER_43_269 ();
 sg13g2_fill_2 FILLER_43_273 ();
 sg13g2_fill_2 FILLER_43_312 ();
 sg13g2_decap_4 FILLER_43_318 ();
 sg13g2_fill_2 FILLER_43_348 ();
 sg13g2_fill_1 FILLER_43_350 ();
 sg13g2_fill_1 FILLER_43_398 ();
 sg13g2_fill_2 FILLER_43_403 ();
 sg13g2_fill_2 FILLER_43_410 ();
 sg13g2_fill_2 FILLER_43_416 ();
 sg13g2_fill_1 FILLER_43_418 ();
 sg13g2_fill_2 FILLER_43_445 ();
 sg13g2_fill_1 FILLER_43_447 ();
 sg13g2_decap_4 FILLER_43_453 ();
 sg13g2_fill_2 FILLER_43_457 ();
 sg13g2_fill_2 FILLER_43_463 ();
 sg13g2_fill_1 FILLER_43_484 ();
 sg13g2_fill_1 FILLER_43_526 ();
 sg13g2_fill_2 FILLER_43_531 ();
 sg13g2_decap_8 FILLER_43_537 ();
 sg13g2_decap_8 FILLER_43_544 ();
 sg13g2_decap_8 FILLER_43_551 ();
 sg13g2_decap_8 FILLER_43_558 ();
 sg13g2_decap_8 FILLER_43_565 ();
 sg13g2_decap_8 FILLER_43_572 ();
 sg13g2_decap_8 FILLER_43_579 ();
 sg13g2_decap_4 FILLER_43_597 ();
 sg13g2_fill_2 FILLER_43_601 ();
 sg13g2_fill_1 FILLER_43_614 ();
 sg13g2_fill_1 FILLER_43_620 ();
 sg13g2_decap_4 FILLER_43_627 ();
 sg13g2_fill_2 FILLER_43_650 ();
 sg13g2_fill_2 FILLER_43_657 ();
 sg13g2_fill_2 FILLER_43_664 ();
 sg13g2_fill_2 FILLER_43_680 ();
 sg13g2_fill_1 FILLER_43_682 ();
 sg13g2_fill_2 FILLER_43_691 ();
 sg13g2_fill_2 FILLER_43_727 ();
 sg13g2_fill_1 FILLER_43_729 ();
 sg13g2_decap_8 FILLER_43_734 ();
 sg13g2_decap_8 FILLER_43_741 ();
 sg13g2_decap_8 FILLER_43_748 ();
 sg13g2_decap_8 FILLER_43_755 ();
 sg13g2_decap_4 FILLER_43_767 ();
 sg13g2_decap_8 FILLER_43_775 ();
 sg13g2_decap_8 FILLER_43_782 ();
 sg13g2_fill_1 FILLER_43_828 ();
 sg13g2_fill_2 FILLER_43_855 ();
 sg13g2_fill_1 FILLER_43_857 ();
 sg13g2_fill_2 FILLER_43_864 ();
 sg13g2_fill_2 FILLER_43_914 ();
 sg13g2_fill_1 FILLER_43_916 ();
 sg13g2_fill_2 FILLER_43_930 ();
 sg13g2_fill_2 FILLER_43_972 ();
 sg13g2_decap_4 FILLER_43_978 ();
 sg13g2_fill_2 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_993 ();
 sg13g2_fill_2 FILLER_43_1000 ();
 sg13g2_fill_1 FILLER_43_1002 ();
 sg13g2_decap_4 FILLER_43_1012 ();
 sg13g2_fill_1 FILLER_43_1016 ();
 sg13g2_decap_8 FILLER_43_1023 ();
 sg13g2_fill_1 FILLER_43_1030 ();
 sg13g2_decap_4 FILLER_43_1039 ();
 sg13g2_fill_1 FILLER_43_1052 ();
 sg13g2_fill_1 FILLER_43_1062 ();
 sg13g2_fill_2 FILLER_43_1115 ();
 sg13g2_fill_1 FILLER_43_1117 ();
 sg13g2_decap_8 FILLER_43_1143 ();
 sg13g2_decap_8 FILLER_43_1154 ();
 sg13g2_fill_1 FILLER_43_1161 ();
 sg13g2_fill_2 FILLER_43_1172 ();
 sg13g2_fill_1 FILLER_43_1184 ();
 sg13g2_fill_2 FILLER_43_1189 ();
 sg13g2_decap_8 FILLER_43_1253 ();
 sg13g2_fill_2 FILLER_43_1260 ();
 sg13g2_fill_1 FILLER_43_1262 ();
 sg13g2_fill_2 FILLER_43_1297 ();
 sg13g2_fill_1 FILLER_43_1299 ();
 sg13g2_fill_2 FILLER_43_1309 ();
 sg13g2_decap_8 FILLER_43_1337 ();
 sg13g2_decap_8 FILLER_43_1344 ();
 sg13g2_decap_8 FILLER_43_1351 ();
 sg13g2_decap_8 FILLER_43_1358 ();
 sg13g2_fill_2 FILLER_43_1365 ();
 sg13g2_fill_1 FILLER_43_1367 ();
 sg13g2_decap_8 FILLER_43_1373 ();
 sg13g2_decap_4 FILLER_43_1380 ();
 sg13g2_fill_2 FILLER_43_1384 ();
 sg13g2_fill_1 FILLER_43_1390 ();
 sg13g2_decap_8 FILLER_43_1443 ();
 sg13g2_decap_4 FILLER_43_1450 ();
 sg13g2_fill_1 FILLER_43_1454 ();
 sg13g2_decap_4 FILLER_43_1459 ();
 sg13g2_fill_2 FILLER_43_1463 ();
 sg13g2_decap_8 FILLER_43_1473 ();
 sg13g2_decap_8 FILLER_43_1480 ();
 sg13g2_decap_4 FILLER_43_1487 ();
 sg13g2_fill_2 FILLER_43_1491 ();
 sg13g2_decap_8 FILLER_43_1540 ();
 sg13g2_decap_8 FILLER_43_1573 ();
 sg13g2_decap_4 FILLER_43_1580 ();
 sg13g2_decap_8 FILLER_43_1706 ();
 sg13g2_decap_8 FILLER_43_1713 ();
 sg13g2_fill_1 FILLER_43_1720 ();
 sg13g2_fill_1 FILLER_43_1726 ();
 sg13g2_fill_2 FILLER_43_1733 ();
 sg13g2_fill_2 FILLER_43_1761 ();
 sg13g2_fill_1 FILLER_43_1770 ();
 sg13g2_fill_2 FILLER_43_1828 ();
 sg13g2_fill_2 FILLER_43_1840 ();
 sg13g2_fill_1 FILLER_43_1842 ();
 sg13g2_decap_4 FILLER_43_1854 ();
 sg13g2_fill_1 FILLER_43_1858 ();
 sg13g2_fill_1 FILLER_43_1864 ();
 sg13g2_fill_1 FILLER_43_1897 ();
 sg13g2_decap_4 FILLER_43_1904 ();
 sg13g2_decap_8 FILLER_43_1916 ();
 sg13g2_decap_8 FILLER_43_1923 ();
 sg13g2_decap_8 FILLER_43_1930 ();
 sg13g2_decap_8 FILLER_43_1941 ();
 sg13g2_fill_2 FILLER_43_1948 ();
 sg13g2_fill_1 FILLER_43_1950 ();
 sg13g2_fill_1 FILLER_43_1957 ();
 sg13g2_decap_4 FILLER_43_1971 ();
 sg13g2_fill_2 FILLER_43_1975 ();
 sg13g2_fill_1 FILLER_43_1981 ();
 sg13g2_fill_1 FILLER_43_1988 ();
 sg13g2_fill_2 FILLER_43_2033 ();
 sg13g2_fill_1 FILLER_43_2035 ();
 sg13g2_fill_1 FILLER_43_2040 ();
 sg13g2_fill_1 FILLER_43_2047 ();
 sg13g2_fill_1 FILLER_43_2053 ();
 sg13g2_fill_1 FILLER_43_2059 ();
 sg13g2_fill_1 FILLER_43_2086 ();
 sg13g2_fill_1 FILLER_43_2091 ();
 sg13g2_fill_1 FILLER_43_2097 ();
 sg13g2_fill_1 FILLER_43_2107 ();
 sg13g2_decap_8 FILLER_43_2134 ();
 sg13g2_fill_1 FILLER_43_2141 ();
 sg13g2_fill_2 FILLER_43_2146 ();
 sg13g2_decap_8 FILLER_43_2174 ();
 sg13g2_decap_4 FILLER_43_2181 ();
 sg13g2_fill_2 FILLER_43_2185 ();
 sg13g2_fill_1 FILLER_43_2194 ();
 sg13g2_decap_8 FILLER_43_2221 ();
 sg13g2_decap_8 FILLER_43_2228 ();
 sg13g2_decap_8 FILLER_43_2235 ();
 sg13g2_decap_4 FILLER_43_2242 ();
 sg13g2_fill_2 FILLER_43_2307 ();
 sg13g2_decap_8 FILLER_43_2313 ();
 sg13g2_decap_4 FILLER_43_2320 ();
 sg13g2_fill_2 FILLER_43_2343 ();
 sg13g2_fill_1 FILLER_43_2349 ();
 sg13g2_fill_2 FILLER_43_2389 ();
 sg13g2_fill_2 FILLER_43_2446 ();
 sg13g2_fill_1 FILLER_43_2448 ();
 sg13g2_decap_8 FILLER_43_2453 ();
 sg13g2_fill_1 FILLER_43_2460 ();
 sg13g2_fill_1 FILLER_43_2467 ();
 sg13g2_fill_2 FILLER_43_2504 ();
 sg13g2_decap_8 FILLER_43_2510 ();
 sg13g2_decap_4 FILLER_43_2517 ();
 sg13g2_fill_1 FILLER_43_2524 ();
 sg13g2_decap_8 FILLER_43_2564 ();
 sg13g2_decap_8 FILLER_43_2571 ();
 sg13g2_decap_8 FILLER_43_2608 ();
 sg13g2_decap_8 FILLER_43_2615 ();
 sg13g2_fill_2 FILLER_43_2627 ();
 sg13g2_fill_1 FILLER_43_2629 ();
 sg13g2_fill_2 FILLER_43_2635 ();
 sg13g2_fill_2 FILLER_43_2668 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_fill_2 FILLER_44_50 ();
 sg13g2_fill_1 FILLER_44_52 ();
 sg13g2_fill_2 FILLER_44_82 ();
 sg13g2_fill_2 FILLER_44_89 ();
 sg13g2_fill_1 FILLER_44_101 ();
 sg13g2_fill_2 FILLER_44_107 ();
 sg13g2_fill_1 FILLER_44_109 ();
 sg13g2_decap_4 FILLER_44_120 ();
 sg13g2_fill_1 FILLER_44_124 ();
 sg13g2_fill_2 FILLER_44_149 ();
 sg13g2_decap_8 FILLER_44_156 ();
 sg13g2_decap_8 FILLER_44_163 ();
 sg13g2_decap_8 FILLER_44_170 ();
 sg13g2_decap_8 FILLER_44_177 ();
 sg13g2_fill_2 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_186 ();
 sg13g2_decap_4 FILLER_44_192 ();
 sg13g2_fill_2 FILLER_44_196 ();
 sg13g2_fill_1 FILLER_44_230 ();
 sg13g2_fill_1 FILLER_44_238 ();
 sg13g2_decap_8 FILLER_44_243 ();
 sg13g2_decap_4 FILLER_44_250 ();
 sg13g2_fill_2 FILLER_44_284 ();
 sg13g2_fill_1 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_300 ();
 sg13g2_fill_2 FILLER_44_307 ();
 sg13g2_fill_2 FILLER_44_318 ();
 sg13g2_decap_8 FILLER_44_335 ();
 sg13g2_fill_1 FILLER_44_342 ();
 sg13g2_decap_8 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_391 ();
 sg13g2_fill_2 FILLER_44_421 ();
 sg13g2_fill_1 FILLER_44_423 ();
 sg13g2_fill_2 FILLER_44_442 ();
 sg13g2_fill_1 FILLER_44_444 ();
 sg13g2_decap_8 FILLER_44_449 ();
 sg13g2_decap_8 FILLER_44_456 ();
 sg13g2_decap_8 FILLER_44_463 ();
 sg13g2_decap_8 FILLER_44_470 ();
 sg13g2_fill_2 FILLER_44_477 ();
 sg13g2_decap_8 FILLER_44_482 ();
 sg13g2_decap_8 FILLER_44_489 ();
 sg13g2_fill_2 FILLER_44_496 ();
 sg13g2_fill_2 FILLER_44_519 ();
 sg13g2_fill_1 FILLER_44_521 ();
 sg13g2_fill_2 FILLER_44_527 ();
 sg13g2_decap_8 FILLER_44_537 ();
 sg13g2_fill_1 FILLER_44_544 ();
 sg13g2_decap_8 FILLER_44_549 ();
 sg13g2_fill_2 FILLER_44_556 ();
 sg13g2_fill_1 FILLER_44_566 ();
 sg13g2_decap_4 FILLER_44_579 ();
 sg13g2_fill_2 FILLER_44_583 ();
 sg13g2_decap_4 FILLER_44_603 ();
 sg13g2_fill_1 FILLER_44_607 ();
 sg13g2_fill_1 FILLER_44_668 ();
 sg13g2_fill_1 FILLER_44_673 ();
 sg13g2_decap_8 FILLER_44_679 ();
 sg13g2_decap_4 FILLER_44_686 ();
 sg13g2_fill_1 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_717 ();
 sg13g2_decap_8 FILLER_44_724 ();
 sg13g2_decap_8 FILLER_44_731 ();
 sg13g2_decap_8 FILLER_44_738 ();
 sg13g2_decap_8 FILLER_44_745 ();
 sg13g2_decap_8 FILLER_44_752 ();
 sg13g2_decap_8 FILLER_44_785 ();
 sg13g2_fill_2 FILLER_44_892 ();
 sg13g2_fill_1 FILLER_44_894 ();
 sg13g2_fill_2 FILLER_44_898 ();
 sg13g2_fill_2 FILLER_44_915 ();
 sg13g2_fill_2 FILLER_44_927 ();
 sg13g2_fill_1 FILLER_44_929 ();
 sg13g2_fill_1 FILLER_44_935 ();
 sg13g2_decap_8 FILLER_44_966 ();
 sg13g2_decap_8 FILLER_44_973 ();
 sg13g2_decap_8 FILLER_44_980 ();
 sg13g2_fill_2 FILLER_44_987 ();
 sg13g2_decap_8 FILLER_44_993 ();
 sg13g2_fill_2 FILLER_44_1000 ();
 sg13g2_fill_1 FILLER_44_1002 ();
 sg13g2_fill_2 FILLER_44_1008 ();
 sg13g2_fill_1 FILLER_44_1010 ();
 sg13g2_decap_4 FILLER_44_1020 ();
 sg13g2_fill_2 FILLER_44_1035 ();
 sg13g2_fill_1 FILLER_44_1037 ();
 sg13g2_decap_4 FILLER_44_1047 ();
 sg13g2_fill_2 FILLER_44_1066 ();
 sg13g2_fill_1 FILLER_44_1132 ();
 sg13g2_fill_1 FILLER_44_1169 ();
 sg13g2_fill_2 FILLER_44_1176 ();
 sg13g2_decap_8 FILLER_44_1190 ();
 sg13g2_decap_4 FILLER_44_1205 ();
 sg13g2_fill_2 FILLER_44_1209 ();
 sg13g2_decap_8 FILLER_44_1230 ();
 sg13g2_decap_8 FILLER_44_1237 ();
 sg13g2_decap_8 FILLER_44_1244 ();
 sg13g2_decap_8 FILLER_44_1251 ();
 sg13g2_decap_8 FILLER_44_1258 ();
 sg13g2_decap_8 FILLER_44_1265 ();
 sg13g2_decap_4 FILLER_44_1275 ();
 sg13g2_fill_2 FILLER_44_1279 ();
 sg13g2_fill_1 FILLER_44_1287 ();
 sg13g2_decap_8 FILLER_44_1292 ();
 sg13g2_fill_1 FILLER_44_1299 ();
 sg13g2_decap_8 FILLER_44_1330 ();
 sg13g2_decap_4 FILLER_44_1337 ();
 sg13g2_fill_1 FILLER_44_1341 ();
 sg13g2_decap_8 FILLER_44_1346 ();
 sg13g2_decap_8 FILLER_44_1353 ();
 sg13g2_decap_8 FILLER_44_1390 ();
 sg13g2_fill_2 FILLER_44_1397 ();
 sg13g2_fill_1 FILLER_44_1399 ();
 sg13g2_decap_8 FILLER_44_1405 ();
 sg13g2_fill_2 FILLER_44_1412 ();
 sg13g2_fill_1 FILLER_44_1419 ();
 sg13g2_decap_8 FILLER_44_1448 ();
 sg13g2_fill_1 FILLER_44_1460 ();
 sg13g2_decap_8 FILLER_44_1487 ();
 sg13g2_decap_8 FILLER_44_1494 ();
 sg13g2_fill_2 FILLER_44_1501 ();
 sg13g2_fill_1 FILLER_44_1503 ();
 sg13g2_decap_4 FILLER_44_1521 ();
 sg13g2_decap_8 FILLER_44_1561 ();
 sg13g2_fill_1 FILLER_44_1568 ();
 sg13g2_fill_2 FILLER_44_1573 ();
 sg13g2_fill_2 FILLER_44_1590 ();
 sg13g2_fill_2 FILLER_44_1597 ();
 sg13g2_fill_1 FILLER_44_1628 ();
 sg13g2_fill_2 FILLER_44_1643 ();
 sg13g2_decap_8 FILLER_44_1695 ();
 sg13g2_decap_8 FILLER_44_1702 ();
 sg13g2_decap_4 FILLER_44_1709 ();
 sg13g2_fill_2 FILLER_44_1713 ();
 sg13g2_decap_8 FILLER_44_1720 ();
 sg13g2_decap_4 FILLER_44_1727 ();
 sg13g2_fill_1 FILLER_44_1731 ();
 sg13g2_fill_2 FILLER_44_1745 ();
 sg13g2_fill_1 FILLER_44_1747 ();
 sg13g2_fill_2 FILLER_44_1753 ();
 sg13g2_decap_8 FILLER_44_1759 ();
 sg13g2_fill_1 FILLER_44_1766 ();
 sg13g2_decap_4 FILLER_44_1847 ();
 sg13g2_fill_2 FILLER_44_1851 ();
 sg13g2_fill_2 FILLER_44_1894 ();
 sg13g2_fill_1 FILLER_44_1901 ();
 sg13g2_decap_8 FILLER_44_1909 ();
 sg13g2_decap_8 FILLER_44_1916 ();
 sg13g2_decap_4 FILLER_44_1923 ();
 sg13g2_fill_2 FILLER_44_1927 ();
 sg13g2_decap_8 FILLER_44_1934 ();
 sg13g2_decap_4 FILLER_44_1946 ();
 sg13g2_fill_1 FILLER_44_1950 ();
 sg13g2_fill_2 FILLER_44_1978 ();
 sg13g2_fill_2 FILLER_44_1983 ();
 sg13g2_decap_8 FILLER_44_2002 ();
 sg13g2_fill_2 FILLER_44_2009 ();
 sg13g2_decap_8 FILLER_44_2021 ();
 sg13g2_decap_8 FILLER_44_2028 ();
 sg13g2_decap_8 FILLER_44_2035 ();
 sg13g2_decap_4 FILLER_44_2042 ();
 sg13g2_fill_2 FILLER_44_2046 ();
 sg13g2_fill_2 FILLER_44_2052 ();
 sg13g2_fill_2 FILLER_44_2093 ();
 sg13g2_fill_2 FILLER_44_2146 ();
 sg13g2_fill_1 FILLER_44_2153 ();
 sg13g2_decap_8 FILLER_44_2180 ();
 sg13g2_decap_8 FILLER_44_2187 ();
 sg13g2_decap_4 FILLER_44_2217 ();
 sg13g2_decap_8 FILLER_44_2251 ();
 sg13g2_fill_2 FILLER_44_2258 ();
 sg13g2_fill_1 FILLER_44_2260 ();
 sg13g2_fill_2 FILLER_44_2273 ();
 sg13g2_fill_1 FILLER_44_2301 ();
 sg13g2_decap_8 FILLER_44_2354 ();
 sg13g2_decap_8 FILLER_44_2361 ();
 sg13g2_fill_2 FILLER_44_2377 ();
 sg13g2_fill_1 FILLER_44_2379 ();
 sg13g2_fill_2 FILLER_44_2416 ();
 sg13g2_fill_1 FILLER_44_2431 ();
 sg13g2_fill_2 FILLER_44_2458 ();
 sg13g2_fill_1 FILLER_44_2460 ();
 sg13g2_fill_2 FILLER_44_2464 ();
 sg13g2_fill_1 FILLER_44_2466 ();
 sg13g2_fill_2 FILLER_44_2471 ();
 sg13g2_fill_1 FILLER_44_2473 ();
 sg13g2_fill_1 FILLER_44_2508 ();
 sg13g2_decap_8 FILLER_44_2513 ();
 sg13g2_fill_1 FILLER_44_2520 ();
 sg13g2_fill_2 FILLER_44_2565 ();
 sg13g2_decap_4 FILLER_44_2654 ();
 sg13g2_fill_1 FILLER_44_2658 ();
 sg13g2_decap_8 FILLER_44_2663 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_fill_1 FILLER_45_61 ();
 sg13g2_fill_1 FILLER_45_85 ();
 sg13g2_fill_2 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_162 ();
 sg13g2_decap_8 FILLER_45_169 ();
 sg13g2_decap_4 FILLER_45_176 ();
 sg13g2_fill_2 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_233 ();
 sg13g2_decap_4 FILLER_45_262 ();
 sg13g2_fill_1 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_277 ();
 sg13g2_fill_1 FILLER_45_286 ();
 sg13g2_decap_4 FILLER_45_321 ();
 sg13g2_fill_1 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_fill_2 FILLER_45_349 ();
 sg13g2_fill_1 FILLER_45_351 ();
 sg13g2_fill_1 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_372 ();
 sg13g2_fill_1 FILLER_45_379 ();
 sg13g2_fill_2 FILLER_45_385 ();
 sg13g2_fill_1 FILLER_45_387 ();
 sg13g2_decap_8 FILLER_45_395 ();
 sg13g2_fill_2 FILLER_45_406 ();
 sg13g2_fill_1 FILLER_45_408 ();
 sg13g2_decap_4 FILLER_45_418 ();
 sg13g2_fill_2 FILLER_45_422 ();
 sg13g2_decap_8 FILLER_45_437 ();
 sg13g2_decap_8 FILLER_45_444 ();
 sg13g2_fill_2 FILLER_45_454 ();
 sg13g2_fill_1 FILLER_45_456 ();
 sg13g2_decap_8 FILLER_45_461 ();
 sg13g2_fill_2 FILLER_45_468 ();
 sg13g2_fill_1 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_551 ();
 sg13g2_decap_4 FILLER_45_558 ();
 sg13g2_fill_2 FILLER_45_566 ();
 sg13g2_fill_1 FILLER_45_578 ();
 sg13g2_fill_2 FILLER_45_584 ();
 sg13g2_fill_1 FILLER_45_586 ();
 sg13g2_fill_1 FILLER_45_591 ();
 sg13g2_fill_1 FILLER_45_597 ();
 sg13g2_fill_2 FILLER_45_602 ();
 sg13g2_fill_2 FILLER_45_611 ();
 sg13g2_fill_2 FILLER_45_618 ();
 sg13g2_fill_1 FILLER_45_620 ();
 sg13g2_fill_1 FILLER_45_634 ();
 sg13g2_decap_4 FILLER_45_644 ();
 sg13g2_fill_1 FILLER_45_648 ();
 sg13g2_decap_4 FILLER_45_658 ();
 sg13g2_fill_2 FILLER_45_667 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_fill_1 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_709 ();
 sg13g2_decap_8 FILLER_45_716 ();
 sg13g2_decap_8 FILLER_45_736 ();
 sg13g2_decap_8 FILLER_45_743 ();
 sg13g2_decap_4 FILLER_45_750 ();
 sg13g2_decap_8 FILLER_45_759 ();
 sg13g2_fill_2 FILLER_45_766 ();
 sg13g2_fill_1 FILLER_45_768 ();
 sg13g2_fill_2 FILLER_45_782 ();
 sg13g2_fill_1 FILLER_45_784 ();
 sg13g2_fill_1 FILLER_45_847 ();
 sg13g2_fill_1 FILLER_45_920 ();
 sg13g2_decap_4 FILLER_45_934 ();
 sg13g2_fill_1 FILLER_45_947 ();
 sg13g2_fill_2 FILLER_45_952 ();
 sg13g2_fill_2 FILLER_45_980 ();
 sg13g2_fill_2 FILLER_45_986 ();
 sg13g2_fill_1 FILLER_45_994 ();
 sg13g2_decap_4 FILLER_45_1025 ();
 sg13g2_decap_4 FILLER_45_1060 ();
 sg13g2_fill_2 FILLER_45_1133 ();
 sg13g2_fill_2 FILLER_45_1167 ();
 sg13g2_fill_2 FILLER_45_1214 ();
 sg13g2_decap_8 FILLER_45_1221 ();
 sg13g2_decap_8 FILLER_45_1228 ();
 sg13g2_fill_1 FILLER_45_1235 ();
 sg13g2_decap_8 FILLER_45_1241 ();
 sg13g2_decap_8 FILLER_45_1248 ();
 sg13g2_decap_8 FILLER_45_1255 ();
 sg13g2_fill_1 FILLER_45_1262 ();
 sg13g2_fill_1 FILLER_45_1271 ();
 sg13g2_decap_8 FILLER_45_1292 ();
 sg13g2_fill_1 FILLER_45_1299 ();
 sg13g2_decap_8 FILLER_45_1317 ();
 sg13g2_decap_4 FILLER_45_1324 ();
 sg13g2_fill_1 FILLER_45_1328 ();
 sg13g2_decap_4 FILLER_45_1371 ();
 sg13g2_fill_2 FILLER_45_1381 ();
 sg13g2_fill_1 FILLER_45_1383 ();
 sg13g2_fill_1 FILLER_45_1389 ();
 sg13g2_decap_4 FILLER_45_1395 ();
 sg13g2_fill_2 FILLER_45_1441 ();
 sg13g2_fill_1 FILLER_45_1443 ();
 sg13g2_decap_4 FILLER_45_1496 ();
 sg13g2_decap_4 FILLER_45_1513 ();
 sg13g2_fill_1 FILLER_45_1517 ();
 sg13g2_decap_8 FILLER_45_1522 ();
 sg13g2_decap_8 FILLER_45_1529 ();
 sg13g2_decap_8 FILLER_45_1536 ();
 sg13g2_decap_8 FILLER_45_1543 ();
 sg13g2_decap_8 FILLER_45_1550 ();
 sg13g2_decap_8 FILLER_45_1557 ();
 sg13g2_decap_8 FILLER_45_1564 ();
 sg13g2_fill_1 FILLER_45_1571 ();
 sg13g2_fill_2 FILLER_45_1581 ();
 sg13g2_decap_8 FILLER_45_1588 ();
 sg13g2_decap_8 FILLER_45_1595 ();
 sg13g2_decap_8 FILLER_45_1602 ();
 sg13g2_decap_4 FILLER_45_1609 ();
 sg13g2_fill_1 FILLER_45_1613 ();
 sg13g2_fill_2 FILLER_45_1630 ();
 sg13g2_fill_1 FILLER_45_1643 ();
 sg13g2_fill_2 FILLER_45_1652 ();
 sg13g2_fill_2 FILLER_45_1718 ();
 sg13g2_fill_2 FILLER_45_1732 ();
 sg13g2_fill_1 FILLER_45_1778 ();
 sg13g2_fill_1 FILLER_45_1794 ();
 sg13g2_fill_2 FILLER_45_1799 ();
 sg13g2_decap_4 FILLER_45_1816 ();
 sg13g2_fill_1 FILLER_45_1820 ();
 sg13g2_fill_1 FILLER_45_1829 ();
 sg13g2_fill_1 FILLER_45_1873 ();
 sg13g2_fill_2 FILLER_45_1901 ();
 sg13g2_decap_8 FILLER_45_1933 ();
 sg13g2_decap_4 FILLER_45_1940 ();
 sg13g2_fill_2 FILLER_45_1944 ();
 sg13g2_fill_2 FILLER_45_1950 ();
 sg13g2_fill_1 FILLER_45_1990 ();
 sg13g2_fill_2 FILLER_45_2006 ();
 sg13g2_fill_1 FILLER_45_2008 ();
 sg13g2_fill_2 FILLER_45_2016 ();
 sg13g2_decap_8 FILLER_45_2024 ();
 sg13g2_decap_8 FILLER_45_2031 ();
 sg13g2_decap_8 FILLER_45_2038 ();
 sg13g2_decap_8 FILLER_45_2045 ();
 sg13g2_decap_4 FILLER_45_2052 ();
 sg13g2_fill_1 FILLER_45_2056 ();
 sg13g2_fill_1 FILLER_45_2062 ();
 sg13g2_fill_1 FILLER_45_2068 ();
 sg13g2_fill_2 FILLER_45_2086 ();
 sg13g2_decap_8 FILLER_45_2104 ();
 sg13g2_decap_8 FILLER_45_2111 ();
 sg13g2_decap_8 FILLER_45_2118 ();
 sg13g2_fill_2 FILLER_45_2125 ();
 sg13g2_fill_1 FILLER_45_2127 ();
 sg13g2_decap_8 FILLER_45_2134 ();
 sg13g2_decap_8 FILLER_45_2141 ();
 sg13g2_decap_8 FILLER_45_2148 ();
 sg13g2_decap_8 FILLER_45_2155 ();
 sg13g2_decap_4 FILLER_45_2162 ();
 sg13g2_fill_2 FILLER_45_2166 ();
 sg13g2_decap_8 FILLER_45_2172 ();
 sg13g2_decap_8 FILLER_45_2179 ();
 sg13g2_fill_1 FILLER_45_2186 ();
 sg13g2_decap_4 FILLER_45_2210 ();
 sg13g2_decap_4 FILLER_45_2240 ();
 sg13g2_fill_1 FILLER_45_2244 ();
 sg13g2_decap_8 FILLER_45_2249 ();
 sg13g2_decap_8 FILLER_45_2256 ();
 sg13g2_decap_8 FILLER_45_2263 ();
 sg13g2_fill_1 FILLER_45_2270 ();
 sg13g2_fill_2 FILLER_45_2277 ();
 sg13g2_fill_1 FILLER_45_2283 ();
 sg13g2_fill_2 FILLER_45_2288 ();
 sg13g2_decap_4 FILLER_45_2294 ();
 sg13g2_decap_8 FILLER_45_2302 ();
 sg13g2_decap_8 FILLER_45_2309 ();
 sg13g2_decap_4 FILLER_45_2316 ();
 sg13g2_fill_2 FILLER_45_2330 ();
 sg13g2_fill_1 FILLER_45_2332 ();
 sg13g2_decap_8 FILLER_45_2337 ();
 sg13g2_decap_8 FILLER_45_2344 ();
 sg13g2_fill_1 FILLER_45_2364 ();
 sg13g2_fill_1 FILLER_45_2382 ();
 sg13g2_fill_1 FILLER_45_2414 ();
 sg13g2_fill_2 FILLER_45_2441 ();
 sg13g2_decap_8 FILLER_45_2461 ();
 sg13g2_fill_2 FILLER_45_2479 ();
 sg13g2_fill_2 FILLER_45_2485 ();
 sg13g2_fill_2 FILLER_45_2491 ();
 sg13g2_fill_1 FILLER_45_2493 ();
 sg13g2_decap_8 FILLER_45_2528 ();
 sg13g2_fill_1 FILLER_45_2535 ();
 sg13g2_decap_4 FILLER_45_2540 ();
 sg13g2_fill_1 FILLER_45_2544 ();
 sg13g2_fill_2 FILLER_45_2549 ();
 sg13g2_fill_1 FILLER_45_2555 ();
 sg13g2_fill_2 FILLER_45_2600 ();
 sg13g2_fill_1 FILLER_45_2602 ();
 sg13g2_decap_8 FILLER_45_2607 ();
 sg13g2_decap_8 FILLER_45_2614 ();
 sg13g2_fill_1 FILLER_45_2621 ();
 sg13g2_decap_4 FILLER_45_2666 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_4 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_110 ();
 sg13g2_fill_1 FILLER_46_117 ();
 sg13g2_decap_8 FILLER_46_122 ();
 sg13g2_fill_1 FILLER_46_129 ();
 sg13g2_decap_8 FILLER_46_152 ();
 sg13g2_decap_4 FILLER_46_159 ();
 sg13g2_fill_2 FILLER_46_163 ();
 sg13g2_decap_4 FILLER_46_245 ();
 sg13g2_decap_8 FILLER_46_254 ();
 sg13g2_fill_1 FILLER_46_267 ();
 sg13g2_fill_2 FILLER_46_277 ();
 sg13g2_fill_1 FILLER_46_294 ();
 sg13g2_decap_4 FILLER_46_330 ();
 sg13g2_fill_1 FILLER_46_360 ();
 sg13g2_fill_1 FILLER_46_371 ();
 sg13g2_fill_2 FILLER_46_376 ();
 sg13g2_fill_2 FILLER_46_404 ();
 sg13g2_decap_4 FILLER_46_410 ();
 sg13g2_fill_1 FILLER_46_414 ();
 sg13g2_decap_8 FILLER_46_419 ();
 sg13g2_fill_2 FILLER_46_426 ();
 sg13g2_fill_1 FILLER_46_433 ();
 sg13g2_fill_1 FILLER_46_443 ();
 sg13g2_fill_2 FILLER_46_456 ();
 sg13g2_fill_1 FILLER_46_458 ();
 sg13g2_decap_4 FILLER_46_504 ();
 sg13g2_fill_2 FILLER_46_508 ();
 sg13g2_fill_2 FILLER_46_527 ();
 sg13g2_decap_8 FILLER_46_534 ();
 sg13g2_decap_4 FILLER_46_541 ();
 sg13g2_fill_1 FILLER_46_545 ();
 sg13g2_decap_4 FILLER_46_549 ();
 sg13g2_fill_2 FILLER_46_553 ();
 sg13g2_decap_8 FILLER_46_562 ();
 sg13g2_decap_8 FILLER_46_569 ();
 sg13g2_fill_2 FILLER_46_576 ();
 sg13g2_fill_1 FILLER_46_578 ();
 sg13g2_decap_4 FILLER_46_584 ();
 sg13g2_fill_1 FILLER_46_588 ();
 sg13g2_decap_4 FILLER_46_594 ();
 sg13g2_fill_2 FILLER_46_598 ();
 sg13g2_decap_4 FILLER_46_606 ();
 sg13g2_fill_1 FILLER_46_620 ();
 sg13g2_decap_4 FILLER_46_627 ();
 sg13g2_decap_8 FILLER_46_635 ();
 sg13g2_fill_1 FILLER_46_642 ();
 sg13g2_fill_1 FILLER_46_651 ();
 sg13g2_fill_1 FILLER_46_670 ();
 sg13g2_decap_4 FILLER_46_682 ();
 sg13g2_fill_2 FILLER_46_686 ();
 sg13g2_decap_4 FILLER_46_716 ();
 sg13g2_decap_8 FILLER_46_724 ();
 sg13g2_decap_8 FILLER_46_731 ();
 sg13g2_decap_8 FILLER_46_738 ();
 sg13g2_decap_8 FILLER_46_745 ();
 sg13g2_decap_8 FILLER_46_752 ();
 sg13g2_fill_2 FILLER_46_759 ();
 sg13g2_decap_8 FILLER_46_765 ();
 sg13g2_fill_1 FILLER_46_772 ();
 sg13g2_decap_8 FILLER_46_778 ();
 sg13g2_decap_8 FILLER_46_785 ();
 sg13g2_decap_8 FILLER_46_797 ();
 sg13g2_fill_1 FILLER_46_804 ();
 sg13g2_decap_4 FILLER_46_815 ();
 sg13g2_fill_1 FILLER_46_819 ();
 sg13g2_fill_2 FILLER_46_824 ();
 sg13g2_fill_1 FILLER_46_826 ();
 sg13g2_fill_2 FILLER_46_837 ();
 sg13g2_fill_2 FILLER_46_843 ();
 sg13g2_fill_1 FILLER_46_888 ();
 sg13g2_decap_4 FILLER_46_898 ();
 sg13g2_fill_1 FILLER_46_902 ();
 sg13g2_decap_8 FILLER_46_942 ();
 sg13g2_fill_1 FILLER_46_949 ();
 sg13g2_decap_8 FILLER_46_959 ();
 sg13g2_fill_2 FILLER_46_1032 ();
 sg13g2_fill_2 FILLER_46_1038 ();
 sg13g2_decap_8 FILLER_46_1071 ();
 sg13g2_decap_4 FILLER_46_1078 ();
 sg13g2_decap_4 FILLER_46_1090 ();
 sg13g2_fill_2 FILLER_46_1112 ();
 sg13g2_fill_1 FILLER_46_1119 ();
 sg13g2_fill_1 FILLER_46_1124 ();
 sg13g2_fill_1 FILLER_46_1133 ();
 sg13g2_fill_1 FILLER_46_1144 ();
 sg13g2_decap_8 FILLER_46_1176 ();
 sg13g2_fill_2 FILLER_46_1183 ();
 sg13g2_decap_4 FILLER_46_1217 ();
 sg13g2_fill_2 FILLER_46_1230 ();
 sg13g2_fill_2 FILLER_46_1269 ();
 sg13g2_decap_4 FILLER_46_1275 ();
 sg13g2_decap_8 FILLER_46_1292 ();
 sg13g2_fill_2 FILLER_46_1299 ();
 sg13g2_fill_1 FILLER_46_1301 ();
 sg13g2_decap_8 FILLER_46_1307 ();
 sg13g2_decap_8 FILLER_46_1314 ();
 sg13g2_fill_1 FILLER_46_1321 ();
 sg13g2_fill_1 FILLER_46_1327 ();
 sg13g2_decap_8 FILLER_46_1332 ();
 sg13g2_fill_2 FILLER_46_1339 ();
 sg13g2_decap_4 FILLER_46_1346 ();
 sg13g2_fill_1 FILLER_46_1350 ();
 sg13g2_fill_2 FILLER_46_1377 ();
 sg13g2_fill_2 FILLER_46_1405 ();
 sg13g2_fill_1 FILLER_46_1407 ();
 sg13g2_fill_2 FILLER_46_1437 ();
 sg13g2_fill_2 FILLER_46_1453 ();
 sg13g2_fill_1 FILLER_46_1459 ();
 sg13g2_fill_2 FILLER_46_1466 ();
 sg13g2_decap_8 FILLER_46_1477 ();
 sg13g2_decap_8 FILLER_46_1484 ();
 sg13g2_fill_2 FILLER_46_1491 ();
 sg13g2_fill_1 FILLER_46_1493 ();
 sg13g2_fill_2 FILLER_46_1520 ();
 sg13g2_fill_1 FILLER_46_1522 ();
 sg13g2_decap_4 FILLER_46_1527 ();
 sg13g2_fill_2 FILLER_46_1531 ();
 sg13g2_fill_2 FILLER_46_1537 ();
 sg13g2_fill_2 FILLER_46_1582 ();
 sg13g2_decap_8 FILLER_46_1610 ();
 sg13g2_decap_8 FILLER_46_1617 ();
 sg13g2_fill_1 FILLER_46_1660 ();
 sg13g2_fill_2 FILLER_46_1666 ();
 sg13g2_fill_2 FILLER_46_1689 ();
 sg13g2_decap_8 FILLER_46_1695 ();
 sg13g2_decap_4 FILLER_46_1702 ();
 sg13g2_fill_2 FILLER_46_1706 ();
 sg13g2_fill_1 FILLER_46_1734 ();
 sg13g2_fill_1 FILLER_46_1807 ();
 sg13g2_decap_4 FILLER_46_1834 ();
 sg13g2_fill_1 FILLER_46_1838 ();
 sg13g2_fill_2 FILLER_46_1862 ();
 sg13g2_fill_1 FILLER_46_1864 ();
 sg13g2_fill_1 FILLER_46_1877 ();
 sg13g2_fill_2 FILLER_46_1883 ();
 sg13g2_fill_1 FILLER_46_1893 ();
 sg13g2_fill_1 FILLER_46_1900 ();
 sg13g2_decap_8 FILLER_46_1906 ();
 sg13g2_fill_1 FILLER_46_1913 ();
 sg13g2_decap_8 FILLER_46_1918 ();
 sg13g2_fill_2 FILLER_46_1925 ();
 sg13g2_fill_1 FILLER_46_1927 ();
 sg13g2_fill_1 FILLER_46_1954 ();
 sg13g2_fill_2 FILLER_46_1961 ();
 sg13g2_fill_1 FILLER_46_1974 ();
 sg13g2_fill_2 FILLER_46_2012 ();
 sg13g2_decap_4 FILLER_46_2028 ();
 sg13g2_fill_1 FILLER_46_2032 ();
 sg13g2_decap_8 FILLER_46_2090 ();
 sg13g2_fill_1 FILLER_46_2097 ();
 sg13g2_decap_8 FILLER_46_2106 ();
 sg13g2_decap_4 FILLER_46_2113 ();
 sg13g2_fill_2 FILLER_46_2117 ();
 sg13g2_decap_4 FILLER_46_2153 ();
 sg13g2_fill_2 FILLER_46_2187 ();
 sg13g2_fill_1 FILLER_46_2189 ();
 sg13g2_decap_8 FILLER_46_2194 ();
 sg13g2_fill_1 FILLER_46_2201 ();
 sg13g2_decap_8 FILLER_46_2208 ();
 sg13g2_decap_8 FILLER_46_2215 ();
 sg13g2_fill_1 FILLER_46_2222 ();
 sg13g2_decap_8 FILLER_46_2229 ();
 sg13g2_fill_2 FILLER_46_2236 ();
 sg13g2_fill_1 FILLER_46_2238 ();
 sg13g2_fill_1 FILLER_46_2243 ();
 sg13g2_fill_1 FILLER_46_2249 ();
 sg13g2_decap_8 FILLER_46_2266 ();
 sg13g2_decap_8 FILLER_46_2273 ();
 sg13g2_decap_8 FILLER_46_2284 ();
 sg13g2_decap_4 FILLER_46_2291 ();
 sg13g2_decap_4 FILLER_46_2298 ();
 sg13g2_fill_1 FILLER_46_2306 ();
 sg13g2_decap_4 FILLER_46_2333 ();
 sg13g2_fill_2 FILLER_46_2337 ();
 sg13g2_decap_4 FILLER_46_2345 ();
 sg13g2_fill_1 FILLER_46_2349 ();
 sg13g2_decap_8 FILLER_46_2354 ();
 sg13g2_fill_2 FILLER_46_2395 ();
 sg13g2_fill_1 FILLER_46_2455 ();
 sg13g2_decap_8 FILLER_46_2462 ();
 sg13g2_decap_4 FILLER_46_2469 ();
 sg13g2_fill_1 FILLER_46_2473 ();
 sg13g2_fill_2 FILLER_46_2483 ();
 sg13g2_decap_8 FILLER_46_2490 ();
 sg13g2_decap_8 FILLER_46_2497 ();
 sg13g2_decap_8 FILLER_46_2504 ();
 sg13g2_decap_8 FILLER_46_2511 ();
 sg13g2_decap_8 FILLER_46_2518 ();
 sg13g2_decap_8 FILLER_46_2525 ();
 sg13g2_decap_8 FILLER_46_2532 ();
 sg13g2_fill_1 FILLER_46_2539 ();
 sg13g2_decap_8 FILLER_46_2550 ();
 sg13g2_decap_8 FILLER_46_2557 ();
 sg13g2_decap_4 FILLER_46_2564 ();
 sg13g2_fill_2 FILLER_46_2568 ();
 sg13g2_fill_1 FILLER_46_2574 ();
 sg13g2_fill_1 FILLER_46_2583 ();
 sg13g2_decap_8 FILLER_46_2597 ();
 sg13g2_decap_8 FILLER_46_2604 ();
 sg13g2_decap_8 FILLER_46_2611 ();
 sg13g2_decap_8 FILLER_46_2618 ();
 sg13g2_fill_2 FILLER_46_2625 ();
 sg13g2_fill_1 FILLER_46_2627 ();
 sg13g2_decap_8 FILLER_46_2651 ();
 sg13g2_decap_8 FILLER_46_2658 ();
 sg13g2_decap_4 FILLER_46_2665 ();
 sg13g2_fill_1 FILLER_46_2669 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_fill_2 FILLER_47_38 ();
 sg13g2_fill_1 FILLER_47_40 ();
 sg13g2_decap_8 FILLER_47_51 ();
 sg13g2_fill_1 FILLER_47_63 ();
 sg13g2_decap_4 FILLER_47_76 ();
 sg13g2_fill_1 FILLER_47_80 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_4 FILLER_47_98 ();
 sg13g2_fill_1 FILLER_47_102 ();
 sg13g2_decap_8 FILLER_47_110 ();
 sg13g2_decap_8 FILLER_47_117 ();
 sg13g2_fill_2 FILLER_47_139 ();
 sg13g2_fill_1 FILLER_47_141 ();
 sg13g2_decap_4 FILLER_47_147 ();
 sg13g2_fill_1 FILLER_47_151 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_decap_8 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_178 ();
 sg13g2_fill_1 FILLER_47_190 ();
 sg13g2_fill_1 FILLER_47_241 ();
 sg13g2_fill_1 FILLER_47_248 ();
 sg13g2_fill_2 FILLER_47_255 ();
 sg13g2_fill_2 FILLER_47_260 ();
 sg13g2_fill_1 FILLER_47_262 ();
 sg13g2_fill_2 FILLER_47_302 ();
 sg13g2_fill_1 FILLER_47_304 ();
 sg13g2_decap_4 FILLER_47_334 ();
 sg13g2_fill_1 FILLER_47_338 ();
 sg13g2_decap_8 FILLER_47_342 ();
 sg13g2_decap_8 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_fill_1 FILLER_47_370 ();
 sg13g2_fill_1 FILLER_47_380 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_fill_2 FILLER_47_440 ();
 sg13g2_fill_2 FILLER_47_481 ();
 sg13g2_fill_1 FILLER_47_483 ();
 sg13g2_fill_2 FILLER_47_487 ();
 sg13g2_decap_4 FILLER_47_515 ();
 sg13g2_fill_2 FILLER_47_528 ();
 sg13g2_decap_8 FILLER_47_540 ();
 sg13g2_decap_8 FILLER_47_547 ();
 sg13g2_decap_8 FILLER_47_554 ();
 sg13g2_fill_1 FILLER_47_561 ();
 sg13g2_fill_2 FILLER_47_577 ();
 sg13g2_fill_1 FILLER_47_579 ();
 sg13g2_decap_8 FILLER_47_589 ();
 sg13g2_decap_4 FILLER_47_607 ();
 sg13g2_fill_1 FILLER_47_611 ();
 sg13g2_fill_2 FILLER_47_626 ();
 sg13g2_fill_2 FILLER_47_657 ();
 sg13g2_fill_2 FILLER_47_666 ();
 sg13g2_fill_1 FILLER_47_697 ();
 sg13g2_decap_4 FILLER_47_729 ();
 sg13g2_fill_2 FILLER_47_733 ();
 sg13g2_decap_4 FILLER_47_753 ();
 sg13g2_fill_2 FILLER_47_757 ();
 sg13g2_fill_2 FILLER_47_790 ();
 sg13g2_fill_1 FILLER_47_792 ();
 sg13g2_fill_1 FILLER_47_802 ();
 sg13g2_decap_8 FILLER_47_807 ();
 sg13g2_fill_1 FILLER_47_814 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_4 FILLER_47_838 ();
 sg13g2_fill_2 FILLER_47_842 ();
 sg13g2_decap_4 FILLER_47_850 ();
 sg13g2_fill_2 FILLER_47_863 ();
 sg13g2_fill_1 FILLER_47_869 ();
 sg13g2_fill_2 FILLER_47_886 ();
 sg13g2_decap_4 FILLER_47_946 ();
 sg13g2_fill_1 FILLER_47_950 ();
 sg13g2_fill_2 FILLER_47_956 ();
 sg13g2_fill_1 FILLER_47_958 ();
 sg13g2_decap_8 FILLER_47_964 ();
 sg13g2_fill_2 FILLER_47_971 ();
 sg13g2_decap_4 FILLER_47_991 ();
 sg13g2_fill_2 FILLER_47_995 ();
 sg13g2_decap_8 FILLER_47_1002 ();
 sg13g2_decap_4 FILLER_47_1013 ();
 sg13g2_fill_1 FILLER_47_1017 ();
 sg13g2_fill_2 FILLER_47_1023 ();
 sg13g2_fill_1 FILLER_47_1025 ();
 sg13g2_decap_4 FILLER_47_1035 ();
 sg13g2_decap_8 FILLER_47_1043 ();
 sg13g2_decap_4 FILLER_47_1050 ();
 sg13g2_fill_2 FILLER_47_1054 ();
 sg13g2_decap_8 FILLER_47_1069 ();
 sg13g2_decap_8 FILLER_47_1076 ();
 sg13g2_fill_1 FILLER_47_1083 ();
 sg13g2_decap_8 FILLER_47_1089 ();
 sg13g2_decap_8 FILLER_47_1096 ();
 sg13g2_decap_8 FILLER_47_1103 ();
 sg13g2_fill_1 FILLER_47_1110 ();
 sg13g2_fill_1 FILLER_47_1169 ();
 sg13g2_decap_4 FILLER_47_1180 ();
 sg13g2_decap_4 FILLER_47_1190 ();
 sg13g2_fill_2 FILLER_47_1194 ();
 sg13g2_decap_4 FILLER_47_1211 ();
 sg13g2_fill_2 FILLER_47_1215 ();
 sg13g2_decap_8 FILLER_47_1243 ();
 sg13g2_fill_2 FILLER_47_1254 ();
 sg13g2_fill_1 FILLER_47_1256 ();
 sg13g2_fill_2 FILLER_47_1286 ();
 sg13g2_decap_4 FILLER_47_1318 ();
 sg13g2_fill_2 FILLER_47_1322 ();
 sg13g2_fill_2 FILLER_47_1355 ();
 sg13g2_decap_4 FILLER_47_1361 ();
 sg13g2_decap_8 FILLER_47_1369 ();
 sg13g2_fill_1 FILLER_47_1376 ();
 sg13g2_decap_4 FILLER_47_1386 ();
 sg13g2_fill_2 FILLER_47_1390 ();
 sg13g2_decap_8 FILLER_47_1397 ();
 sg13g2_fill_2 FILLER_47_1413 ();
 sg13g2_fill_2 FILLER_47_1420 ();
 sg13g2_fill_1 FILLER_47_1422 ();
 sg13g2_fill_1 FILLER_47_1427 ();
 sg13g2_decap_8 FILLER_47_1448 ();
 sg13g2_decap_8 FILLER_47_1455 ();
 sg13g2_decap_8 FILLER_47_1462 ();
 sg13g2_decap_8 FILLER_47_1469 ();
 sg13g2_decap_8 FILLER_47_1476 ();
 sg13g2_decap_8 FILLER_47_1483 ();
 sg13g2_decap_8 FILLER_47_1490 ();
 sg13g2_decap_8 FILLER_47_1497 ();
 sg13g2_fill_2 FILLER_47_1504 ();
 sg13g2_decap_4 FILLER_47_1519 ();
 sg13g2_fill_2 FILLER_47_1523 ();
 sg13g2_fill_2 FILLER_47_1533 ();
 sg13g2_fill_2 FILLER_47_1569 ();
 sg13g2_decap_8 FILLER_47_1576 ();
 sg13g2_decap_8 FILLER_47_1599 ();
 sg13g2_decap_8 FILLER_47_1606 ();
 sg13g2_decap_8 FILLER_47_1613 ();
 sg13g2_decap_8 FILLER_47_1620 ();
 sg13g2_decap_8 FILLER_47_1640 ();
 sg13g2_decap_8 FILLER_47_1647 ();
 sg13g2_decap_4 FILLER_47_1660 ();
 sg13g2_decap_4 FILLER_47_1716 ();
 sg13g2_fill_2 FILLER_47_1720 ();
 sg13g2_fill_2 FILLER_47_1726 ();
 sg13g2_decap_8 FILLER_47_1796 ();
 sg13g2_decap_8 FILLER_47_1803 ();
 sg13g2_decap_8 FILLER_47_1810 ();
 sg13g2_decap_8 FILLER_47_1817 ();
 sg13g2_decap_8 FILLER_47_1824 ();
 sg13g2_fill_1 FILLER_47_1831 ();
 sg13g2_decap_4 FILLER_47_1872 ();
 sg13g2_fill_1 FILLER_47_1897 ();
 sg13g2_decap_8 FILLER_47_1907 ();
 sg13g2_decap_4 FILLER_47_1914 ();
 sg13g2_fill_2 FILLER_47_1918 ();
 sg13g2_fill_1 FILLER_47_1948 ();
 sg13g2_fill_2 FILLER_47_1969 ();
 sg13g2_fill_2 FILLER_47_1981 ();
 sg13g2_fill_1 FILLER_47_1991 ();
 sg13g2_fill_1 FILLER_47_2030 ();
 sg13g2_fill_2 FILLER_47_2040 ();
 sg13g2_fill_1 FILLER_47_2042 ();
 sg13g2_decap_8 FILLER_47_2047 ();
 sg13g2_decap_4 FILLER_47_2054 ();
 sg13g2_fill_2 FILLER_47_2077 ();
 sg13g2_fill_2 FILLER_47_2093 ();
 sg13g2_fill_1 FILLER_47_2100 ();
 sg13g2_decap_8 FILLER_47_2173 ();
 sg13g2_decap_8 FILLER_47_2180 ();
 sg13g2_decap_8 FILLER_47_2187 ();
 sg13g2_fill_2 FILLER_47_2194 ();
 sg13g2_decap_8 FILLER_47_2209 ();
 sg13g2_decap_8 FILLER_47_2216 ();
 sg13g2_fill_2 FILLER_47_2229 ();
 sg13g2_fill_1 FILLER_47_2231 ();
 sg13g2_decap_8 FILLER_47_2240 ();
 sg13g2_decap_8 FILLER_47_2247 ();
 sg13g2_decap_8 FILLER_47_2254 ();
 sg13g2_fill_2 FILLER_47_2261 ();
 sg13g2_fill_1 FILLER_47_2294 ();
 sg13g2_fill_1 FILLER_47_2301 ();
 sg13g2_fill_2 FILLER_47_2328 ();
 sg13g2_decap_8 FILLER_47_2334 ();
 sg13g2_fill_2 FILLER_47_2341 ();
 sg13g2_decap_8 FILLER_47_2347 ();
 sg13g2_fill_1 FILLER_47_2410 ();
 sg13g2_fill_2 FILLER_47_2415 ();
 sg13g2_fill_2 FILLER_47_2473 ();
 sg13g2_fill_2 FILLER_47_2501 ();
 sg13g2_fill_1 FILLER_47_2503 ();
 sg13g2_fill_1 FILLER_47_2540 ();
 sg13g2_fill_2 FILLER_47_2553 ();
 sg13g2_fill_1 FILLER_47_2555 ();
 sg13g2_decap_8 FILLER_47_2563 ();
 sg13g2_decap_8 FILLER_47_2570 ();
 sg13g2_decap_8 FILLER_47_2577 ();
 sg13g2_fill_2 FILLER_47_2584 ();
 sg13g2_fill_1 FILLER_47_2586 ();
 sg13g2_decap_4 FILLER_47_2621 ();
 sg13g2_fill_2 FILLER_47_2667 ();
 sg13g2_fill_1 FILLER_47_2669 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_fill_1 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_34 ();
 sg13g2_decap_4 FILLER_48_55 ();
 sg13g2_fill_1 FILLER_48_59 ();
 sg13g2_decap_8 FILLER_48_72 ();
 sg13g2_fill_1 FILLER_48_79 ();
 sg13g2_decap_4 FILLER_48_94 ();
 sg13g2_fill_1 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_109 ();
 sg13g2_decap_8 FILLER_48_116 ();
 sg13g2_decap_8 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_130 ();
 sg13g2_fill_1 FILLER_48_137 ();
 sg13g2_fill_2 FILLER_48_146 ();
 sg13g2_decap_4 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_203 ();
 sg13g2_decap_4 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_291 ();
 sg13g2_fill_2 FILLER_48_295 ();
 sg13g2_fill_1 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_fill_1 FILLER_48_371 ();
 sg13g2_fill_2 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_48_383 ();
 sg13g2_fill_1 FILLER_48_428 ();
 sg13g2_decap_4 FILLER_48_433 ();
 sg13g2_decap_8 FILLER_48_446 ();
 sg13g2_fill_2 FILLER_48_467 ();
 sg13g2_fill_1 FILLER_48_520 ();
 sg13g2_decap_4 FILLER_48_550 ();
 sg13g2_fill_1 FILLER_48_554 ();
 sg13g2_decap_4 FILLER_48_559 ();
 sg13g2_decap_4 FILLER_48_585 ();
 sg13g2_fill_1 FILLER_48_598 ();
 sg13g2_fill_1 FILLER_48_609 ();
 sg13g2_fill_1 FILLER_48_614 ();
 sg13g2_decap_4 FILLER_48_626 ();
 sg13g2_fill_2 FILLER_48_630 ();
 sg13g2_fill_2 FILLER_48_640 ();
 sg13g2_fill_1 FILLER_48_642 ();
 sg13g2_fill_1 FILLER_48_652 ();
 sg13g2_fill_2 FILLER_48_662 ();
 sg13g2_fill_1 FILLER_48_664 ();
 sg13g2_fill_2 FILLER_48_680 ();
 sg13g2_fill_2 FILLER_48_687 ();
 sg13g2_fill_2 FILLER_48_702 ();
 sg13g2_decap_8 FILLER_48_708 ();
 sg13g2_decap_8 FILLER_48_715 ();
 sg13g2_decap_8 FILLER_48_722 ();
 sg13g2_decap_8 FILLER_48_729 ();
 sg13g2_decap_8 FILLER_48_736 ();
 sg13g2_fill_1 FILLER_48_743 ();
 sg13g2_fill_2 FILLER_48_775 ();
 sg13g2_decap_8 FILLER_48_821 ();
 sg13g2_fill_2 FILLER_48_828 ();
 sg13g2_fill_1 FILLER_48_830 ();
 sg13g2_fill_1 FILLER_48_871 ();
 sg13g2_fill_2 FILLER_48_906 ();
 sg13g2_decap_8 FILLER_48_946 ();
 sg13g2_decap_8 FILLER_48_953 ();
 sg13g2_decap_8 FILLER_48_960 ();
 sg13g2_decap_8 FILLER_48_967 ();
 sg13g2_fill_2 FILLER_48_1009 ();
 sg13g2_fill_2 FILLER_48_1014 ();
 sg13g2_fill_1 FILLER_48_1042 ();
 sg13g2_decap_8 FILLER_48_1095 ();
 sg13g2_fill_2 FILLER_48_1102 ();
 sg13g2_fill_1 FILLER_48_1104 ();
 sg13g2_decap_8 FILLER_48_1113 ();
 sg13g2_fill_1 FILLER_48_1120 ();
 sg13g2_fill_1 FILLER_48_1187 ();
 sg13g2_decap_4 FILLER_48_1201 ();
 sg13g2_decap_8 FILLER_48_1209 ();
 sg13g2_decap_4 FILLER_48_1216 ();
 sg13g2_decap_8 FILLER_48_1224 ();
 sg13g2_decap_8 FILLER_48_1231 ();
 sg13g2_fill_2 FILLER_48_1238 ();
 sg13g2_fill_2 FILLER_48_1250 ();
 sg13g2_fill_1 FILLER_48_1252 ();
 sg13g2_fill_1 FILLER_48_1263 ();
 sg13g2_fill_1 FILLER_48_1277 ();
 sg13g2_fill_1 FILLER_48_1283 ();
 sg13g2_decap_8 FILLER_48_1316 ();
 sg13g2_fill_1 FILLER_48_1323 ();
 sg13g2_decap_4 FILLER_48_1329 ();
 sg13g2_fill_2 FILLER_48_1333 ();
 sg13g2_decap_8 FILLER_48_1339 ();
 sg13g2_decap_8 FILLER_48_1346 ();
 sg13g2_decap_8 FILLER_48_1353 ();
 sg13g2_decap_8 FILLER_48_1360 ();
 sg13g2_decap_8 FILLER_48_1380 ();
 sg13g2_fill_2 FILLER_48_1387 ();
 sg13g2_decap_8 FILLER_48_1416 ();
 sg13g2_fill_2 FILLER_48_1423 ();
 sg13g2_fill_1 FILLER_48_1425 ();
 sg13g2_decap_8 FILLER_48_1486 ();
 sg13g2_decap_4 FILLER_48_1493 ();
 sg13g2_fill_1 FILLER_48_1497 ();
 sg13g2_decap_8 FILLER_48_1548 ();
 sg13g2_decap_8 FILLER_48_1555 ();
 sg13g2_decap_8 FILLER_48_1562 ();
 sg13g2_fill_2 FILLER_48_1569 ();
 sg13g2_fill_1 FILLER_48_1571 ();
 sg13g2_decap_8 FILLER_48_1581 ();
 sg13g2_fill_2 FILLER_48_1592 ();
 sg13g2_fill_1 FILLER_48_1594 ();
 sg13g2_decap_4 FILLER_48_1652 ();
 sg13g2_fill_2 FILLER_48_1667 ();
 sg13g2_decap_8 FILLER_48_1673 ();
 sg13g2_decap_8 FILLER_48_1680 ();
 sg13g2_decap_8 FILLER_48_1687 ();
 sg13g2_decap_8 FILLER_48_1694 ();
 sg13g2_decap_4 FILLER_48_1701 ();
 sg13g2_fill_1 FILLER_48_1705 ();
 sg13g2_decap_4 FILLER_48_1715 ();
 sg13g2_fill_1 FILLER_48_1719 ();
 sg13g2_decap_8 FILLER_48_1732 ();
 sg13g2_fill_2 FILLER_48_1739 ();
 sg13g2_fill_2 FILLER_48_1767 ();
 sg13g2_fill_1 FILLER_48_1769 ();
 sg13g2_decap_8 FILLER_48_1790 ();
 sg13g2_decap_8 FILLER_48_1797 ();
 sg13g2_decap_8 FILLER_48_1808 ();
 sg13g2_decap_4 FILLER_48_1815 ();
 sg13g2_fill_1 FILLER_48_1819 ();
 sg13g2_decap_8 FILLER_48_1830 ();
 sg13g2_decap_8 FILLER_48_1837 ();
 sg13g2_decap_8 FILLER_48_1847 ();
 sg13g2_decap_8 FILLER_48_1857 ();
 sg13g2_fill_1 FILLER_48_1895 ();
 sg13g2_fill_1 FILLER_48_1931 ();
 sg13g2_fill_2 FILLER_48_1935 ();
 sg13g2_fill_1 FILLER_48_1937 ();
 sg13g2_decap_4 FILLER_48_1975 ();
 sg13g2_fill_1 FILLER_48_1979 ();
 sg13g2_decap_8 FILLER_48_2019 ();
 sg13g2_decap_4 FILLER_48_2026 ();
 sg13g2_fill_2 FILLER_48_2030 ();
 sg13g2_fill_2 FILLER_48_2068 ();
 sg13g2_decap_8 FILLER_48_2082 ();
 sg13g2_decap_8 FILLER_48_2089 ();
 sg13g2_fill_1 FILLER_48_2096 ();
 sg13g2_fill_1 FILLER_48_2123 ();
 sg13g2_fill_1 FILLER_48_2129 ();
 sg13g2_fill_1 FILLER_48_2174 ();
 sg13g2_decap_8 FILLER_48_2180 ();
 sg13g2_fill_1 FILLER_48_2187 ();
 sg13g2_decap_4 FILLER_48_2197 ();
 sg13g2_fill_1 FILLER_48_2201 ();
 sg13g2_fill_2 FILLER_48_2258 ();
 sg13g2_fill_1 FILLER_48_2260 ();
 sg13g2_fill_2 FILLER_48_2265 ();
 sg13g2_fill_1 FILLER_48_2267 ();
 sg13g2_decap_4 FILLER_48_2294 ();
 sg13g2_fill_2 FILLER_48_2302 ();
 sg13g2_fill_1 FILLER_48_2304 ();
 sg13g2_decap_4 FILLER_48_2362 ();
 sg13g2_fill_2 FILLER_48_2366 ();
 sg13g2_fill_2 FILLER_48_2373 ();
 sg13g2_fill_1 FILLER_48_2375 ();
 sg13g2_decap_8 FILLER_48_2406 ();
 sg13g2_decap_8 FILLER_48_2413 ();
 sg13g2_fill_2 FILLER_48_2428 ();
 sg13g2_decap_8 FILLER_48_2434 ();
 sg13g2_fill_2 FILLER_48_2441 ();
 sg13g2_fill_1 FILLER_48_2443 ();
 sg13g2_fill_1 FILLER_48_2504 ();
 sg13g2_fill_1 FILLER_48_2622 ();
 sg13g2_fill_1 FILLER_48_2631 ();
 sg13g2_fill_1 FILLER_48_2636 ();
 sg13g2_fill_2 FILLER_48_2668 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_19 ();
 sg13g2_fill_2 FILLER_49_26 ();
 sg13g2_fill_1 FILLER_49_28 ();
 sg13g2_fill_2 FILLER_49_81 ();
 sg13g2_fill_1 FILLER_49_83 ();
 sg13g2_decap_4 FILLER_49_110 ();
 sg13g2_fill_2 FILLER_49_114 ();
 sg13g2_decap_4 FILLER_49_124 ();
 sg13g2_fill_2 FILLER_49_128 ();
 sg13g2_decap_4 FILLER_49_156 ();
 sg13g2_decap_8 FILLER_49_170 ();
 sg13g2_fill_2 FILLER_49_177 ();
 sg13g2_fill_1 FILLER_49_179 ();
 sg13g2_fill_1 FILLER_49_219 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_fill_2 FILLER_49_238 ();
 sg13g2_fill_1 FILLER_49_240 ();
 sg13g2_decap_4 FILLER_49_252 ();
 sg13g2_fill_2 FILLER_49_256 ();
 sg13g2_fill_2 FILLER_49_266 ();
 sg13g2_fill_1 FILLER_49_271 ();
 sg13g2_decap_8 FILLER_49_279 ();
 sg13g2_decap_8 FILLER_49_286 ();
 sg13g2_fill_1 FILLER_49_293 ();
 sg13g2_decap_8 FILLER_49_299 ();
 sg13g2_fill_1 FILLER_49_306 ();
 sg13g2_decap_4 FILLER_49_311 ();
 sg13g2_decap_4 FILLER_49_318 ();
 sg13g2_decap_8 FILLER_49_334 ();
 sg13g2_fill_2 FILLER_49_351 ();
 sg13g2_decap_8 FILLER_49_366 ();
 sg13g2_fill_2 FILLER_49_373 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_4 FILLER_49_399 ();
 sg13g2_fill_1 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_415 ();
 sg13g2_decap_8 FILLER_49_422 ();
 sg13g2_fill_2 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_440 ();
 sg13g2_decap_8 FILLER_49_447 ();
 sg13g2_decap_8 FILLER_49_454 ();
 sg13g2_fill_2 FILLER_49_465 ();
 sg13g2_fill_1 FILLER_49_467 ();
 sg13g2_decap_8 FILLER_49_471 ();
 sg13g2_decap_4 FILLER_49_478 ();
 sg13g2_fill_1 FILLER_49_482 ();
 sg13g2_fill_2 FILLER_49_503 ();
 sg13g2_decap_4 FILLER_49_519 ();
 sg13g2_decap_4 FILLER_49_528 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_4 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_566 ();
 sg13g2_decap_4 FILLER_49_573 ();
 sg13g2_fill_2 FILLER_49_581 ();
 sg13g2_fill_1 FILLER_49_583 ();
 sg13g2_decap_8 FILLER_49_600 ();
 sg13g2_decap_8 FILLER_49_607 ();
 sg13g2_decap_4 FILLER_49_614 ();
 sg13g2_fill_2 FILLER_49_634 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_fill_2 FILLER_49_660 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_4 FILLER_49_683 ();
 sg13g2_fill_1 FILLER_49_687 ();
 sg13g2_decap_8 FILLER_49_707 ();
 sg13g2_decap_4 FILLER_49_714 ();
 sg13g2_fill_2 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_787 ();
 sg13g2_decap_4 FILLER_49_794 ();
 sg13g2_decap_8 FILLER_49_827 ();
 sg13g2_decap_4 FILLER_49_834 ();
 sg13g2_decap_4 FILLER_49_870 ();
 sg13g2_fill_1 FILLER_49_874 ();
 sg13g2_fill_2 FILLER_49_888 ();
 sg13g2_fill_1 FILLER_49_902 ();
 sg13g2_decap_4 FILLER_49_952 ();
 sg13g2_fill_1 FILLER_49_956 ();
 sg13g2_decap_8 FILLER_49_961 ();
 sg13g2_decap_8 FILLER_49_968 ();
 sg13g2_decap_4 FILLER_49_975 ();
 sg13g2_fill_1 FILLER_49_979 ();
 sg13g2_decap_8 FILLER_49_985 ();
 sg13g2_decap_4 FILLER_49_992 ();
 sg13g2_fill_2 FILLER_49_996 ();
 sg13g2_fill_2 FILLER_49_1008 ();
 sg13g2_fill_1 FILLER_49_1075 ();
 sg13g2_decap_4 FILLER_49_1080 ();
 sg13g2_decap_8 FILLER_49_1120 ();
 sg13g2_decap_8 FILLER_49_1127 ();
 sg13g2_decap_8 FILLER_49_1134 ();
 sg13g2_decap_4 FILLER_49_1141 ();
 sg13g2_fill_1 FILLER_49_1145 ();
 sg13g2_decap_4 FILLER_49_1155 ();
 sg13g2_fill_1 FILLER_49_1159 ();
 sg13g2_decap_8 FILLER_49_1211 ();
 sg13g2_fill_1 FILLER_49_1218 ();
 sg13g2_decap_8 FILLER_49_1233 ();
 sg13g2_decap_8 FILLER_49_1240 ();
 sg13g2_decap_8 FILLER_49_1247 ();
 sg13g2_fill_2 FILLER_49_1254 ();
 sg13g2_fill_1 FILLER_49_1256 ();
 sg13g2_fill_1 FILLER_49_1270 ();
 sg13g2_fill_1 FILLER_49_1302 ();
 sg13g2_decap_8 FILLER_49_1345 ();
 sg13g2_decap_4 FILLER_49_1352 ();
 sg13g2_fill_2 FILLER_49_1356 ();
 sg13g2_decap_4 FILLER_49_1388 ();
 sg13g2_decap_4 FILLER_49_1418 ();
 sg13g2_fill_2 FILLER_49_1422 ();
 sg13g2_decap_8 FILLER_49_1433 ();
 sg13g2_decap_8 FILLER_49_1440 ();
 sg13g2_decap_8 FILLER_49_1447 ();
 sg13g2_fill_1 FILLER_49_1454 ();
 sg13g2_decap_8 FILLER_49_1492 ();
 sg13g2_decap_4 FILLER_49_1499 ();
 sg13g2_decap_8 FILLER_49_1507 ();
 sg13g2_decap_4 FILLER_49_1514 ();
 sg13g2_fill_1 FILLER_49_1522 ();
 sg13g2_decap_8 FILLER_49_1558 ();
 sg13g2_decap_8 FILLER_49_1565 ();
 sg13g2_decap_8 FILLER_49_1572 ();
 sg13g2_decap_4 FILLER_49_1579 ();
 sg13g2_fill_1 FILLER_49_1583 ();
 sg13g2_fill_1 FILLER_49_1590 ();
 sg13g2_decap_4 FILLER_49_1660 ();
 sg13g2_fill_1 FILLER_49_1664 ();
 sg13g2_decap_4 FILLER_49_1670 ();
 sg13g2_fill_2 FILLER_49_1674 ();
 sg13g2_fill_2 FILLER_49_1679 ();
 sg13g2_fill_2 FILLER_49_1707 ();
 sg13g2_decap_8 FILLER_49_1735 ();
 sg13g2_decap_4 FILLER_49_1742 ();
 sg13g2_fill_1 FILLER_49_1746 ();
 sg13g2_fill_2 FILLER_49_1750 ();
 sg13g2_decap_4 FILLER_49_1759 ();
 sg13g2_fill_1 FILLER_49_1763 ();
 sg13g2_fill_1 FILLER_49_1768 ();
 sg13g2_fill_1 FILLER_49_1774 ();
 sg13g2_fill_1 FILLER_49_1780 ();
 sg13g2_fill_2 FILLER_49_1786 ();
 sg13g2_fill_1 FILLER_49_1814 ();
 sg13g2_decap_4 FILLER_49_1828 ();
 sg13g2_fill_2 FILLER_49_1838 ();
 sg13g2_fill_1 FILLER_49_1840 ();
 sg13g2_fill_2 FILLER_49_1849 ();
 sg13g2_decap_8 FILLER_49_1862 ();
 sg13g2_decap_8 FILLER_49_1869 ();
 sg13g2_decap_4 FILLER_49_1876 ();
 sg13g2_fill_2 FILLER_49_1880 ();
 sg13g2_decap_4 FILLER_49_1887 ();
 sg13g2_fill_2 FILLER_49_1891 ();
 sg13g2_fill_2 FILLER_49_1904 ();
 sg13g2_decap_4 FILLER_49_1910 ();
 sg13g2_fill_2 FILLER_49_1914 ();
 sg13g2_fill_1 FILLER_49_1975 ();
 sg13g2_fill_1 FILLER_49_1988 ();
 sg13g2_fill_1 FILLER_49_2002 ();
 sg13g2_decap_8 FILLER_49_2011 ();
 sg13g2_fill_1 FILLER_49_2018 ();
 sg13g2_decap_8 FILLER_49_2049 ();
 sg13g2_fill_1 FILLER_49_2056 ();
 sg13g2_decap_8 FILLER_49_2063 ();
 sg13g2_decap_8 FILLER_49_2070 ();
 sg13g2_decap_8 FILLER_49_2077 ();
 sg13g2_decap_8 FILLER_49_2084 ();
 sg13g2_fill_1 FILLER_49_2091 ();
 sg13g2_decap_4 FILLER_49_2128 ();
 sg13g2_fill_1 FILLER_49_2132 ();
 sg13g2_fill_2 FILLER_49_2178 ();
 sg13g2_decap_8 FILLER_49_2190 ();
 sg13g2_decap_8 FILLER_49_2197 ();
 sg13g2_fill_2 FILLER_49_2204 ();
 sg13g2_decap_8 FILLER_49_2211 ();
 sg13g2_decap_8 FILLER_49_2218 ();
 sg13g2_decap_8 FILLER_49_2225 ();
 sg13g2_decap_8 FILLER_49_2232 ();
 sg13g2_fill_2 FILLER_49_2239 ();
 sg13g2_fill_1 FILLER_49_2245 ();
 sg13g2_fill_1 FILLER_49_2252 ();
 sg13g2_fill_1 FILLER_49_2268 ();
 sg13g2_fill_2 FILLER_49_2273 ();
 sg13g2_fill_2 FILLER_49_2279 ();
 sg13g2_fill_1 FILLER_49_2281 ();
 sg13g2_decap_8 FILLER_49_2294 ();
 sg13g2_decap_4 FILLER_49_2301 ();
 sg13g2_decap_8 FILLER_49_2317 ();
 sg13g2_fill_2 FILLER_49_2324 ();
 sg13g2_fill_1 FILLER_49_2393 ();
 sg13g2_decap_8 FILLER_49_2398 ();
 sg13g2_decap_8 FILLER_49_2405 ();
 sg13g2_decap_8 FILLER_49_2412 ();
 sg13g2_decap_8 FILLER_49_2419 ();
 sg13g2_fill_1 FILLER_49_2426 ();
 sg13g2_decap_8 FILLER_49_2434 ();
 sg13g2_decap_8 FILLER_49_2441 ();
 sg13g2_fill_2 FILLER_49_2452 ();
 sg13g2_decap_8 FILLER_49_2458 ();
 sg13g2_decap_4 FILLER_49_2465 ();
 sg13g2_fill_1 FILLER_49_2469 ();
 sg13g2_fill_1 FILLER_49_2534 ();
 sg13g2_fill_2 FILLER_49_2584 ();
 sg13g2_decap_8 FILLER_49_2614 ();
 sg13g2_decap_4 FILLER_49_2621 ();
 sg13g2_fill_2 FILLER_49_2625 ();
 sg13g2_decap_4 FILLER_49_2665 ();
 sg13g2_fill_1 FILLER_49_2669 ();
 sg13g2_fill_1 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_31 ();
 sg13g2_decap_4 FILLER_50_64 ();
 sg13g2_fill_2 FILLER_50_91 ();
 sg13g2_fill_1 FILLER_50_93 ();
 sg13g2_fill_2 FILLER_50_104 ();
 sg13g2_fill_2 FILLER_50_113 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_decap_8 FILLER_50_194 ();
 sg13g2_decap_4 FILLER_50_201 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_220 ();
 sg13g2_decap_8 FILLER_50_227 ();
 sg13g2_decap_8 FILLER_50_234 ();
 sg13g2_decap_4 FILLER_50_241 ();
 sg13g2_decap_8 FILLER_50_249 ();
 sg13g2_decap_8 FILLER_50_256 ();
 sg13g2_decap_8 FILLER_50_263 ();
 sg13g2_fill_2 FILLER_50_270 ();
 sg13g2_fill_1 FILLER_50_272 ();
 sg13g2_fill_1 FILLER_50_415 ();
 sg13g2_decap_8 FILLER_50_421 ();
 sg13g2_decap_8 FILLER_50_428 ();
 sg13g2_decap_8 FILLER_50_435 ();
 sg13g2_decap_8 FILLER_50_442 ();
 sg13g2_decap_8 FILLER_50_449 ();
 sg13g2_fill_2 FILLER_50_456 ();
 sg13g2_fill_1 FILLER_50_458 ();
 sg13g2_decap_8 FILLER_50_472 ();
 sg13g2_decap_8 FILLER_50_479 ();
 sg13g2_fill_2 FILLER_50_486 ();
 sg13g2_fill_1 FILLER_50_488 ();
 sg13g2_decap_8 FILLER_50_500 ();
 sg13g2_decap_8 FILLER_50_507 ();
 sg13g2_decap_4 FILLER_50_514 ();
 sg13g2_decap_8 FILLER_50_547 ();
 sg13g2_decap_8 FILLER_50_554 ();
 sg13g2_decap_8 FILLER_50_565 ();
 sg13g2_fill_2 FILLER_50_572 ();
 sg13g2_fill_1 FILLER_50_591 ();
 sg13g2_fill_2 FILLER_50_602 ();
 sg13g2_decap_8 FILLER_50_616 ();
 sg13g2_decap_8 FILLER_50_623 ();
 sg13g2_fill_2 FILLER_50_630 ();
 sg13g2_decap_8 FILLER_50_636 ();
 sg13g2_decap_4 FILLER_50_643 ();
 sg13g2_fill_1 FILLER_50_647 ();
 sg13g2_fill_2 FILLER_50_653 ();
 sg13g2_decap_8 FILLER_50_659 ();
 sg13g2_decap_4 FILLER_50_666 ();
 sg13g2_fill_2 FILLER_50_670 ();
 sg13g2_decap_8 FILLER_50_678 ();
 sg13g2_fill_1 FILLER_50_685 ();
 sg13g2_fill_1 FILLER_50_690 ();
 sg13g2_fill_1 FILLER_50_696 ();
 sg13g2_fill_1 FILLER_50_701 ();
 sg13g2_decap_8 FILLER_50_707 ();
 sg13g2_decap_8 FILLER_50_719 ();
 sg13g2_fill_1 FILLER_50_731 ();
 sg13g2_decap_8 FILLER_50_766 ();
 sg13g2_decap_4 FILLER_50_773 ();
 sg13g2_fill_1 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_786 ();
 sg13g2_fill_2 FILLER_50_793 ();
 sg13g2_decap_4 FILLER_50_800 ();
 sg13g2_decap_8 FILLER_50_845 ();
 sg13g2_decap_4 FILLER_50_852 ();
 sg13g2_fill_1 FILLER_50_856 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_fill_2 FILLER_50_868 ();
 sg13g2_fill_1 FILLER_50_908 ();
 sg13g2_fill_1 FILLER_50_920 ();
 sg13g2_decap_8 FILLER_50_962 ();
 sg13g2_fill_2 FILLER_50_969 ();
 sg13g2_fill_1 FILLER_50_971 ();
 sg13g2_fill_2 FILLER_50_998 ();
 sg13g2_fill_1 FILLER_50_1000 ();
 sg13g2_fill_2 FILLER_50_1007 ();
 sg13g2_decap_4 FILLER_50_1042 ();
 sg13g2_fill_1 FILLER_50_1046 ();
 sg13g2_fill_2 FILLER_50_1057 ();
 sg13g2_decap_4 FILLER_50_1082 ();
 sg13g2_fill_1 FILLER_50_1120 ();
 sg13g2_fill_2 FILLER_50_1131 ();
 sg13g2_fill_1 FILLER_50_1133 ();
 sg13g2_decap_8 FILLER_50_1139 ();
 sg13g2_decap_4 FILLER_50_1146 ();
 sg13g2_fill_1 FILLER_50_1150 ();
 sg13g2_fill_2 FILLER_50_1163 ();
 sg13g2_fill_2 FILLER_50_1170 ();
 sg13g2_decap_8 FILLER_50_1206 ();
 sg13g2_fill_2 FILLER_50_1213 ();
 sg13g2_fill_1 FILLER_50_1215 ();
 sg13g2_decap_8 FILLER_50_1242 ();
 sg13g2_fill_2 FILLER_50_1253 ();
 sg13g2_decap_8 FILLER_50_1260 ();
 sg13g2_decap_8 FILLER_50_1267 ();
 sg13g2_fill_2 FILLER_50_1287 ();
 sg13g2_decap_4 FILLER_50_1304 ();
 sg13g2_fill_2 FILLER_50_1308 ();
 sg13g2_decap_8 FILLER_50_1319 ();
 sg13g2_decap_4 FILLER_50_1326 ();
 sg13g2_fill_1 FILLER_50_1330 ();
 sg13g2_fill_1 FILLER_50_1340 ();
 sg13g2_fill_1 FILLER_50_1433 ();
 sg13g2_fill_1 FILLER_50_1465 ();
 sg13g2_fill_2 FILLER_50_1470 ();
 sg13g2_decap_8 FILLER_50_1476 ();
 sg13g2_decap_8 FILLER_50_1483 ();
 sg13g2_fill_2 FILLER_50_1503 ();
 sg13g2_decap_4 FILLER_50_1548 ();
 sg13g2_fill_1 FILLER_50_1552 ();
 sg13g2_fill_1 FILLER_50_1556 ();
 sg13g2_fill_2 FILLER_50_1561 ();
 sg13g2_fill_1 FILLER_50_1563 ();
 sg13g2_fill_1 FILLER_50_1597 ();
 sg13g2_fill_1 FILLER_50_1602 ();
 sg13g2_fill_2 FILLER_50_1607 ();
 sg13g2_fill_1 FILLER_50_1609 ();
 sg13g2_decap_4 FILLER_50_1614 ();
 sg13g2_fill_1 FILLER_50_1618 ();
 sg13g2_decap_4 FILLER_50_1624 ();
 sg13g2_fill_2 FILLER_50_1674 ();
 sg13g2_fill_2 FILLER_50_1684 ();
 sg13g2_fill_1 FILLER_50_1686 ();
 sg13g2_decap_8 FILLER_50_1691 ();
 sg13g2_fill_1 FILLER_50_1698 ();
 sg13g2_decap_8 FILLER_50_1706 ();
 sg13g2_fill_2 FILLER_50_1713 ();
 sg13g2_decap_4 FILLER_50_1720 ();
 sg13g2_fill_2 FILLER_50_1724 ();
 sg13g2_fill_1 FILLER_50_1739 ();
 sg13g2_decap_8 FILLER_50_1776 ();
 sg13g2_fill_2 FILLER_50_1828 ();
 sg13g2_fill_1 FILLER_50_1846 ();
 sg13g2_fill_2 FILLER_50_1862 ();
 sg13g2_decap_8 FILLER_50_1871 ();
 sg13g2_decap_8 FILLER_50_1884 ();
 sg13g2_fill_1 FILLER_50_1891 ();
 sg13g2_decap_4 FILLER_50_1897 ();
 sg13g2_fill_2 FILLER_50_1901 ();
 sg13g2_fill_1 FILLER_50_1958 ();
 sg13g2_fill_1 FILLER_50_1967 ();
 sg13g2_fill_2 FILLER_50_1974 ();
 sg13g2_fill_2 FILLER_50_1981 ();
 sg13g2_fill_1 FILLER_50_2007 ();
 sg13g2_decap_4 FILLER_50_2036 ();
 sg13g2_fill_1 FILLER_50_2044 ();
 sg13g2_decap_8 FILLER_50_2070 ();
 sg13g2_decap_8 FILLER_50_2077 ();
 sg13g2_decap_8 FILLER_50_2084 ();
 sg13g2_decap_8 FILLER_50_2099 ();
 sg13g2_fill_1 FILLER_50_2106 ();
 sg13g2_decap_8 FILLER_50_2111 ();
 sg13g2_decap_8 FILLER_50_2118 ();
 sg13g2_fill_2 FILLER_50_2125 ();
 sg13g2_decap_8 FILLER_50_2133 ();
 sg13g2_fill_2 FILLER_50_2140 ();
 sg13g2_decap_8 FILLER_50_2229 ();
 sg13g2_decap_8 FILLER_50_2236 ();
 sg13g2_fill_2 FILLER_50_2243 ();
 sg13g2_fill_1 FILLER_50_2245 ();
 sg13g2_decap_4 FILLER_50_2252 ();
 sg13g2_decap_4 FILLER_50_2282 ();
 sg13g2_fill_2 FILLER_50_2286 ();
 sg13g2_decap_8 FILLER_50_2294 ();
 sg13g2_fill_2 FILLER_50_2301 ();
 sg13g2_decap_4 FILLER_50_2333 ();
 sg13g2_decap_8 FILLER_50_2341 ();
 sg13g2_fill_1 FILLER_50_2348 ();
 sg13g2_decap_8 FILLER_50_2353 ();
 sg13g2_fill_1 FILLER_50_2360 ();
 sg13g2_fill_1 FILLER_50_2365 ();
 sg13g2_decap_8 FILLER_50_2374 ();
 sg13g2_decap_8 FILLER_50_2381 ();
 sg13g2_fill_1 FILLER_50_2388 ();
 sg13g2_decap_8 FILLER_50_2393 ();
 sg13g2_fill_1 FILLER_50_2400 ();
 sg13g2_decap_8 FILLER_50_2463 ();
 sg13g2_decap_4 FILLER_50_2470 ();
 sg13g2_fill_2 FILLER_50_2474 ();
 sg13g2_fill_2 FILLER_50_2480 ();
 sg13g2_fill_1 FILLER_50_2482 ();
 sg13g2_fill_1 FILLER_50_2487 ();
 sg13g2_decap_8 FILLER_50_2504 ();
 sg13g2_decap_8 FILLER_50_2511 ();
 sg13g2_decap_8 FILLER_50_2518 ();
 sg13g2_decap_4 FILLER_50_2525 ();
 sg13g2_decap_8 FILLER_50_2563 ();
 sg13g2_decap_8 FILLER_50_2570 ();
 sg13g2_decap_4 FILLER_50_2577 ();
 sg13g2_fill_2 FILLER_50_2581 ();
 sg13g2_decap_4 FILLER_50_2596 ();
 sg13g2_decap_8 FILLER_50_2604 ();
 sg13g2_decap_8 FILLER_50_2611 ();
 sg13g2_decap_8 FILLER_50_2618 ();
 sg13g2_decap_4 FILLER_50_2625 ();
 sg13g2_fill_1 FILLER_50_2629 ();
 sg13g2_decap_8 FILLER_50_2634 ();
 sg13g2_decap_8 FILLER_50_2641 ();
 sg13g2_decap_8 FILLER_50_2648 ();
 sg13g2_decap_8 FILLER_50_2655 ();
 sg13g2_decap_8 FILLER_50_2662 ();
 sg13g2_fill_1 FILLER_50_2669 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_4 FILLER_51_14 ();
 sg13g2_fill_1 FILLER_51_18 ();
 sg13g2_fill_1 FILLER_51_59 ();
 sg13g2_decap_4 FILLER_51_70 ();
 sg13g2_fill_2 FILLER_51_74 ();
 sg13g2_decap_8 FILLER_51_81 ();
 sg13g2_decap_8 FILLER_51_88 ();
 sg13g2_decap_8 FILLER_51_95 ();
 sg13g2_decap_8 FILLER_51_102 ();
 sg13g2_fill_2 FILLER_51_109 ();
 sg13g2_fill_1 FILLER_51_111 ();
 sg13g2_fill_2 FILLER_51_127 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_decap_4 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_180 ();
 sg13g2_decap_4 FILLER_51_217 ();
 sg13g2_fill_1 FILLER_51_221 ();
 sg13g2_decap_8 FILLER_51_226 ();
 sg13g2_decap_8 FILLER_51_233 ();
 sg13g2_decap_8 FILLER_51_240 ();
 sg13g2_decap_8 FILLER_51_247 ();
 sg13g2_decap_8 FILLER_51_254 ();
 sg13g2_decap_4 FILLER_51_261 ();
 sg13g2_fill_2 FILLER_51_265 ();
 sg13g2_fill_2 FILLER_51_271 ();
 sg13g2_fill_1 FILLER_51_273 ();
 sg13g2_decap_8 FILLER_51_278 ();
 sg13g2_decap_4 FILLER_51_285 ();
 sg13g2_fill_2 FILLER_51_289 ();
 sg13g2_decap_8 FILLER_51_295 ();
 sg13g2_fill_2 FILLER_51_307 ();
 sg13g2_decap_8 FILLER_51_319 ();
 sg13g2_decap_4 FILLER_51_330 ();
 sg13g2_fill_2 FILLER_51_334 ();
 sg13g2_fill_1 FILLER_51_343 ();
 sg13g2_fill_1 FILLER_51_350 ();
 sg13g2_fill_1 FILLER_51_358 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_fill_1 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_409 ();
 sg13g2_decap_4 FILLER_51_416 ();
 sg13g2_fill_1 FILLER_51_420 ();
 sg13g2_fill_2 FILLER_51_425 ();
 sg13g2_decap_4 FILLER_51_436 ();
 sg13g2_fill_1 FILLER_51_440 ();
 sg13g2_fill_1 FILLER_51_444 ();
 sg13g2_fill_2 FILLER_51_448 ();
 sg13g2_fill_2 FILLER_51_457 ();
 sg13g2_decap_4 FILLER_51_478 ();
 sg13g2_fill_2 FILLER_51_482 ();
 sg13g2_fill_1 FILLER_51_518 ();
 sg13g2_decap_8 FILLER_51_528 ();
 sg13g2_decap_8 FILLER_51_535 ();
 sg13g2_decap_4 FILLER_51_542 ();
 sg13g2_decap_8 FILLER_51_550 ();
 sg13g2_fill_2 FILLER_51_557 ();
 sg13g2_decap_8 FILLER_51_569 ();
 sg13g2_decap_4 FILLER_51_576 ();
 sg13g2_decap_8 FILLER_51_623 ();
 sg13g2_decap_4 FILLER_51_630 ();
 sg13g2_fill_1 FILLER_51_634 ();
 sg13g2_decap_8 FILLER_51_639 ();
 sg13g2_fill_2 FILLER_51_646 ();
 sg13g2_fill_1 FILLER_51_648 ();
 sg13g2_fill_1 FILLER_51_664 ();
 sg13g2_fill_1 FILLER_51_673 ();
 sg13g2_fill_2 FILLER_51_678 ();
 sg13g2_decap_8 FILLER_51_688 ();
 sg13g2_decap_4 FILLER_51_698 ();
 sg13g2_fill_2 FILLER_51_702 ();
 sg13g2_decap_8 FILLER_51_708 ();
 sg13g2_decap_4 FILLER_51_715 ();
 sg13g2_fill_1 FILLER_51_719 ();
 sg13g2_fill_1 FILLER_51_751 ();
 sg13g2_fill_1 FILLER_51_809 ();
 sg13g2_fill_1 FILLER_51_816 ();
 sg13g2_decap_8 FILLER_51_821 ();
 sg13g2_fill_2 FILLER_51_828 ();
 sg13g2_fill_2 FILLER_51_835 ();
 sg13g2_fill_1 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_843 ();
 sg13g2_fill_1 FILLER_51_850 ();
 sg13g2_decap_4 FILLER_51_882 ();
 sg13g2_fill_1 FILLER_51_886 ();
 sg13g2_fill_2 FILLER_51_892 ();
 sg13g2_fill_1 FILLER_51_920 ();
 sg13g2_fill_1 FILLER_51_952 ();
 sg13g2_fill_1 FILLER_51_959 ();
 sg13g2_decap_4 FILLER_51_966 ();
 sg13g2_fill_1 FILLER_51_970 ();
 sg13g2_decap_4 FILLER_51_1040 ();
 sg13g2_fill_1 FILLER_51_1044 ();
 sg13g2_decap_8 FILLER_51_1074 ();
 sg13g2_decap_8 FILLER_51_1081 ();
 sg13g2_decap_8 FILLER_51_1088 ();
 sg13g2_decap_8 FILLER_51_1095 ();
 sg13g2_fill_2 FILLER_51_1102 ();
 sg13g2_decap_4 FILLER_51_1130 ();
 sg13g2_fill_2 FILLER_51_1134 ();
 sg13g2_decap_8 FILLER_51_1162 ();
 sg13g2_decap_8 FILLER_51_1169 ();
 sg13g2_decap_8 FILLER_51_1176 ();
 sg13g2_fill_1 FILLER_51_1183 ();
 sg13g2_decap_8 FILLER_51_1188 ();
 sg13g2_decap_8 FILLER_51_1195 ();
 sg13g2_fill_2 FILLER_51_1202 ();
 sg13g2_fill_1 FILLER_51_1204 ();
 sg13g2_fill_1 FILLER_51_1214 ();
 sg13g2_fill_1 FILLER_51_1241 ();
 sg13g2_fill_2 FILLER_51_1248 ();
 sg13g2_fill_1 FILLER_51_1253 ();
 sg13g2_fill_2 FILLER_51_1312 ();
 sg13g2_fill_1 FILLER_51_1314 ();
 sg13g2_decap_4 FILLER_51_1346 ();
 sg13g2_fill_1 FILLER_51_1350 ();
 sg13g2_decap_4 FILLER_51_1355 ();
 sg13g2_decap_8 FILLER_51_1365 ();
 sg13g2_fill_2 FILLER_51_1416 ();
 sg13g2_fill_1 FILLER_51_1418 ();
 sg13g2_fill_1 FILLER_51_1445 ();
 sg13g2_decap_8 FILLER_51_1472 ();
 sg13g2_fill_1 FILLER_51_1479 ();
 sg13g2_decap_4 FILLER_51_1486 ();
 sg13g2_decap_4 FILLER_51_1539 ();
 sg13g2_fill_1 FILLER_51_1543 ();
 sg13g2_fill_1 FILLER_51_1587 ();
 sg13g2_fill_2 FILLER_51_1605 ();
 sg13g2_fill_2 FILLER_51_1610 ();
 sg13g2_fill_1 FILLER_51_1612 ();
 sg13g2_fill_2 FILLER_51_1622 ();
 sg13g2_fill_2 FILLER_51_1633 ();
 sg13g2_fill_1 FILLER_51_1635 ();
 sg13g2_fill_2 FILLER_51_1659 ();
 sg13g2_fill_1 FILLER_51_1661 ();
 sg13g2_decap_8 FILLER_51_1669 ();
 sg13g2_fill_2 FILLER_51_1707 ();
 sg13g2_decap_8 FILLER_51_1748 ();
 sg13g2_decap_4 FILLER_51_1755 ();
 sg13g2_fill_2 FILLER_51_1759 ();
 sg13g2_fill_2 FILLER_51_1766 ();
 sg13g2_decap_4 FILLER_51_1772 ();
 sg13g2_fill_2 FILLER_51_1776 ();
 sg13g2_fill_2 FILLER_51_1782 ();
 sg13g2_fill_1 FILLER_51_1788 ();
 sg13g2_decap_8 FILLER_51_1800 ();
 sg13g2_fill_1 FILLER_51_1827 ();
 sg13g2_fill_2 FILLER_51_1833 ();
 sg13g2_fill_1 FILLER_51_1835 ();
 sg13g2_decap_4 FILLER_51_1874 ();
 sg13g2_fill_2 FILLER_51_1878 ();
 sg13g2_fill_1 FILLER_51_1884 ();
 sg13g2_fill_2 FILLER_51_1898 ();
 sg13g2_fill_2 FILLER_51_1904 ();
 sg13g2_fill_1 FILLER_51_1906 ();
 sg13g2_fill_1 FILLER_51_1938 ();
 sg13g2_decap_4 FILLER_51_1947 ();
 sg13g2_fill_1 FILLER_51_1998 ();
 sg13g2_decap_8 FILLER_51_2007 ();
 sg13g2_fill_1 FILLER_51_2014 ();
 sg13g2_decap_8 FILLER_51_2041 ();
 sg13g2_decap_8 FILLER_51_2048 ();
 sg13g2_fill_2 FILLER_51_2055 ();
 sg13g2_decap_8 FILLER_51_2062 ();
 sg13g2_decap_8 FILLER_51_2069 ();
 sg13g2_fill_2 FILLER_51_2076 ();
 sg13g2_fill_1 FILLER_51_2078 ();
 sg13g2_decap_4 FILLER_51_2082 ();
 sg13g2_fill_2 FILLER_51_2086 ();
 sg13g2_decap_8 FILLER_51_2126 ();
 sg13g2_decap_4 FILLER_51_2133 ();
 sg13g2_fill_2 FILLER_51_2137 ();
 sg13g2_fill_2 FILLER_51_2143 ();
 sg13g2_fill_1 FILLER_51_2145 ();
 sg13g2_decap_8 FILLER_51_2172 ();
 sg13g2_decap_8 FILLER_51_2179 ();
 sg13g2_decap_8 FILLER_51_2186 ();
 sg13g2_fill_2 FILLER_51_2229 ();
 sg13g2_fill_1 FILLER_51_2231 ();
 sg13g2_fill_2 FILLER_51_2251 ();
 sg13g2_decap_4 FILLER_51_2293 ();
 sg13g2_fill_1 FILLER_51_2297 ();
 sg13g2_decap_8 FILLER_51_2332 ();
 sg13g2_decap_8 FILLER_51_2339 ();
 sg13g2_decap_8 FILLER_51_2346 ();
 sg13g2_decap_8 FILLER_51_2353 ();
 sg13g2_decap_4 FILLER_51_2360 ();
 sg13g2_fill_1 FILLER_51_2364 ();
 sg13g2_decap_8 FILLER_51_2371 ();
 sg13g2_decap_8 FILLER_51_2378 ();
 sg13g2_decap_8 FILLER_51_2385 ();
 sg13g2_decap_8 FILLER_51_2392 ();
 sg13g2_fill_2 FILLER_51_2399 ();
 sg13g2_fill_1 FILLER_51_2401 ();
 sg13g2_decap_8 FILLER_51_2428 ();
 sg13g2_decap_8 FILLER_51_2435 ();
 sg13g2_fill_2 FILLER_51_2442 ();
 sg13g2_fill_1 FILLER_51_2444 ();
 sg13g2_decap_8 FILLER_51_2449 ();
 sg13g2_decap_4 FILLER_51_2456 ();
 sg13g2_fill_2 FILLER_51_2460 ();
 sg13g2_decap_8 FILLER_51_2498 ();
 sg13g2_decap_8 FILLER_51_2505 ();
 sg13g2_decap_4 FILLER_51_2512 ();
 sg13g2_decap_8 FILLER_51_2520 ();
 sg13g2_decap_8 FILLER_51_2527 ();
 sg13g2_fill_2 FILLER_51_2534 ();
 sg13g2_fill_2 FILLER_51_2544 ();
 sg13g2_fill_1 FILLER_51_2546 ();
 sg13g2_decap_4 FILLER_51_2580 ();
 sg13g2_fill_2 FILLER_51_2584 ();
 sg13g2_fill_2 FILLER_51_2589 ();
 sg13g2_fill_1 FILLER_51_2591 ();
 sg13g2_decap_8 FILLER_51_2622 ();
 sg13g2_decap_8 FILLER_51_2629 ();
 sg13g2_decap_8 FILLER_51_2636 ();
 sg13g2_decap_8 FILLER_51_2643 ();
 sg13g2_decap_8 FILLER_51_2650 ();
 sg13g2_decap_8 FILLER_51_2657 ();
 sg13g2_decap_4 FILLER_51_2664 ();
 sg13g2_fill_2 FILLER_51_2668 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_fill_1 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_39 ();
 sg13g2_fill_1 FILLER_52_60 ();
 sg13g2_decap_8 FILLER_52_73 ();
 sg13g2_decap_8 FILLER_52_80 ();
 sg13g2_decap_4 FILLER_52_87 ();
 sg13g2_fill_2 FILLER_52_91 ();
 sg13g2_decap_4 FILLER_52_103 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_4 FILLER_52_161 ();
 sg13g2_fill_1 FILLER_52_165 ();
 sg13g2_decap_8 FILLER_52_179 ();
 sg13g2_decap_8 FILLER_52_186 ();
 sg13g2_decap_4 FILLER_52_193 ();
 sg13g2_decap_8 FILLER_52_202 ();
 sg13g2_decap_8 FILLER_52_209 ();
 sg13g2_decap_8 FILLER_52_216 ();
 sg13g2_decap_8 FILLER_52_223 ();
 sg13g2_decap_8 FILLER_52_230 ();
 sg13g2_fill_1 FILLER_52_237 ();
 sg13g2_decap_4 FILLER_52_247 ();
 sg13g2_decap_8 FILLER_52_255 ();
 sg13g2_decap_8 FILLER_52_262 ();
 sg13g2_decap_4 FILLER_52_269 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_4 FILLER_52_301 ();
 sg13g2_fill_2 FILLER_52_315 ();
 sg13g2_fill_1 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_325 ();
 sg13g2_fill_2 FILLER_52_333 ();
 sg13g2_decap_8 FILLER_52_383 ();
 sg13g2_fill_2 FILLER_52_390 ();
 sg13g2_fill_1 FILLER_52_395 ();
 sg13g2_decap_4 FILLER_52_419 ();
 sg13g2_fill_1 FILLER_52_423 ();
 sg13g2_decap_8 FILLER_52_480 ();
 sg13g2_decap_4 FILLER_52_487 ();
 sg13g2_fill_1 FILLER_52_495 ();
 sg13g2_fill_1 FILLER_52_520 ();
 sg13g2_decap_8 FILLER_52_526 ();
 sg13g2_decap_8 FILLER_52_533 ();
 sg13g2_fill_2 FILLER_52_540 ();
 sg13g2_fill_2 FILLER_52_562 ();
 sg13g2_fill_1 FILLER_52_564 ();
 sg13g2_decap_8 FILLER_52_570 ();
 sg13g2_fill_1 FILLER_52_577 ();
 sg13g2_fill_2 FILLER_52_583 ();
 sg13g2_fill_1 FILLER_52_585 ();
 sg13g2_fill_1 FILLER_52_594 ();
 sg13g2_fill_1 FILLER_52_600 ();
 sg13g2_fill_2 FILLER_52_608 ();
 sg13g2_fill_2 FILLER_52_621 ();
 sg13g2_fill_2 FILLER_52_643 ();
 sg13g2_decap_8 FILLER_52_648 ();
 sg13g2_decap_8 FILLER_52_655 ();
 sg13g2_decap_4 FILLER_52_662 ();
 sg13g2_fill_2 FILLER_52_666 ();
 sg13g2_fill_2 FILLER_52_678 ();
 sg13g2_fill_1 FILLER_52_680 ();
 sg13g2_decap_4 FILLER_52_685 ();
 sg13g2_fill_2 FILLER_52_689 ();
 sg13g2_decap_4 FILLER_52_709 ();
 sg13g2_fill_2 FILLER_52_713 ();
 sg13g2_decap_8 FILLER_52_741 ();
 sg13g2_fill_2 FILLER_52_748 ();
 sg13g2_fill_1 FILLER_52_750 ();
 sg13g2_fill_2 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_fill_1 FILLER_52_791 ();
 sg13g2_decap_4 FILLER_52_802 ();
 sg13g2_fill_2 FILLER_52_812 ();
 sg13g2_fill_1 FILLER_52_814 ();
 sg13g2_decap_4 FILLER_52_819 ();
 sg13g2_fill_1 FILLER_52_855 ();
 sg13g2_decap_8 FILLER_52_862 ();
 sg13g2_decap_8 FILLER_52_869 ();
 sg13g2_fill_1 FILLER_52_881 ();
 sg13g2_decap_8 FILLER_52_891 ();
 sg13g2_decap_4 FILLER_52_898 ();
 sg13g2_fill_1 FILLER_52_902 ();
 sg13g2_fill_2 FILLER_52_906 ();
 sg13g2_fill_1 FILLER_52_908 ();
 sg13g2_fill_1 FILLER_52_961 ();
 sg13g2_fill_2 FILLER_52_967 ();
 sg13g2_fill_2 FILLER_52_998 ();
 sg13g2_fill_1 FILLER_52_1008 ();
 sg13g2_decap_8 FILLER_52_1038 ();
 sg13g2_decap_8 FILLER_52_1045 ();
 sg13g2_decap_8 FILLER_52_1052 ();
 sg13g2_decap_8 FILLER_52_1064 ();
 sg13g2_decap_8 FILLER_52_1071 ();
 sg13g2_decap_8 FILLER_52_1078 ();
 sg13g2_decap_8 FILLER_52_1085 ();
 sg13g2_decap_8 FILLER_52_1092 ();
 sg13g2_fill_2 FILLER_52_1099 ();
 sg13g2_decap_8 FILLER_52_1114 ();
 sg13g2_decap_4 FILLER_52_1121 ();
 sg13g2_decap_8 FILLER_52_1140 ();
 sg13g2_decap_8 FILLER_52_1147 ();
 sg13g2_decap_8 FILLER_52_1154 ();
 sg13g2_decap_8 FILLER_52_1161 ();
 sg13g2_decap_4 FILLER_52_1168 ();
 sg13g2_fill_2 FILLER_52_1172 ();
 sg13g2_decap_8 FILLER_52_1178 ();
 sg13g2_decap_8 FILLER_52_1185 ();
 sg13g2_decap_4 FILLER_52_1192 ();
 sg13g2_fill_2 FILLER_52_1233 ();
 sg13g2_fill_2 FILLER_52_1240 ();
 sg13g2_fill_1 FILLER_52_1242 ();
 sg13g2_decap_4 FILLER_52_1262 ();
 sg13g2_fill_2 FILLER_52_1266 ();
 sg13g2_fill_2 FILLER_52_1301 ();
 sg13g2_decap_4 FILLER_52_1312 ();
 sg13g2_decap_8 FILLER_52_1321 ();
 sg13g2_fill_1 FILLER_52_1328 ();
 sg13g2_fill_1 FILLER_52_1333 ();
 sg13g2_decap_8 FILLER_52_1364 ();
 sg13g2_decap_8 FILLER_52_1371 ();
 sg13g2_fill_1 FILLER_52_1378 ();
 sg13g2_decap_8 FILLER_52_1388 ();
 sg13g2_fill_2 FILLER_52_1395 ();
 sg13g2_fill_1 FILLER_52_1397 ();
 sg13g2_decap_4 FILLER_52_1424 ();
 sg13g2_decap_8 FILLER_52_1433 ();
 sg13g2_decap_4 FILLER_52_1440 ();
 sg13g2_decap_4 FILLER_52_1453 ();
 sg13g2_fill_2 FILLER_52_1457 ();
 sg13g2_decap_8 FILLER_52_1464 ();
 sg13g2_decap_4 FILLER_52_1471 ();
 sg13g2_fill_1 FILLER_52_1475 ();
 sg13g2_decap_4 FILLER_52_1502 ();
 sg13g2_fill_1 FILLER_52_1506 ();
 sg13g2_decap_4 FILLER_52_1511 ();
 sg13g2_fill_1 FILLER_52_1530 ();
 sg13g2_fill_1 FILLER_52_1557 ();
 sg13g2_decap_4 FILLER_52_1615 ();
 sg13g2_fill_2 FILLER_52_1662 ();
 sg13g2_fill_1 FILLER_52_1664 ();
 sg13g2_fill_1 FILLER_52_1695 ();
 sg13g2_decap_8 FILLER_52_1700 ();
 sg13g2_decap_8 FILLER_52_1707 ();
 sg13g2_fill_1 FILLER_52_1714 ();
 sg13g2_decap_4 FILLER_52_1724 ();
 sg13g2_fill_2 FILLER_52_1728 ();
 sg13g2_decap_8 FILLER_52_1734 ();
 sg13g2_decap_8 FILLER_52_1741 ();
 sg13g2_decap_8 FILLER_52_1748 ();
 sg13g2_decap_4 FILLER_52_1755 ();
 sg13g2_fill_2 FILLER_52_1759 ();
 sg13g2_decap_8 FILLER_52_1787 ();
 sg13g2_decap_8 FILLER_52_1794 ();
 sg13g2_decap_4 FILLER_52_1801 ();
 sg13g2_fill_1 FILLER_52_1813 ();
 sg13g2_fill_1 FILLER_52_1851 ();
 sg13g2_decap_8 FILLER_52_1856 ();
 sg13g2_fill_1 FILLER_52_1863 ();
 sg13g2_decap_8 FILLER_52_1868 ();
 sg13g2_fill_1 FILLER_52_1875 ();
 sg13g2_fill_1 FILLER_52_1884 ();
 sg13g2_decap_8 FILLER_52_1911 ();
 sg13g2_fill_1 FILLER_52_1918 ();
 sg13g2_decap_4 FILLER_52_1923 ();
 sg13g2_decap_8 FILLER_52_1930 ();
 sg13g2_fill_2 FILLER_52_1937 ();
 sg13g2_fill_1 FILLER_52_1939 ();
 sg13g2_fill_2 FILLER_52_1953 ();
 sg13g2_fill_1 FILLER_52_1955 ();
 sg13g2_fill_1 FILLER_52_1999 ();
 sg13g2_fill_1 FILLER_52_2004 ();
 sg13g2_fill_1 FILLER_52_2036 ();
 sg13g2_decap_4 FILLER_52_2063 ();
 sg13g2_fill_1 FILLER_52_2067 ();
 sg13g2_decap_8 FILLER_52_2072 ();
 sg13g2_decap_4 FILLER_52_2079 ();
 sg13g2_fill_2 FILLER_52_2091 ();
 sg13g2_decap_8 FILLER_52_2120 ();
 sg13g2_decap_4 FILLER_52_2135 ();
 sg13g2_decap_8 FILLER_52_2144 ();
 sg13g2_decap_8 FILLER_52_2151 ();
 sg13g2_decap_8 FILLER_52_2158 ();
 sg13g2_decap_8 FILLER_52_2165 ();
 sg13g2_decap_8 FILLER_52_2172 ();
 sg13g2_decap_8 FILLER_52_2179 ();
 sg13g2_fill_1 FILLER_52_2186 ();
 sg13g2_fill_2 FILLER_52_2196 ();
 sg13g2_fill_1 FILLER_52_2240 ();
 sg13g2_fill_2 FILLER_52_2249 ();
 sg13g2_fill_2 FILLER_52_2257 ();
 sg13g2_fill_1 FILLER_52_2284 ();
 sg13g2_decap_8 FILLER_52_2291 ();
 sg13g2_fill_2 FILLER_52_2298 ();
 sg13g2_fill_1 FILLER_52_2300 ();
 sg13g2_decap_8 FILLER_52_2305 ();
 sg13g2_fill_1 FILLER_52_2316 ();
 sg13g2_fill_2 FILLER_52_2343 ();
 sg13g2_decap_8 FILLER_52_2421 ();
 sg13g2_decap_4 FILLER_52_2432 ();
 sg13g2_fill_2 FILLER_52_2436 ();
 sg13g2_decap_8 FILLER_52_2494 ();
 sg13g2_decap_8 FILLER_52_2501 ();
 sg13g2_fill_2 FILLER_52_2508 ();
 sg13g2_fill_1 FILLER_52_2510 ();
 sg13g2_fill_2 FILLER_52_2522 ();
 sg13g2_fill_2 FILLER_52_2538 ();
 sg13g2_decap_4 FILLER_52_2590 ();
 sg13g2_fill_2 FILLER_52_2594 ();
 sg13g2_fill_1 FILLER_52_2600 ();
 sg13g2_decap_4 FILLER_52_2631 ();
 sg13g2_fill_1 FILLER_52_2635 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_1 FILLER_53_2 ();
 sg13g2_decap_8 FILLER_53_33 ();
 sg13g2_decap_8 FILLER_53_40 ();
 sg13g2_decap_8 FILLER_53_47 ();
 sg13g2_decap_8 FILLER_53_54 ();
 sg13g2_fill_1 FILLER_53_71 ();
 sg13g2_fill_2 FILLER_53_77 ();
 sg13g2_fill_2 FILLER_53_105 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_1 FILLER_53_113 ();
 sg13g2_fill_2 FILLER_53_119 ();
 sg13g2_decap_4 FILLER_53_126 ();
 sg13g2_fill_2 FILLER_53_130 ();
 sg13g2_decap_8 FILLER_53_137 ();
 sg13g2_decap_4 FILLER_53_144 ();
 sg13g2_decap_8 FILLER_53_162 ();
 sg13g2_decap_4 FILLER_53_169 ();
 sg13g2_fill_1 FILLER_53_194 ();
 sg13g2_fill_1 FILLER_53_199 ();
 sg13g2_fill_2 FILLER_53_204 ();
 sg13g2_fill_1 FILLER_53_206 ();
 sg13g2_decap_8 FILLER_53_283 ();
 sg13g2_decap_8 FILLER_53_290 ();
 sg13g2_decap_8 FILLER_53_297 ();
 sg13g2_fill_2 FILLER_53_304 ();
 sg13g2_fill_1 FILLER_53_306 ();
 sg13g2_fill_2 FILLER_53_392 ();
 sg13g2_fill_1 FILLER_53_413 ();
 sg13g2_fill_1 FILLER_53_421 ();
 sg13g2_fill_1 FILLER_53_436 ();
 sg13g2_fill_2 FILLER_53_478 ();
 sg13g2_fill_1 FILLER_53_480 ();
 sg13g2_fill_2 FILLER_53_524 ();
 sg13g2_decap_8 FILLER_53_544 ();
 sg13g2_fill_2 FILLER_53_551 ();
 sg13g2_fill_1 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_566 ();
 sg13g2_decap_4 FILLER_53_573 ();
 sg13g2_fill_1 FILLER_53_654 ();
 sg13g2_decap_4 FILLER_53_673 ();
 sg13g2_decap_8 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_712 ();
 sg13g2_decap_8 FILLER_53_719 ();
 sg13g2_fill_2 FILLER_53_726 ();
 sg13g2_fill_1 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_739 ();
 sg13g2_fill_1 FILLER_53_746 ();
 sg13g2_fill_1 FILLER_53_752 ();
 sg13g2_decap_4 FILLER_53_758 ();
 sg13g2_decap_8 FILLER_53_825 ();
 sg13g2_decap_8 FILLER_53_836 ();
 sg13g2_fill_1 FILLER_53_912 ();
 sg13g2_fill_2 FILLER_53_935 ();
 sg13g2_fill_1 FILLER_53_937 ();
 sg13g2_fill_2 FILLER_53_941 ();
 sg13g2_fill_2 FILLER_53_962 ();
 sg13g2_decap_8 FILLER_53_1003 ();
 sg13g2_decap_4 FILLER_53_1015 ();
 sg13g2_fill_2 FILLER_53_1019 ();
 sg13g2_decap_8 FILLER_53_1025 ();
 sg13g2_decap_8 FILLER_53_1032 ();
 sg13g2_decap_8 FILLER_53_1039 ();
 sg13g2_decap_8 FILLER_53_1046 ();
 sg13g2_decap_8 FILLER_53_1053 ();
 sg13g2_decap_8 FILLER_53_1060 ();
 sg13g2_decap_8 FILLER_53_1067 ();
 sg13g2_decap_8 FILLER_53_1074 ();
 sg13g2_decap_8 FILLER_53_1081 ();
 sg13g2_decap_8 FILLER_53_1088 ();
 sg13g2_decap_8 FILLER_53_1095 ();
 sg13g2_decap_4 FILLER_53_1102 ();
 sg13g2_decap_8 FILLER_53_1133 ();
 sg13g2_decap_8 FILLER_53_1140 ();
 sg13g2_decap_8 FILLER_53_1147 ();
 sg13g2_decap_8 FILLER_53_1154 ();
 sg13g2_fill_2 FILLER_53_1161 ();
 sg13g2_fill_1 FILLER_53_1163 ();
 sg13g2_decap_8 FILLER_53_1168 ();
 sg13g2_decap_4 FILLER_53_1175 ();
 sg13g2_decap_8 FILLER_53_1184 ();
 sg13g2_decap_8 FILLER_53_1191 ();
 sg13g2_decap_4 FILLER_53_1198 ();
 sg13g2_fill_2 FILLER_53_1202 ();
 sg13g2_fill_2 FILLER_53_1234 ();
 sg13g2_fill_2 FILLER_53_1296 ();
 sg13g2_decap_4 FILLER_53_1324 ();
 sg13g2_fill_2 FILLER_53_1328 ();
 sg13g2_decap_8 FILLER_53_1361 ();
 sg13g2_decap_4 FILLER_53_1368 ();
 sg13g2_fill_1 FILLER_53_1372 ();
 sg13g2_decap_8 FILLER_53_1413 ();
 sg13g2_decap_4 FILLER_53_1429 ();
 sg13g2_fill_1 FILLER_53_1433 ();
 sg13g2_decap_4 FILLER_53_1442 ();
 sg13g2_fill_2 FILLER_53_1446 ();
 sg13g2_decap_8 FILLER_53_1451 ();
 sg13g2_fill_1 FILLER_53_1492 ();
 sg13g2_fill_2 FILLER_53_1497 ();
 sg13g2_fill_1 FILLER_53_1499 ();
 sg13g2_fill_1 FILLER_53_1593 ();
 sg13g2_decap_8 FILLER_53_1611 ();
 sg13g2_decap_8 FILLER_53_1630 ();
 sg13g2_decap_4 FILLER_53_1637 ();
 sg13g2_fill_1 FILLER_53_1641 ();
 sg13g2_fill_1 FILLER_53_1658 ();
 sg13g2_fill_1 FILLER_53_1696 ();
 sg13g2_decap_8 FILLER_53_1702 ();
 sg13g2_decap_8 FILLER_53_1709 ();
 sg13g2_fill_1 FILLER_53_1730 ();
 sg13g2_decap_8 FILLER_53_1735 ();
 sg13g2_decap_8 FILLER_53_1742 ();
 sg13g2_decap_4 FILLER_53_1749 ();
 sg13g2_fill_2 FILLER_53_1753 ();
 sg13g2_decap_8 FILLER_53_1760 ();
 sg13g2_decap_8 FILLER_53_1767 ();
 sg13g2_decap_8 FILLER_53_1774 ();
 sg13g2_decap_4 FILLER_53_1781 ();
 sg13g2_fill_1 FILLER_53_1785 ();
 sg13g2_decap_8 FILLER_53_1794 ();
 sg13g2_fill_1 FILLER_53_1801 ();
 sg13g2_decap_4 FILLER_53_1872 ();
 sg13g2_fill_2 FILLER_53_1876 ();
 sg13g2_fill_1 FILLER_53_1887 ();
 sg13g2_decap_8 FILLER_53_1897 ();
 sg13g2_decap_8 FILLER_53_1904 ();
 sg13g2_decap_8 FILLER_53_1911 ();
 sg13g2_decap_8 FILLER_53_1918 ();
 sg13g2_fill_2 FILLER_53_1925 ();
 sg13g2_fill_2 FILLER_53_1932 ();
 sg13g2_fill_1 FILLER_53_1949 ();
 sg13g2_decap_8 FILLER_53_1955 ();
 sg13g2_decap_8 FILLER_53_1962 ();
 sg13g2_decap_8 FILLER_53_1969 ();
 sg13g2_decap_8 FILLER_53_1976 ();
 sg13g2_decap_8 FILLER_53_1983 ();
 sg13g2_decap_8 FILLER_53_1990 ();
 sg13g2_fill_2 FILLER_53_1997 ();
 sg13g2_decap_8 FILLER_53_2012 ();
 sg13g2_fill_2 FILLER_53_2019 ();
 sg13g2_fill_1 FILLER_53_2021 ();
 sg13g2_fill_1 FILLER_53_2037 ();
 sg13g2_decap_4 FILLER_53_2042 ();
 sg13g2_fill_2 FILLER_53_2046 ();
 sg13g2_fill_1 FILLER_53_2052 ();
 sg13g2_fill_2 FILLER_53_2083 ();
 sg13g2_decap_4 FILLER_53_2133 ();
 sg13g2_fill_2 FILLER_53_2137 ();
 sg13g2_decap_8 FILLER_53_2143 ();
 sg13g2_decap_8 FILLER_53_2150 ();
 sg13g2_fill_2 FILLER_53_2157 ();
 sg13g2_fill_1 FILLER_53_2159 ();
 sg13g2_fill_2 FILLER_53_2169 ();
 sg13g2_fill_1 FILLER_53_2171 ();
 sg13g2_fill_2 FILLER_53_2198 ();
 sg13g2_decap_4 FILLER_53_2230 ();
 sg13g2_fill_2 FILLER_53_2234 ();
 sg13g2_fill_1 FILLER_53_2242 ();
 sg13g2_fill_1 FILLER_53_2255 ();
 sg13g2_fill_2 FILLER_53_2287 ();
 sg13g2_fill_1 FILLER_53_2289 ();
 sg13g2_decap_8 FILLER_53_2333 ();
 sg13g2_decap_8 FILLER_53_2346 ();
 sg13g2_fill_2 FILLER_53_2353 ();
 sg13g2_fill_1 FILLER_53_2355 ();
 sg13g2_decap_8 FILLER_53_2360 ();
 sg13g2_decap_8 FILLER_53_2367 ();
 sg13g2_fill_1 FILLER_53_2374 ();
 sg13g2_decap_8 FILLER_53_2405 ();
 sg13g2_decap_8 FILLER_53_2412 ();
 sg13g2_decap_8 FILLER_53_2419 ();
 sg13g2_fill_2 FILLER_53_2426 ();
 sg13g2_fill_1 FILLER_53_2468 ();
 sg13g2_decap_4 FILLER_53_2490 ();
 sg13g2_fill_2 FILLER_53_2494 ();
 sg13g2_fill_2 FILLER_53_2551 ();
 sg13g2_fill_1 FILLER_53_2553 ();
 sg13g2_decap_8 FILLER_53_2559 ();
 sg13g2_decap_4 FILLER_53_2566 ();
 sg13g2_fill_2 FILLER_53_2580 ();
 sg13g2_fill_1 FILLER_53_2629 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_17 ();
 sg13g2_fill_2 FILLER_54_24 ();
 sg13g2_fill_1 FILLER_54_26 ();
 sg13g2_fill_1 FILLER_54_30 ();
 sg13g2_fill_1 FILLER_54_35 ();
 sg13g2_fill_1 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_47 ();
 sg13g2_fill_1 FILLER_54_53 ();
 sg13g2_decap_4 FILLER_54_64 ();
 sg13g2_decap_8 FILLER_54_75 ();
 sg13g2_decap_8 FILLER_54_82 ();
 sg13g2_decap_8 FILLER_54_89 ();
 sg13g2_decap_8 FILLER_54_96 ();
 sg13g2_decap_4 FILLER_54_103 ();
 sg13g2_fill_1 FILLER_54_107 ();
 sg13g2_decap_4 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_fill_2 FILLER_54_128 ();
 sg13g2_fill_2 FILLER_54_139 ();
 sg13g2_fill_2 FILLER_54_146 ();
 sg13g2_fill_1 FILLER_54_152 ();
 sg13g2_fill_1 FILLER_54_156 ();
 sg13g2_fill_1 FILLER_54_162 ();
 sg13g2_fill_1 FILLER_54_172 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_fill_2 FILLER_54_184 ();
 sg13g2_fill_1 FILLER_54_191 ();
 sg13g2_decap_4 FILLER_54_197 ();
 sg13g2_fill_2 FILLER_54_201 ();
 sg13g2_fill_1 FILLER_54_207 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_decap_4 FILLER_54_220 ();
 sg13g2_decap_8 FILLER_54_280 ();
 sg13g2_decap_8 FILLER_54_287 ();
 sg13g2_decap_8 FILLER_54_294 ();
 sg13g2_decap_4 FILLER_54_301 ();
 sg13g2_fill_1 FILLER_54_323 ();
 sg13g2_fill_2 FILLER_54_333 ();
 sg13g2_fill_2 FILLER_54_363 ();
 sg13g2_fill_1 FILLER_54_365 ();
 sg13g2_fill_1 FILLER_54_371 ();
 sg13g2_fill_2 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_54_379 ();
 sg13g2_decap_4 FILLER_54_387 ();
 sg13g2_fill_2 FILLER_54_429 ();
 sg13g2_fill_1 FILLER_54_431 ();
 sg13g2_fill_2 FILLER_54_441 ();
 sg13g2_fill_2 FILLER_54_456 ();
 sg13g2_fill_2 FILLER_54_476 ();
 sg13g2_fill_1 FILLER_54_486 ();
 sg13g2_decap_8 FILLER_54_543 ();
 sg13g2_decap_8 FILLER_54_557 ();
 sg13g2_decap_8 FILLER_54_564 ();
 sg13g2_fill_2 FILLER_54_571 ();
 sg13g2_fill_1 FILLER_54_573 ();
 sg13g2_fill_2 FILLER_54_652 ();
 sg13g2_fill_1 FILLER_54_654 ();
 sg13g2_decap_4 FILLER_54_673 ();
 sg13g2_decap_4 FILLER_54_686 ();
 sg13g2_fill_2 FILLER_54_690 ();
 sg13g2_decap_8 FILLER_54_702 ();
 sg13g2_decap_4 FILLER_54_709 ();
 sg13g2_decap_8 FILLER_54_724 ();
 sg13g2_decap_8 FILLER_54_735 ();
 sg13g2_decap_8 FILLER_54_742 ();
 sg13g2_fill_2 FILLER_54_749 ();
 sg13g2_fill_2 FILLER_54_760 ();
 sg13g2_fill_1 FILLER_54_762 ();
 sg13g2_decap_8 FILLER_54_819 ();
 sg13g2_fill_1 FILLER_54_826 ();
 sg13g2_fill_2 FILLER_54_832 ();
 sg13g2_fill_1 FILLER_54_834 ();
 sg13g2_decap_4 FILLER_54_849 ();
 sg13g2_fill_1 FILLER_54_853 ();
 sg13g2_fill_2 FILLER_54_858 ();
 sg13g2_decap_4 FILLER_54_865 ();
 sg13g2_decap_8 FILLER_54_873 ();
 sg13g2_fill_2 FILLER_54_880 ();
 sg13g2_fill_2 FILLER_54_887 ();
 sg13g2_decap_8 FILLER_54_897 ();
 sg13g2_decap_8 FILLER_54_904 ();
 sg13g2_decap_8 FILLER_54_911 ();
 sg13g2_decap_8 FILLER_54_918 ();
 sg13g2_fill_2 FILLER_54_925 ();
 sg13g2_fill_1 FILLER_54_927 ();
 sg13g2_fill_1 FILLER_54_937 ();
 sg13g2_fill_1 FILLER_54_948 ();
 sg13g2_decap_8 FILLER_54_953 ();
 sg13g2_fill_1 FILLER_54_960 ();
 sg13g2_decap_4 FILLER_54_964 ();
 sg13g2_fill_2 FILLER_54_968 ();
 sg13g2_fill_1 FILLER_54_979 ();
 sg13g2_decap_8 FILLER_54_984 ();
 sg13g2_decap_8 FILLER_54_991 ();
 sg13g2_fill_1 FILLER_54_998 ();
 sg13g2_fill_2 FILLER_54_1011 ();
 sg13g2_fill_1 FILLER_54_1013 ();
 sg13g2_fill_2 FILLER_54_1040 ();
 sg13g2_fill_2 FILLER_54_1076 ();
 sg13g2_fill_1 FILLER_54_1078 ();
 sg13g2_fill_2 FILLER_54_1083 ();
 sg13g2_fill_1 FILLER_54_1090 ();
 sg13g2_decap_8 FILLER_54_1095 ();
 sg13g2_fill_2 FILLER_54_1128 ();
 sg13g2_fill_1 FILLER_54_1130 ();
 sg13g2_decap_8 FILLER_54_1137 ();
 sg13g2_fill_2 FILLER_54_1144 ();
 sg13g2_fill_1 FILLER_54_1146 ();
 sg13g2_decap_8 FILLER_54_1185 ();
 sg13g2_decap_8 FILLER_54_1192 ();
 sg13g2_decap_8 FILLER_54_1199 ();
 sg13g2_decap_4 FILLER_54_1206 ();
 sg13g2_fill_1 FILLER_54_1210 ();
 sg13g2_decap_8 FILLER_54_1214 ();
 sg13g2_fill_2 FILLER_54_1221 ();
 sg13g2_fill_1 FILLER_54_1223 ();
 sg13g2_fill_1 FILLER_54_1229 ();
 sg13g2_fill_2 FILLER_54_1234 ();
 sg13g2_fill_1 FILLER_54_1236 ();
 sg13g2_fill_1 FILLER_54_1263 ();
 sg13g2_decap_8 FILLER_54_1286 ();
 sg13g2_decap_8 FILLER_54_1293 ();
 sg13g2_fill_1 FILLER_54_1300 ();
 sg13g2_decap_8 FILLER_54_1332 ();
 sg13g2_decap_8 FILLER_54_1339 ();
 sg13g2_fill_2 FILLER_54_1346 ();
 sg13g2_fill_1 FILLER_54_1348 ();
 sg13g2_decap_8 FILLER_54_1375 ();
 sg13g2_decap_8 FILLER_54_1382 ();
 sg13g2_decap_8 FILLER_54_1389 ();
 sg13g2_decap_8 FILLER_54_1396 ();
 sg13g2_fill_2 FILLER_54_1403 ();
 sg13g2_fill_1 FILLER_54_1405 ();
 sg13g2_decap_4 FILLER_54_1416 ();
 sg13g2_fill_2 FILLER_54_1420 ();
 sg13g2_fill_1 FILLER_54_1453 ();
 sg13g2_decap_8 FILLER_54_1458 ();
 sg13g2_decap_8 FILLER_54_1465 ();
 sg13g2_fill_2 FILLER_54_1472 ();
 sg13g2_decap_8 FILLER_54_1485 ();
 sg13g2_decap_4 FILLER_54_1492 ();
 sg13g2_fill_2 FILLER_54_1496 ();
 sg13g2_fill_1 FILLER_54_1502 ();
 sg13g2_fill_2 FILLER_54_1508 ();
 sg13g2_fill_2 FILLER_54_1618 ();
 sg13g2_fill_1 FILLER_54_1620 ();
 sg13g2_decap_4 FILLER_54_1628 ();
 sg13g2_fill_2 FILLER_54_1640 ();
 sg13g2_fill_2 FILLER_54_1653 ();
 sg13g2_fill_1 FILLER_54_1688 ();
 sg13g2_decap_8 FILLER_54_1710 ();
 sg13g2_fill_1 FILLER_54_1717 ();
 sg13g2_decap_4 FILLER_54_1748 ();
 sg13g2_fill_2 FILLER_54_1752 ();
 sg13g2_decap_8 FILLER_54_1758 ();
 sg13g2_decap_4 FILLER_54_1782 ();
 sg13g2_fill_1 FILLER_54_1792 ();
 sg13g2_fill_1 FILLER_54_1819 ();
 sg13g2_decap_8 FILLER_54_1875 ();
 sg13g2_fill_2 FILLER_54_1885 ();
 sg13g2_fill_1 FILLER_54_1887 ();
 sg13g2_decap_8 FILLER_54_1896 ();
 sg13g2_decap_8 FILLER_54_1903 ();
 sg13g2_decap_8 FILLER_54_1910 ();
 sg13g2_decap_8 FILLER_54_1917 ();
 sg13g2_decap_8 FILLER_54_1924 ();
 sg13g2_decap_8 FILLER_54_1931 ();
 sg13g2_decap_8 FILLER_54_1938 ();
 sg13g2_decap_4 FILLER_54_1945 ();
 sg13g2_decap_8 FILLER_54_1966 ();
 sg13g2_decap_8 FILLER_54_1973 ();
 sg13g2_decap_8 FILLER_54_1985 ();
 sg13g2_decap_4 FILLER_54_1992 ();
 sg13g2_decap_8 FILLER_54_2005 ();
 sg13g2_decap_8 FILLER_54_2012 ();
 sg13g2_fill_1 FILLER_54_2019 ();
 sg13g2_decap_8 FILLER_54_2024 ();
 sg13g2_decap_8 FILLER_54_2031 ();
 sg13g2_decap_8 FILLER_54_2038 ();
 sg13g2_decap_4 FILLER_54_2045 ();
 sg13g2_fill_2 FILLER_54_2049 ();
 sg13g2_fill_2 FILLER_54_2056 ();
 sg13g2_fill_1 FILLER_54_2058 ();
 sg13g2_fill_1 FILLER_54_2063 ();
 sg13g2_fill_1 FILLER_54_2093 ();
 sg13g2_fill_1 FILLER_54_2126 ();
 sg13g2_decap_8 FILLER_54_2132 ();
 sg13g2_fill_2 FILLER_54_2139 ();
 sg13g2_fill_1 FILLER_54_2172 ();
 sg13g2_fill_1 FILLER_54_2178 ();
 sg13g2_fill_1 FILLER_54_2205 ();
 sg13g2_fill_2 FILLER_54_2244 ();
 sg13g2_fill_2 FILLER_54_2255 ();
 sg13g2_fill_2 FILLER_54_2265 ();
 sg13g2_fill_1 FILLER_54_2267 ();
 sg13g2_fill_1 FILLER_54_2278 ();
 sg13g2_fill_2 FILLER_54_2306 ();
 sg13g2_decap_4 FILLER_54_2312 ();
 sg13g2_fill_1 FILLER_54_2316 ();
 sg13g2_decap_8 FILLER_54_2347 ();
 sg13g2_decap_8 FILLER_54_2354 ();
 sg13g2_decap_8 FILLER_54_2361 ();
 sg13g2_decap_4 FILLER_54_2368 ();
 sg13g2_fill_2 FILLER_54_2372 ();
 sg13g2_fill_1 FILLER_54_2378 ();
 sg13g2_fill_2 FILLER_54_2383 ();
 sg13g2_fill_2 FILLER_54_2389 ();
 sg13g2_decap_8 FILLER_54_2395 ();
 sg13g2_decap_8 FILLER_54_2402 ();
 sg13g2_decap_8 FILLER_54_2409 ();
 sg13g2_decap_8 FILLER_54_2416 ();
 sg13g2_decap_8 FILLER_54_2423 ();
 sg13g2_decap_8 FILLER_54_2430 ();
 sg13g2_fill_1 FILLER_54_2475 ();
 sg13g2_fill_2 FILLER_54_2482 ();
 sg13g2_fill_1 FILLER_54_2484 ();
 sg13g2_fill_2 FILLER_54_2505 ();
 sg13g2_fill_1 FILLER_54_2507 ();
 sg13g2_fill_2 FILLER_54_2534 ();
 sg13g2_fill_1 FILLER_54_2536 ();
 sg13g2_fill_1 FILLER_54_2540 ();
 sg13g2_decap_4 FILLER_54_2550 ();
 sg13g2_decap_8 FILLER_54_2558 ();
 sg13g2_decap_8 FILLER_54_2565 ();
 sg13g2_decap_8 FILLER_54_2572 ();
 sg13g2_decap_8 FILLER_54_2579 ();
 sg13g2_decap_4 FILLER_54_2586 ();
 sg13g2_fill_1 FILLER_54_2590 ();
 sg13g2_fill_2 FILLER_54_2617 ();
 sg13g2_fill_2 FILLER_54_2632 ();
 sg13g2_fill_1 FILLER_54_2634 ();
 sg13g2_fill_2 FILLER_54_2648 ();
 sg13g2_fill_1 FILLER_54_2650 ();
 sg13g2_decap_8 FILLER_54_2655 ();
 sg13g2_decap_8 FILLER_54_2662 ();
 sg13g2_fill_1 FILLER_54_2669 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_4 FILLER_55_24 ();
 sg13g2_fill_2 FILLER_55_28 ();
 sg13g2_fill_1 FILLER_55_51 ();
 sg13g2_fill_2 FILLER_55_72 ();
 sg13g2_decap_8 FILLER_55_92 ();
 sg13g2_decap_8 FILLER_55_99 ();
 sg13g2_decap_8 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_113 ();
 sg13g2_fill_1 FILLER_55_115 ();
 sg13g2_decap_8 FILLER_55_120 ();
 sg13g2_decap_4 FILLER_55_127 ();
 sg13g2_fill_1 FILLER_55_131 ();
 sg13g2_fill_2 FILLER_55_141 ();
 sg13g2_fill_1 FILLER_55_143 ();
 sg13g2_fill_2 FILLER_55_148 ();
 sg13g2_fill_2 FILLER_55_160 ();
 sg13g2_decap_4 FILLER_55_166 ();
 sg13g2_fill_2 FILLER_55_170 ();
 sg13g2_decap_4 FILLER_55_176 ();
 sg13g2_fill_2 FILLER_55_180 ();
 sg13g2_decap_4 FILLER_55_190 ();
 sg13g2_fill_2 FILLER_55_194 ();
 sg13g2_decap_8 FILLER_55_200 ();
 sg13g2_fill_1 FILLER_55_207 ();
 sg13g2_decap_8 FILLER_55_234 ();
 sg13g2_fill_2 FILLER_55_277 ();
 sg13g2_fill_1 FILLER_55_279 ();
 sg13g2_decap_8 FILLER_55_288 ();
 sg13g2_decap_8 FILLER_55_295 ();
 sg13g2_decap_8 FILLER_55_302 ();
 sg13g2_fill_2 FILLER_55_309 ();
 sg13g2_fill_1 FILLER_55_311 ();
 sg13g2_fill_2 FILLER_55_315 ();
 sg13g2_fill_1 FILLER_55_317 ();
 sg13g2_decap_4 FILLER_55_323 ();
 sg13g2_fill_1 FILLER_55_327 ();
 sg13g2_decap_8 FILLER_55_333 ();
 sg13g2_fill_2 FILLER_55_340 ();
 sg13g2_fill_1 FILLER_55_342 ();
 sg13g2_decap_8 FILLER_55_353 ();
 sg13g2_decap_8 FILLER_55_360 ();
 sg13g2_fill_2 FILLER_55_367 ();
 sg13g2_fill_2 FILLER_55_400 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_fill_2 FILLER_55_413 ();
 sg13g2_fill_1 FILLER_55_415 ();
 sg13g2_decap_8 FILLER_55_421 ();
 sg13g2_decap_4 FILLER_55_428 ();
 sg13g2_fill_1 FILLER_55_432 ();
 sg13g2_fill_2 FILLER_55_443 ();
 sg13g2_fill_1 FILLER_55_445 ();
 sg13g2_fill_2 FILLER_55_460 ();
 sg13g2_fill_2 FILLER_55_477 ();
 sg13g2_fill_1 FILLER_55_484 ();
 sg13g2_decap_4 FILLER_55_513 ();
 sg13g2_fill_2 FILLER_55_517 ();
 sg13g2_fill_2 FILLER_55_522 ();
 sg13g2_fill_1 FILLER_55_524 ();
 sg13g2_fill_1 FILLER_55_533 ();
 sg13g2_decap_8 FILLER_55_542 ();
 sg13g2_decap_4 FILLER_55_549 ();
 sg13g2_fill_1 FILLER_55_553 ();
 sg13g2_decap_4 FILLER_55_559 ();
 sg13g2_fill_2 FILLER_55_563 ();
 sg13g2_fill_1 FILLER_55_584 ();
 sg13g2_fill_1 FILLER_55_589 ();
 sg13g2_fill_1 FILLER_55_613 ();
 sg13g2_fill_2 FILLER_55_635 ();
 sg13g2_decap_8 FILLER_55_684 ();
 sg13g2_decap_4 FILLER_55_710 ();
 sg13g2_fill_1 FILLER_55_714 ();
 sg13g2_decap_8 FILLER_55_723 ();
 sg13g2_decap_8 FILLER_55_730 ();
 sg13g2_decap_8 FILLER_55_767 ();
 sg13g2_fill_1 FILLER_55_774 ();
 sg13g2_fill_1 FILLER_55_793 ();
 sg13g2_fill_2 FILLER_55_799 ();
 sg13g2_fill_1 FILLER_55_801 ();
 sg13g2_fill_2 FILLER_55_811 ();
 sg13g2_fill_1 FILLER_55_839 ();
 sg13g2_fill_1 FILLER_55_845 ();
 sg13g2_decap_8 FILLER_55_881 ();
 sg13g2_fill_2 FILLER_55_888 ();
 sg13g2_fill_2 FILLER_55_899 ();
 sg13g2_fill_1 FILLER_55_901 ();
 sg13g2_decap_8 FILLER_55_907 ();
 sg13g2_fill_2 FILLER_55_914 ();
 sg13g2_decap_4 FILLER_55_921 ();
 sg13g2_fill_1 FILLER_55_925 ();
 sg13g2_decap_8 FILLER_55_930 ();
 sg13g2_decap_8 FILLER_55_937 ();
 sg13g2_decap_4 FILLER_55_957 ();
 sg13g2_decap_4 FILLER_55_966 ();
 sg13g2_fill_1 FILLER_55_970 ();
 sg13g2_fill_1 FILLER_55_997 ();
 sg13g2_fill_2 FILLER_55_1016 ();
 sg13g2_fill_2 FILLER_55_1050 ();
 sg13g2_fill_1 FILLER_55_1057 ();
 sg13g2_fill_2 FILLER_55_1140 ();
 sg13g2_fill_1 FILLER_55_1146 ();
 sg13g2_fill_2 FILLER_55_1173 ();
 sg13g2_fill_1 FILLER_55_1175 ();
 sg13g2_decap_4 FILLER_55_1202 ();
 sg13g2_fill_2 FILLER_55_1206 ();
 sg13g2_fill_1 FILLER_55_1216 ();
 sg13g2_fill_2 FILLER_55_1242 ();
 sg13g2_fill_2 FILLER_55_1263 ();
 sg13g2_decap_8 FILLER_55_1292 ();
 sg13g2_fill_1 FILLER_55_1299 ();
 sg13g2_fill_1 FILLER_55_1311 ();
 sg13g2_decap_8 FILLER_55_1316 ();
 sg13g2_decap_8 FILLER_55_1323 ();
 sg13g2_decap_8 FILLER_55_1330 ();
 sg13g2_decap_8 FILLER_55_1337 ();
 sg13g2_decap_4 FILLER_55_1344 ();
 sg13g2_fill_2 FILLER_55_1348 ();
 sg13g2_decap_8 FILLER_55_1359 ();
 sg13g2_decap_8 FILLER_55_1366 ();
 sg13g2_decap_8 FILLER_55_1373 ();
 sg13g2_decap_8 FILLER_55_1380 ();
 sg13g2_decap_8 FILLER_55_1387 ();
 sg13g2_fill_2 FILLER_55_1415 ();
 sg13g2_decap_8 FILLER_55_1421 ();
 sg13g2_fill_2 FILLER_55_1428 ();
 sg13g2_fill_1 FILLER_55_1442 ();
 sg13g2_decap_8 FILLER_55_1475 ();
 sg13g2_decap_8 FILLER_55_1482 ();
 sg13g2_decap_4 FILLER_55_1489 ();
 sg13g2_fill_2 FILLER_55_1523 ();
 sg13g2_fill_2 FILLER_55_1539 ();
 sg13g2_decap_8 FILLER_55_1558 ();
 sg13g2_decap_4 FILLER_55_1565 ();
 sg13g2_fill_1 FILLER_55_1609 ();
 sg13g2_fill_2 FILLER_55_1615 ();
 sg13g2_fill_2 FILLER_55_1694 ();
 sg13g2_decap_8 FILLER_55_1710 ();
 sg13g2_fill_2 FILLER_55_1717 ();
 sg13g2_fill_1 FILLER_55_1719 ();
 sg13g2_fill_2 FILLER_55_1751 ();
 sg13g2_decap_8 FILLER_55_1784 ();
 sg13g2_decap_8 FILLER_55_1791 ();
 sg13g2_decap_4 FILLER_55_1798 ();
 sg13g2_fill_2 FILLER_55_1802 ();
 sg13g2_fill_2 FILLER_55_1838 ();
 sg13g2_fill_2 FILLER_55_1847 ();
 sg13g2_fill_1 FILLER_55_1859 ();
 sg13g2_fill_1 FILLER_55_1891 ();
 sg13g2_decap_8 FILLER_55_1924 ();
 sg13g2_decap_8 FILLER_55_1931 ();
 sg13g2_decap_8 FILLER_55_1938 ();
 sg13g2_fill_1 FILLER_55_1945 ();
 sg13g2_decap_8 FILLER_55_1950 ();
 sg13g2_decap_8 FILLER_55_1957 ();
 sg13g2_fill_1 FILLER_55_1964 ();
 sg13g2_fill_2 FILLER_55_1970 ();
 sg13g2_fill_1 FILLER_55_1979 ();
 sg13g2_decap_8 FILLER_55_2011 ();
 sg13g2_decap_8 FILLER_55_2018 ();
 sg13g2_decap_4 FILLER_55_2025 ();
 sg13g2_decap_4 FILLER_55_2045 ();
 sg13g2_fill_1 FILLER_55_2049 ();
 sg13g2_fill_2 FILLER_55_2099 ();
 sg13g2_fill_2 FILLER_55_2111 ();
 sg13g2_fill_1 FILLER_55_2117 ();
 sg13g2_fill_1 FILLER_55_2136 ();
 sg13g2_fill_2 FILLER_55_2169 ();
 sg13g2_fill_1 FILLER_55_2171 ();
 sg13g2_decap_8 FILLER_55_2176 ();
 sg13g2_decap_8 FILLER_55_2183 ();
 sg13g2_decap_8 FILLER_55_2190 ();
 sg13g2_fill_2 FILLER_55_2197 ();
 sg13g2_fill_1 FILLER_55_2199 ();
 sg13g2_decap_4 FILLER_55_2250 ();
 sg13g2_fill_1 FILLER_55_2254 ();
 sg13g2_fill_2 FILLER_55_2291 ();
 sg13g2_decap_8 FILLER_55_2319 ();
 sg13g2_fill_1 FILLER_55_2326 ();
 sg13g2_decap_8 FILLER_55_2331 ();
 sg13g2_decap_8 FILLER_55_2338 ();
 sg13g2_decap_8 FILLER_55_2345 ();
 sg13g2_fill_2 FILLER_55_2352 ();
 sg13g2_decap_4 FILLER_55_2384 ();
 sg13g2_decap_8 FILLER_55_2392 ();
 sg13g2_fill_2 FILLER_55_2399 ();
 sg13g2_decap_4 FILLER_55_2405 ();
 sg13g2_fill_1 FILLER_55_2409 ();
 sg13g2_decap_8 FILLER_55_2440 ();
 sg13g2_decap_8 FILLER_55_2447 ();
 sg13g2_fill_2 FILLER_55_2454 ();
 sg13g2_fill_1 FILLER_55_2456 ();
 sg13g2_decap_8 FILLER_55_2460 ();
 sg13g2_fill_1 FILLER_55_2471 ();
 sg13g2_fill_2 FILLER_55_2476 ();
 sg13g2_fill_1 FILLER_55_2483 ();
 sg13g2_fill_2 FILLER_55_2493 ();
 sg13g2_fill_1 FILLER_55_2495 ();
 sg13g2_fill_1 FILLER_55_2499 ();
 sg13g2_fill_1 FILLER_55_2530 ();
 sg13g2_fill_1 FILLER_55_2536 ();
 sg13g2_decap_8 FILLER_55_2576 ();
 sg13g2_decap_8 FILLER_55_2583 ();
 sg13g2_decap_4 FILLER_55_2590 ();
 sg13g2_fill_1 FILLER_55_2594 ();
 sg13g2_fill_2 FILLER_55_2599 ();
 sg13g2_decap_8 FILLER_55_2605 ();
 sg13g2_decap_8 FILLER_55_2612 ();
 sg13g2_decap_8 FILLER_55_2619 ();
 sg13g2_decap_4 FILLER_55_2631 ();
 sg13g2_fill_1 FILLER_55_2635 ();
 sg13g2_decap_4 FILLER_55_2666 ();
 sg13g2_fill_2 FILLER_56_0 ();
 sg13g2_fill_2 FILLER_56_28 ();
 sg13g2_fill_1 FILLER_56_30 ();
 sg13g2_fill_1 FILLER_56_35 ();
 sg13g2_fill_1 FILLER_56_55 ();
 sg13g2_fill_1 FILLER_56_60 ();
 sg13g2_fill_1 FILLER_56_65 ();
 sg13g2_decap_4 FILLER_56_76 ();
 sg13g2_fill_1 FILLER_56_80 ();
 sg13g2_decap_4 FILLER_56_86 ();
 sg13g2_decap_8 FILLER_56_94 ();
 sg13g2_decap_8 FILLER_56_101 ();
 sg13g2_fill_2 FILLER_56_108 ();
 sg13g2_fill_1 FILLER_56_110 ();
 sg13g2_decap_4 FILLER_56_129 ();
 sg13g2_decap_4 FILLER_56_138 ();
 sg13g2_decap_8 FILLER_56_151 ();
 sg13g2_decap_8 FILLER_56_158 ();
 sg13g2_fill_2 FILLER_56_165 ();
 sg13g2_decap_8 FILLER_56_177 ();
 sg13g2_decap_8 FILLER_56_184 ();
 sg13g2_decap_8 FILLER_56_191 ();
 sg13g2_decap_4 FILLER_56_198 ();
 sg13g2_fill_2 FILLER_56_202 ();
 sg13g2_fill_2 FILLER_56_230 ();
 sg13g2_decap_8 FILLER_56_236 ();
 sg13g2_decap_8 FILLER_56_243 ();
 sg13g2_decap_8 FILLER_56_250 ();
 sg13g2_decap_8 FILLER_56_257 ();
 sg13g2_decap_4 FILLER_56_264 ();
 sg13g2_fill_2 FILLER_56_268 ();
 sg13g2_decap_8 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_319 ();
 sg13g2_fill_1 FILLER_56_321 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_335 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_347 ();
 sg13g2_decap_4 FILLER_56_354 ();
 sg13g2_fill_1 FILLER_56_358 ();
 sg13g2_fill_1 FILLER_56_391 ();
 sg13g2_fill_1 FILLER_56_397 ();
 sg13g2_fill_2 FILLER_56_408 ();
 sg13g2_decap_8 FILLER_56_416 ();
 sg13g2_decap_8 FILLER_56_423 ();
 sg13g2_fill_2 FILLER_56_430 ();
 sg13g2_fill_1 FILLER_56_432 ();
 sg13g2_fill_1 FILLER_56_438 ();
 sg13g2_fill_2 FILLER_56_442 ();
 sg13g2_decap_8 FILLER_56_447 ();
 sg13g2_decap_8 FILLER_56_454 ();
 sg13g2_fill_2 FILLER_56_461 ();
 sg13g2_fill_2 FILLER_56_468 ();
 sg13g2_fill_1 FILLER_56_470 ();
 sg13g2_fill_2 FILLER_56_486 ();
 sg13g2_fill_1 FILLER_56_493 ();
 sg13g2_fill_2 FILLER_56_511 ();
 sg13g2_fill_1 FILLER_56_513 ();
 sg13g2_decap_8 FILLER_56_540 ();
 sg13g2_decap_8 FILLER_56_547 ();
 sg13g2_decap_8 FILLER_56_558 ();
 sg13g2_decap_8 FILLER_56_565 ();
 sg13g2_decap_4 FILLER_56_572 ();
 sg13g2_fill_1 FILLER_56_605 ();
 sg13g2_decap_4 FILLER_56_660 ();
 sg13g2_fill_2 FILLER_56_664 ();
 sg13g2_fill_1 FILLER_56_671 ();
 sg13g2_fill_1 FILLER_56_680 ();
 sg13g2_fill_1 FILLER_56_697 ();
 sg13g2_fill_1 FILLER_56_712 ();
 sg13g2_decap_8 FILLER_56_724 ();
 sg13g2_decap_8 FILLER_56_731 ();
 sg13g2_decap_8 FILLER_56_738 ();
 sg13g2_decap_8 FILLER_56_745 ();
 sg13g2_decap_8 FILLER_56_752 ();
 sg13g2_decap_8 FILLER_56_759 ();
 sg13g2_decap_8 FILLER_56_766 ();
 sg13g2_fill_2 FILLER_56_773 ();
 sg13g2_decap_4 FILLER_56_810 ();
 sg13g2_fill_1 FILLER_56_814 ();
 sg13g2_fill_2 FILLER_56_819 ();
 sg13g2_fill_1 FILLER_56_821 ();
 sg13g2_decap_8 FILLER_56_831 ();
 sg13g2_decap_8 FILLER_56_838 ();
 sg13g2_decap_8 FILLER_56_845 ();
 sg13g2_fill_2 FILLER_56_852 ();
 sg13g2_decap_4 FILLER_56_911 ();
 sg13g2_fill_1 FILLER_56_945 ();
 sg13g2_fill_2 FILLER_56_950 ();
 sg13g2_fill_1 FILLER_56_952 ();
 sg13g2_fill_2 FILLER_56_957 ();
 sg13g2_decap_8 FILLER_56_977 ();
 sg13g2_fill_2 FILLER_56_984 ();
 sg13g2_fill_1 FILLER_56_986 ();
 sg13g2_fill_2 FILLER_56_990 ();
 sg13g2_fill_2 FILLER_56_1018 ();
 sg13g2_fill_1 FILLER_56_1020 ();
 sg13g2_fill_2 FILLER_56_1031 ();
 sg13g2_decap_8 FILLER_56_1074 ();
 sg13g2_fill_2 FILLER_56_1081 ();
 sg13g2_decap_8 FILLER_56_1137 ();
 sg13g2_fill_1 FILLER_56_1144 ();
 sg13g2_decap_4 FILLER_56_1159 ();
 sg13g2_fill_1 FILLER_56_1163 ();
 sg13g2_fill_2 FILLER_56_1168 ();
 sg13g2_fill_1 FILLER_56_1170 ();
 sg13g2_fill_2 FILLER_56_1176 ();
 sg13g2_fill_1 FILLER_56_1178 ();
 sg13g2_fill_2 FILLER_56_1184 ();
 sg13g2_fill_2 FILLER_56_1212 ();
 sg13g2_fill_1 FILLER_56_1214 ();
 sg13g2_fill_2 FILLER_56_1266 ();
 sg13g2_decap_8 FILLER_56_1294 ();
 sg13g2_decap_8 FILLER_56_1301 ();
 sg13g2_decap_8 FILLER_56_1308 ();
 sg13g2_decap_8 FILLER_56_1315 ();
 sg13g2_decap_8 FILLER_56_1322 ();
 sg13g2_fill_2 FILLER_56_1329 ();
 sg13g2_decap_8 FILLER_56_1340 ();
 sg13g2_decap_8 FILLER_56_1347 ();
 sg13g2_decap_4 FILLER_56_1354 ();
 sg13g2_fill_1 FILLER_56_1393 ();
 sg13g2_decap_8 FILLER_56_1467 ();
 sg13g2_decap_8 FILLER_56_1474 ();
 sg13g2_decap_8 FILLER_56_1481 ();
 sg13g2_fill_2 FILLER_56_1488 ();
 sg13g2_decap_8 FILLER_56_1495 ();
 sg13g2_decap_8 FILLER_56_1502 ();
 sg13g2_fill_2 FILLER_56_1509 ();
 sg13g2_decap_8 FILLER_56_1514 ();
 sg13g2_fill_2 FILLER_56_1521 ();
 sg13g2_fill_1 FILLER_56_1523 ();
 sg13g2_fill_2 FILLER_56_1528 ();
 sg13g2_fill_1 FILLER_56_1543 ();
 sg13g2_fill_2 FILLER_56_1593 ();
 sg13g2_fill_2 FILLER_56_1599 ();
 sg13g2_fill_2 FILLER_56_1614 ();
 sg13g2_fill_1 FILLER_56_1616 ();
 sg13g2_decap_4 FILLER_56_1621 ();
 sg13g2_fill_2 FILLER_56_1634 ();
 sg13g2_fill_1 FILLER_56_1636 ();
 sg13g2_decap_4 FILLER_56_1667 ();
 sg13g2_fill_1 FILLER_56_1671 ();
 sg13g2_fill_2 FILLER_56_1677 ();
 sg13g2_fill_1 FILLER_56_1679 ();
 sg13g2_fill_2 FILLER_56_1744 ();
 sg13g2_fill_1 FILLER_56_1746 ();
 sg13g2_decap_8 FILLER_56_1752 ();
 sg13g2_decap_8 FILLER_56_1759 ();
 sg13g2_decap_8 FILLER_56_1766 ();
 sg13g2_decap_4 FILLER_56_1777 ();
 sg13g2_fill_2 FILLER_56_1781 ();
 sg13g2_decap_4 FILLER_56_1788 ();
 sg13g2_fill_1 FILLER_56_1792 ();
 sg13g2_decap_8 FILLER_56_1801 ();
 sg13g2_fill_2 FILLER_56_1844 ();
 sg13g2_fill_2 FILLER_56_1860 ();
 sg13g2_fill_1 FILLER_56_1881 ();
 sg13g2_decap_4 FILLER_56_1898 ();
 sg13g2_fill_2 FILLER_56_1902 ();
 sg13g2_decap_4 FILLER_56_1913 ();
 sg13g2_fill_1 FILLER_56_1925 ();
 sg13g2_decap_4 FILLER_56_1965 ();
 sg13g2_fill_1 FILLER_56_1969 ();
 sg13g2_fill_1 FILLER_56_2008 ();
 sg13g2_decap_8 FILLER_56_2088 ();
 sg13g2_decap_4 FILLER_56_2095 ();
 sg13g2_fill_2 FILLER_56_2099 ();
 sg13g2_decap_8 FILLER_56_2110 ();
 sg13g2_decap_8 FILLER_56_2117 ();
 sg13g2_decap_8 FILLER_56_2129 ();
 sg13g2_decap_8 FILLER_56_2136 ();
 sg13g2_decap_4 FILLER_56_2143 ();
 sg13g2_fill_1 FILLER_56_2147 ();
 sg13g2_fill_2 FILLER_56_2158 ();
 sg13g2_fill_2 FILLER_56_2166 ();
 sg13g2_fill_1 FILLER_56_2172 ();
 sg13g2_decap_8 FILLER_56_2204 ();
 sg13g2_fill_2 FILLER_56_2211 ();
 sg13g2_decap_8 FILLER_56_2244 ();
 sg13g2_decap_8 FILLER_56_2251 ();
 sg13g2_decap_4 FILLER_56_2258 ();
 sg13g2_fill_1 FILLER_56_2262 ();
 sg13g2_fill_1 FILLER_56_2286 ();
 sg13g2_fill_2 FILLER_56_2293 ();
 sg13g2_fill_1 FILLER_56_2295 ();
 sg13g2_decap_8 FILLER_56_2313 ();
 sg13g2_fill_1 FILLER_56_2320 ();
 sg13g2_decap_8 FILLER_56_2355 ();
 sg13g2_fill_2 FILLER_56_2362 ();
 sg13g2_fill_1 FILLER_56_2364 ();
 sg13g2_fill_2 FILLER_56_2369 ();
 sg13g2_fill_1 FILLER_56_2371 ();
 sg13g2_fill_2 FILLER_56_2449 ();
 sg13g2_fill_1 FILLER_56_2451 ();
 sg13g2_fill_1 FILLER_56_2456 ();
 sg13g2_fill_2 FILLER_56_2460 ();
 sg13g2_fill_2 FILLER_56_2505 ();
 sg13g2_fill_2 FILLER_56_2511 ();
 sg13g2_fill_1 FILLER_56_2513 ();
 sg13g2_fill_1 FILLER_56_2518 ();
 sg13g2_decap_8 FILLER_56_2553 ();
 sg13g2_fill_2 FILLER_56_2560 ();
 sg13g2_decap_4 FILLER_56_2588 ();
 sg13g2_fill_1 FILLER_56_2592 ();
 sg13g2_fill_1 FILLER_56_2597 ();
 sg13g2_decap_8 FILLER_56_2628 ();
 sg13g2_decap_4 FILLER_56_2635 ();
 sg13g2_fill_1 FILLER_56_2639 ();
 sg13g2_decap_8 FILLER_56_2648 ();
 sg13g2_fill_2 FILLER_56_2655 ();
 sg13g2_fill_1 FILLER_56_2657 ();
 sg13g2_decap_8 FILLER_56_2662 ();
 sg13g2_fill_1 FILLER_56_2669 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_fill_2 FILLER_57_7 ();
 sg13g2_fill_1 FILLER_57_9 ();
 sg13g2_decap_4 FILLER_57_20 ();
 sg13g2_fill_1 FILLER_57_24 ();
 sg13g2_decap_4 FILLER_57_32 ();
 sg13g2_fill_1 FILLER_57_36 ();
 sg13g2_fill_2 FILLER_57_82 ();
 sg13g2_fill_1 FILLER_57_84 ();
 sg13g2_fill_2 FILLER_57_100 ();
 sg13g2_fill_2 FILLER_57_141 ();
 sg13g2_decap_4 FILLER_57_153 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_fill_1 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_187 ();
 sg13g2_decap_4 FILLER_57_194 ();
 sg13g2_fill_2 FILLER_57_198 ();
 sg13g2_fill_2 FILLER_57_210 ();
 sg13g2_fill_1 FILLER_57_212 ();
 sg13g2_decap_4 FILLER_57_227 ();
 sg13g2_decap_8 FILLER_57_241 ();
 sg13g2_decap_8 FILLER_57_248 ();
 sg13g2_fill_2 FILLER_57_255 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_4 FILLER_57_287 ();
 sg13g2_fill_2 FILLER_57_291 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_2 FILLER_57_349 ();
 sg13g2_decap_8 FILLER_57_356 ();
 sg13g2_fill_1 FILLER_57_363 ();
 sg13g2_decap_4 FILLER_57_400 ();
 sg13g2_decap_4 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_414 ();
 sg13g2_decap_4 FILLER_57_421 ();
 sg13g2_fill_2 FILLER_57_483 ();
 sg13g2_fill_1 FILLER_57_485 ();
 sg13g2_fill_2 FILLER_57_495 ();
 sg13g2_fill_1 FILLER_57_497 ();
 sg13g2_fill_1 FILLER_57_502 ();
 sg13g2_fill_2 FILLER_57_507 ();
 sg13g2_decap_4 FILLER_57_513 ();
 sg13g2_decap_4 FILLER_57_529 ();
 sg13g2_decap_4 FILLER_57_545 ();
 sg13g2_fill_1 FILLER_57_549 ();
 sg13g2_decap_8 FILLER_57_555 ();
 sg13g2_decap_8 FILLER_57_562 ();
 sg13g2_decap_4 FILLER_57_569 ();
 sg13g2_fill_1 FILLER_57_573 ();
 sg13g2_fill_2 FILLER_57_594 ();
 sg13g2_fill_2 FILLER_57_606 ();
 sg13g2_fill_2 FILLER_57_612 ();
 sg13g2_fill_1 FILLER_57_632 ();
 sg13g2_fill_1 FILLER_57_642 ();
 sg13g2_decap_4 FILLER_57_651 ();
 sg13g2_fill_2 FILLER_57_655 ();
 sg13g2_decap_4 FILLER_57_662 ();
 sg13g2_fill_1 FILLER_57_666 ();
 sg13g2_fill_2 FILLER_57_698 ();
 sg13g2_fill_1 FILLER_57_704 ();
 sg13g2_fill_2 FILLER_57_709 ();
 sg13g2_fill_1 FILLER_57_711 ();
 sg13g2_decap_8 FILLER_57_717 ();
 sg13g2_decap_8 FILLER_57_724 ();
 sg13g2_decap_8 FILLER_57_731 ();
 sg13g2_fill_1 FILLER_57_738 ();
 sg13g2_decap_8 FILLER_57_774 ();
 sg13g2_decap_4 FILLER_57_781 ();
 sg13g2_fill_1 FILLER_57_785 ();
 sg13g2_decap_4 FILLER_57_794 ();
 sg13g2_fill_1 FILLER_57_803 ();
 sg13g2_fill_1 FILLER_57_830 ();
 sg13g2_decap_8 FILLER_57_837 ();
 sg13g2_decap_8 FILLER_57_844 ();
 sg13g2_fill_1 FILLER_57_879 ();
 sg13g2_decap_4 FILLER_57_906 ();
 sg13g2_fill_2 FILLER_57_910 ();
 sg13g2_decap_8 FILLER_57_972 ();
 sg13g2_decap_8 FILLER_57_979 ();
 sg13g2_fill_1 FILLER_57_986 ();
 sg13g2_fill_1 FILLER_57_992 ();
 sg13g2_fill_1 FILLER_57_1017 ();
 sg13g2_decap_4 FILLER_57_1028 ();
 sg13g2_fill_2 FILLER_57_1032 ();
 sg13g2_fill_2 FILLER_57_1039 ();
 sg13g2_fill_1 FILLER_57_1041 ();
 sg13g2_decap_8 FILLER_57_1046 ();
 sg13g2_fill_1 FILLER_57_1053 ();
 sg13g2_decap_8 FILLER_57_1059 ();
 sg13g2_decap_4 FILLER_57_1066 ();
 sg13g2_fill_2 FILLER_57_1070 ();
 sg13g2_decap_8 FILLER_57_1078 ();
 sg13g2_fill_1 FILLER_57_1085 ();
 sg13g2_fill_2 FILLER_57_1108 ();
 sg13g2_fill_2 FILLER_57_1118 ();
 sg13g2_decap_4 FILLER_57_1130 ();
 sg13g2_decap_8 FILLER_57_1137 ();
 sg13g2_fill_1 FILLER_57_1144 ();
 sg13g2_decap_8 FILLER_57_1150 ();
 sg13g2_decap_4 FILLER_57_1157 ();
 sg13g2_fill_2 FILLER_57_1161 ();
 sg13g2_decap_8 FILLER_57_1167 ();
 sg13g2_decap_8 FILLER_57_1174 ();
 sg13g2_fill_2 FILLER_57_1181 ();
 sg13g2_decap_8 FILLER_57_1187 ();
 sg13g2_decap_4 FILLER_57_1194 ();
 sg13g2_fill_2 FILLER_57_1211 ();
 sg13g2_fill_1 FILLER_57_1218 ();
 sg13g2_fill_2 FILLER_57_1229 ();
 sg13g2_fill_2 FILLER_57_1269 ();
 sg13g2_decap_8 FILLER_57_1297 ();
 sg13g2_decap_8 FILLER_57_1304 ();
 sg13g2_fill_2 FILLER_57_1311 ();
 sg13g2_decap_8 FILLER_57_1318 ();
 sg13g2_fill_1 FILLER_57_1325 ();
 sg13g2_decap_4 FILLER_57_1330 ();
 sg13g2_fill_2 FILLER_57_1360 ();
 sg13g2_decap_8 FILLER_57_1393 ();
 sg13g2_decap_4 FILLER_57_1400 ();
 sg13g2_fill_1 FILLER_57_1404 ();
 sg13g2_fill_1 FILLER_57_1414 ();
 sg13g2_decap_4 FILLER_57_1420 ();
 sg13g2_fill_1 FILLER_57_1437 ();
 sg13g2_decap_8 FILLER_57_1450 ();
 sg13g2_decap_4 FILLER_57_1457 ();
 sg13g2_fill_1 FILLER_57_1461 ();
 sg13g2_decap_4 FILLER_57_1467 ();
 sg13g2_fill_1 FILLER_57_1475 ();
 sg13g2_decap_8 FILLER_57_1480 ();
 sg13g2_decap_4 FILLER_57_1487 ();
 sg13g2_fill_2 FILLER_57_1491 ();
 sg13g2_decap_4 FILLER_57_1498 ();
 sg13g2_fill_2 FILLER_57_1502 ();
 sg13g2_fill_2 FILLER_57_1509 ();
 sg13g2_fill_1 FILLER_57_1516 ();
 sg13g2_decap_8 FILLER_57_1543 ();
 sg13g2_fill_2 FILLER_57_1550 ();
 sg13g2_fill_1 FILLER_57_1552 ();
 sg13g2_decap_4 FILLER_57_1561 ();
 sg13g2_fill_2 FILLER_57_1565 ();
 sg13g2_decap_8 FILLER_57_1597 ();
 sg13g2_decap_8 FILLER_57_1604 ();
 sg13g2_fill_2 FILLER_57_1611 ();
 sg13g2_fill_2 FILLER_57_1631 ();
 sg13g2_fill_1 FILLER_57_1633 ();
 sg13g2_decap_8 FILLER_57_1664 ();
 sg13g2_fill_2 FILLER_57_1671 ();
 sg13g2_fill_2 FILLER_57_1680 ();
 sg13g2_fill_1 FILLER_57_1682 ();
 sg13g2_decap_8 FILLER_57_1695 ();
 sg13g2_fill_1 FILLER_57_1702 ();
 sg13g2_fill_1 FILLER_57_1706 ();
 sg13g2_fill_2 FILLER_57_1712 ();
 sg13g2_fill_1 FILLER_57_1714 ();
 sg13g2_decap_4 FILLER_57_1731 ();
 sg13g2_fill_1 FILLER_57_1735 ();
 sg13g2_decap_8 FILLER_57_1744 ();
 sg13g2_decap_4 FILLER_57_1799 ();
 sg13g2_fill_2 FILLER_57_1803 ();
 sg13g2_fill_1 FILLER_57_1816 ();
 sg13g2_fill_1 FILLER_57_1830 ();
 sg13g2_fill_1 FILLER_57_1847 ();
 sg13g2_decap_8 FILLER_57_1908 ();
 sg13g2_fill_2 FILLER_57_1915 ();
 sg13g2_decap_8 FILLER_57_1933 ();
 sg13g2_decap_4 FILLER_57_1945 ();
 sg13g2_decap_4 FILLER_57_1970 ();
 sg13g2_fill_2 FILLER_57_1974 ();
 sg13g2_fill_1 FILLER_57_1987 ();
 sg13g2_decap_8 FILLER_57_1994 ();
 sg13g2_decap_4 FILLER_57_2001 ();
 sg13g2_fill_1 FILLER_57_2005 ();
 sg13g2_fill_2 FILLER_57_2061 ();
 sg13g2_fill_1 FILLER_57_2072 ();
 sg13g2_fill_2 FILLER_57_2087 ();
 sg13g2_fill_1 FILLER_57_2089 ();
 sg13g2_fill_1 FILLER_57_2093 ();
 sg13g2_fill_1 FILLER_57_2104 ();
 sg13g2_fill_1 FILLER_57_2115 ();
 sg13g2_fill_2 FILLER_57_2132 ();
 sg13g2_fill_2 FILLER_57_2139 ();
 sg13g2_fill_2 FILLER_57_2145 ();
 sg13g2_decap_8 FILLER_57_2152 ();
 sg13g2_fill_2 FILLER_57_2159 ();
 sg13g2_fill_1 FILLER_57_2161 ();
 sg13g2_fill_1 FILLER_57_2172 ();
 sg13g2_fill_2 FILLER_57_2199 ();
 sg13g2_fill_1 FILLER_57_2201 ();
 sg13g2_decap_8 FILLER_57_2211 ();
 sg13g2_decap_8 FILLER_57_2218 ();
 sg13g2_decap_8 FILLER_57_2251 ();
 sg13g2_decap_8 FILLER_57_2258 ();
 sg13g2_fill_2 FILLER_57_2265 ();
 sg13g2_fill_1 FILLER_57_2267 ();
 sg13g2_fill_1 FILLER_57_2302 ();
 sg13g2_decap_8 FILLER_57_2311 ();
 sg13g2_fill_1 FILLER_57_2318 ();
 sg13g2_decap_8 FILLER_57_2323 ();
 sg13g2_fill_1 FILLER_57_2330 ();
 sg13g2_decap_4 FILLER_57_2335 ();
 sg13g2_fill_1 FILLER_57_2339 ();
 sg13g2_decap_8 FILLER_57_2366 ();
 sg13g2_decap_8 FILLER_57_2373 ();
 sg13g2_fill_2 FILLER_57_2380 ();
 sg13g2_fill_1 FILLER_57_2382 ();
 sg13g2_fill_1 FILLER_57_2400 ();
 sg13g2_fill_2 FILLER_57_2420 ();
 sg13g2_fill_1 FILLER_57_2492 ();
 sg13g2_fill_2 FILLER_57_2497 ();
 sg13g2_fill_1 FILLER_57_2499 ();
 sg13g2_fill_2 FILLER_57_2526 ();
 sg13g2_fill_1 FILLER_57_2528 ();
 sg13g2_fill_1 FILLER_57_2541 ();
 sg13g2_decap_4 FILLER_57_2546 ();
 sg13g2_decap_8 FILLER_57_2620 ();
 sg13g2_fill_1 FILLER_57_2639 ();
 sg13g2_decap_8 FILLER_57_2651 ();
 sg13g2_decap_8 FILLER_57_2658 ();
 sg13g2_decap_4 FILLER_57_2665 ();
 sg13g2_fill_1 FILLER_57_2669 ();
 sg13g2_fill_2 FILLER_58_0 ();
 sg13g2_decap_4 FILLER_58_40 ();
 sg13g2_fill_1 FILLER_58_44 ();
 sg13g2_fill_2 FILLER_58_75 ();
 sg13g2_fill_1 FILLER_58_77 ();
 sg13g2_decap_4 FILLER_58_98 ();
 sg13g2_fill_1 FILLER_58_132 ();
 sg13g2_fill_1 FILLER_58_143 ();
 sg13g2_fill_2 FILLER_58_167 ();
 sg13g2_fill_1 FILLER_58_169 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_decap_4 FILLER_58_248 ();
 sg13g2_fill_1 FILLER_58_252 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_decap_8 FILLER_58_302 ();
 sg13g2_decap_4 FILLER_58_309 ();
 sg13g2_decap_4 FILLER_58_351 ();
 sg13g2_fill_2 FILLER_58_355 ();
 sg13g2_decap_4 FILLER_58_364 ();
 sg13g2_fill_1 FILLER_58_368 ();
 sg13g2_fill_2 FILLER_58_396 ();
 sg13g2_fill_1 FILLER_58_398 ();
 sg13g2_fill_2 FILLER_58_470 ();
 sg13g2_fill_1 FILLER_58_472 ();
 sg13g2_decap_8 FILLER_58_480 ();
 sg13g2_decap_4 FILLER_58_487 ();
 sg13g2_fill_1 FILLER_58_495 ();
 sg13g2_decap_8 FILLER_58_515 ();
 sg13g2_decap_8 FILLER_58_522 ();
 sg13g2_fill_1 FILLER_58_529 ();
 sg13g2_decap_8 FILLER_58_564 ();
 sg13g2_decap_8 FILLER_58_571 ();
 sg13g2_fill_2 FILLER_58_640 ();
 sg13g2_decap_4 FILLER_58_647 ();
 sg13g2_fill_2 FILLER_58_656 ();
 sg13g2_fill_1 FILLER_58_658 ();
 sg13g2_fill_2 FILLER_58_662 ();
 sg13g2_fill_1 FILLER_58_664 ();
 sg13g2_decap_4 FILLER_58_674 ();
 sg13g2_fill_1 FILLER_58_678 ();
 sg13g2_fill_1 FILLER_58_690 ();
 sg13g2_decap_8 FILLER_58_706 ();
 sg13g2_decap_8 FILLER_58_713 ();
 sg13g2_decap_8 FILLER_58_720 ();
 sg13g2_fill_2 FILLER_58_727 ();
 sg13g2_fill_1 FILLER_58_729 ();
 sg13g2_decap_4 FILLER_58_738 ();
 sg13g2_decap_8 FILLER_58_747 ();
 sg13g2_decap_4 FILLER_58_754 ();
 sg13g2_fill_1 FILLER_58_758 ();
 sg13g2_decap_8 FILLER_58_764 ();
 sg13g2_decap_8 FILLER_58_776 ();
 sg13g2_fill_2 FILLER_58_783 ();
 sg13g2_fill_1 FILLER_58_785 ();
 sg13g2_decap_4 FILLER_58_791 ();
 sg13g2_fill_2 FILLER_58_795 ();
 sg13g2_fill_1 FILLER_58_801 ();
 sg13g2_fill_1 FILLER_58_834 ();
 sg13g2_decap_8 FILLER_58_841 ();
 sg13g2_decap_8 FILLER_58_848 ();
 sg13g2_fill_2 FILLER_58_855 ();
 sg13g2_fill_2 FILLER_58_883 ();
 sg13g2_fill_1 FILLER_58_909 ();
 sg13g2_fill_1 FILLER_58_915 ();
 sg13g2_fill_1 FILLER_58_924 ();
 sg13g2_fill_2 FILLER_58_936 ();
 sg13g2_fill_1 FILLER_58_949 ();
 sg13g2_fill_1 FILLER_58_955 ();
 sg13g2_fill_1 FILLER_58_982 ();
 sg13g2_decap_8 FILLER_58_1015 ();
 sg13g2_decap_8 FILLER_58_1027 ();
 sg13g2_decap_8 FILLER_58_1034 ();
 sg13g2_decap_4 FILLER_58_1041 ();
 sg13g2_fill_2 FILLER_58_1045 ();
 sg13g2_decap_4 FILLER_58_1073 ();
 sg13g2_fill_1 FILLER_58_1077 ();
 sg13g2_decap_8 FILLER_58_1083 ();
 sg13g2_fill_2 FILLER_58_1090 ();
 sg13g2_fill_1 FILLER_58_1092 ();
 sg13g2_fill_1 FILLER_58_1128 ();
 sg13g2_decap_4 FILLER_58_1194 ();
 sg13g2_fill_1 FILLER_58_1198 ();
 sg13g2_fill_2 FILLER_58_1228 ();
 sg13g2_fill_2 FILLER_58_1262 ();
 sg13g2_fill_1 FILLER_58_1264 ();
 sg13g2_decap_8 FILLER_58_1287 ();
 sg13g2_decap_4 FILLER_58_1294 ();
 sg13g2_fill_1 FILLER_58_1302 ();
 sg13g2_fill_1 FILLER_58_1309 ();
 sg13g2_fill_1 FILLER_58_1314 ();
 sg13g2_fill_1 FILLER_58_1341 ();
 sg13g2_fill_1 FILLER_58_1350 ();
 sg13g2_fill_2 FILLER_58_1356 ();
 sg13g2_fill_2 FILLER_58_1363 ();
 sg13g2_fill_1 FILLER_58_1365 ();
 sg13g2_fill_1 FILLER_58_1371 ();
 sg13g2_fill_2 FILLER_58_1376 ();
 sg13g2_fill_1 FILLER_58_1378 ();
 sg13g2_fill_2 FILLER_58_1463 ();
 sg13g2_decap_8 FILLER_58_1491 ();
 sg13g2_decap_8 FILLER_58_1498 ();
 sg13g2_decap_8 FILLER_58_1505 ();
 sg13g2_decap_8 FILLER_58_1512 ();
 sg13g2_decap_8 FILLER_58_1519 ();
 sg13g2_decap_8 FILLER_58_1526 ();
 sg13g2_decap_8 FILLER_58_1533 ();
 sg13g2_decap_4 FILLER_58_1540 ();
 sg13g2_fill_1 FILLER_58_1552 ();
 sg13g2_decap_8 FILLER_58_1557 ();
 sg13g2_decap_8 FILLER_58_1564 ();
 sg13g2_fill_2 FILLER_58_1571 ();
 sg13g2_decap_4 FILLER_58_1611 ();
 sg13g2_decap_8 FILLER_58_1653 ();
 sg13g2_fill_2 FILLER_58_1660 ();
 sg13g2_fill_1 FILLER_58_1662 ();
 sg13g2_decap_8 FILLER_58_1668 ();
 sg13g2_fill_2 FILLER_58_1675 ();
 sg13g2_fill_1 FILLER_58_1702 ();
 sg13g2_fill_2 FILLER_58_1713 ();
 sg13g2_fill_1 FILLER_58_1715 ();
 sg13g2_fill_2 FILLER_58_1746 ();
 sg13g2_decap_4 FILLER_58_1757 ();
 sg13g2_decap_4 FILLER_58_1787 ();
 sg13g2_fill_2 FILLER_58_1826 ();
 sg13g2_fill_1 FILLER_58_1842 ();
 sg13g2_fill_1 FILLER_58_1851 ();
 sg13g2_fill_1 FILLER_58_1878 ();
 sg13g2_decap_8 FILLER_58_1883 ();
 sg13g2_fill_2 FILLER_58_1895 ();
 sg13g2_decap_4 FILLER_58_1900 ();
 sg13g2_fill_1 FILLER_58_1904 ();
 sg13g2_decap_4 FILLER_58_1940 ();
 sg13g2_fill_2 FILLER_58_1976 ();
 sg13g2_fill_1 FILLER_58_1978 ();
 sg13g2_fill_2 FILLER_58_1988 ();
 sg13g2_fill_2 FILLER_58_1999 ();
 sg13g2_decap_8 FILLER_58_2016 ();
 sg13g2_fill_2 FILLER_58_2023 ();
 sg13g2_fill_1 FILLER_58_2025 ();
 sg13g2_fill_1 FILLER_58_2029 ();
 sg13g2_fill_2 FILLER_58_2033 ();
 sg13g2_fill_1 FILLER_58_2035 ();
 sg13g2_decap_4 FILLER_58_2040 ();
 sg13g2_fill_2 FILLER_58_2064 ();
 sg13g2_fill_2 FILLER_58_2080 ();
 sg13g2_fill_1 FILLER_58_2100 ();
 sg13g2_fill_2 FILLER_58_2158 ();
 sg13g2_fill_1 FILLER_58_2209 ();
 sg13g2_decap_8 FILLER_58_2214 ();
 sg13g2_decap_8 FILLER_58_2221 ();
 sg13g2_fill_2 FILLER_58_2228 ();
 sg13g2_fill_1 FILLER_58_2230 ();
 sg13g2_fill_1 FILLER_58_2235 ();
 sg13g2_fill_2 FILLER_58_2250 ();
 sg13g2_fill_1 FILLER_58_2252 ();
 sg13g2_fill_1 FILLER_58_2259 ();
 sg13g2_decap_8 FILLER_58_2264 ();
 sg13g2_decap_8 FILLER_58_2271 ();
 sg13g2_decap_8 FILLER_58_2278 ();
 sg13g2_decap_8 FILLER_58_2298 ();
 sg13g2_fill_1 FILLER_58_2305 ();
 sg13g2_fill_2 FILLER_58_2316 ();
 sg13g2_fill_2 FILLER_58_2344 ();
 sg13g2_fill_1 FILLER_58_2346 ();
 sg13g2_fill_2 FILLER_58_2351 ();
 sg13g2_fill_1 FILLER_58_2353 ();
 sg13g2_fill_2 FILLER_58_2380 ();
 sg13g2_decap_8 FILLER_58_2386 ();
 sg13g2_decap_4 FILLER_58_2393 ();
 sg13g2_fill_1 FILLER_58_2397 ();
 sg13g2_fill_2 FILLER_58_2430 ();
 sg13g2_fill_1 FILLER_58_2432 ();
 sg13g2_fill_2 FILLER_58_2446 ();
 sg13g2_fill_1 FILLER_58_2456 ();
 sg13g2_decap_8 FILLER_58_2476 ();
 sg13g2_decap_8 FILLER_58_2483 ();
 sg13g2_decap_8 FILLER_58_2490 ();
 sg13g2_decap_4 FILLER_58_2497 ();
 sg13g2_fill_1 FILLER_58_2501 ();
 sg13g2_decap_8 FILLER_58_2506 ();
 sg13g2_fill_2 FILLER_58_2513 ();
 sg13g2_fill_2 FILLER_58_2545 ();
 sg13g2_fill_1 FILLER_58_2547 ();
 sg13g2_decap_4 FILLER_58_2565 ();
 sg13g2_decap_8 FILLER_58_2577 ();
 sg13g2_decap_8 FILLER_58_2584 ();
 sg13g2_decap_8 FILLER_58_2604 ();
 sg13g2_decap_8 FILLER_58_2611 ();
 sg13g2_fill_2 FILLER_58_2618 ();
 sg13g2_decap_8 FILLER_58_2659 ();
 sg13g2_decap_4 FILLER_58_2666 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_fill_2 FILLER_59_31 ();
 sg13g2_fill_2 FILLER_59_53 ();
 sg13g2_fill_1 FILLER_59_65 ();
 sg13g2_decap_8 FILLER_59_76 ();
 sg13g2_fill_2 FILLER_59_98 ();
 sg13g2_fill_1 FILLER_59_105 ();
 sg13g2_fill_2 FILLER_59_133 ();
 sg13g2_fill_2 FILLER_59_157 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_2 FILLER_59_164 ();
 sg13g2_decap_4 FILLER_59_184 ();
 sg13g2_fill_2 FILLER_59_188 ();
 sg13g2_fill_2 FILLER_59_195 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_decap_4 FILLER_59_208 ();
 sg13g2_fill_2 FILLER_59_212 ();
 sg13g2_decap_4 FILLER_59_240 ();
 sg13g2_decap_8 FILLER_59_270 ();
 sg13g2_decap_8 FILLER_59_277 ();
 sg13g2_decap_8 FILLER_59_294 ();
 sg13g2_decap_4 FILLER_59_301 ();
 sg13g2_fill_2 FILLER_59_305 ();
 sg13g2_fill_2 FILLER_59_331 ();
 sg13g2_fill_2 FILLER_59_338 ();
 sg13g2_decap_4 FILLER_59_366 ();
 sg13g2_fill_2 FILLER_59_370 ();
 sg13g2_fill_2 FILLER_59_377 ();
 sg13g2_fill_1 FILLER_59_379 ();
 sg13g2_decap_8 FILLER_59_390 ();
 sg13g2_decap_8 FILLER_59_397 ();
 sg13g2_decap_4 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_412 ();
 sg13g2_fill_2 FILLER_59_421 ();
 sg13g2_fill_2 FILLER_59_436 ();
 sg13g2_fill_1 FILLER_59_443 ();
 sg13g2_decap_4 FILLER_59_464 ();
 sg13g2_fill_1 FILLER_59_468 ();
 sg13g2_fill_2 FILLER_59_505 ();
 sg13g2_decap_8 FILLER_59_515 ();
 sg13g2_decap_8 FILLER_59_522 ();
 sg13g2_fill_1 FILLER_59_529 ();
 sg13g2_decap_8 FILLER_59_534 ();
 sg13g2_decap_8 FILLER_59_541 ();
 sg13g2_decap_4 FILLER_59_548 ();
 sg13g2_fill_1 FILLER_59_552 ();
 sg13g2_decap_8 FILLER_59_584 ();
 sg13g2_decap_8 FILLER_59_591 ();
 sg13g2_decap_4 FILLER_59_598 ();
 sg13g2_fill_1 FILLER_59_602 ();
 sg13g2_decap_8 FILLER_59_610 ();
 sg13g2_fill_2 FILLER_59_617 ();
 sg13g2_fill_1 FILLER_59_619 ();
 sg13g2_decap_4 FILLER_59_637 ();
 sg13g2_decap_4 FILLER_59_646 ();
 sg13g2_fill_2 FILLER_59_650 ();
 sg13g2_decap_8 FILLER_59_660 ();
 sg13g2_fill_2 FILLER_59_667 ();
 sg13g2_fill_1 FILLER_59_669 ();
 sg13g2_decap_8 FILLER_59_707 ();
 sg13g2_decap_8 FILLER_59_714 ();
 sg13g2_fill_2 FILLER_59_721 ();
 sg13g2_fill_2 FILLER_59_758 ();
 sg13g2_decap_8 FILLER_59_786 ();
 sg13g2_fill_2 FILLER_59_793 ();
 sg13g2_fill_2 FILLER_59_800 ();
 sg13g2_fill_2 FILLER_59_833 ();
 sg13g2_decap_8 FILLER_59_841 ();
 sg13g2_decap_8 FILLER_59_848 ();
 sg13g2_decap_8 FILLER_59_855 ();
 sg13g2_decap_4 FILLER_59_862 ();
 sg13g2_fill_2 FILLER_59_866 ();
 sg13g2_decap_8 FILLER_59_876 ();
 sg13g2_fill_2 FILLER_59_883 ();
 sg13g2_fill_1 FILLER_59_929 ();
 sg13g2_decap_4 FILLER_59_939 ();
 sg13g2_fill_1 FILLER_59_943 ();
 sg13g2_fill_1 FILLER_59_949 ();
 sg13g2_decap_4 FILLER_59_954 ();
 sg13g2_fill_2 FILLER_59_958 ();
 sg13g2_decap_8 FILLER_59_963 ();
 sg13g2_fill_1 FILLER_59_970 ();
 sg13g2_fill_2 FILLER_59_976 ();
 sg13g2_fill_1 FILLER_59_1012 ();
 sg13g2_fill_2 FILLER_59_1017 ();
 sg13g2_decap_4 FILLER_59_1023 ();
 sg13g2_fill_2 FILLER_59_1027 ();
 sg13g2_fill_1 FILLER_59_1099 ();
 sg13g2_fill_2 FILLER_59_1164 ();
 sg13g2_decap_4 FILLER_59_1171 ();
 sg13g2_fill_1 FILLER_59_1175 ();
 sg13g2_fill_1 FILLER_59_1186 ();
 sg13g2_decap_4 FILLER_59_1199 ();
 sg13g2_decap_4 FILLER_59_1258 ();
 sg13g2_decap_8 FILLER_59_1319 ();
 sg13g2_fill_2 FILLER_59_1326 ();
 sg13g2_fill_2 FILLER_59_1332 ();
 sg13g2_fill_1 FILLER_59_1334 ();
 sg13g2_decap_8 FILLER_59_1365 ();
 sg13g2_fill_1 FILLER_59_1372 ();
 sg13g2_fill_2 FILLER_59_1382 ();
 sg13g2_fill_1 FILLER_59_1394 ();
 sg13g2_fill_2 FILLER_59_1404 ();
 sg13g2_decap_4 FILLER_59_1411 ();
 sg13g2_fill_2 FILLER_59_1415 ();
 sg13g2_fill_1 FILLER_59_1421 ();
 sg13g2_decap_4 FILLER_59_1453 ();
 sg13g2_fill_1 FILLER_59_1457 ();
 sg13g2_decap_8 FILLER_59_1495 ();
 sg13g2_decap_8 FILLER_59_1502 ();
 sg13g2_decap_4 FILLER_59_1509 ();
 sg13g2_fill_1 FILLER_59_1513 ();
 sg13g2_decap_4 FILLER_59_1532 ();
 sg13g2_fill_1 FILLER_59_1536 ();
 sg13g2_fill_1 FILLER_59_1542 ();
 sg13g2_fill_2 FILLER_59_1574 ();
 sg13g2_decap_4 FILLER_59_1580 ();
 sg13g2_fill_1 FILLER_59_1610 ();
 sg13g2_decap_4 FILLER_59_1642 ();
 sg13g2_fill_1 FILLER_59_1646 ();
 sg13g2_fill_2 FILLER_59_1751 ();
 sg13g2_fill_1 FILLER_59_1758 ();
 sg13g2_decap_8 FILLER_59_1768 ();
 sg13g2_decap_8 FILLER_59_1775 ();
 sg13g2_decap_8 FILLER_59_1782 ();
 sg13g2_decap_8 FILLER_59_1789 ();
 sg13g2_fill_2 FILLER_59_1796 ();
 sg13g2_decap_8 FILLER_59_1802 ();
 sg13g2_decap_4 FILLER_59_1809 ();
 sg13g2_fill_1 FILLER_59_1813 ();
 sg13g2_fill_2 FILLER_59_1821 ();
 sg13g2_fill_2 FILLER_59_1847 ();
 sg13g2_fill_2 FILLER_59_1854 ();
 sg13g2_fill_2 FILLER_59_1862 ();
 sg13g2_fill_2 FILLER_59_1876 ();
 sg13g2_decap_4 FILLER_59_1886 ();
 sg13g2_fill_2 FILLER_59_1890 ();
 sg13g2_fill_2 FILLER_59_1908 ();
 sg13g2_decap_4 FILLER_59_1915 ();
 sg13g2_fill_1 FILLER_59_1919 ();
 sg13g2_fill_1 FILLER_59_1939 ();
 sg13g2_fill_2 FILLER_59_1961 ();
 sg13g2_fill_1 FILLER_59_1963 ();
 sg13g2_fill_2 FILLER_59_1968 ();
 sg13g2_decap_8 FILLER_59_1975 ();
 sg13g2_decap_8 FILLER_59_1991 ();
 sg13g2_decap_8 FILLER_59_1998 ();
 sg13g2_fill_1 FILLER_59_2005 ();
 sg13g2_decap_8 FILLER_59_2014 ();
 sg13g2_decap_4 FILLER_59_2021 ();
 sg13g2_fill_1 FILLER_59_2025 ();
 sg13g2_decap_8 FILLER_59_2042 ();
 sg13g2_fill_2 FILLER_59_2049 ();
 sg13g2_fill_1 FILLER_59_2051 ();
 sg13g2_decap_8 FILLER_59_2056 ();
 sg13g2_fill_1 FILLER_59_2072 ();
 sg13g2_decap_8 FILLER_59_2079 ();
 sg13g2_decap_4 FILLER_59_2086 ();
 sg13g2_decap_4 FILLER_59_2093 ();
 sg13g2_fill_1 FILLER_59_2097 ();
 sg13g2_decap_8 FILLER_59_2102 ();
 sg13g2_fill_2 FILLER_59_2109 ();
 sg13g2_fill_2 FILLER_59_2123 ();
 sg13g2_fill_1 FILLER_59_2125 ();
 sg13g2_decap_4 FILLER_59_2206 ();
 sg13g2_fill_2 FILLER_59_2250 ();
 sg13g2_fill_2 FILLER_59_2278 ();
 sg13g2_fill_1 FILLER_59_2280 ();
 sg13g2_fill_1 FILLER_59_2311 ();
 sg13g2_decap_8 FILLER_59_2342 ();
 sg13g2_fill_2 FILLER_59_2349 ();
 sg13g2_fill_1 FILLER_59_2351 ();
 sg13g2_decap_4 FILLER_59_2356 ();
 sg13g2_fill_2 FILLER_59_2360 ();
 sg13g2_fill_1 FILLER_59_2374 ();
 sg13g2_decap_8 FILLER_59_2430 ();
 sg13g2_decap_8 FILLER_59_2437 ();
 sg13g2_decap_8 FILLER_59_2444 ();
 sg13g2_decap_4 FILLER_59_2451 ();
 sg13g2_fill_2 FILLER_59_2455 ();
 sg13g2_decap_8 FILLER_59_2460 ();
 sg13g2_decap_8 FILLER_59_2473 ();
 sg13g2_decap_4 FILLER_59_2480 ();
 sg13g2_fill_2 FILLER_59_2484 ();
 sg13g2_decap_4 FILLER_59_2498 ();
 sg13g2_fill_1 FILLER_59_2502 ();
 sg13g2_decap_4 FILLER_59_2529 ();
 sg13g2_fill_1 FILLER_59_2533 ();
 sg13g2_decap_4 FILLER_59_2540 ();
 sg13g2_fill_2 FILLER_59_2544 ();
 sg13g2_decap_8 FILLER_59_2572 ();
 sg13g2_decap_8 FILLER_59_2579 ();
 sg13g2_decap_8 FILLER_59_2586 ();
 sg13g2_fill_1 FILLER_59_2593 ();
 sg13g2_decap_8 FILLER_59_2604 ();
 sg13g2_decap_8 FILLER_59_2611 ();
 sg13g2_fill_2 FILLER_59_2618 ();
 sg13g2_decap_4 FILLER_59_2624 ();
 sg13g2_fill_1 FILLER_59_2633 ();
 sg13g2_decap_4 FILLER_59_2638 ();
 sg13g2_fill_2 FILLER_59_2668 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_18 ();
 sg13g2_fill_1 FILLER_60_67 ();
 sg13g2_fill_2 FILLER_60_78 ();
 sg13g2_fill_1 FILLER_60_85 ();
 sg13g2_fill_2 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_127 ();
 sg13g2_decap_8 FILLER_60_142 ();
 sg13g2_fill_2 FILLER_60_149 ();
 sg13g2_fill_2 FILLER_60_164 ();
 sg13g2_decap_8 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_219 ();
 sg13g2_fill_2 FILLER_60_230 ();
 sg13g2_fill_1 FILLER_60_232 ();
 sg13g2_decap_8 FILLER_60_253 ();
 sg13g2_decap_4 FILLER_60_260 ();
 sg13g2_fill_2 FILLER_60_264 ();
 sg13g2_fill_2 FILLER_60_303 ();
 sg13g2_fill_2 FILLER_60_320 ();
 sg13g2_decap_8 FILLER_60_329 ();
 sg13g2_fill_2 FILLER_60_336 ();
 sg13g2_fill_1 FILLER_60_338 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_375 ();
 sg13g2_fill_1 FILLER_60_399 ();
 sg13g2_fill_2 FILLER_60_405 ();
 sg13g2_fill_1 FILLER_60_407 ();
 sg13g2_fill_1 FILLER_60_420 ();
 sg13g2_fill_1 FILLER_60_426 ();
 sg13g2_fill_1 FILLER_60_432 ();
 sg13g2_fill_2 FILLER_60_443 ();
 sg13g2_decap_8 FILLER_60_458 ();
 sg13g2_decap_4 FILLER_60_465 ();
 sg13g2_fill_1 FILLER_60_469 ();
 sg13g2_decap_8 FILLER_60_477 ();
 sg13g2_fill_2 FILLER_60_484 ();
 sg13g2_decap_4 FILLER_60_520 ();
 sg13g2_fill_1 FILLER_60_524 ();
 sg13g2_fill_2 FILLER_60_530 ();
 sg13g2_fill_1 FILLER_60_532 ();
 sg13g2_decap_8 FILLER_60_546 ();
 sg13g2_decap_8 FILLER_60_553 ();
 sg13g2_decap_8 FILLER_60_560 ();
 sg13g2_decap_8 FILLER_60_567 ();
 sg13g2_decap_8 FILLER_60_574 ();
 sg13g2_fill_2 FILLER_60_581 ();
 sg13g2_fill_1 FILLER_60_583 ();
 sg13g2_fill_1 FILLER_60_593 ();
 sg13g2_fill_1 FILLER_60_600 ();
 sg13g2_decap_8 FILLER_60_609 ();
 sg13g2_decap_4 FILLER_60_616 ();
 sg13g2_fill_1 FILLER_60_620 ();
 sg13g2_fill_2 FILLER_60_639 ();
 sg13g2_decap_8 FILLER_60_658 ();
 sg13g2_decap_8 FILLER_60_665 ();
 sg13g2_decap_4 FILLER_60_672 ();
 sg13g2_fill_2 FILLER_60_676 ();
 sg13g2_fill_1 FILLER_60_682 ();
 sg13g2_fill_1 FILLER_60_688 ();
 sg13g2_fill_1 FILLER_60_694 ();
 sg13g2_decap_8 FILLER_60_700 ();
 sg13g2_decap_8 FILLER_60_707 ();
 sg13g2_decap_4 FILLER_60_714 ();
 sg13g2_fill_1 FILLER_60_718 ();
 sg13g2_decap_8 FILLER_60_745 ();
 sg13g2_decap_8 FILLER_60_752 ();
 sg13g2_decap_8 FILLER_60_759 ();
 sg13g2_decap_4 FILLER_60_766 ();
 sg13g2_fill_2 FILLER_60_775 ();
 sg13g2_decap_8 FILLER_60_807 ();
 sg13g2_fill_2 FILLER_60_814 ();
 sg13g2_fill_1 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_843 ();
 sg13g2_decap_8 FILLER_60_850 ();
 sg13g2_fill_1 FILLER_60_857 ();
 sg13g2_fill_2 FILLER_60_890 ();
 sg13g2_fill_2 FILLER_60_910 ();
 sg13g2_fill_1 FILLER_60_912 ();
 sg13g2_fill_2 FILLER_60_922 ();
 sg13g2_fill_2 FILLER_60_994 ();
 sg13g2_fill_1 FILLER_60_996 ();
 sg13g2_fill_2 FILLER_60_1001 ();
 sg13g2_fill_1 FILLER_60_1008 ();
 sg13g2_fill_2 FILLER_60_1035 ();
 sg13g2_fill_2 FILLER_60_1041 ();
 sg13g2_fill_1 FILLER_60_1053 ();
 sg13g2_decap_4 FILLER_60_1058 ();
 sg13g2_fill_1 FILLER_60_1071 ();
 sg13g2_decap_8 FILLER_60_1078 ();
 sg13g2_fill_1 FILLER_60_1098 ();
 sg13g2_fill_1 FILLER_60_1103 ();
 sg13g2_fill_1 FILLER_60_1112 ();
 sg13g2_fill_1 FILLER_60_1118 ();
 sg13g2_fill_1 FILLER_60_1140 ();
 sg13g2_decap_8 FILLER_60_1146 ();
 sg13g2_decap_8 FILLER_60_1153 ();
 sg13g2_fill_2 FILLER_60_1160 ();
 sg13g2_decap_4 FILLER_60_1168 ();
 sg13g2_fill_1 FILLER_60_1172 ();
 sg13g2_decap_8 FILLER_60_1198 ();
 sg13g2_fill_1 FILLER_60_1205 ();
 sg13g2_fill_1 FILLER_60_1232 ();
 sg13g2_fill_2 FILLER_60_1239 ();
 sg13g2_fill_2 FILLER_60_1244 ();
 sg13g2_fill_1 FILLER_60_1246 ();
 sg13g2_fill_1 FILLER_60_1253 ();
 sg13g2_decap_4 FILLER_60_1260 ();
 sg13g2_decap_8 FILLER_60_1272 ();
 sg13g2_decap_4 FILLER_60_1279 ();
 sg13g2_fill_1 FILLER_60_1283 ();
 sg13g2_decap_8 FILLER_60_1293 ();
 sg13g2_decap_4 FILLER_60_1300 ();
 sg13g2_fill_1 FILLER_60_1304 ();
 sg13g2_fill_2 FILLER_60_1311 ();
 sg13g2_fill_1 FILLER_60_1313 ();
 sg13g2_decap_4 FILLER_60_1340 ();
 sg13g2_fill_2 FILLER_60_1344 ();
 sg13g2_decap_8 FILLER_60_1367 ();
 sg13g2_decap_8 FILLER_60_1374 ();
 sg13g2_fill_2 FILLER_60_1381 ();
 sg13g2_decap_8 FILLER_60_1396 ();
 sg13g2_decap_8 FILLER_60_1403 ();
 sg13g2_decap_4 FILLER_60_1410 ();
 sg13g2_fill_2 FILLER_60_1418 ();
 sg13g2_fill_1 FILLER_60_1425 ();
 sg13g2_decap_8 FILLER_60_1432 ();
 sg13g2_decap_8 FILLER_60_1439 ();
 sg13g2_fill_2 FILLER_60_1446 ();
 sg13g2_fill_1 FILLER_60_1448 ();
 sg13g2_decap_8 FILLER_60_1481 ();
 sg13g2_decap_8 FILLER_60_1488 ();
 sg13g2_decap_4 FILLER_60_1495 ();
 sg13g2_fill_1 FILLER_60_1499 ();
 sg13g2_decap_8 FILLER_60_1516 ();
 sg13g2_decap_4 FILLER_60_1523 ();
 sg13g2_decap_8 FILLER_60_1558 ();
 sg13g2_decap_8 FILLER_60_1565 ();
 sg13g2_fill_2 FILLER_60_1572 ();
 sg13g2_fill_1 FILLER_60_1574 ();
 sg13g2_fill_1 FILLER_60_1580 ();
 sg13g2_decap_4 FILLER_60_1611 ();
 sg13g2_decap_4 FILLER_60_1623 ();
 sg13g2_decap_4 FILLER_60_1636 ();
 sg13g2_decap_8 FILLER_60_1644 ();
 sg13g2_decap_4 FILLER_60_1659 ();
 sg13g2_fill_2 FILLER_60_1681 ();
 sg13g2_fill_1 FILLER_60_1683 ();
 sg13g2_decap_8 FILLER_60_1688 ();
 sg13g2_fill_1 FILLER_60_1695 ();
 sg13g2_decap_4 FILLER_60_1704 ();
 sg13g2_fill_1 FILLER_60_1708 ();
 sg13g2_fill_2 FILLER_60_1745 ();
 sg13g2_fill_2 FILLER_60_1762 ();
 sg13g2_fill_2 FILLER_60_1769 ();
 sg13g2_decap_8 FILLER_60_1801 ();
 sg13g2_decap_8 FILLER_60_1808 ();
 sg13g2_decap_8 FILLER_60_1815 ();
 sg13g2_fill_1 FILLER_60_1822 ();
 sg13g2_fill_1 FILLER_60_1827 ();
 sg13g2_fill_1 FILLER_60_1858 ();
 sg13g2_decap_8 FILLER_60_1884 ();
 sg13g2_fill_2 FILLER_60_1917 ();
 sg13g2_fill_1 FILLER_60_1919 ();
 sg13g2_fill_2 FILLER_60_1928 ();
 sg13g2_fill_1 FILLER_60_1930 ();
 sg13g2_decap_4 FILLER_60_1999 ();
 sg13g2_fill_2 FILLER_60_2003 ();
 sg13g2_decap_4 FILLER_60_2010 ();
 sg13g2_fill_1 FILLER_60_2014 ();
 sg13g2_fill_2 FILLER_60_2024 ();
 sg13g2_fill_1 FILLER_60_2033 ();
 sg13g2_decap_8 FILLER_60_2038 ();
 sg13g2_decap_8 FILLER_60_2045 ();
 sg13g2_decap_4 FILLER_60_2056 ();
 sg13g2_fill_1 FILLER_60_2060 ();
 sg13g2_fill_1 FILLER_60_2124 ();
 sg13g2_decap_8 FILLER_60_2154 ();
 sg13g2_decap_4 FILLER_60_2161 ();
 sg13g2_fill_1 FILLER_60_2165 ();
 sg13g2_decap_8 FILLER_60_2225 ();
 sg13g2_decap_8 FILLER_60_2232 ();
 sg13g2_decap_8 FILLER_60_2239 ();
 sg13g2_decap_8 FILLER_60_2246 ();
 sg13g2_decap_8 FILLER_60_2253 ();
 sg13g2_decap_4 FILLER_60_2260 ();
 sg13g2_fill_2 FILLER_60_2264 ();
 sg13g2_decap_8 FILLER_60_2310 ();
 sg13g2_decap_8 FILLER_60_2317 ();
 sg13g2_decap_8 FILLER_60_2324 ();
 sg13g2_decap_8 FILLER_60_2335 ();
 sg13g2_decap_8 FILLER_60_2342 ();
 sg13g2_decap_8 FILLER_60_2349 ();
 sg13g2_fill_2 FILLER_60_2356 ();
 sg13g2_fill_1 FILLER_60_2358 ();
 sg13g2_fill_2 FILLER_60_2363 ();
 sg13g2_decap_4 FILLER_60_2369 ();
 sg13g2_fill_1 FILLER_60_2373 ();
 sg13g2_fill_2 FILLER_60_2426 ();
 sg13g2_fill_1 FILLER_60_2428 ();
 sg13g2_decap_8 FILLER_60_2459 ();
 sg13g2_decap_4 FILLER_60_2466 ();
 sg13g2_fill_2 FILLER_60_2470 ();
 sg13g2_decap_8 FILLER_60_2482 ();
 sg13g2_decap_8 FILLER_60_2489 ();
 sg13g2_decap_4 FILLER_60_2496 ();
 sg13g2_fill_1 FILLER_60_2500 ();
 sg13g2_decap_8 FILLER_60_2531 ();
 sg13g2_fill_1 FILLER_60_2538 ();
 sg13g2_decap_4 FILLER_60_2543 ();
 sg13g2_fill_2 FILLER_60_2551 ();
 sg13g2_fill_1 FILLER_60_2553 ();
 sg13g2_decap_4 FILLER_60_2564 ();
 sg13g2_decap_4 FILLER_60_2572 ();
 sg13g2_fill_1 FILLER_60_2580 ();
 sg13g2_decap_8 FILLER_60_2585 ();
 sg13g2_decap_8 FILLER_60_2592 ();
 sg13g2_decap_8 FILLER_60_2599 ();
 sg13g2_decap_8 FILLER_60_2606 ();
 sg13g2_decap_8 FILLER_60_2613 ();
 sg13g2_decap_4 FILLER_60_2620 ();
 sg13g2_fill_2 FILLER_60_2624 ();
 sg13g2_decap_4 FILLER_60_2666 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_fill_2 FILLER_61_7 ();
 sg13g2_fill_2 FILLER_61_45 ();
 sg13g2_fill_1 FILLER_61_47 ();
 sg13g2_fill_1 FILLER_61_53 ();
 sg13g2_fill_2 FILLER_61_64 ();
 sg13g2_decap_4 FILLER_61_76 ();
 sg13g2_fill_2 FILLER_61_80 ();
 sg13g2_decap_4 FILLER_61_87 ();
 sg13g2_fill_2 FILLER_61_91 ();
 sg13g2_decap_4 FILLER_61_103 ();
 sg13g2_decap_4 FILLER_61_120 ();
 sg13g2_fill_2 FILLER_61_124 ();
 sg13g2_decap_8 FILLER_61_153 ();
 sg13g2_decap_8 FILLER_61_164 ();
 sg13g2_fill_2 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_173 ();
 sg13g2_decap_4 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_201 ();
 sg13g2_decap_4 FILLER_61_208 ();
 sg13g2_fill_2 FILLER_61_238 ();
 sg13g2_decap_8 FILLER_61_245 ();
 sg13g2_decap_8 FILLER_61_252 ();
 sg13g2_decap_8 FILLER_61_259 ();
 sg13g2_fill_1 FILLER_61_266 ();
 sg13g2_fill_2 FILLER_61_315 ();
 sg13g2_decap_8 FILLER_61_321 ();
 sg13g2_fill_2 FILLER_61_328 ();
 sg13g2_fill_1 FILLER_61_330 ();
 sg13g2_decap_8 FILLER_61_334 ();
 sg13g2_fill_2 FILLER_61_341 ();
 sg13g2_fill_1 FILLER_61_385 ();
 sg13g2_fill_1 FILLER_61_412 ();
 sg13g2_fill_1 FILLER_61_444 ();
 sg13g2_fill_2 FILLER_61_450 ();
 sg13g2_fill_1 FILLER_61_452 ();
 sg13g2_fill_1 FILLER_61_511 ();
 sg13g2_decap_4 FILLER_61_517 ();
 sg13g2_decap_8 FILLER_61_560 ();
 sg13g2_decap_8 FILLER_61_567 ();
 sg13g2_decap_8 FILLER_61_574 ();
 sg13g2_fill_1 FILLER_61_581 ();
 sg13g2_fill_2 FILLER_61_595 ();
 sg13g2_decap_4 FILLER_61_604 ();
 sg13g2_fill_1 FILLER_61_613 ();
 sg13g2_fill_1 FILLER_61_618 ();
 sg13g2_fill_2 FILLER_61_632 ();
 sg13g2_fill_1 FILLER_61_634 ();
 sg13g2_fill_2 FILLER_61_640 ();
 sg13g2_fill_1 FILLER_61_642 ();
 sg13g2_decap_8 FILLER_61_660 ();
 sg13g2_fill_2 FILLER_61_667 ();
 sg13g2_fill_1 FILLER_61_674 ();
 sg13g2_decap_8 FILLER_61_681 ();
 sg13g2_decap_8 FILLER_61_688 ();
 sg13g2_decap_8 FILLER_61_695 ();
 sg13g2_decap_4 FILLER_61_702 ();
 sg13g2_decap_8 FILLER_61_712 ();
 sg13g2_decap_8 FILLER_61_719 ();
 sg13g2_decap_8 FILLER_61_726 ();
 sg13g2_fill_1 FILLER_61_733 ();
 sg13g2_fill_2 FILLER_61_748 ();
 sg13g2_fill_1 FILLER_61_750 ();
 sg13g2_decap_4 FILLER_61_755 ();
 sg13g2_fill_1 FILLER_61_759 ();
 sg13g2_decap_8 FILLER_61_794 ();
 sg13g2_decap_8 FILLER_61_806 ();
 sg13g2_decap_8 FILLER_61_813 ();
 sg13g2_fill_1 FILLER_61_820 ();
 sg13g2_decap_8 FILLER_61_839 ();
 sg13g2_fill_1 FILLER_61_846 ();
 sg13g2_fill_1 FILLER_61_856 ();
 sg13g2_fill_2 FILLER_61_894 ();
 sg13g2_fill_1 FILLER_61_896 ();
 sg13g2_decap_8 FILLER_61_913 ();
 sg13g2_decap_8 FILLER_61_970 ();
 sg13g2_decap_8 FILLER_61_977 ();
 sg13g2_decap_4 FILLER_61_984 ();
 sg13g2_decap_8 FILLER_61_993 ();
 sg13g2_decap_8 FILLER_61_1056 ();
 sg13g2_fill_1 FILLER_61_1063 ();
 sg13g2_decap_8 FILLER_61_1082 ();
 sg13g2_fill_2 FILLER_61_1093 ();
 sg13g2_fill_1 FILLER_61_1095 ();
 sg13g2_fill_2 FILLER_61_1108 ();
 sg13g2_decap_8 FILLER_61_1119 ();
 sg13g2_decap_4 FILLER_61_1126 ();
 sg13g2_fill_1 FILLER_61_1130 ();
 sg13g2_fill_1 FILLER_61_1134 ();
 sg13g2_decap_8 FILLER_61_1142 ();
 sg13g2_decap_8 FILLER_61_1149 ();
 sg13g2_decap_4 FILLER_61_1156 ();
 sg13g2_fill_2 FILLER_61_1172 ();
 sg13g2_fill_1 FILLER_61_1174 ();
 sg13g2_fill_1 FILLER_61_1190 ();
 sg13g2_fill_2 FILLER_61_1195 ();
 sg13g2_decap_4 FILLER_61_1203 ();
 sg13g2_fill_2 FILLER_61_1207 ();
 sg13g2_fill_2 FILLER_61_1235 ();
 sg13g2_fill_1 FILLER_61_1237 ();
 sg13g2_decap_8 FILLER_61_1243 ();
 sg13g2_decap_8 FILLER_61_1256 ();
 sg13g2_decap_8 FILLER_61_1263 ();
 sg13g2_fill_2 FILLER_61_1270 ();
 sg13g2_fill_1 FILLER_61_1272 ();
 sg13g2_decap_8 FILLER_61_1281 ();
 sg13g2_fill_2 FILLER_61_1288 ();
 sg13g2_fill_1 FILLER_61_1290 ();
 sg13g2_decap_4 FILLER_61_1321 ();
 sg13g2_fill_2 FILLER_61_1330 ();
 sg13g2_decap_8 FILLER_61_1338 ();
 sg13g2_decap_8 FILLER_61_1345 ();
 sg13g2_decap_4 FILLER_61_1352 ();
 sg13g2_fill_2 FILLER_61_1361 ();
 sg13g2_decap_8 FILLER_61_1420 ();
 sg13g2_decap_4 FILLER_61_1427 ();
 sg13g2_fill_1 FILLER_61_1431 ();
 sg13g2_decap_8 FILLER_61_1478 ();
 sg13g2_fill_2 FILLER_61_1485 ();
 sg13g2_fill_2 FILLER_61_1493 ();
 sg13g2_fill_2 FILLER_61_1532 ();
 sg13g2_decap_8 FILLER_61_1560 ();
 sg13g2_decap_8 FILLER_61_1589 ();
 sg13g2_fill_1 FILLER_61_1596 ();
 sg13g2_decap_8 FILLER_61_1602 ();
 sg13g2_decap_4 FILLER_61_1609 ();
 sg13g2_fill_2 FILLER_61_1613 ();
 sg13g2_fill_2 FILLER_61_1649 ();
 sg13g2_fill_1 FILLER_61_1651 ();
 sg13g2_fill_2 FILLER_61_1670 ();
 sg13g2_decap_4 FILLER_61_1683 ();
 sg13g2_fill_2 FILLER_61_1687 ();
 sg13g2_decap_4 FILLER_61_1696 ();
 sg13g2_fill_1 FILLER_61_1700 ();
 sg13g2_fill_2 FILLER_61_1713 ();
 sg13g2_fill_1 FILLER_61_1715 ();
 sg13g2_decap_8 FILLER_61_1725 ();
 sg13g2_decap_8 FILLER_61_1732 ();
 sg13g2_decap_8 FILLER_61_1739 ();
 sg13g2_decap_4 FILLER_61_1746 ();
 sg13g2_fill_1 FILLER_61_1750 ();
 sg13g2_decap_8 FILLER_61_1781 ();
 sg13g2_decap_4 FILLER_61_1788 ();
 sg13g2_decap_8 FILLER_61_1798 ();
 sg13g2_decap_8 FILLER_61_1810 ();
 sg13g2_decap_8 FILLER_61_1817 ();
 sg13g2_decap_8 FILLER_61_1824 ();
 sg13g2_fill_2 FILLER_61_1837 ();
 sg13g2_fill_1 FILLER_61_1847 ();
 sg13g2_fill_1 FILLER_61_1866 ();
 sg13g2_decap_8 FILLER_61_1889 ();
 sg13g2_fill_1 FILLER_61_1896 ();
 sg13g2_decap_8 FILLER_61_1911 ();
 sg13g2_fill_1 FILLER_61_1923 ();
 sg13g2_decap_4 FILLER_61_1950 ();
 sg13g2_fill_1 FILLER_61_1954 ();
 sg13g2_fill_1 FILLER_61_1960 ();
 sg13g2_fill_2 FILLER_61_1968 ();
 sg13g2_fill_2 FILLER_61_1980 ();
 sg13g2_fill_2 FILLER_61_1991 ();
 sg13g2_fill_2 FILLER_61_2012 ();
 sg13g2_fill_2 FILLER_61_2019 ();
 sg13g2_fill_2 FILLER_61_2047 ();
 sg13g2_fill_1 FILLER_61_2049 ();
 sg13g2_decap_4 FILLER_61_2167 ();
 sg13g2_fill_1 FILLER_61_2171 ();
 sg13g2_decap_8 FILLER_61_2176 ();
 sg13g2_decap_8 FILLER_61_2183 ();
 sg13g2_decap_8 FILLER_61_2190 ();
 sg13g2_fill_1 FILLER_61_2197 ();
 sg13g2_decap_4 FILLER_61_2209 ();
 sg13g2_decap_8 FILLER_61_2218 ();
 sg13g2_fill_1 FILLER_61_2225 ();
 sg13g2_decap_8 FILLER_61_2232 ();
 sg13g2_fill_1 FILLER_61_2239 ();
 sg13g2_fill_1 FILLER_61_2266 ();
 sg13g2_fill_1 FILLER_61_2271 ();
 sg13g2_fill_1 FILLER_61_2277 ();
 sg13g2_decap_8 FILLER_61_2310 ();
 sg13g2_decap_4 FILLER_61_2317 ();
 sg13g2_fill_2 FILLER_61_2321 ();
 sg13g2_decap_8 FILLER_61_2327 ();
 sg13g2_decap_8 FILLER_61_2334 ();
 sg13g2_decap_8 FILLER_61_2371 ();
 sg13g2_decap_4 FILLER_61_2378 ();
 sg13g2_decap_4 FILLER_61_2395 ();
 sg13g2_fill_2 FILLER_61_2399 ();
 sg13g2_fill_1 FILLER_61_2405 ();
 sg13g2_fill_1 FILLER_61_2410 ();
 sg13g2_decap_8 FILLER_61_2453 ();
 sg13g2_decap_8 FILLER_61_2460 ();
 sg13g2_decap_4 FILLER_61_2475 ();
 sg13g2_fill_2 FILLER_61_2479 ();
 sg13g2_fill_2 FILLER_61_2516 ();
 sg13g2_fill_1 FILLER_61_2518 ();
 sg13g2_decap_4 FILLER_61_2549 ();
 sg13g2_fill_2 FILLER_61_2591 ();
 sg13g2_fill_1 FILLER_61_2629 ();
 sg13g2_fill_1 FILLER_61_2642 ();
 sg13g2_decap_8 FILLER_61_2662 ();
 sg13g2_fill_1 FILLER_61_2669 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_4 FILLER_62_28 ();
 sg13g2_fill_1 FILLER_62_32 ();
 sg13g2_decap_8 FILLER_62_37 ();
 sg13g2_fill_2 FILLER_62_44 ();
 sg13g2_fill_1 FILLER_62_61 ();
 sg13g2_fill_1 FILLER_62_82 ();
 sg13g2_fill_2 FILLER_62_103 ();
 sg13g2_fill_1 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_115 ();
 sg13g2_decap_8 FILLER_62_122 ();
 sg13g2_fill_2 FILLER_62_137 ();
 sg13g2_fill_1 FILLER_62_139 ();
 sg13g2_fill_1 FILLER_62_145 ();
 sg13g2_decap_8 FILLER_62_151 ();
 sg13g2_decap_8 FILLER_62_158 ();
 sg13g2_decap_8 FILLER_62_165 ();
 sg13g2_decap_8 FILLER_62_172 ();
 sg13g2_decap_8 FILLER_62_179 ();
 sg13g2_fill_2 FILLER_62_186 ();
 sg13g2_decap_8 FILLER_62_201 ();
 sg13g2_decap_8 FILLER_62_208 ();
 sg13g2_fill_2 FILLER_62_215 ();
 sg13g2_fill_1 FILLER_62_217 ();
 sg13g2_fill_1 FILLER_62_223 ();
 sg13g2_fill_2 FILLER_62_236 ();
 sg13g2_fill_2 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_248 ();
 sg13g2_fill_2 FILLER_62_259 ();
 sg13g2_fill_1 FILLER_62_261 ();
 sg13g2_fill_2 FILLER_62_288 ();
 sg13g2_decap_8 FILLER_62_316 ();
 sg13g2_fill_2 FILLER_62_323 ();
 sg13g2_fill_1 FILLER_62_325 ();
 sg13g2_decap_8 FILLER_62_352 ();
 sg13g2_decap_4 FILLER_62_359 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_decap_8 FILLER_62_367 ();
 sg13g2_fill_2 FILLER_62_374 ();
 sg13g2_fill_2 FILLER_62_393 ();
 sg13g2_fill_2 FILLER_62_423 ();
 sg13g2_fill_2 FILLER_62_451 ();
 sg13g2_decap_8 FILLER_62_461 ();
 sg13g2_decap_8 FILLER_62_468 ();
 sg13g2_decap_8 FILLER_62_475 ();
 sg13g2_fill_1 FILLER_62_482 ();
 sg13g2_fill_2 FILLER_62_507 ();
 sg13g2_decap_8 FILLER_62_535 ();
 sg13g2_fill_2 FILLER_62_542 ();
 sg13g2_fill_1 FILLER_62_544 ();
 sg13g2_decap_4 FILLER_62_555 ();
 sg13g2_fill_1 FILLER_62_563 ();
 sg13g2_decap_4 FILLER_62_568 ();
 sg13g2_decap_8 FILLER_62_577 ();
 sg13g2_decap_8 FILLER_62_589 ();
 sg13g2_fill_1 FILLER_62_596 ();
 sg13g2_decap_4 FILLER_62_650 ();
 sg13g2_decap_4 FILLER_62_658 ();
 sg13g2_fill_1 FILLER_62_667 ();
 sg13g2_decap_8 FILLER_62_716 ();
 sg13g2_fill_1 FILLER_62_723 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_fill_2 FILLER_62_735 ();
 sg13g2_decap_4 FILLER_62_763 ();
 sg13g2_fill_1 FILLER_62_767 ();
 sg13g2_decap_8 FILLER_62_794 ();
 sg13g2_decap_8 FILLER_62_813 ();
 sg13g2_decap_8 FILLER_62_820 ();
 sg13g2_fill_2 FILLER_62_827 ();
 sg13g2_fill_1 FILLER_62_829 ();
 sg13g2_fill_2 FILLER_62_834 ();
 sg13g2_fill_1 FILLER_62_836 ();
 sg13g2_fill_1 FILLER_62_858 ();
 sg13g2_decap_8 FILLER_62_912 ();
 sg13g2_decap_8 FILLER_62_919 ();
 sg13g2_decap_4 FILLER_62_978 ();
 sg13g2_fill_1 FILLER_62_982 ();
 sg13g2_fill_2 FILLER_62_999 ();
 sg13g2_fill_1 FILLER_62_1001 ();
 sg13g2_fill_2 FILLER_62_1016 ();
 sg13g2_fill_1 FILLER_62_1032 ();
 sg13g2_fill_1 FILLER_62_1045 ();
 sg13g2_fill_2 FILLER_62_1076 ();
 sg13g2_fill_2 FILLER_62_1114 ();
 sg13g2_fill_2 FILLER_62_1177 ();
 sg13g2_fill_1 FILLER_62_1179 ();
 sg13g2_decap_4 FILLER_62_1211 ();
 sg13g2_fill_2 FILLER_62_1220 ();
 sg13g2_fill_1 FILLER_62_1222 ();
 sg13g2_fill_1 FILLER_62_1258 ();
 sg13g2_fill_2 FILLER_62_1285 ();
 sg13g2_fill_1 FILLER_62_1287 ();
 sg13g2_decap_8 FILLER_62_1292 ();
 sg13g2_fill_2 FILLER_62_1304 ();
 sg13g2_decap_4 FILLER_62_1310 ();
 sg13g2_decap_8 FILLER_62_1319 ();
 sg13g2_decap_8 FILLER_62_1326 ();
 sg13g2_decap_8 FILLER_62_1333 ();
 sg13g2_fill_2 FILLER_62_1340 ();
 sg13g2_fill_2 FILLER_62_1356 ();
 sg13g2_fill_1 FILLER_62_1358 ();
 sg13g2_decap_8 FILLER_62_1385 ();
 sg13g2_decap_4 FILLER_62_1392 ();
 sg13g2_fill_1 FILLER_62_1396 ();
 sg13g2_decap_4 FILLER_62_1411 ();
 sg13g2_decap_4 FILLER_62_1441 ();
 sg13g2_decap_4 FILLER_62_1450 ();
 sg13g2_decap_8 FILLER_62_1458 ();
 sg13g2_decap_8 FILLER_62_1470 ();
 sg13g2_fill_2 FILLER_62_1477 ();
 sg13g2_fill_1 FILLER_62_1483 ();
 sg13g2_fill_1 FILLER_62_1546 ();
 sg13g2_decap_4 FILLER_62_1573 ();
 sg13g2_fill_1 FILLER_62_1577 ();
 sg13g2_fill_2 FILLER_62_1608 ();
 sg13g2_decap_8 FILLER_62_1640 ();
 sg13g2_fill_1 FILLER_62_1703 ();
 sg13g2_fill_2 FILLER_62_1749 ();
 sg13g2_decap_8 FILLER_62_1765 ();
 sg13g2_decap_4 FILLER_62_1772 ();
 sg13g2_decap_8 FILLER_62_1780 ();
 sg13g2_decap_8 FILLER_62_1787 ();
 sg13g2_decap_8 FILLER_62_1794 ();
 sg13g2_decap_8 FILLER_62_1801 ();
 sg13g2_fill_2 FILLER_62_1833 ();
 sg13g2_fill_1 FILLER_62_1861 ();
 sg13g2_fill_1 FILLER_62_1866 ();
 sg13g2_fill_2 FILLER_62_1871 ();
 sg13g2_fill_1 FILLER_62_1873 ();
 sg13g2_decap_4 FILLER_62_1892 ();
 sg13g2_decap_8 FILLER_62_1902 ();
 sg13g2_fill_2 FILLER_62_1909 ();
 sg13g2_fill_1 FILLER_62_1911 ();
 sg13g2_fill_2 FILLER_62_1940 ();
 sg13g2_fill_1 FILLER_62_1942 ();
 sg13g2_fill_1 FILLER_62_1960 ();
 sg13g2_fill_1 FILLER_62_1966 ();
 sg13g2_fill_1 FILLER_62_1972 ();
 sg13g2_fill_2 FILLER_62_2050 ();
 sg13g2_fill_1 FILLER_62_2102 ();
 sg13g2_fill_2 FILLER_62_2121 ();
 sg13g2_decap_8 FILLER_62_2140 ();
 sg13g2_fill_2 FILLER_62_2147 ();
 sg13g2_fill_2 FILLER_62_2168 ();
 sg13g2_fill_1 FILLER_62_2170 ();
 sg13g2_decap_4 FILLER_62_2176 ();
 sg13g2_fill_1 FILLER_62_2186 ();
 sg13g2_fill_2 FILLER_62_2213 ();
 sg13g2_fill_2 FILLER_62_2241 ();
 sg13g2_decap_4 FILLER_62_2268 ();
 sg13g2_fill_2 FILLER_62_2272 ();
 sg13g2_decap_8 FILLER_62_2280 ();
 sg13g2_decap_8 FILLER_62_2287 ();
 sg13g2_fill_2 FILLER_62_2294 ();
 sg13g2_decap_8 FILLER_62_2299 ();
 sg13g2_fill_2 FILLER_62_2306 ();
 sg13g2_fill_1 FILLER_62_2308 ();
 sg13g2_fill_2 FILLER_62_2315 ();
 sg13g2_fill_2 FILLER_62_2323 ();
 sg13g2_fill_1 FILLER_62_2325 ();
 sg13g2_decap_8 FILLER_62_2378 ();
 sg13g2_decap_8 FILLER_62_2385 ();
 sg13g2_decap_8 FILLER_62_2392 ();
 sg13g2_decap_8 FILLER_62_2399 ();
 sg13g2_decap_8 FILLER_62_2406 ();
 sg13g2_fill_2 FILLER_62_2413 ();
 sg13g2_fill_1 FILLER_62_2415 ();
 sg13g2_fill_2 FILLER_62_2464 ();
 sg13g2_fill_1 FILLER_62_2466 ();
 sg13g2_fill_2 FILLER_62_2470 ();
 sg13g2_fill_1 FILLER_62_2472 ();
 sg13g2_decap_4 FILLER_62_2477 ();
 sg13g2_fill_1 FILLER_62_2481 ();
 sg13g2_fill_2 FILLER_62_2494 ();
 sg13g2_fill_1 FILLER_62_2496 ();
 sg13g2_fill_2 FILLER_62_2501 ();
 sg13g2_decap_8 FILLER_62_2507 ();
 sg13g2_decap_8 FILLER_62_2514 ();
 sg13g2_decap_4 FILLER_62_2521 ();
 sg13g2_fill_2 FILLER_62_2525 ();
 sg13g2_fill_2 FILLER_62_2553 ();
 sg13g2_fill_1 FILLER_62_2555 ();
 sg13g2_fill_2 FILLER_62_2627 ();
 sg13g2_decap_8 FILLER_62_2637 ();
 sg13g2_decap_8 FILLER_62_2644 ();
 sg13g2_decap_8 FILLER_62_2651 ();
 sg13g2_decap_8 FILLER_62_2658 ();
 sg13g2_decap_4 FILLER_62_2665 ();
 sg13g2_fill_1 FILLER_62_2669 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_4 FILLER_63_14 ();
 sg13g2_decap_4 FILLER_63_28 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_decap_8 FILLER_63_38 ();
 sg13g2_decap_8 FILLER_63_45 ();
 sg13g2_decap_4 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_56 ();
 sg13g2_fill_2 FILLER_63_87 ();
 sg13g2_fill_1 FILLER_63_99 ();
 sg13g2_fill_1 FILLER_63_104 ();
 sg13g2_fill_1 FILLER_63_110 ();
 sg13g2_fill_2 FILLER_63_121 ();
 sg13g2_decap_8 FILLER_63_128 ();
 sg13g2_fill_2 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_137 ();
 sg13g2_decap_8 FILLER_63_142 ();
 sg13g2_decap_8 FILLER_63_149 ();
 sg13g2_decap_4 FILLER_63_171 ();
 sg13g2_decap_4 FILLER_63_185 ();
 sg13g2_fill_2 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_230 ();
 sg13g2_decap_8 FILLER_63_236 ();
 sg13g2_decap_8 FILLER_63_243 ();
 sg13g2_decap_8 FILLER_63_250 ();
 sg13g2_decap_8 FILLER_63_257 ();
 sg13g2_decap_4 FILLER_63_264 ();
 sg13g2_decap_8 FILLER_63_304 ();
 sg13g2_decap_8 FILLER_63_311 ();
 sg13g2_decap_8 FILLER_63_318 ();
 sg13g2_decap_8 FILLER_63_325 ();
 sg13g2_decap_8 FILLER_63_332 ();
 sg13g2_decap_8 FILLER_63_339 ();
 sg13g2_decap_8 FILLER_63_346 ();
 sg13g2_decap_8 FILLER_63_353 ();
 sg13g2_decap_8 FILLER_63_360 ();
 sg13g2_decap_8 FILLER_63_367 ();
 sg13g2_decap_4 FILLER_63_378 ();
 sg13g2_fill_1 FILLER_63_390 ();
 sg13g2_fill_2 FILLER_63_424 ();
 sg13g2_fill_1 FILLER_63_444 ();
 sg13g2_fill_2 FILLER_63_459 ();
 sg13g2_decap_8 FILLER_63_466 ();
 sg13g2_decap_8 FILLER_63_473 ();
 sg13g2_fill_2 FILLER_63_480 ();
 sg13g2_decap_8 FILLER_63_518 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_fill_2 FILLER_63_539 ();
 sg13g2_fill_1 FILLER_63_541 ();
 sg13g2_decap_8 FILLER_63_594 ();
 sg13g2_decap_4 FILLER_63_601 ();
 sg13g2_fill_2 FILLER_63_609 ();
 sg13g2_decap_4 FILLER_63_636 ();
 sg13g2_fill_1 FILLER_63_640 ();
 sg13g2_decap_8 FILLER_63_661 ();
 sg13g2_decap_8 FILLER_63_668 ();
 sg13g2_fill_2 FILLER_63_675 ();
 sg13g2_fill_1 FILLER_63_677 ();
 sg13g2_fill_2 FILLER_63_704 ();
 sg13g2_decap_8 FILLER_63_732 ();
 sg13g2_decap_8 FILLER_63_748 ();
 sg13g2_decap_8 FILLER_63_755 ();
 sg13g2_fill_1 FILLER_63_762 ();
 sg13g2_fill_1 FILLER_63_772 ();
 sg13g2_fill_2 FILLER_63_808 ();
 sg13g2_decap_8 FILLER_63_816 ();
 sg13g2_fill_2 FILLER_63_823 ();
 sg13g2_fill_2 FILLER_63_830 ();
 sg13g2_fill_1 FILLER_63_832 ();
 sg13g2_fill_1 FILLER_63_873 ();
 sg13g2_fill_1 FILLER_63_909 ();
 sg13g2_fill_1 FILLER_63_936 ();
 sg13g2_fill_2 FILLER_63_968 ();
 sg13g2_fill_2 FILLER_63_1054 ();
 sg13g2_fill_1 FILLER_63_1056 ();
 sg13g2_fill_2 FILLER_63_1060 ();
 sg13g2_fill_1 FILLER_63_1062 ();
 sg13g2_decap_8 FILLER_63_1072 ();
 sg13g2_decap_4 FILLER_63_1079 ();
 sg13g2_fill_2 FILLER_63_1083 ();
 sg13g2_decap_8 FILLER_63_1121 ();
 sg13g2_fill_2 FILLER_63_1128 ();
 sg13g2_fill_1 FILLER_63_1130 ();
 sg13g2_fill_1 FILLER_63_1157 ();
 sg13g2_fill_1 FILLER_63_1164 ();
 sg13g2_fill_1 FILLER_63_1174 ();
 sg13g2_decap_8 FILLER_63_1214 ();
 sg13g2_decap_8 FILLER_63_1221 ();
 sg13g2_fill_2 FILLER_63_1228 ();
 sg13g2_fill_1 FILLER_63_1230 ();
 sg13g2_decap_4 FILLER_63_1236 ();
 sg13g2_decap_8 FILLER_63_1278 ();
 sg13g2_decap_8 FILLER_63_1285 ();
 sg13g2_decap_8 FILLER_63_1292 ();
 sg13g2_decap_8 FILLER_63_1299 ();
 sg13g2_decap_8 FILLER_63_1306 ();
 sg13g2_fill_2 FILLER_63_1313 ();
 sg13g2_fill_1 FILLER_63_1315 ();
 sg13g2_fill_2 FILLER_63_1342 ();
 sg13g2_fill_1 FILLER_63_1344 ();
 sg13g2_decap_8 FILLER_63_1371 ();
 sg13g2_decap_4 FILLER_63_1378 ();
 sg13g2_fill_1 FILLER_63_1382 ();
 sg13g2_decap_8 FILLER_63_1389 ();
 sg13g2_decap_4 FILLER_63_1396 ();
 sg13g2_decap_8 FILLER_63_1419 ();
 sg13g2_decap_8 FILLER_63_1426 ();
 sg13g2_decap_8 FILLER_63_1442 ();
 sg13g2_decap_8 FILLER_63_1449 ();
 sg13g2_decap_4 FILLER_63_1456 ();
 sg13g2_fill_2 FILLER_63_1494 ();
 sg13g2_fill_2 FILLER_63_1509 ();
 sg13g2_decap_8 FILLER_63_1562 ();
 sg13g2_decap_8 FILLER_63_1569 ();
 sg13g2_decap_8 FILLER_63_1576 ();
 sg13g2_decap_8 FILLER_63_1583 ();
 sg13g2_decap_8 FILLER_63_1590 ();
 sg13g2_decap_8 FILLER_63_1597 ();
 sg13g2_decap_8 FILLER_63_1604 ();
 sg13g2_fill_2 FILLER_63_1611 ();
 sg13g2_fill_1 FILLER_63_1613 ();
 sg13g2_decap_8 FILLER_63_1629 ();
 sg13g2_fill_1 FILLER_63_1636 ();
 sg13g2_decap_8 FILLER_63_1658 ();
 sg13g2_fill_2 FILLER_63_1665 ();
 sg13g2_decap_4 FILLER_63_1670 ();
 sg13g2_fill_2 FILLER_63_1713 ();
 sg13g2_fill_1 FILLER_63_1715 ();
 sg13g2_fill_2 FILLER_63_1721 ();
 sg13g2_fill_2 FILLER_63_1733 ();
 sg13g2_fill_1 FILLER_63_1735 ();
 sg13g2_decap_4 FILLER_63_1754 ();
 sg13g2_decap_4 FILLER_63_1763 ();
 sg13g2_fill_1 FILLER_63_1767 ();
 sg13g2_decap_8 FILLER_63_1794 ();
 sg13g2_fill_1 FILLER_63_1801 ();
 sg13g2_decap_4 FILLER_63_1833 ();
 sg13g2_decap_4 FILLER_63_1845 ();
 sg13g2_fill_1 FILLER_63_1849 ();
 sg13g2_fill_2 FILLER_63_1854 ();
 sg13g2_decap_4 FILLER_63_1876 ();
 sg13g2_decap_8 FILLER_63_1892 ();
 sg13g2_fill_1 FILLER_63_1899 ();
 sg13g2_decap_8 FILLER_63_1905 ();
 sg13g2_fill_2 FILLER_63_1917 ();
 sg13g2_fill_2 FILLER_63_1945 ();
 sg13g2_fill_1 FILLER_63_1947 ();
 sg13g2_fill_1 FILLER_63_1954 ();
 sg13g2_fill_2 FILLER_63_1964 ();
 sg13g2_decap_4 FILLER_63_1977 ();
 sg13g2_fill_2 FILLER_63_1981 ();
 sg13g2_decap_8 FILLER_63_2015 ();
 sg13g2_decap_8 FILLER_63_2022 ();
 sg13g2_decap_4 FILLER_63_2029 ();
 sg13g2_fill_2 FILLER_63_2033 ();
 sg13g2_decap_4 FILLER_63_2061 ();
 sg13g2_fill_2 FILLER_63_2100 ();
 sg13g2_fill_1 FILLER_63_2102 ();
 sg13g2_fill_2 FILLER_63_2109 ();
 sg13g2_fill_1 FILLER_63_2111 ();
 sg13g2_decap_4 FILLER_63_2152 ();
 sg13g2_fill_2 FILLER_63_2164 ();
 sg13g2_fill_2 FILLER_63_2170 ();
 sg13g2_fill_1 FILLER_63_2172 ();
 sg13g2_fill_1 FILLER_63_2178 ();
 sg13g2_fill_2 FILLER_63_2183 ();
 sg13g2_fill_1 FILLER_63_2251 ();
 sg13g2_decap_8 FILLER_63_2267 ();
 sg13g2_decap_4 FILLER_63_2274 ();
 sg13g2_fill_1 FILLER_63_2278 ();
 sg13g2_fill_2 FILLER_63_2287 ();
 sg13g2_fill_1 FILLER_63_2289 ();
 sg13g2_fill_2 FILLER_63_2299 ();
 sg13g2_decap_8 FILLER_63_2341 ();
 sg13g2_fill_1 FILLER_63_2348 ();
 sg13g2_decap_4 FILLER_63_2357 ();
 sg13g2_fill_2 FILLER_63_2361 ();
 sg13g2_decap_8 FILLER_63_2367 ();
 sg13g2_decap_4 FILLER_63_2374 ();
 sg13g2_decap_8 FILLER_63_2384 ();
 sg13g2_decap_8 FILLER_63_2508 ();
 sg13g2_fill_1 FILLER_63_2515 ();
 sg13g2_decap_8 FILLER_63_2553 ();
 sg13g2_decap_8 FILLER_63_2560 ();
 sg13g2_decap_8 FILLER_63_2567 ();
 sg13g2_decap_8 FILLER_63_2574 ();
 sg13g2_decap_8 FILLER_63_2581 ();
 sg13g2_fill_1 FILLER_63_2588 ();
 sg13g2_decap_8 FILLER_63_2593 ();
 sg13g2_fill_1 FILLER_63_2604 ();
 sg13g2_fill_2 FILLER_63_2609 ();
 sg13g2_fill_2 FILLER_63_2616 ();
 sg13g2_fill_2 FILLER_63_2626 ();
 sg13g2_decap_8 FILLER_63_2633 ();
 sg13g2_decap_8 FILLER_63_2640 ();
 sg13g2_decap_8 FILLER_63_2647 ();
 sg13g2_decap_8 FILLER_63_2654 ();
 sg13g2_decap_8 FILLER_63_2661 ();
 sg13g2_fill_2 FILLER_63_2668 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_fill_2 FILLER_64_18 ();
 sg13g2_decap_8 FILLER_64_50 ();
 sg13g2_fill_2 FILLER_64_57 ();
 sg13g2_fill_1 FILLER_64_59 ();
 sg13g2_decap_4 FILLER_64_80 ();
 sg13g2_decap_8 FILLER_64_94 ();
 sg13g2_fill_2 FILLER_64_101 ();
 sg13g2_fill_1 FILLER_64_103 ();
 sg13g2_decap_4 FILLER_64_109 ();
 sg13g2_fill_1 FILLER_64_113 ();
 sg13g2_decap_8 FILLER_64_133 ();
 sg13g2_decap_4 FILLER_64_149 ();
 sg13g2_fill_2 FILLER_64_153 ();
 sg13g2_decap_4 FILLER_64_167 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_decap_4 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_202 ();
 sg13g2_fill_2 FILLER_64_208 ();
 sg13g2_fill_1 FILLER_64_210 ();
 sg13g2_decap_8 FILLER_64_247 ();
 sg13g2_decap_8 FILLER_64_254 ();
 sg13g2_decap_8 FILLER_64_261 ();
 sg13g2_decap_8 FILLER_64_268 ();
 sg13g2_decap_8 FILLER_64_275 ();
 sg13g2_decap_8 FILLER_64_282 ();
 sg13g2_decap_8 FILLER_64_299 ();
 sg13g2_decap_8 FILLER_64_306 ();
 sg13g2_decap_8 FILLER_64_313 ();
 sg13g2_decap_8 FILLER_64_320 ();
 sg13g2_decap_8 FILLER_64_327 ();
 sg13g2_decap_8 FILLER_64_334 ();
 sg13g2_decap_4 FILLER_64_341 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_fill_2 FILLER_64_381 ();
 sg13g2_fill_1 FILLER_64_383 ();
 sg13g2_fill_2 FILLER_64_392 ();
 sg13g2_decap_8 FILLER_64_448 ();
 sg13g2_fill_1 FILLER_64_455 ();
 sg13g2_decap_4 FILLER_64_460 ();
 sg13g2_fill_1 FILLER_64_464 ();
 sg13g2_fill_1 FILLER_64_468 ();
 sg13g2_fill_1 FILLER_64_476 ();
 sg13g2_fill_2 FILLER_64_481 ();
 sg13g2_decap_8 FILLER_64_493 ();
 sg13g2_decap_4 FILLER_64_500 ();
 sg13g2_fill_2 FILLER_64_504 ();
 sg13g2_fill_1 FILLER_64_511 ();
 sg13g2_decap_4 FILLER_64_518 ();
 sg13g2_decap_8 FILLER_64_525 ();
 sg13g2_decap_8 FILLER_64_532 ();
 sg13g2_decap_8 FILLER_64_539 ();
 sg13g2_decap_8 FILLER_64_546 ();
 sg13g2_decap_4 FILLER_64_553 ();
 sg13g2_decap_8 FILLER_64_587 ();
 sg13g2_decap_8 FILLER_64_594 ();
 sg13g2_decap_8 FILLER_64_601 ();
 sg13g2_fill_2 FILLER_64_608 ();
 sg13g2_fill_1 FILLER_64_610 ();
 sg13g2_decap_4 FILLER_64_618 ();
 sg13g2_fill_2 FILLER_64_625 ();
 sg13g2_fill_1 FILLER_64_627 ();
 sg13g2_decap_8 FILLER_64_675 ();
 sg13g2_decap_8 FILLER_64_682 ();
 sg13g2_decap_4 FILLER_64_689 ();
 sg13g2_fill_1 FILLER_64_723 ();
 sg13g2_fill_2 FILLER_64_776 ();
 sg13g2_fill_1 FILLER_64_778 ();
 sg13g2_fill_2 FILLER_64_784 ();
 sg13g2_decap_4 FILLER_64_816 ();
 sg13g2_fill_2 FILLER_64_820 ();
 sg13g2_fill_1 FILLER_64_857 ();
 sg13g2_fill_2 FILLER_64_874 ();
 sg13g2_fill_2 FILLER_64_885 ();
 sg13g2_decap_8 FILLER_64_893 ();
 sg13g2_fill_1 FILLER_64_900 ();
 sg13g2_decap_8 FILLER_64_907 ();
 sg13g2_decap_8 FILLER_64_914 ();
 sg13g2_decap_8 FILLER_64_921 ();
 sg13g2_fill_1 FILLER_64_931 ();
 sg13g2_decap_8 FILLER_64_949 ();
 sg13g2_decap_8 FILLER_64_956 ();
 sg13g2_fill_2 FILLER_64_966 ();
 sg13g2_fill_1 FILLER_64_968 ();
 sg13g2_fill_1 FILLER_64_998 ();
 sg13g2_fill_1 FILLER_64_1039 ();
 sg13g2_decap_4 FILLER_64_1053 ();
 sg13g2_fill_1 FILLER_64_1062 ();
 sg13g2_decap_8 FILLER_64_1073 ();
 sg13g2_fill_1 FILLER_64_1080 ();
 sg13g2_fill_1 FILLER_64_1120 ();
 sg13g2_fill_2 FILLER_64_1156 ();
 sg13g2_decap_4 FILLER_64_1172 ();
 sg13g2_fill_1 FILLER_64_1176 ();
 sg13g2_decap_4 FILLER_64_1207 ();
 sg13g2_fill_2 FILLER_64_1211 ();
 sg13g2_fill_2 FILLER_64_1239 ();
 sg13g2_fill_1 FILLER_64_1241 ();
 sg13g2_decap_8 FILLER_64_1246 ();
 sg13g2_decap_4 FILLER_64_1253 ();
 sg13g2_decap_8 FILLER_64_1285 ();
 sg13g2_decap_8 FILLER_64_1292 ();
 sg13g2_decap_8 FILLER_64_1299 ();
 sg13g2_decap_8 FILLER_64_1306 ();
 sg13g2_fill_2 FILLER_64_1313 ();
 sg13g2_decap_8 FILLER_64_1324 ();
 sg13g2_decap_8 FILLER_64_1331 ();
 sg13g2_decap_8 FILLER_64_1338 ();
 sg13g2_fill_2 FILLER_64_1350 ();
 sg13g2_decap_8 FILLER_64_1389 ();
 sg13g2_decap_8 FILLER_64_1396 ();
 sg13g2_decap_4 FILLER_64_1408 ();
 sg13g2_fill_1 FILLER_64_1412 ();
 sg13g2_decap_4 FILLER_64_1427 ();
 sg13g2_fill_2 FILLER_64_1431 ();
 sg13g2_decap_4 FILLER_64_1468 ();
 sg13g2_fill_1 FILLER_64_1495 ();
 sg13g2_fill_1 FILLER_64_1522 ();
 sg13g2_fill_1 FILLER_64_1530 ();
 sg13g2_fill_1 FILLER_64_1548 ();
 sg13g2_decap_4 FILLER_64_1553 ();
 sg13g2_decap_8 FILLER_64_1583 ();
 sg13g2_decap_8 FILLER_64_1590 ();
 sg13g2_decap_4 FILLER_64_1597 ();
 sg13g2_fill_1 FILLER_64_1601 ();
 sg13g2_decap_4 FILLER_64_1623 ();
 sg13g2_fill_2 FILLER_64_1627 ();
 sg13g2_decap_8 FILLER_64_1638 ();
 sg13g2_fill_1 FILLER_64_1645 ();
 sg13g2_decap_8 FILLER_64_1649 ();
 sg13g2_decap_4 FILLER_64_1656 ();
 sg13g2_fill_1 FILLER_64_1673 ();
 sg13g2_fill_2 FILLER_64_1715 ();
 sg13g2_fill_2 FILLER_64_1757 ();
 sg13g2_fill_2 FILLER_64_1789 ();
 sg13g2_fill_2 FILLER_64_1822 ();
 sg13g2_fill_2 FILLER_64_1827 ();
 sg13g2_fill_1 FILLER_64_1829 ();
 sg13g2_fill_1 FILLER_64_1850 ();
 sg13g2_fill_2 FILLER_64_1855 ();
 sg13g2_fill_1 FILLER_64_1857 ();
 sg13g2_fill_2 FILLER_64_1870 ();
 sg13g2_decap_8 FILLER_64_1877 ();
 sg13g2_decap_4 FILLER_64_1884 ();
 sg13g2_fill_2 FILLER_64_1888 ();
 sg13g2_fill_1 FILLER_64_1918 ();
 sg13g2_fill_1 FILLER_64_1928 ();
 sg13g2_fill_1 FILLER_64_1935 ();
 sg13g2_decap_4 FILLER_64_1941 ();
 sg13g2_fill_1 FILLER_64_1945 ();
 sg13g2_decap_8 FILLER_64_1955 ();
 sg13g2_decap_8 FILLER_64_1962 ();
 sg13g2_decap_8 FILLER_64_1969 ();
 sg13g2_decap_4 FILLER_64_1976 ();
 sg13g2_fill_1 FILLER_64_1980 ();
 sg13g2_fill_1 FILLER_64_2005 ();
 sg13g2_decap_8 FILLER_64_2010 ();
 sg13g2_decap_8 FILLER_64_2017 ();
 sg13g2_decap_4 FILLER_64_2027 ();
 sg13g2_decap_4 FILLER_64_2036 ();
 sg13g2_fill_2 FILLER_64_2050 ();
 sg13g2_fill_2 FILLER_64_2058 ();
 sg13g2_fill_2 FILLER_64_2066 ();
 sg13g2_fill_1 FILLER_64_2068 ();
 sg13g2_fill_2 FILLER_64_2072 ();
 sg13g2_fill_1 FILLER_64_2074 ();
 sg13g2_decap_4 FILLER_64_2090 ();
 sg13g2_decap_8 FILLER_64_2098 ();
 sg13g2_decap_8 FILLER_64_2105 ();
 sg13g2_decap_4 FILLER_64_2112 ();
 sg13g2_fill_1 FILLER_64_2116 ();
 sg13g2_fill_1 FILLER_64_2146 ();
 sg13g2_fill_2 FILLER_64_2159 ();
 sg13g2_fill_1 FILLER_64_2161 ();
 sg13g2_decap_4 FILLER_64_2188 ();
 sg13g2_fill_2 FILLER_64_2192 ();
 sg13g2_decap_8 FILLER_64_2198 ();
 sg13g2_fill_1 FILLER_64_2205 ();
 sg13g2_fill_2 FILLER_64_2211 ();
 sg13g2_fill_1 FILLER_64_2244 ();
 sg13g2_fill_1 FILLER_64_2254 ();
 sg13g2_fill_2 FILLER_64_2281 ();
 sg13g2_fill_1 FILLER_64_2283 ();
 sg13g2_decap_4 FILLER_64_2290 ();
 sg13g2_fill_2 FILLER_64_2294 ();
 sg13g2_decap_8 FILLER_64_2308 ();
 sg13g2_decap_4 FILLER_64_2315 ();
 sg13g2_fill_1 FILLER_64_2319 ();
 sg13g2_fill_2 FILLER_64_2324 ();
 sg13g2_decap_8 FILLER_64_2360 ();
 sg13g2_decap_8 FILLER_64_2367 ();
 sg13g2_decap_8 FILLER_64_2374 ();
 sg13g2_fill_2 FILLER_64_2381 ();
 sg13g2_fill_1 FILLER_64_2383 ();
 sg13g2_decap_8 FILLER_64_2418 ();
 sg13g2_decap_8 FILLER_64_2425 ();
 sg13g2_decap_4 FILLER_64_2432 ();
 sg13g2_fill_1 FILLER_64_2440 ();
 sg13g2_fill_2 FILLER_64_2470 ();
 sg13g2_fill_1 FILLER_64_2476 ();
 sg13g2_fill_1 FILLER_64_2509 ();
 sg13g2_fill_2 FILLER_64_2514 ();
 sg13g2_fill_2 FILLER_64_2528 ();
 sg13g2_fill_2 FILLER_64_2534 ();
 sg13g2_fill_2 FILLER_64_2540 ();
 sg13g2_decap_8 FILLER_64_2546 ();
 sg13g2_decap_4 FILLER_64_2553 ();
 sg13g2_fill_2 FILLER_64_2557 ();
 sg13g2_fill_2 FILLER_64_2610 ();
 sg13g2_decap_8 FILLER_64_2638 ();
 sg13g2_fill_1 FILLER_64_2645 ();
 sg13g2_decap_8 FILLER_64_2659 ();
 sg13g2_decap_4 FILLER_64_2666 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_fill_2 FILLER_65_14 ();
 sg13g2_decap_4 FILLER_65_46 ();
 sg13g2_fill_2 FILLER_65_50 ();
 sg13g2_decap_4 FILLER_65_62 ();
 sg13g2_fill_2 FILLER_65_189 ();
 sg13g2_fill_1 FILLER_65_191 ();
 sg13g2_decap_8 FILLER_65_202 ();
 sg13g2_fill_1 FILLER_65_209 ();
 sg13g2_fill_2 FILLER_65_220 ();
 sg13g2_decap_8 FILLER_65_227 ();
 sg13g2_decap_4 FILLER_65_234 ();
 sg13g2_fill_1 FILLER_65_238 ();
 sg13g2_decap_4 FILLER_65_249 ();
 sg13g2_decap_4 FILLER_65_279 ();
 sg13g2_fill_1 FILLER_65_283 ();
 sg13g2_decap_8 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_decap_4 FILLER_65_331 ();
 sg13g2_fill_2 FILLER_65_335 ();
 sg13g2_fill_1 FILLER_65_340 ();
 sg13g2_decap_8 FILLER_65_347 ();
 sg13g2_fill_2 FILLER_65_354 ();
 sg13g2_decap_8 FILLER_65_359 ();
 sg13g2_fill_2 FILLER_65_366 ();
 sg13g2_fill_1 FILLER_65_368 ();
 sg13g2_decap_8 FILLER_65_374 ();
 sg13g2_decap_8 FILLER_65_381 ();
 sg13g2_decap_8 FILLER_65_388 ();
 sg13g2_decap_4 FILLER_65_395 ();
 sg13g2_fill_1 FILLER_65_399 ();
 sg13g2_decap_4 FILLER_65_408 ();
 sg13g2_fill_2 FILLER_65_412 ();
 sg13g2_fill_2 FILLER_65_419 ();
 sg13g2_decap_8 FILLER_65_443 ();
 sg13g2_decap_4 FILLER_65_450 ();
 sg13g2_decap_8 FILLER_65_459 ();
 sg13g2_decap_8 FILLER_65_466 ();
 sg13g2_fill_2 FILLER_65_473 ();
 sg13g2_fill_1 FILLER_65_475 ();
 sg13g2_fill_2 FILLER_65_479 ();
 sg13g2_fill_2 FILLER_65_507 ();
 sg13g2_fill_1 FILLER_65_514 ();
 sg13g2_decap_4 FILLER_65_593 ();
 sg13g2_fill_2 FILLER_65_597 ();
 sg13g2_fill_1 FILLER_65_604 ();
 sg13g2_fill_2 FILLER_65_611 ();
 sg13g2_fill_1 FILLER_65_613 ();
 sg13g2_fill_2 FILLER_65_619 ();
 sg13g2_fill_1 FILLER_65_621 ();
 sg13g2_decap_4 FILLER_65_674 ();
 sg13g2_fill_1 FILLER_65_678 ();
 sg13g2_decap_8 FILLER_65_687 ();
 sg13g2_decap_8 FILLER_65_694 ();
 sg13g2_decap_8 FILLER_65_701 ();
 sg13g2_decap_4 FILLER_65_708 ();
 sg13g2_fill_2 FILLER_65_712 ();
 sg13g2_decap_8 FILLER_65_724 ();
 sg13g2_decap_8 FILLER_65_731 ();
 sg13g2_decap_8 FILLER_65_738 ();
 sg13g2_fill_2 FILLER_65_745 ();
 sg13g2_fill_2 FILLER_65_752 ();
 sg13g2_decap_8 FILLER_65_759 ();
 sg13g2_decap_8 FILLER_65_766 ();
 sg13g2_decap_8 FILLER_65_773 ();
 sg13g2_decap_4 FILLER_65_780 ();
 sg13g2_fill_1 FILLER_65_793 ();
 sg13g2_fill_1 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_808 ();
 sg13g2_fill_1 FILLER_65_841 ();
 sg13g2_fill_2 FILLER_65_872 ();
 sg13g2_fill_2 FILLER_65_882 ();
 sg13g2_decap_8 FILLER_65_892 ();
 sg13g2_fill_2 FILLER_65_899 ();
 sg13g2_decap_8 FILLER_65_905 ();
 sg13g2_decap_8 FILLER_65_912 ();
 sg13g2_decap_4 FILLER_65_919 ();
 sg13g2_fill_1 FILLER_65_923 ();
 sg13g2_fill_2 FILLER_65_952 ();
 sg13g2_fill_1 FILLER_65_954 ();
 sg13g2_fill_2 FILLER_65_959 ();
 sg13g2_fill_2 FILLER_65_993 ();
 sg13g2_fill_1 FILLER_65_1000 ();
 sg13g2_decap_8 FILLER_65_1006 ();
 sg13g2_decap_8 FILLER_65_1013 ();
 sg13g2_fill_1 FILLER_65_1020 ();
 sg13g2_fill_1 FILLER_65_1024 ();
 sg13g2_fill_1 FILLER_65_1028 ();
 sg13g2_fill_2 FILLER_65_1063 ();
 sg13g2_fill_1 FILLER_65_1065 ();
 sg13g2_fill_1 FILLER_65_1128 ();
 sg13g2_decap_8 FILLER_65_1181 ();
 sg13g2_fill_2 FILLER_65_1188 ();
 sg13g2_fill_2 FILLER_65_1205 ();
 sg13g2_decap_4 FILLER_65_1215 ();
 sg13g2_decap_8 FILLER_65_1223 ();
 sg13g2_fill_1 FILLER_65_1230 ();
 sg13g2_fill_1 FILLER_65_1282 ();
 sg13g2_fill_1 FILLER_65_1291 ();
 sg13g2_fill_1 FILLER_65_1297 ();
 sg13g2_decap_8 FILLER_65_1304 ();
 sg13g2_fill_1 FILLER_65_1311 ();
 sg13g2_decap_8 FILLER_65_1338 ();
 sg13g2_fill_1 FILLER_65_1345 ();
 sg13g2_fill_2 FILLER_65_1385 ();
 sg13g2_decap_4 FILLER_65_1413 ();
 sg13g2_decap_4 FILLER_65_1443 ();
 sg13g2_decap_8 FILLER_65_1453 ();
 sg13g2_decap_8 FILLER_65_1460 ();
 sg13g2_fill_2 FILLER_65_1467 ();
 sg13g2_fill_1 FILLER_65_1469 ();
 sg13g2_fill_2 FILLER_65_1486 ();
 sg13g2_fill_2 FILLER_65_1494 ();
 sg13g2_fill_1 FILLER_65_1514 ();
 sg13g2_fill_2 FILLER_65_1520 ();
 sg13g2_fill_2 FILLER_65_1542 ();
 sg13g2_fill_2 FILLER_65_1570 ();
 sg13g2_fill_1 FILLER_65_1572 ();
 sg13g2_decap_8 FILLER_65_1581 ();
 sg13g2_fill_1 FILLER_65_1588 ();
 sg13g2_fill_2 FILLER_65_1628 ();
 sg13g2_fill_2 FILLER_65_1635 ();
 sg13g2_fill_1 FILLER_65_1637 ();
 sg13g2_fill_2 FILLER_65_1725 ();
 sg13g2_fill_1 FILLER_65_1758 ();
 sg13g2_fill_2 FILLER_65_1772 ();
 sg13g2_decap_8 FILLER_65_1800 ();
 sg13g2_decap_8 FILLER_65_1807 ();
 sg13g2_fill_2 FILLER_65_1819 ();
 sg13g2_fill_1 FILLER_65_1821 ();
 sg13g2_decap_8 FILLER_65_1834 ();
 sg13g2_fill_2 FILLER_65_1841 ();
 sg13g2_fill_1 FILLER_65_1843 ();
 sg13g2_fill_2 FILLER_65_1881 ();
 sg13g2_fill_1 FILLER_65_1883 ();
 sg13g2_fill_2 FILLER_65_1887 ();
 sg13g2_fill_2 FILLER_65_1895 ();
 sg13g2_fill_1 FILLER_65_1897 ();
 sg13g2_decap_8 FILLER_65_1904 ();
 sg13g2_decap_4 FILLER_65_1911 ();
 sg13g2_decap_4 FILLER_65_1931 ();
 sg13g2_decap_4 FILLER_65_1941 ();
 sg13g2_fill_2 FILLER_65_1945 ();
 sg13g2_fill_2 FILLER_65_1970 ();
 sg13g2_fill_1 FILLER_65_1972 ();
 sg13g2_fill_2 FILLER_65_1979 ();
 sg13g2_decap_4 FILLER_65_1986 ();
 sg13g2_decap_4 FILLER_65_1994 ();
 sg13g2_decap_8 FILLER_65_2004 ();
 sg13g2_decap_8 FILLER_65_2027 ();
 sg13g2_fill_1 FILLER_65_2060 ();
 sg13g2_fill_1 FILLER_65_2086 ();
 sg13g2_fill_2 FILLER_65_2097 ();
 sg13g2_fill_2 FILLER_65_2105 ();
 sg13g2_decap_8 FILLER_65_2113 ();
 sg13g2_decap_4 FILLER_65_2120 ();
 sg13g2_fill_1 FILLER_65_2124 ();
 sg13g2_decap_8 FILLER_65_2138 ();
 sg13g2_fill_2 FILLER_65_2145 ();
 sg13g2_decap_8 FILLER_65_2165 ();
 sg13g2_fill_1 FILLER_65_2172 ();
 sg13g2_decap_8 FILLER_65_2181 ();
 sg13g2_decap_4 FILLER_65_2188 ();
 sg13g2_fill_1 FILLER_65_2192 ();
 sg13g2_decap_8 FILLER_65_2198 ();
 sg13g2_decap_4 FILLER_65_2205 ();
 sg13g2_fill_2 FILLER_65_2209 ();
 sg13g2_fill_1 FILLER_65_2220 ();
 sg13g2_decap_8 FILLER_65_2338 ();
 sg13g2_decap_8 FILLER_65_2345 ();
 sg13g2_decap_8 FILLER_65_2352 ();
 sg13g2_decap_8 FILLER_65_2389 ();
 sg13g2_fill_2 FILLER_65_2396 ();
 sg13g2_fill_2 FILLER_65_2402 ();
 sg13g2_fill_1 FILLER_65_2404 ();
 sg13g2_fill_1 FILLER_65_2411 ();
 sg13g2_decap_8 FILLER_65_2429 ();
 sg13g2_decap_4 FILLER_65_2436 ();
 sg13g2_fill_1 FILLER_65_2440 ();
 sg13g2_decap_8 FILLER_65_2445 ();
 sg13g2_decap_8 FILLER_65_2452 ();
 sg13g2_decap_4 FILLER_65_2459 ();
 sg13g2_decap_4 FILLER_65_2557 ();
 sg13g2_fill_2 FILLER_65_2561 ();
 sg13g2_decap_8 FILLER_65_2599 ();
 sg13g2_decap_8 FILLER_65_2637 ();
 sg13g2_decap_8 FILLER_65_2644 ();
 sg13g2_decap_8 FILLER_65_2651 ();
 sg13g2_decap_8 FILLER_65_2658 ();
 sg13g2_decap_4 FILLER_65_2665 ();
 sg13g2_fill_1 FILLER_65_2669 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_fill_2 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_40 ();
 sg13g2_decap_8 FILLER_66_47 ();
 sg13g2_decap_8 FILLER_66_54 ();
 sg13g2_decap_8 FILLER_66_61 ();
 sg13g2_fill_1 FILLER_66_68 ();
 sg13g2_fill_2 FILLER_66_98 ();
 sg13g2_fill_2 FILLER_66_136 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_1 FILLER_66_151 ();
 sg13g2_fill_2 FILLER_66_157 ();
 sg13g2_fill_1 FILLER_66_159 ();
 sg13g2_decap_4 FILLER_66_164 ();
 sg13g2_decap_4 FILLER_66_172 ();
 sg13g2_fill_2 FILLER_66_176 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_decap_4 FILLER_66_204 ();
 sg13g2_fill_1 FILLER_66_208 ();
 sg13g2_fill_2 FILLER_66_219 ();
 sg13g2_fill_2 FILLER_66_296 ();
 sg13g2_fill_1 FILLER_66_298 ();
 sg13g2_decap_4 FILLER_66_325 ();
 sg13g2_decap_8 FILLER_66_355 ();
 sg13g2_fill_2 FILLER_66_362 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_371 ();
 sg13g2_fill_2 FILLER_66_378 ();
 sg13g2_decap_8 FILLER_66_383 ();
 sg13g2_decap_8 FILLER_66_390 ();
 sg13g2_decap_8 FILLER_66_397 ();
 sg13g2_decap_8 FILLER_66_404 ();
 sg13g2_decap_4 FILLER_66_411 ();
 sg13g2_fill_2 FILLER_66_441 ();
 sg13g2_fill_2 FILLER_66_449 ();
 sg13g2_fill_1 FILLER_66_451 ();
 sg13g2_fill_1 FILLER_66_458 ();
 sg13g2_fill_2 FILLER_66_463 ();
 sg13g2_fill_1 FILLER_66_470 ();
 sg13g2_fill_1 FILLER_66_477 ();
 sg13g2_fill_2 FILLER_66_504 ();
 sg13g2_fill_2 FILLER_66_522 ();
 sg13g2_decap_8 FILLER_66_528 ();
 sg13g2_decap_8 FILLER_66_535 ();
 sg13g2_decap_8 FILLER_66_542 ();
 sg13g2_decap_8 FILLER_66_549 ();
 sg13g2_fill_2 FILLER_66_556 ();
 sg13g2_fill_2 FILLER_66_565 ();
 sg13g2_fill_1 FILLER_66_575 ();
 sg13g2_fill_2 FILLER_66_615 ();
 sg13g2_fill_2 FILLER_66_630 ();
 sg13g2_fill_1 FILLER_66_636 ();
 sg13g2_decap_8 FILLER_66_677 ();
 sg13g2_fill_2 FILLER_66_684 ();
 sg13g2_decap_8 FILLER_66_691 ();
 sg13g2_decap_8 FILLER_66_698 ();
 sg13g2_fill_1 FILLER_66_705 ();
 sg13g2_decap_4 FILLER_66_723 ();
 sg13g2_fill_2 FILLER_66_727 ();
 sg13g2_decap_4 FILLER_66_734 ();
 sg13g2_decap_8 FILLER_66_742 ();
 sg13g2_fill_1 FILLER_66_749 ();
 sg13g2_fill_1 FILLER_66_799 ();
 sg13g2_decap_4 FILLER_66_826 ();
 sg13g2_fill_2 FILLER_66_830 ();
 sg13g2_decap_8 FILLER_66_838 ();
 sg13g2_fill_1 FILLER_66_845 ();
 sg13g2_decap_8 FILLER_66_941 ();
 sg13g2_decap_8 FILLER_66_948 ();
 sg13g2_decap_8 FILLER_66_973 ();
 sg13g2_decap_8 FILLER_66_980 ();
 sg13g2_fill_2 FILLER_66_987 ();
 sg13g2_fill_1 FILLER_66_994 ();
 sg13g2_fill_1 FILLER_66_1006 ();
 sg13g2_fill_2 FILLER_66_1018 ();
 sg13g2_fill_1 FILLER_66_1020 ();
 sg13g2_decap_8 FILLER_66_1027 ();
 sg13g2_fill_2 FILLER_66_1034 ();
 sg13g2_fill_1 FILLER_66_1041 ();
 sg13g2_fill_2 FILLER_66_1050 ();
 sg13g2_fill_1 FILLER_66_1052 ();
 sg13g2_fill_1 FILLER_66_1062 ();
 sg13g2_fill_2 FILLER_66_1102 ();
 sg13g2_fill_1 FILLER_66_1109 ();
 sg13g2_fill_2 FILLER_66_1168 ();
 sg13g2_fill_2 FILLER_66_1175 ();
 sg13g2_fill_1 FILLER_66_1177 ();
 sg13g2_decap_8 FILLER_66_1182 ();
 sg13g2_decap_4 FILLER_66_1189 ();
 sg13g2_fill_2 FILLER_66_1193 ();
 sg13g2_fill_1 FILLER_66_1253 ();
 sg13g2_fill_2 FILLER_66_1267 ();
 sg13g2_decap_4 FILLER_66_1304 ();
 sg13g2_fill_2 FILLER_66_1379 ();
 sg13g2_decap_8 FILLER_66_1411 ();
 sg13g2_decap_8 FILLER_66_1418 ();
 sg13g2_decap_4 FILLER_66_1425 ();
 sg13g2_fill_2 FILLER_66_1429 ();
 sg13g2_decap_8 FILLER_66_1460 ();
 sg13g2_decap_8 FILLER_66_1548 ();
 sg13g2_fill_1 FILLER_66_1555 ();
 sg13g2_fill_2 FILLER_66_1559 ();
 sg13g2_decap_8 FILLER_66_1569 ();
 sg13g2_fill_1 FILLER_66_1576 ();
 sg13g2_decap_8 FILLER_66_1582 ();
 sg13g2_fill_1 FILLER_66_1589 ();
 sg13g2_decap_8 FILLER_66_1595 ();
 sg13g2_decap_8 FILLER_66_1602 ();
 sg13g2_decap_8 FILLER_66_1609 ();
 sg13g2_fill_1 FILLER_66_1616 ();
 sg13g2_fill_1 FILLER_66_1657 ();
 sg13g2_fill_2 FILLER_66_1665 ();
 sg13g2_fill_1 FILLER_66_1678 ();
 sg13g2_fill_1 FILLER_66_1708 ();
 sg13g2_decap_8 FILLER_66_1716 ();
 sg13g2_fill_2 FILLER_66_1763 ();
 sg13g2_fill_1 FILLER_66_1765 ();
 sg13g2_decap_8 FILLER_66_1790 ();
 sg13g2_decap_8 FILLER_66_1797 ();
 sg13g2_decap_4 FILLER_66_1804 ();
 sg13g2_decap_8 FILLER_66_1813 ();
 sg13g2_decap_4 FILLER_66_1820 ();
 sg13g2_fill_2 FILLER_66_1824 ();
 sg13g2_decap_8 FILLER_66_1832 ();
 sg13g2_fill_2 FILLER_66_1839 ();
 sg13g2_fill_1 FILLER_66_1841 ();
 sg13g2_decap_4 FILLER_66_1845 ();
 sg13g2_fill_1 FILLER_66_1849 ();
 sg13g2_decap_8 FILLER_66_1855 ();
 sg13g2_fill_2 FILLER_66_1882 ();
 sg13g2_fill_2 FILLER_66_1890 ();
 sg13g2_decap_4 FILLER_66_1928 ();
 sg13g2_fill_1 FILLER_66_1951 ();
 sg13g2_fill_2 FILLER_66_1955 ();
 sg13g2_fill_2 FILLER_66_2001 ();
 sg13g2_fill_1 FILLER_66_2003 ();
 sg13g2_fill_2 FILLER_66_2010 ();
 sg13g2_decap_4 FILLER_66_2043 ();
 sg13g2_fill_2 FILLER_66_2047 ();
 sg13g2_fill_1 FILLER_66_2055 ();
 sg13g2_fill_2 FILLER_66_2082 ();
 sg13g2_fill_2 FILLER_66_2094 ();
 sg13g2_fill_1 FILLER_66_2096 ();
 sg13g2_fill_2 FILLER_66_2123 ();
 sg13g2_fill_1 FILLER_66_2125 ();
 sg13g2_fill_1 FILLER_66_2130 ();
 sg13g2_decap_4 FILLER_66_2162 ();
 sg13g2_fill_1 FILLER_66_2166 ();
 sg13g2_decap_8 FILLER_66_2211 ();
 sg13g2_fill_2 FILLER_66_2218 ();
 sg13g2_fill_1 FILLER_66_2220 ();
 sg13g2_decap_8 FILLER_66_2227 ();
 sg13g2_decap_8 FILLER_66_2234 ();
 sg13g2_decap_8 FILLER_66_2241 ();
 sg13g2_decap_4 FILLER_66_2248 ();
 sg13g2_fill_1 FILLER_66_2262 ();
 sg13g2_fill_2 FILLER_66_2273 ();
 sg13g2_fill_1 FILLER_66_2275 ();
 sg13g2_decap_8 FILLER_66_2305 ();
 sg13g2_decap_4 FILLER_66_2312 ();
 sg13g2_fill_2 FILLER_66_2321 ();
 sg13g2_decap_8 FILLER_66_2327 ();
 sg13g2_decap_8 FILLER_66_2334 ();
 sg13g2_fill_2 FILLER_66_2375 ();
 sg13g2_fill_1 FILLER_66_2377 ();
 sg13g2_fill_2 FILLER_66_2430 ();
 sg13g2_fill_2 FILLER_66_2491 ();
 sg13g2_fill_1 FILLER_66_2493 ();
 sg13g2_fill_1 FILLER_66_2498 ();
 sg13g2_fill_2 FILLER_66_2525 ();
 sg13g2_decap_8 FILLER_66_2553 ();
 sg13g2_decap_8 FILLER_66_2560 ();
 sg13g2_decap_8 FILLER_66_2588 ();
 sg13g2_decap_8 FILLER_66_2595 ();
 sg13g2_fill_2 FILLER_66_2602 ();
 sg13g2_decap_8 FILLER_66_2620 ();
 sg13g2_decap_8 FILLER_66_2627 ();
 sg13g2_decap_8 FILLER_66_2634 ();
 sg13g2_decap_8 FILLER_66_2641 ();
 sg13g2_decap_8 FILLER_66_2648 ();
 sg13g2_decap_8 FILLER_66_2655 ();
 sg13g2_decap_8 FILLER_66_2662 ();
 sg13g2_fill_1 FILLER_66_2669 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_4 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_11 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_fill_2 FILLER_67_56 ();
 sg13g2_fill_1 FILLER_67_92 ();
 sg13g2_fill_2 FILLER_67_102 ();
 sg13g2_fill_1 FILLER_67_134 ();
 sg13g2_fill_2 FILLER_67_139 ();
 sg13g2_fill_1 FILLER_67_141 ();
 sg13g2_fill_1 FILLER_67_146 ();
 sg13g2_decap_8 FILLER_67_151 ();
 sg13g2_fill_1 FILLER_67_158 ();
 sg13g2_fill_2 FILLER_67_166 ();
 sg13g2_decap_8 FILLER_67_201 ();
 sg13g2_fill_2 FILLER_67_208 ();
 sg13g2_fill_1 FILLER_67_210 ();
 sg13g2_fill_1 FILLER_67_221 ();
 sg13g2_decap_8 FILLER_67_243 ();
 sg13g2_decap_8 FILLER_67_250 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_decap_8 FILLER_67_310 ();
 sg13g2_decap_4 FILLER_67_317 ();
 sg13g2_fill_2 FILLER_67_331 ();
 sg13g2_fill_2 FILLER_67_339 ();
 sg13g2_decap_8 FILLER_67_347 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_fill_1 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_398 ();
 sg13g2_decap_8 FILLER_67_405 ();
 sg13g2_decap_8 FILLER_67_412 ();
 sg13g2_fill_1 FILLER_67_424 ();
 sg13g2_fill_2 FILLER_67_456 ();
 sg13g2_fill_1 FILLER_67_464 ();
 sg13g2_fill_1 FILLER_67_475 ();
 sg13g2_fill_1 FILLER_67_484 ();
 sg13g2_decap_8 FILLER_67_503 ();
 sg13g2_decap_8 FILLER_67_510 ();
 sg13g2_decap_8 FILLER_67_517 ();
 sg13g2_decap_8 FILLER_67_524 ();
 sg13g2_decap_8 FILLER_67_531 ();
 sg13g2_decap_8 FILLER_67_538 ();
 sg13g2_fill_2 FILLER_67_545 ();
 sg13g2_fill_1 FILLER_67_547 ();
 sg13g2_decap_8 FILLER_67_585 ();
 sg13g2_fill_1 FILLER_67_592 ();
 sg13g2_fill_2 FILLER_67_642 ();
 sg13g2_fill_2 FILLER_67_648 ();
 sg13g2_fill_1 FILLER_67_660 ();
 sg13g2_decap_8 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_691 ();
 sg13g2_decap_4 FILLER_67_698 ();
 sg13g2_fill_1 FILLER_67_702 ();
 sg13g2_decap_4 FILLER_67_708 ();
 sg13g2_fill_2 FILLER_67_712 ();
 sg13g2_fill_2 FILLER_67_740 ();
 sg13g2_fill_1 FILLER_67_742 ();
 sg13g2_fill_1 FILLER_67_769 ();
 sg13g2_decap_8 FILLER_67_774 ();
 sg13g2_decap_4 FILLER_67_781 ();
 sg13g2_fill_1 FILLER_67_785 ();
 sg13g2_decap_8 FILLER_67_801 ();
 sg13g2_decap_4 FILLER_67_808 ();
 sg13g2_fill_2 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_4 FILLER_67_833 ();
 sg13g2_fill_2 FILLER_67_857 ();
 sg13g2_fill_2 FILLER_67_873 ();
 sg13g2_fill_2 FILLER_67_878 ();
 sg13g2_fill_2 FILLER_67_886 ();
 sg13g2_decap_8 FILLER_67_892 ();
 sg13g2_decap_4 FILLER_67_899 ();
 sg13g2_fill_1 FILLER_67_903 ();
 sg13g2_fill_1 FILLER_67_914 ();
 sg13g2_fill_2 FILLER_67_919 ();
 sg13g2_decap_4 FILLER_67_932 ();
 sg13g2_fill_1 FILLER_67_960 ();
 sg13g2_fill_1 FILLER_67_967 ();
 sg13g2_decap_4 FILLER_67_989 ();
 sg13g2_fill_2 FILLER_67_993 ();
 sg13g2_decap_8 FILLER_67_1004 ();
 sg13g2_decap_4 FILLER_67_1011 ();
 sg13g2_decap_8 FILLER_67_1027 ();
 sg13g2_decap_8 FILLER_67_1034 ();
 sg13g2_decap_4 FILLER_67_1041 ();
 sg13g2_fill_1 FILLER_67_1045 ();
 sg13g2_fill_1 FILLER_67_1118 ();
 sg13g2_decap_8 FILLER_67_1125 ();
 sg13g2_decap_8 FILLER_67_1141 ();
 sg13g2_decap_8 FILLER_67_1148 ();
 sg13g2_fill_2 FILLER_67_1155 ();
 sg13g2_fill_2 FILLER_67_1203 ();
 sg13g2_fill_2 FILLER_67_1213 ();
 sg13g2_fill_1 FILLER_67_1215 ();
 sg13g2_fill_1 FILLER_67_1221 ();
 sg13g2_decap_4 FILLER_67_1228 ();
 sg13g2_fill_1 FILLER_67_1232 ();
 sg13g2_fill_1 FILLER_67_1243 ();
 sg13g2_fill_2 FILLER_67_1270 ();
 sg13g2_decap_8 FILLER_67_1306 ();
 sg13g2_decap_4 FILLER_67_1313 ();
 sg13g2_fill_1 FILLER_67_1322 ();
 sg13g2_decap_4 FILLER_67_1327 ();
 sg13g2_decap_8 FILLER_67_1340 ();
 sg13g2_fill_2 FILLER_67_1347 ();
 sg13g2_fill_1 FILLER_67_1354 ();
 sg13g2_fill_2 FILLER_67_1359 ();
 sg13g2_fill_1 FILLER_67_1366 ();
 sg13g2_fill_1 FILLER_67_1388 ();
 sg13g2_decap_4 FILLER_67_1411 ();
 sg13g2_fill_2 FILLER_67_1415 ();
 sg13g2_decap_8 FILLER_67_1422 ();
 sg13g2_fill_2 FILLER_67_1429 ();
 sg13g2_decap_8 FILLER_67_1436 ();
 sg13g2_fill_1 FILLER_67_1443 ();
 sg13g2_decap_8 FILLER_67_1454 ();
 sg13g2_decap_8 FILLER_67_1461 ();
 sg13g2_fill_2 FILLER_67_1468 ();
 sg13g2_fill_2 FILLER_67_1479 ();
 sg13g2_fill_2 FILLER_67_1520 ();
 sg13g2_decap_8 FILLER_67_1528 ();
 sg13g2_fill_2 FILLER_67_1535 ();
 sg13g2_decap_8 FILLER_67_1540 ();
 sg13g2_fill_1 FILLER_67_1547 ();
 sg13g2_fill_2 FILLER_67_1551 ();
 sg13g2_decap_8 FILLER_67_1565 ();
 sg13g2_decap_8 FILLER_67_1572 ();
 sg13g2_fill_1 FILLER_67_1579 ();
 sg13g2_decap_4 FILLER_67_1588 ();
 sg13g2_decap_8 FILLER_67_1627 ();
 sg13g2_fill_2 FILLER_67_1634 ();
 sg13g2_fill_1 FILLER_67_1636 ();
 sg13g2_fill_2 FILLER_67_1642 ();
 sg13g2_fill_1 FILLER_67_1644 ();
 sg13g2_decap_8 FILLER_67_1653 ();
 sg13g2_decap_4 FILLER_67_1660 ();
 sg13g2_fill_1 FILLER_67_1664 ();
 sg13g2_fill_1 FILLER_67_1674 ();
 sg13g2_fill_2 FILLER_67_1701 ();
 sg13g2_decap_8 FILLER_67_1708 ();
 sg13g2_decap_8 FILLER_67_1715 ();
 sg13g2_fill_1 FILLER_67_1722 ();
 sg13g2_fill_1 FILLER_67_1728 ();
 sg13g2_decap_8 FILLER_67_1735 ();
 sg13g2_decap_8 FILLER_67_1742 ();
 sg13g2_fill_2 FILLER_67_1749 ();
 sg13g2_decap_4 FILLER_67_1760 ();
 sg13g2_fill_2 FILLER_67_1764 ();
 sg13g2_decap_8 FILLER_67_1801 ();
 sg13g2_fill_1 FILLER_67_1808 ();
 sg13g2_fill_1 FILLER_67_1835 ();
 sg13g2_fill_1 FILLER_67_1839 ();
 sg13g2_fill_1 FILLER_67_1873 ();
 sg13g2_fill_1 FILLER_67_1880 ();
 sg13g2_fill_2 FILLER_67_1919 ();
 sg13g2_decap_8 FILLER_67_1927 ();
 sg13g2_decap_8 FILLER_67_1934 ();
 sg13g2_fill_2 FILLER_67_1950 ();
 sg13g2_fill_1 FILLER_67_1958 ();
 sg13g2_fill_2 FILLER_67_1979 ();
 sg13g2_fill_1 FILLER_67_2012 ();
 sg13g2_fill_1 FILLER_67_2016 ();
 sg13g2_decap_8 FILLER_67_2043 ();
 sg13g2_decap_8 FILLER_67_2050 ();
 sg13g2_fill_1 FILLER_67_2057 ();
 sg13g2_decap_4 FILLER_67_2064 ();
 sg13g2_fill_1 FILLER_67_2068 ();
 sg13g2_fill_2 FILLER_67_2078 ();
 sg13g2_decap_4 FILLER_67_2093 ();
 sg13g2_decap_8 FILLER_67_2140 ();
 sg13g2_decap_8 FILLER_67_2147 ();
 sg13g2_decap_4 FILLER_67_2158 ();
 sg13g2_fill_2 FILLER_67_2172 ();
 sg13g2_fill_1 FILLER_67_2174 ();
 sg13g2_fill_1 FILLER_67_2181 ();
 sg13g2_decap_8 FILLER_67_2191 ();
 sg13g2_decap_4 FILLER_67_2198 ();
 sg13g2_fill_2 FILLER_67_2237 ();
 sg13g2_fill_1 FILLER_67_2239 ();
 sg13g2_decap_8 FILLER_67_2244 ();
 sg13g2_fill_1 FILLER_67_2251 ();
 sg13g2_fill_1 FILLER_67_2296 ();
 sg13g2_fill_1 FILLER_67_2305 ();
 sg13g2_fill_2 FILLER_67_2312 ();
 sg13g2_fill_2 FILLER_67_2320 ();
 sg13g2_fill_1 FILLER_67_2375 ();
 sg13g2_fill_1 FILLER_67_2381 ();
 sg13g2_fill_1 FILLER_67_2386 ();
 sg13g2_fill_1 FILLER_67_2391 ();
 sg13g2_fill_2 FILLER_67_2397 ();
 sg13g2_fill_1 FILLER_67_2455 ();
 sg13g2_fill_2 FILLER_67_2473 ();
 sg13g2_fill_2 FILLER_67_2488 ();
 sg13g2_decap_4 FILLER_67_2494 ();
 sg13g2_fill_1 FILLER_67_2507 ();
 sg13g2_fill_2 FILLER_67_2525 ();
 sg13g2_fill_1 FILLER_67_2527 ();
 sg13g2_decap_4 FILLER_67_2532 ();
 sg13g2_decap_4 FILLER_67_2540 ();
 sg13g2_decap_8 FILLER_67_2548 ();
 sg13g2_decap_8 FILLER_67_2555 ();
 sg13g2_decap_8 FILLER_67_2562 ();
 sg13g2_fill_2 FILLER_67_2569 ();
 sg13g2_decap_8 FILLER_67_2575 ();
 sg13g2_decap_8 FILLER_67_2582 ();
 sg13g2_decap_8 FILLER_67_2623 ();
 sg13g2_decap_8 FILLER_67_2630 ();
 sg13g2_decap_8 FILLER_67_2637 ();
 sg13g2_decap_8 FILLER_67_2644 ();
 sg13g2_decap_8 FILLER_67_2655 ();
 sg13g2_decap_8 FILLER_67_2662 ();
 sg13g2_fill_1 FILLER_67_2669 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_4 FILLER_68_21 ();
 sg13g2_fill_2 FILLER_68_25 ();
 sg13g2_decap_4 FILLER_68_56 ();
 sg13g2_fill_1 FILLER_68_78 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_171 ();
 sg13g2_decap_8 FILLER_68_178 ();
 sg13g2_decap_8 FILLER_68_185 ();
 sg13g2_decap_8 FILLER_68_192 ();
 sg13g2_decap_8 FILLER_68_199 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_decap_8 FILLER_68_213 ();
 sg13g2_decap_8 FILLER_68_220 ();
 sg13g2_decap_4 FILLER_68_227 ();
 sg13g2_fill_1 FILLER_68_231 ();
 sg13g2_decap_8 FILLER_68_247 ();
 sg13g2_decap_8 FILLER_68_254 ();
 sg13g2_decap_8 FILLER_68_261 ();
 sg13g2_decap_8 FILLER_68_268 ();
 sg13g2_decap_8 FILLER_68_275 ();
 sg13g2_decap_8 FILLER_68_282 ();
 sg13g2_decap_8 FILLER_68_289 ();
 sg13g2_decap_4 FILLER_68_296 ();
 sg13g2_fill_1 FILLER_68_300 ();
 sg13g2_fill_1 FILLER_68_314 ();
 sg13g2_decap_8 FILLER_68_394 ();
 sg13g2_decap_8 FILLER_68_409 ();
 sg13g2_decap_8 FILLER_68_416 ();
 sg13g2_fill_1 FILLER_68_423 ();
 sg13g2_fill_2 FILLER_68_433 ();
 sg13g2_fill_1 FILLER_68_445 ();
 sg13g2_decap_4 FILLER_68_455 ();
 sg13g2_fill_1 FILLER_68_459 ();
 sg13g2_fill_2 FILLER_68_464 ();
 sg13g2_fill_1 FILLER_68_466 ();
 sg13g2_fill_2 FILLER_68_496 ();
 sg13g2_fill_1 FILLER_68_498 ();
 sg13g2_decap_8 FILLER_68_525 ();
 sg13g2_decap_8 FILLER_68_532 ();
 sg13g2_decap_8 FILLER_68_539 ();
 sg13g2_fill_2 FILLER_68_554 ();
 sg13g2_fill_1 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_598 ();
 sg13g2_decap_4 FILLER_68_615 ();
 sg13g2_fill_1 FILLER_68_619 ();
 sg13g2_fill_1 FILLER_68_633 ();
 sg13g2_fill_2 FILLER_68_644 ();
 sg13g2_decap_8 FILLER_68_651 ();
 sg13g2_decap_8 FILLER_68_658 ();
 sg13g2_decap_8 FILLER_68_665 ();
 sg13g2_decap_8 FILLER_68_672 ();
 sg13g2_fill_1 FILLER_68_679 ();
 sg13g2_decap_8 FILLER_68_710 ();
 sg13g2_fill_2 FILLER_68_717 ();
 sg13g2_fill_1 FILLER_68_719 ();
 sg13g2_fill_1 FILLER_68_728 ();
 sg13g2_fill_1 FILLER_68_764 ();
 sg13g2_fill_1 FILLER_68_812 ();
 sg13g2_decap_8 FILLER_68_822 ();
 sg13g2_decap_4 FILLER_68_829 ();
 sg13g2_fill_1 FILLER_68_833 ();
 sg13g2_fill_1 FILLER_68_874 ();
 sg13g2_fill_2 FILLER_68_878 ();
 sg13g2_decap_8 FILLER_68_892 ();
 sg13g2_fill_2 FILLER_68_899 ();
 sg13g2_fill_1 FILLER_68_901 ();
 sg13g2_decap_8 FILLER_68_908 ();
 sg13g2_fill_1 FILLER_68_915 ();
 sg13g2_fill_2 FILLER_68_924 ();
 sg13g2_fill_1 FILLER_68_926 ();
 sg13g2_fill_2 FILLER_68_966 ();
 sg13g2_fill_2 FILLER_68_977 ();
 sg13g2_decap_4 FILLER_68_992 ();
 sg13g2_decap_8 FILLER_68_1032 ();
 sg13g2_decap_4 FILLER_68_1039 ();
 sg13g2_fill_2 FILLER_68_1043 ();
 sg13g2_fill_1 FILLER_68_1071 ();
 sg13g2_fill_2 FILLER_68_1100 ();
 sg13g2_decap_4 FILLER_68_1109 ();
 sg13g2_fill_2 FILLER_68_1118 ();
 sg13g2_fill_1 FILLER_68_1132 ();
 sg13g2_decap_4 FILLER_68_1159 ();
 sg13g2_decap_4 FILLER_68_1189 ();
 sg13g2_fill_1 FILLER_68_1193 ();
 sg13g2_decap_8 FILLER_68_1198 ();
 sg13g2_decap_8 FILLER_68_1205 ();
 sg13g2_decap_4 FILLER_68_1212 ();
 sg13g2_decap_8 FILLER_68_1225 ();
 sg13g2_decap_8 FILLER_68_1232 ();
 sg13g2_decap_8 FILLER_68_1239 ();
 sg13g2_fill_1 FILLER_68_1246 ();
 sg13g2_fill_2 FILLER_68_1252 ();
 sg13g2_fill_2 FILLER_68_1270 ();
 sg13g2_fill_2 FILLER_68_1305 ();
 sg13g2_fill_1 FILLER_68_1307 ();
 sg13g2_decap_8 FILLER_68_1320 ();
 sg13g2_decap_8 FILLER_68_1327 ();
 sg13g2_decap_8 FILLER_68_1346 ();
 sg13g2_decap_8 FILLER_68_1353 ();
 sg13g2_decap_8 FILLER_68_1360 ();
 sg13g2_decap_8 FILLER_68_1367 ();
 sg13g2_fill_2 FILLER_68_1374 ();
 sg13g2_fill_1 FILLER_68_1376 ();
 sg13g2_decap_8 FILLER_68_1410 ();
 sg13g2_decap_4 FILLER_68_1417 ();
 sg13g2_fill_2 FILLER_68_1421 ();
 sg13g2_fill_2 FILLER_68_1461 ();
 sg13g2_fill_1 FILLER_68_1463 ();
 sg13g2_decap_8 FILLER_68_1507 ();
 sg13g2_decap_4 FILLER_68_1514 ();
 sg13g2_fill_1 FILLER_68_1527 ();
 sg13g2_fill_2 FILLER_68_1534 ();
 sg13g2_fill_1 FILLER_68_1536 ();
 sg13g2_decap_4 FILLER_68_1574 ();
 sg13g2_fill_2 FILLER_68_1578 ();
 sg13g2_decap_8 FILLER_68_1584 ();
 sg13g2_decap_8 FILLER_68_1591 ();
 sg13g2_decap_4 FILLER_68_1598 ();
 sg13g2_decap_4 FILLER_68_1605 ();
 sg13g2_fill_2 FILLER_68_1609 ();
 sg13g2_decap_4 FILLER_68_1645 ();
 sg13g2_fill_2 FILLER_68_1659 ();
 sg13g2_fill_2 FILLER_68_1665 ();
 sg13g2_fill_1 FILLER_68_1667 ();
 sg13g2_fill_2 FILLER_68_1671 ();
 sg13g2_decap_4 FILLER_68_1699 ();
 sg13g2_decap_8 FILLER_68_1734 ();
 sg13g2_decap_8 FILLER_68_1741 ();
 sg13g2_decap_8 FILLER_68_1748 ();
 sg13g2_fill_1 FILLER_68_1755 ();
 sg13g2_decap_4 FILLER_68_1760 ();
 sg13g2_decap_4 FILLER_68_1769 ();
 sg13g2_fill_2 FILLER_68_1773 ();
 sg13g2_decap_4 FILLER_68_1779 ();
 sg13g2_fill_2 FILLER_68_1783 ();
 sg13g2_fill_2 FILLER_68_1789 ();
 sg13g2_decap_8 FILLER_68_1797 ();
 sg13g2_decap_8 FILLER_68_1804 ();
 sg13g2_decap_4 FILLER_68_1811 ();
 sg13g2_fill_2 FILLER_68_1815 ();
 sg13g2_decap_8 FILLER_68_1820 ();
 sg13g2_fill_1 FILLER_68_1827 ();
 sg13g2_fill_2 FILLER_68_1845 ();
 sg13g2_decap_8 FILLER_68_1924 ();
 sg13g2_fill_1 FILLER_68_1931 ();
 sg13g2_decap_8 FILLER_68_1958 ();
 sg13g2_fill_2 FILLER_68_1971 ();
 sg13g2_decap_8 FILLER_68_2022 ();
 sg13g2_decap_8 FILLER_68_2029 ();
 sg13g2_decap_8 FILLER_68_2036 ();
 sg13g2_decap_8 FILLER_68_2043 ();
 sg13g2_decap_8 FILLER_68_2050 ();
 sg13g2_decap_8 FILLER_68_2057 ();
 sg13g2_decap_4 FILLER_68_2064 ();
 sg13g2_decap_4 FILLER_68_2078 ();
 sg13g2_decap_4 FILLER_68_2118 ();
 sg13g2_fill_1 FILLER_68_2122 ();
 sg13g2_fill_1 FILLER_68_2128 ();
 sg13g2_fill_1 FILLER_68_2133 ();
 sg13g2_fill_1 FILLER_68_2139 ();
 sg13g2_fill_2 FILLER_68_2144 ();
 sg13g2_fill_1 FILLER_68_2181 ();
 sg13g2_fill_2 FILLER_68_2203 ();
 sg13g2_fill_1 FILLER_68_2205 ();
 sg13g2_decap_4 FILLER_68_2248 ();
 sg13g2_fill_1 FILLER_68_2252 ();
 sg13g2_fill_2 FILLER_68_2265 ();
 sg13g2_decap_8 FILLER_68_2280 ();
 sg13g2_fill_2 FILLER_68_2287 ();
 sg13g2_fill_1 FILLER_68_2289 ();
 sg13g2_decap_4 FILLER_68_2296 ();
 sg13g2_fill_1 FILLER_68_2300 ();
 sg13g2_decap_8 FILLER_68_2306 ();
 sg13g2_fill_2 FILLER_68_2313 ();
 sg13g2_fill_2 FILLER_68_2319 ();
 sg13g2_decap_4 FILLER_68_2355 ();
 sg13g2_decap_4 FILLER_68_2363 ();
 sg13g2_decap_8 FILLER_68_2373 ();
 sg13g2_decap_8 FILLER_68_2380 ();
 sg13g2_decap_8 FILLER_68_2387 ();
 sg13g2_decap_8 FILLER_68_2394 ();
 sg13g2_decap_4 FILLER_68_2401 ();
 sg13g2_fill_1 FILLER_68_2405 ();
 sg13g2_decap_8 FILLER_68_2414 ();
 sg13g2_fill_2 FILLER_68_2421 ();
 sg13g2_fill_1 FILLER_68_2423 ();
 sg13g2_fill_1 FILLER_68_2434 ();
 sg13g2_fill_1 FILLER_68_2439 ();
 sg13g2_decap_4 FILLER_68_2454 ();
 sg13g2_fill_1 FILLER_68_2458 ();
 sg13g2_decap_8 FILLER_68_2474 ();
 sg13g2_decap_4 FILLER_68_2481 ();
 sg13g2_fill_2 FILLER_68_2500 ();
 sg13g2_fill_1 FILLER_68_2502 ();
 sg13g2_fill_2 FILLER_68_2559 ();
 sg13g2_decap_8 FILLER_68_2587 ();
 sg13g2_decap_8 FILLER_68_2594 ();
 sg13g2_fill_1 FILLER_68_2601 ();
 sg13g2_decap_8 FILLER_68_2618 ();
 sg13g2_decap_8 FILLER_68_2625 ();
 sg13g2_decap_4 FILLER_68_2666 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_4 FILLER_69_21 ();
 sg13g2_fill_2 FILLER_69_25 ();
 sg13g2_fill_1 FILLER_69_80 ();
 sg13g2_fill_2 FILLER_69_86 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_fill_1 FILLER_69_94 ();
 sg13g2_fill_2 FILLER_69_105 ();
 sg13g2_decap_4 FILLER_69_119 ();
 sg13g2_fill_2 FILLER_69_123 ();
 sg13g2_fill_1 FILLER_69_146 ();
 sg13g2_fill_1 FILLER_69_154 ();
 sg13g2_fill_1 FILLER_69_161 ();
 sg13g2_fill_1 FILLER_69_181 ();
 sg13g2_decap_8 FILLER_69_187 ();
 sg13g2_decap_8 FILLER_69_194 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_decap_8 FILLER_69_215 ();
 sg13g2_decap_8 FILLER_69_222 ();
 sg13g2_fill_1 FILLER_69_229 ();
 sg13g2_fill_2 FILLER_69_235 ();
 sg13g2_fill_1 FILLER_69_237 ();
 sg13g2_fill_2 FILLER_69_243 ();
 sg13g2_decap_8 FILLER_69_250 ();
 sg13g2_decap_8 FILLER_69_257 ();
 sg13g2_decap_8 FILLER_69_264 ();
 sg13g2_decap_8 FILLER_69_271 ();
 sg13g2_decap_4 FILLER_69_278 ();
 sg13g2_fill_2 FILLER_69_282 ();
 sg13g2_fill_2 FILLER_69_304 ();
 sg13g2_decap_4 FILLER_69_332 ();
 sg13g2_decap_4 FILLER_69_339 ();
 sg13g2_decap_8 FILLER_69_349 ();
 sg13g2_fill_2 FILLER_69_356 ();
 sg13g2_decap_8 FILLER_69_398 ();
 sg13g2_fill_1 FILLER_69_405 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_414 ();
 sg13g2_fill_2 FILLER_69_421 ();
 sg13g2_decap_8 FILLER_69_427 ();
 sg13g2_fill_1 FILLER_69_434 ();
 sg13g2_decap_4 FILLER_69_439 ();
 sg13g2_fill_1 FILLER_69_443 ();
 sg13g2_fill_1 FILLER_69_451 ();
 sg13g2_fill_1 FILLER_69_456 ();
 sg13g2_decap_4 FILLER_69_462 ();
 sg13g2_fill_2 FILLER_69_471 ();
 sg13g2_fill_2 FILLER_69_492 ();
 sg13g2_fill_2 FILLER_69_499 ();
 sg13g2_fill_1 FILLER_69_501 ();
 sg13g2_decap_8 FILLER_69_528 ();
 sg13g2_decap_8 FILLER_69_535 ();
 sg13g2_decap_8 FILLER_69_542 ();
 sg13g2_fill_1 FILLER_69_549 ();
 sg13g2_fill_1 FILLER_69_581 ();
 sg13g2_decap_4 FILLER_69_596 ();
 sg13g2_fill_1 FILLER_69_600 ();
 sg13g2_fill_1 FILLER_69_630 ();
 sg13g2_decap_8 FILLER_69_660 ();
 sg13g2_decap_8 FILLER_69_667 ();
 sg13g2_fill_2 FILLER_69_674 ();
 sg13g2_fill_1 FILLER_69_676 ();
 sg13g2_decap_4 FILLER_69_703 ();
 sg13g2_fill_2 FILLER_69_738 ();
 sg13g2_fill_1 FILLER_69_744 ();
 sg13g2_decap_8 FILLER_69_834 ();
 sg13g2_fill_2 FILLER_69_852 ();
 sg13g2_fill_1 FILLER_69_871 ();
 sg13g2_fill_1 FILLER_69_887 ();
 sg13g2_fill_2 FILLER_69_891 ();
 sg13g2_decap_4 FILLER_69_922 ();
 sg13g2_fill_2 FILLER_69_926 ();
 sg13g2_fill_2 FILLER_69_961 ();
 sg13g2_fill_2 FILLER_69_985 ();
 sg13g2_decap_8 FILLER_69_1005 ();
 sg13g2_fill_2 FILLER_69_1039 ();
 sg13g2_decap_4 FILLER_69_1051 ();
 sg13g2_fill_1 FILLER_69_1055 ();
 sg13g2_fill_1 FILLER_69_1071 ();
 sg13g2_decap_4 FILLER_69_1081 ();
 sg13g2_fill_2 FILLER_69_1085 ();
 sg13g2_fill_2 FILLER_69_1096 ();
 sg13g2_fill_1 FILLER_69_1098 ();
 sg13g2_fill_1 FILLER_69_1129 ();
 sg13g2_decap_8 FILLER_69_1139 ();
 sg13g2_decap_8 FILLER_69_1146 ();
 sg13g2_decap_4 FILLER_69_1153 ();
 sg13g2_fill_2 FILLER_69_1157 ();
 sg13g2_fill_2 FILLER_69_1176 ();
 sg13g2_fill_1 FILLER_69_1178 ();
 sg13g2_decap_8 FILLER_69_1205 ();
 sg13g2_decap_4 FILLER_69_1212 ();
 sg13g2_fill_2 FILLER_69_1216 ();
 sg13g2_decap_8 FILLER_69_1222 ();
 sg13g2_fill_2 FILLER_69_1229 ();
 sg13g2_fill_1 FILLER_69_1231 ();
 sg13g2_decap_8 FILLER_69_1237 ();
 sg13g2_fill_2 FILLER_69_1254 ();
 sg13g2_fill_2 FILLER_69_1261 ();
 sg13g2_fill_1 FILLER_69_1279 ();
 sg13g2_fill_2 FILLER_69_1302 ();
 sg13g2_fill_1 FILLER_69_1339 ();
 sg13g2_decap_8 FILLER_69_1352 ();
 sg13g2_fill_2 FILLER_69_1359 ();
 sg13g2_decap_4 FILLER_69_1366 ();
 sg13g2_fill_1 FILLER_69_1370 ();
 sg13g2_fill_1 FILLER_69_1379 ();
 sg13g2_decap_4 FILLER_69_1415 ();
 sg13g2_fill_1 FILLER_69_1419 ();
 sg13g2_decap_8 FILLER_69_1426 ();
 sg13g2_fill_2 FILLER_69_1433 ();
 sg13g2_fill_1 FILLER_69_1435 ();
 sg13g2_decap_4 FILLER_69_1441 ();
 sg13g2_fill_1 FILLER_69_1449 ();
 sg13g2_fill_1 FILLER_69_1486 ();
 sg13g2_fill_2 FILLER_69_1516 ();
 sg13g2_fill_1 FILLER_69_1583 ();
 sg13g2_decap_8 FILLER_69_1588 ();
 sg13g2_decap_4 FILLER_69_1595 ();
 sg13g2_fill_2 FILLER_69_1623 ();
 sg13g2_fill_1 FILLER_69_1625 ();
 sg13g2_fill_1 FILLER_69_1664 ();
 sg13g2_fill_2 FILLER_69_1678 ();
 sg13g2_fill_1 FILLER_69_1680 ();
 sg13g2_decap_8 FILLER_69_1685 ();
 sg13g2_fill_1 FILLER_69_1692 ();
 sg13g2_decap_4 FILLER_69_1698 ();
 sg13g2_fill_1 FILLER_69_1702 ();
 sg13g2_decap_4 FILLER_69_1716 ();
 sg13g2_fill_2 FILLER_69_1724 ();
 sg13g2_decap_4 FILLER_69_1734 ();
 sg13g2_fill_2 FILLER_69_1738 ();
 sg13g2_decap_8 FILLER_69_1744 ();
 sg13g2_decap_4 FILLER_69_1751 ();
 sg13g2_fill_1 FILLER_69_1755 ();
 sg13g2_fill_1 FILLER_69_1764 ();
 sg13g2_decap_8 FILLER_69_1804 ();
 sg13g2_fill_1 FILLER_69_1826 ();
 sg13g2_fill_1 FILLER_69_1839 ();
 sg13g2_fill_2 FILLER_69_1879 ();
 sg13g2_fill_1 FILLER_69_1892 ();
 sg13g2_decap_8 FILLER_69_1917 ();
 sg13g2_decap_8 FILLER_69_1924 ();
 sg13g2_decap_8 FILLER_69_1931 ();
 sg13g2_decap_8 FILLER_69_1938 ();
 sg13g2_decap_4 FILLER_69_1945 ();
 sg13g2_fill_2 FILLER_69_1961 ();
 sg13g2_fill_2 FILLER_69_1981 ();
 sg13g2_fill_1 FILLER_69_1983 ();
 sg13g2_fill_2 FILLER_69_2003 ();
 sg13g2_fill_2 FILLER_69_2011 ();
 sg13g2_decap_8 FILLER_69_2021 ();
 sg13g2_decap_8 FILLER_69_2028 ();
 sg13g2_decap_4 FILLER_69_2035 ();
 sg13g2_decap_8 FILLER_69_2045 ();
 sg13g2_fill_1 FILLER_69_2052 ();
 sg13g2_decap_8 FILLER_69_2062 ();
 sg13g2_decap_4 FILLER_69_2069 ();
 sg13g2_decap_4 FILLER_69_2084 ();
 sg13g2_fill_2 FILLER_69_2092 ();
 sg13g2_fill_1 FILLER_69_2102 ();
 sg13g2_decap_8 FILLER_69_2111 ();
 sg13g2_decap_8 FILLER_69_2118 ();
 sg13g2_decap_8 FILLER_69_2151 ();
 sg13g2_decap_8 FILLER_69_2158 ();
 sg13g2_decap_8 FILLER_69_2165 ();
 sg13g2_fill_2 FILLER_69_2172 ();
 sg13g2_fill_1 FILLER_69_2174 ();
 sg13g2_fill_1 FILLER_69_2181 ();
 sg13g2_fill_2 FILLER_69_2185 ();
 sg13g2_fill_1 FILLER_69_2187 ();
 sg13g2_decap_8 FILLER_69_2194 ();
 sg13g2_fill_2 FILLER_69_2201 ();
 sg13g2_fill_1 FILLER_69_2212 ();
 sg13g2_decap_8 FILLER_69_2218 ();
 sg13g2_decap_4 FILLER_69_2225 ();
 sg13g2_decap_4 FILLER_69_2261 ();
 sg13g2_fill_2 FILLER_69_2265 ();
 sg13g2_decap_8 FILLER_69_2275 ();
 sg13g2_decap_8 FILLER_69_2282 ();
 sg13g2_fill_2 FILLER_69_2289 ();
 sg13g2_fill_1 FILLER_69_2291 ();
 sg13g2_decap_8 FILLER_69_2298 ();
 sg13g2_decap_8 FILLER_69_2305 ();
 sg13g2_decap_8 FILLER_69_2312 ();
 sg13g2_decap_4 FILLER_69_2319 ();
 sg13g2_decap_8 FILLER_69_2353 ();
 sg13g2_decap_8 FILLER_69_2360 ();
 sg13g2_decap_8 FILLER_69_2408 ();
 sg13g2_fill_2 FILLER_69_2415 ();
 sg13g2_fill_1 FILLER_69_2417 ();
 sg13g2_decap_4 FILLER_69_2428 ();
 sg13g2_decap_4 FILLER_69_2465 ();
 sg13g2_fill_2 FILLER_69_2564 ();
 sg13g2_fill_2 FILLER_69_2570 ();
 sg13g2_fill_1 FILLER_69_2572 ();
 sg13g2_decap_8 FILLER_69_2590 ();
 sg13g2_fill_2 FILLER_69_2597 ();
 sg13g2_decap_8 FILLER_69_2612 ();
 sg13g2_fill_2 FILLER_69_2619 ();
 sg13g2_fill_1 FILLER_69_2621 ();
 sg13g2_fill_2 FILLER_69_2660 ();
 sg13g2_decap_4 FILLER_69_2666 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_35 ();
 sg13g2_fill_2 FILLER_70_51 ();
 sg13g2_fill_2 FILLER_70_64 ();
 sg13g2_fill_1 FILLER_70_66 ();
 sg13g2_fill_2 FILLER_70_112 ();
 sg13g2_fill_1 FILLER_70_114 ();
 sg13g2_fill_2 FILLER_70_120 ();
 sg13g2_fill_1 FILLER_70_122 ();
 sg13g2_decap_8 FILLER_70_128 ();
 sg13g2_decap_4 FILLER_70_135 ();
 sg13g2_decap_8 FILLER_70_144 ();
 sg13g2_fill_1 FILLER_70_151 ();
 sg13g2_decap_8 FILLER_70_155 ();
 sg13g2_fill_2 FILLER_70_167 ();
 sg13g2_decap_4 FILLER_70_184 ();
 sg13g2_decap_8 FILLER_70_192 ();
 sg13g2_decap_8 FILLER_70_199 ();
 sg13g2_decap_4 FILLER_70_206 ();
 sg13g2_fill_2 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_220 ();
 sg13g2_decap_8 FILLER_70_227 ();
 sg13g2_decap_4 FILLER_70_254 ();
 sg13g2_fill_2 FILLER_70_294 ();
 sg13g2_fill_1 FILLER_70_296 ();
 sg13g2_decap_8 FILLER_70_323 ();
 sg13g2_decap_8 FILLER_70_330 ();
 sg13g2_decap_4 FILLER_70_337 ();
 sg13g2_fill_2 FILLER_70_341 ();
 sg13g2_fill_2 FILLER_70_436 ();
 sg13g2_fill_2 FILLER_70_442 ();
 sg13g2_fill_1 FILLER_70_444 ();
 sg13g2_fill_1 FILLER_70_455 ();
 sg13g2_fill_2 FILLER_70_459 ();
 sg13g2_fill_1 FILLER_70_461 ();
 sg13g2_fill_2 FILLER_70_466 ();
 sg13g2_fill_1 FILLER_70_468 ();
 sg13g2_fill_2 FILLER_70_474 ();
 sg13g2_fill_1 FILLER_70_476 ();
 sg13g2_fill_1 FILLER_70_491 ();
 sg13g2_fill_2 FILLER_70_523 ();
 sg13g2_fill_1 FILLER_70_525 ();
 sg13g2_fill_1 FILLER_70_557 ();
 sg13g2_fill_1 FILLER_70_570 ();
 sg13g2_decap_8 FILLER_70_597 ();
 sg13g2_decap_8 FILLER_70_604 ();
 sg13g2_decap_8 FILLER_70_611 ();
 sg13g2_fill_2 FILLER_70_622 ();
 sg13g2_fill_1 FILLER_70_649 ();
 sg13g2_decap_8 FILLER_70_654 ();
 sg13g2_decap_8 FILLER_70_661 ();
 sg13g2_decap_8 FILLER_70_668 ();
 sg13g2_decap_8 FILLER_70_675 ();
 sg13g2_decap_4 FILLER_70_682 ();
 sg13g2_fill_2 FILLER_70_686 ();
 sg13g2_fill_2 FILLER_70_697 ();
 sg13g2_decap_8 FILLER_70_712 ();
 sg13g2_decap_8 FILLER_70_719 ();
 sg13g2_fill_2 FILLER_70_726 ();
 sg13g2_fill_1 FILLER_70_754 ();
 sg13g2_fill_1 FILLER_70_773 ();
 sg13g2_fill_1 FILLER_70_843 ();
 sg13g2_fill_1 FILLER_70_875 ();
 sg13g2_fill_2 FILLER_70_888 ();
 sg13g2_decap_8 FILLER_70_933 ();
 sg13g2_decap_8 FILLER_70_940 ();
 sg13g2_fill_1 FILLER_70_947 ();
 sg13g2_fill_2 FILLER_70_980 ();
 sg13g2_fill_2 FILLER_70_991 ();
 sg13g2_fill_2 FILLER_70_997 ();
 sg13g2_fill_2 FILLER_70_1025 ();
 sg13g2_decap_8 FILLER_70_1053 ();
 sg13g2_decap_8 FILLER_70_1060 ();
 sg13g2_decap_8 FILLER_70_1067 ();
 sg13g2_decap_8 FILLER_70_1074 ();
 sg13g2_decap_8 FILLER_70_1081 ();
 sg13g2_decap_4 FILLER_70_1088 ();
 sg13g2_fill_2 FILLER_70_1092 ();
 sg13g2_decap_8 FILLER_70_1099 ();
 sg13g2_fill_1 FILLER_70_1106 ();
 sg13g2_fill_1 FILLER_70_1115 ();
 sg13g2_decap_8 FILLER_70_1142 ();
 sg13g2_decap_8 FILLER_70_1149 ();
 sg13g2_decap_8 FILLER_70_1156 ();
 sg13g2_decap_8 FILLER_70_1163 ();
 sg13g2_fill_2 FILLER_70_1182 ();
 sg13g2_fill_1 FILLER_70_1184 ();
 sg13g2_decap_8 FILLER_70_1215 ();
 sg13g2_fill_2 FILLER_70_1222 ();
 sg13g2_fill_2 FILLER_70_1258 ();
 sg13g2_fill_1 FILLER_70_1260 ();
 sg13g2_decap_8 FILLER_70_1267 ();
 sg13g2_fill_1 FILLER_70_1274 ();
 sg13g2_decap_8 FILLER_70_1279 ();
 sg13g2_fill_2 FILLER_70_1286 ();
 sg13g2_decap_8 FILLER_70_1294 ();
 sg13g2_fill_1 FILLER_70_1301 ();
 sg13g2_decap_8 FILLER_70_1342 ();
 sg13g2_decap_8 FILLER_70_1349 ();
 sg13g2_decap_4 FILLER_70_1356 ();
 sg13g2_fill_2 FILLER_70_1360 ();
 sg13g2_fill_2 FILLER_70_1366 ();
 sg13g2_fill_1 FILLER_70_1376 ();
 sg13g2_decap_8 FILLER_70_1393 ();
 sg13g2_decap_4 FILLER_70_1400 ();
 sg13g2_fill_1 FILLER_70_1404 ();
 sg13g2_fill_1 FILLER_70_1436 ();
 sg13g2_fill_1 FILLER_70_1441 ();
 sg13g2_fill_1 FILLER_70_1468 ();
 sg13g2_fill_1 FILLER_70_1475 ();
 sg13g2_fill_2 FILLER_70_1481 ();
 sg13g2_decap_4 FILLER_70_1487 ();
 sg13g2_fill_1 FILLER_70_1491 ();
 sg13g2_decap_8 FILLER_70_1502 ();
 sg13g2_decap_8 FILLER_70_1509 ();
 sg13g2_fill_2 FILLER_70_1516 ();
 sg13g2_decap_8 FILLER_70_1589 ();
 sg13g2_decap_8 FILLER_70_1596 ();
 sg13g2_fill_2 FILLER_70_1603 ();
 sg13g2_fill_1 FILLER_70_1605 ();
 sg13g2_fill_2 FILLER_70_1614 ();
 sg13g2_decap_4 FILLER_70_1630 ();
 sg13g2_fill_2 FILLER_70_1634 ();
 sg13g2_decap_8 FILLER_70_1676 ();
 sg13g2_decap_8 FILLER_70_1683 ();
 sg13g2_fill_2 FILLER_70_1690 ();
 sg13g2_fill_2 FILLER_70_1700 ();
 sg13g2_fill_1 FILLER_70_1702 ();
 sg13g2_decap_8 FILLER_70_1733 ();
 sg13g2_fill_1 FILLER_70_1757 ();
 sg13g2_decap_8 FILLER_70_1784 ();
 sg13g2_fill_1 FILLER_70_1794 ();
 sg13g2_fill_1 FILLER_70_1812 ();
 sg13g2_fill_1 FILLER_70_1858 ();
 sg13g2_fill_2 FILLER_70_1875 ();
 sg13g2_fill_2 FILLER_70_1915 ();
 sg13g2_fill_2 FILLER_70_1936 ();
 sg13g2_decap_8 FILLER_70_1946 ();
 sg13g2_decap_8 FILLER_70_1953 ();
 sg13g2_decap_4 FILLER_70_1960 ();
 sg13g2_fill_2 FILLER_70_1970 ();
 sg13g2_decap_8 FILLER_70_1980 ();
 sg13g2_fill_2 FILLER_70_1993 ();
 sg13g2_fill_1 FILLER_70_2041 ();
 sg13g2_decap_4 FILLER_70_2056 ();
 sg13g2_fill_2 FILLER_70_2060 ();
 sg13g2_fill_2 FILLER_70_2073 ();
 sg13g2_fill_1 FILLER_70_2075 ();
 sg13g2_fill_1 FILLER_70_2080 ();
 sg13g2_fill_2 FILLER_70_2091 ();
 sg13g2_fill_1 FILLER_70_2093 ();
 sg13g2_decap_8 FILLER_70_2104 ();
 sg13g2_decap_8 FILLER_70_2111 ();
 sg13g2_decap_8 FILLER_70_2118 ();
 sg13g2_decap_8 FILLER_70_2125 ();
 sg13g2_fill_1 FILLER_70_2132 ();
 sg13g2_decap_4 FILLER_70_2153 ();
 sg13g2_fill_1 FILLER_70_2170 ();
 sg13g2_fill_1 FILLER_70_2185 ();
 sg13g2_decap_8 FILLER_70_2196 ();
 sg13g2_fill_2 FILLER_70_2203 ();
 sg13g2_fill_1 FILLER_70_2231 ();
 sg13g2_fill_1 FILLER_70_2240 ();
 sg13g2_decap_8 FILLER_70_2251 ();
 sg13g2_decap_4 FILLER_70_2258 ();
 sg13g2_fill_1 FILLER_70_2262 ();
 sg13g2_fill_2 FILLER_70_2275 ();
 sg13g2_fill_2 FILLER_70_2287 ();
 sg13g2_fill_2 FILLER_70_2307 ();
 sg13g2_fill_1 FILLER_70_2309 ();
 sg13g2_decap_8 FILLER_70_2314 ();
 sg13g2_decap_4 FILLER_70_2321 ();
 sg13g2_decap_8 FILLER_70_2342 ();
 sg13g2_decap_8 FILLER_70_2349 ();
 sg13g2_decap_4 FILLER_70_2356 ();
 sg13g2_fill_2 FILLER_70_2360 ();
 sg13g2_decap_8 FILLER_70_2424 ();
 sg13g2_decap_4 FILLER_70_2439 ();
 sg13g2_fill_1 FILLER_70_2443 ();
 sg13g2_fill_2 FILLER_70_2459 ();
 sg13g2_fill_1 FILLER_70_2461 ();
 sg13g2_fill_2 FILLER_70_2469 ();
 sg13g2_fill_1 FILLER_70_2471 ();
 sg13g2_decap_8 FILLER_70_2478 ();
 sg13g2_decap_8 FILLER_70_2514 ();
 sg13g2_decap_4 FILLER_70_2521 ();
 sg13g2_decap_4 FILLER_70_2528 ();
 sg13g2_fill_1 FILLER_70_2532 ();
 sg13g2_fill_2 FILLER_70_2541 ();
 sg13g2_decap_8 FILLER_70_2547 ();
 sg13g2_fill_1 FILLER_70_2554 ();
 sg13g2_decap_4 FILLER_70_2585 ();
 sg13g2_decap_4 FILLER_70_2593 ();
 sg13g2_decap_8 FILLER_70_2602 ();
 sg13g2_decap_4 FILLER_70_2609 ();
 sg13g2_fill_2 FILLER_70_2613 ();
 sg13g2_fill_1 FILLER_70_2649 ();
 sg13g2_fill_2 FILLER_70_2667 ();
 sg13g2_fill_1 FILLER_70_2669 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_32 ();
 sg13g2_fill_2 FILLER_71_39 ();
 sg13g2_fill_1 FILLER_71_67 ();
 sg13g2_decap_4 FILLER_71_77 ();
 sg13g2_fill_1 FILLER_71_101 ();
 sg13g2_fill_2 FILLER_71_112 ();
 sg13g2_fill_1 FILLER_71_119 ();
 sg13g2_fill_2 FILLER_71_130 ();
 sg13g2_decap_4 FILLER_71_163 ();
 sg13g2_decap_4 FILLER_71_203 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_decap_4 FILLER_71_270 ();
 sg13g2_fill_1 FILLER_71_274 ();
 sg13g2_decap_8 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_292 ();
 sg13g2_decap_8 FILLER_71_299 ();
 sg13g2_decap_8 FILLER_71_306 ();
 sg13g2_decap_8 FILLER_71_313 ();
 sg13g2_decap_8 FILLER_71_320 ();
 sg13g2_decap_8 FILLER_71_327 ();
 sg13g2_decap_8 FILLER_71_334 ();
 sg13g2_decap_8 FILLER_71_341 ();
 sg13g2_decap_8 FILLER_71_348 ();
 sg13g2_decap_8 FILLER_71_355 ();
 sg13g2_fill_1 FILLER_71_377 ();
 sg13g2_fill_1 FILLER_71_382 ();
 sg13g2_fill_1 FILLER_71_399 ();
 sg13g2_decap_8 FILLER_71_409 ();
 sg13g2_fill_1 FILLER_71_481 ();
 sg13g2_fill_1 FILLER_71_487 ();
 sg13g2_decap_8 FILLER_71_497 ();
 sg13g2_decap_8 FILLER_71_504 ();
 sg13g2_decap_8 FILLER_71_511 ();
 sg13g2_decap_8 FILLER_71_518 ();
 sg13g2_decap_8 FILLER_71_525 ();
 sg13g2_decap_4 FILLER_71_532 ();
 sg13g2_fill_1 FILLER_71_536 ();
 sg13g2_fill_1 FILLER_71_542 ();
 sg13g2_fill_1 FILLER_71_549 ();
 sg13g2_fill_2 FILLER_71_560 ();
 sg13g2_decap_8 FILLER_71_598 ();
 sg13g2_fill_1 FILLER_71_605 ();
 sg13g2_decap_4 FILLER_71_616 ();
 sg13g2_decap_4 FILLER_71_624 ();
 sg13g2_decap_8 FILLER_71_654 ();
 sg13g2_decap_8 FILLER_71_661 ();
 sg13g2_decap_4 FILLER_71_668 ();
 sg13g2_fill_1 FILLER_71_698 ();
 sg13g2_decap_4 FILLER_71_712 ();
 sg13g2_decap_8 FILLER_71_742 ();
 sg13g2_decap_4 FILLER_71_749 ();
 sg13g2_fill_2 FILLER_71_753 ();
 sg13g2_decap_8 FILLER_71_764 ();
 sg13g2_fill_2 FILLER_71_771 ();
 sg13g2_fill_1 FILLER_71_773 ();
 sg13g2_decap_4 FILLER_71_840 ();
 sg13g2_fill_1 FILLER_71_856 ();
 sg13g2_fill_2 FILLER_71_862 ();
 sg13g2_fill_2 FILLER_71_925 ();
 sg13g2_fill_1 FILLER_71_927 ();
 sg13g2_fill_1 FILLER_71_966 ();
 sg13g2_decap_4 FILLER_71_1010 ();
 sg13g2_fill_2 FILLER_71_1019 ();
 sg13g2_decap_8 FILLER_71_1095 ();
 sg13g2_fill_2 FILLER_71_1102 ();
 sg13g2_decap_8 FILLER_71_1130 ();
 sg13g2_decap_8 FILLER_71_1137 ();
 sg13g2_decap_4 FILLER_71_1144 ();
 sg13g2_decap_8 FILLER_71_1151 ();
 sg13g2_decap_4 FILLER_71_1158 ();
 sg13g2_fill_2 FILLER_71_1162 ();
 sg13g2_fill_2 FILLER_71_1187 ();
 sg13g2_decap_4 FILLER_71_1192 ();
 sg13g2_fill_1 FILLER_71_1196 ();
 sg13g2_decap_8 FILLER_71_1206 ();
 sg13g2_fill_2 FILLER_71_1213 ();
 sg13g2_decap_4 FILLER_71_1230 ();
 sg13g2_fill_2 FILLER_71_1234 ();
 sg13g2_fill_2 FILLER_71_1262 ();
 sg13g2_fill_1 FILLER_71_1264 ();
 sg13g2_decap_4 FILLER_71_1275 ();
 sg13g2_fill_1 FILLER_71_1279 ();
 sg13g2_fill_2 FILLER_71_1284 ();
 sg13g2_fill_1 FILLER_71_1295 ();
 sg13g2_decap_8 FILLER_71_1326 ();
 sg13g2_fill_1 FILLER_71_1359 ();
 sg13g2_fill_2 FILLER_71_1364 ();
 sg13g2_fill_1 FILLER_71_1366 ();
 sg13g2_fill_2 FILLER_71_1397 ();
 sg13g2_fill_1 FILLER_71_1399 ();
 sg13g2_decap_8 FILLER_71_1504 ();
 sg13g2_fill_1 FILLER_71_1511 ();
 sg13g2_fill_1 FILLER_71_1517 ();
 sg13g2_fill_1 FILLER_71_1537 ();
 sg13g2_fill_1 FILLER_71_1609 ();
 sg13g2_fill_1 FILLER_71_1639 ();
 sg13g2_decap_4 FILLER_71_1667 ();
 sg13g2_fill_2 FILLER_71_1671 ();
 sg13g2_fill_2 FILLER_71_1722 ();
 sg13g2_fill_2 FILLER_71_1729 ();
 sg13g2_fill_2 FILLER_71_1790 ();
 sg13g2_fill_2 FILLER_71_1833 ();
 sg13g2_fill_1 FILLER_71_1843 ();
 sg13g2_fill_2 FILLER_71_1857 ();
 sg13g2_decap_8 FILLER_71_1875 ();
 sg13g2_decap_4 FILLER_71_1882 ();
 sg13g2_fill_1 FILLER_71_1917 ();
 sg13g2_fill_1 FILLER_71_1963 ();
 sg13g2_fill_1 FILLER_71_1988 ();
 sg13g2_fill_2 FILLER_71_2039 ();
 sg13g2_fill_1 FILLER_71_2051 ();
 sg13g2_fill_2 FILLER_71_2078 ();
 sg13g2_fill_1 FILLER_71_2080 ();
 sg13g2_decap_8 FILLER_71_2115 ();
 sg13g2_fill_1 FILLER_71_2122 ();
 sg13g2_fill_1 FILLER_71_2139 ();
 sg13g2_decap_8 FILLER_71_2155 ();
 sg13g2_decap_8 FILLER_71_2162 ();
 sg13g2_decap_4 FILLER_71_2169 ();
 sg13g2_fill_1 FILLER_71_2173 ();
 sg13g2_decap_4 FILLER_71_2178 ();
 sg13g2_fill_1 FILLER_71_2182 ();
 sg13g2_decap_8 FILLER_71_2264 ();
 sg13g2_fill_1 FILLER_71_2271 ();
 sg13g2_fill_2 FILLER_71_2283 ();
 sg13g2_fill_1 FILLER_71_2285 ();
 sg13g2_fill_2 FILLER_71_2297 ();
 sg13g2_fill_1 FILLER_71_2303 ();
 sg13g2_fill_2 FILLER_71_2336 ();
 sg13g2_fill_1 FILLER_71_2338 ();
 sg13g2_fill_2 FILLER_71_2343 ();
 sg13g2_decap_4 FILLER_71_2350 ();
 sg13g2_fill_1 FILLER_71_2354 ();
 sg13g2_decap_8 FILLER_71_2368 ();
 sg13g2_fill_1 FILLER_71_2375 ();
 sg13g2_fill_1 FILLER_71_2380 ();
 sg13g2_fill_2 FILLER_71_2385 ();
 sg13g2_fill_1 FILLER_71_2421 ();
 sg13g2_fill_1 FILLER_71_2454 ();
 sg13g2_decap_8 FILLER_71_2518 ();
 sg13g2_decap_8 FILLER_71_2531 ();
 sg13g2_fill_2 FILLER_71_2538 ();
 sg13g2_decap_8 FILLER_71_2570 ();
 sg13g2_decap_4 FILLER_71_2577 ();
 sg13g2_fill_2 FILLER_71_2581 ();
 sg13g2_decap_8 FILLER_71_2609 ();
 sg13g2_decap_4 FILLER_71_2616 ();
 sg13g2_fill_1 FILLER_71_2656 ();
 sg13g2_decap_8 FILLER_71_2661 ();
 sg13g2_fill_2 FILLER_71_2668 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_73 ();
 sg13g2_fill_2 FILLER_72_79 ();
 sg13g2_fill_1 FILLER_72_81 ();
 sg13g2_decap_8 FILLER_72_102 ();
 sg13g2_decap_8 FILLER_72_109 ();
 sg13g2_decap_8 FILLER_72_116 ();
 sg13g2_decap_4 FILLER_72_123 ();
 sg13g2_fill_1 FILLER_72_161 ();
 sg13g2_fill_1 FILLER_72_172 ();
 sg13g2_fill_1 FILLER_72_199 ();
 sg13g2_decap_8 FILLER_72_226 ();
 sg13g2_fill_1 FILLER_72_233 ();
 sg13g2_fill_2 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_fill_1 FILLER_72_322 ();
 sg13g2_fill_2 FILLER_72_349 ();
 sg13g2_fill_1 FILLER_72_351 ();
 sg13g2_decap_4 FILLER_72_357 ();
 sg13g2_fill_2 FILLER_72_361 ();
 sg13g2_fill_1 FILLER_72_371 ();
 sg13g2_decap_4 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_385 ();
 sg13g2_fill_2 FILLER_72_402 ();
 sg13g2_fill_1 FILLER_72_409 ();
 sg13g2_fill_1 FILLER_72_435 ();
 sg13g2_fill_2 FILLER_72_457 ();
 sg13g2_fill_1 FILLER_72_459 ();
 sg13g2_fill_1 FILLER_72_465 ();
 sg13g2_fill_2 FILLER_72_489 ();
 sg13g2_fill_1 FILLER_72_491 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_504 ();
 sg13g2_decap_8 FILLER_72_511 ();
 sg13g2_decap_8 FILLER_72_518 ();
 sg13g2_decap_4 FILLER_72_577 ();
 sg13g2_fill_2 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_623 ();
 sg13g2_decap_4 FILLER_72_630 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_4 FILLER_72_679 ();
 sg13g2_fill_1 FILLER_72_683 ();
 sg13g2_fill_1 FILLER_72_701 ();
 sg13g2_decap_4 FILLER_72_712 ();
 sg13g2_fill_1 FILLER_72_720 ();
 sg13g2_fill_1 FILLER_72_733 ();
 sg13g2_fill_1 FILLER_72_775 ();
 sg13g2_fill_2 FILLER_72_792 ();
 sg13g2_fill_1 FILLER_72_808 ();
 sg13g2_decap_8 FILLER_72_829 ();
 sg13g2_fill_2 FILLER_72_891 ();
 sg13g2_decap_4 FILLER_72_930 ();
 sg13g2_fill_1 FILLER_72_934 ();
 sg13g2_decap_8 FILLER_72_939 ();
 sg13g2_fill_2 FILLER_72_946 ();
 sg13g2_fill_2 FILLER_72_957 ();
 sg13g2_fill_2 FILLER_72_968 ();
 sg13g2_decap_8 FILLER_72_974 ();
 sg13g2_decap_8 FILLER_72_981 ();
 sg13g2_decap_8 FILLER_72_988 ();
 sg13g2_decap_8 FILLER_72_995 ();
 sg13g2_fill_1 FILLER_72_1002 ();
 sg13g2_fill_2 FILLER_72_1021 ();
 sg13g2_fill_1 FILLER_72_1023 ();
 sg13g2_decap_8 FILLER_72_1033 ();
 sg13g2_fill_2 FILLER_72_1045 ();
 sg13g2_fill_2 FILLER_72_1051 ();
 sg13g2_fill_2 FILLER_72_1057 ();
 sg13g2_fill_1 FILLER_72_1059 ();
 sg13g2_fill_2 FILLER_72_1091 ();
 sg13g2_fill_2 FILLER_72_1119 ();
 sg13g2_decap_8 FILLER_72_1127 ();
 sg13g2_fill_1 FILLER_72_1134 ();
 sg13g2_fill_2 FILLER_72_1195 ();
 sg13g2_fill_1 FILLER_72_1203 ();
 sg13g2_decap_8 FILLER_72_1240 ();
 sg13g2_fill_1 FILLER_72_1265 ();
 sg13g2_decap_8 FILLER_72_1292 ();
 sg13g2_decap_8 FILLER_72_1308 ();
 sg13g2_fill_1 FILLER_72_1315 ();
 sg13g2_fill_2 FILLER_72_1342 ();
 sg13g2_fill_1 FILLER_72_1344 ();
 sg13g2_decap_8 FILLER_72_1349 ();
 sg13g2_decap_4 FILLER_72_1356 ();
 sg13g2_decap_8 FILLER_72_1396 ();
 sg13g2_fill_2 FILLER_72_1403 ();
 sg13g2_fill_1 FILLER_72_1410 ();
 sg13g2_fill_2 FILLER_72_1415 ();
 sg13g2_decap_8 FILLER_72_1421 ();
 sg13g2_fill_2 FILLER_72_1433 ();
 sg13g2_decap_8 FILLER_72_1474 ();
 sg13g2_decap_8 FILLER_72_1481 ();
 sg13g2_fill_2 FILLER_72_1488 ();
 sg13g2_fill_1 FILLER_72_1525 ();
 sg13g2_fill_1 FILLER_72_1561 ();
 sg13g2_fill_2 FILLER_72_1617 ();
 sg13g2_decap_8 FILLER_72_1645 ();
 sg13g2_decap_4 FILLER_72_1652 ();
 sg13g2_fill_2 FILLER_72_1662 ();
 sg13g2_fill_1 FILLER_72_1664 ();
 sg13g2_decap_8 FILLER_72_1713 ();
 sg13g2_fill_2 FILLER_72_1720 ();
 sg13g2_fill_1 FILLER_72_1753 ();
 sg13g2_decap_8 FILLER_72_1775 ();
 sg13g2_fill_1 FILLER_72_1782 ();
 sg13g2_fill_2 FILLER_72_1809 ();
 sg13g2_fill_2 FILLER_72_1853 ();
 sg13g2_fill_1 FILLER_72_1869 ();
 sg13g2_fill_2 FILLER_72_1894 ();
 sg13g2_fill_1 FILLER_72_1908 ();
 sg13g2_fill_1 FILLER_72_1922 ();
 sg13g2_decap_4 FILLER_72_1940 ();
 sg13g2_fill_1 FILLER_72_1944 ();
 sg13g2_fill_1 FILLER_72_2000 ();
 sg13g2_fill_1 FILLER_72_2030 ();
 sg13g2_fill_1 FILLER_72_2057 ();
 sg13g2_decap_4 FILLER_72_2084 ();
 sg13g2_fill_1 FILLER_72_2088 ();
 sg13g2_fill_1 FILLER_72_2093 ();
 sg13g2_decap_8 FILLER_72_2120 ();
 sg13g2_decap_8 FILLER_72_2127 ();
 sg13g2_fill_2 FILLER_72_2134 ();
 sg13g2_fill_1 FILLER_72_2136 ();
 sg13g2_decap_4 FILLER_72_2142 ();
 sg13g2_fill_1 FILLER_72_2146 ();
 sg13g2_decap_8 FILLER_72_2173 ();
 sg13g2_decap_8 FILLER_72_2180 ();
 sg13g2_decap_8 FILLER_72_2187 ();
 sg13g2_decap_8 FILLER_72_2194 ();
 sg13g2_decap_8 FILLER_72_2201 ();
 sg13g2_decap_4 FILLER_72_2208 ();
 sg13g2_decap_8 FILLER_72_2242 ();
 sg13g2_decap_8 FILLER_72_2249 ();
 sg13g2_fill_2 FILLER_72_2262 ();
 sg13g2_decap_4 FILLER_72_2269 ();
 sg13g2_fill_1 FILLER_72_2273 ();
 sg13g2_decap_8 FILLER_72_2300 ();
 sg13g2_decap_8 FILLER_72_2307 ();
 sg13g2_decap_8 FILLER_72_2314 ();
 sg13g2_decap_8 FILLER_72_2321 ();
 sg13g2_decap_8 FILLER_72_2328 ();
 sg13g2_decap_4 FILLER_72_2335 ();
 sg13g2_decap_4 FILLER_72_2369 ();
 sg13g2_decap_8 FILLER_72_2377 ();
 sg13g2_decap_8 FILLER_72_2384 ();
 sg13g2_fill_2 FILLER_72_2391 ();
 sg13g2_fill_1 FILLER_72_2400 ();
 sg13g2_fill_1 FILLER_72_2405 ();
 sg13g2_fill_1 FILLER_72_2410 ();
 sg13g2_fill_1 FILLER_72_2415 ();
 sg13g2_fill_2 FILLER_72_2446 ();
 sg13g2_fill_2 FILLER_72_2480 ();
 sg13g2_decap_4 FILLER_72_2498 ();
 sg13g2_decap_8 FILLER_72_2506 ();
 sg13g2_decap_8 FILLER_72_2513 ();
 sg13g2_fill_2 FILLER_72_2523 ();
 sg13g2_fill_1 FILLER_72_2525 ();
 sg13g2_decap_4 FILLER_72_2532 ();
 sg13g2_decap_8 FILLER_72_2566 ();
 sg13g2_decap_8 FILLER_72_2573 ();
 sg13g2_fill_1 FILLER_72_2580 ();
 sg13g2_decap_8 FILLER_72_2606 ();
 sg13g2_decap_8 FILLER_72_2613 ();
 sg13g2_decap_8 FILLER_72_2620 ();
 sg13g2_fill_2 FILLER_72_2627 ();
 sg13g2_fill_2 FILLER_72_2633 ();
 sg13g2_fill_1 FILLER_72_2635 ();
 sg13g2_decap_8 FILLER_72_2655 ();
 sg13g2_decap_8 FILLER_72_2662 ();
 sg13g2_fill_1 FILLER_72_2669 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_4 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_11 ();
 sg13g2_fill_2 FILLER_73_23 ();
 sg13g2_fill_1 FILLER_73_25 ();
 sg13g2_fill_2 FILLER_73_33 ();
 sg13g2_fill_1 FILLER_73_35 ();
 sg13g2_fill_1 FILLER_73_94 ();
 sg13g2_fill_2 FILLER_73_105 ();
 sg13g2_decap_8 FILLER_73_120 ();
 sg13g2_decap_8 FILLER_73_127 ();
 sg13g2_decap_8 FILLER_73_134 ();
 sg13g2_decap_8 FILLER_73_141 ();
 sg13g2_decap_8 FILLER_73_148 ();
 sg13g2_decap_8 FILLER_73_155 ();
 sg13g2_decap_8 FILLER_73_162 ();
 sg13g2_fill_2 FILLER_73_169 ();
 sg13g2_fill_1 FILLER_73_171 ();
 sg13g2_decap_8 FILLER_73_196 ();
 sg13g2_decap_8 FILLER_73_203 ();
 sg13g2_decap_8 FILLER_73_210 ();
 sg13g2_fill_2 FILLER_73_217 ();
 sg13g2_fill_1 FILLER_73_219 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_decap_8 FILLER_73_277 ();
 sg13g2_decap_8 FILLER_73_284 ();
 sg13g2_decap_8 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_298 ();
 sg13g2_decap_4 FILLER_73_305 ();
 sg13g2_fill_2 FILLER_73_309 ();
 sg13g2_decap_8 FILLER_73_321 ();
 sg13g2_decap_4 FILLER_73_328 ();
 sg13g2_fill_2 FILLER_73_332 ();
 sg13g2_fill_2 FILLER_73_365 ();
 sg13g2_decap_8 FILLER_73_405 ();
 sg13g2_fill_2 FILLER_73_424 ();
 sg13g2_fill_2 FILLER_73_482 ();
 sg13g2_fill_1 FILLER_73_484 ();
 sg13g2_fill_1 FILLER_73_490 ();
 sg13g2_fill_2 FILLER_73_496 ();
 sg13g2_fill_1 FILLER_73_537 ();
 sg13g2_fill_1 FILLER_73_549 ();
 sg13g2_fill_2 FILLER_73_555 ();
 sg13g2_fill_1 FILLER_73_557 ();
 sg13g2_decap_8 FILLER_73_563 ();
 sg13g2_fill_2 FILLER_73_570 ();
 sg13g2_fill_1 FILLER_73_572 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_fill_2 FILLER_73_599 ();
 sg13g2_decap_4 FILLER_73_605 ();
 sg13g2_fill_2 FILLER_73_613 ();
 sg13g2_fill_1 FILLER_73_615 ();
 sg13g2_fill_2 FILLER_73_662 ();
 sg13g2_fill_1 FILLER_73_664 ();
 sg13g2_fill_1 FILLER_73_730 ();
 sg13g2_decap_8 FILLER_73_749 ();
 sg13g2_decap_4 FILLER_73_756 ();
 sg13g2_fill_2 FILLER_73_760 ();
 sg13g2_fill_1 FILLER_73_788 ();
 sg13g2_fill_2 FILLER_73_803 ();
 sg13g2_fill_2 FILLER_73_810 ();
 sg13g2_decap_8 FILLER_73_838 ();
 sg13g2_decap_4 FILLER_73_845 ();
 sg13g2_fill_1 FILLER_73_849 ();
 sg13g2_fill_2 FILLER_73_879 ();
 sg13g2_fill_1 FILLER_73_887 ();
 sg13g2_fill_1 FILLER_73_897 ();
 sg13g2_fill_2 FILLER_73_909 ();
 sg13g2_decap_8 FILLER_73_973 ();
 sg13g2_fill_2 FILLER_73_980 ();
 sg13g2_fill_1 FILLER_73_982 ();
 sg13g2_fill_2 FILLER_73_989 ();
 sg13g2_fill_1 FILLER_73_991 ();
 sg13g2_fill_2 FILLER_73_1049 ();
 sg13g2_fill_1 FILLER_73_1051 ();
 sg13g2_fill_2 FILLER_73_1087 ();
 sg13g2_fill_1 FILLER_73_1089 ();
 sg13g2_fill_2 FILLER_73_1094 ();
 sg13g2_fill_1 FILLER_73_1096 ();
 sg13g2_decap_8 FILLER_73_1102 ();
 sg13g2_decap_4 FILLER_73_1109 ();
 sg13g2_fill_2 FILLER_73_1113 ();
 sg13g2_decap_4 FILLER_73_1119 ();
 sg13g2_fill_1 FILLER_73_1164 ();
 sg13g2_fill_2 FILLER_73_1172 ();
 sg13g2_fill_2 FILLER_73_1178 ();
 sg13g2_fill_2 FILLER_73_1223 ();
 sg13g2_fill_1 FILLER_73_1225 ();
 sg13g2_decap_8 FILLER_73_1232 ();
 sg13g2_fill_2 FILLER_73_1239 ();
 sg13g2_fill_2 FILLER_73_1267 ();
 sg13g2_fill_1 FILLER_73_1287 ();
 sg13g2_fill_2 FILLER_73_1296 ();
 sg13g2_fill_1 FILLER_73_1298 ();
 sg13g2_decap_4 FILLER_73_1340 ();
 sg13g2_fill_2 FILLER_73_1349 ();
 sg13g2_decap_4 FILLER_73_1362 ();
 sg13g2_fill_2 FILLER_73_1366 ();
 sg13g2_fill_1 FILLER_73_1405 ();
 sg13g2_decap_8 FILLER_73_1410 ();
 sg13g2_decap_8 FILLER_73_1417 ();
 sg13g2_decap_8 FILLER_73_1424 ();
 sg13g2_fill_2 FILLER_73_1431 ();
 sg13g2_fill_2 FILLER_73_1464 ();
 sg13g2_fill_2 FILLER_73_1497 ();
 sg13g2_fill_1 FILLER_73_1525 ();
 sg13g2_fill_2 FILLER_73_1530 ();
 sg13g2_fill_1 FILLER_73_1541 ();
 sg13g2_fill_1 FILLER_73_1558 ();
 sg13g2_fill_2 FILLER_73_1606 ();
 sg13g2_fill_1 FILLER_73_1660 ();
 sg13g2_decap_4 FILLER_73_1665 ();
 sg13g2_fill_2 FILLER_73_1669 ();
 sg13g2_fill_2 FILLER_73_1676 ();
 sg13g2_decap_4 FILLER_73_1688 ();
 sg13g2_fill_1 FILLER_73_1692 ();
 sg13g2_decap_8 FILLER_73_1697 ();
 sg13g2_decap_8 FILLER_73_1704 ();
 sg13g2_fill_1 FILLER_73_1711 ();
 sg13g2_fill_1 FILLER_73_1717 ();
 sg13g2_fill_1 FILLER_73_1748 ();
 sg13g2_fill_2 FILLER_73_1768 ();
 sg13g2_decap_8 FILLER_73_1777 ();
 sg13g2_decap_8 FILLER_73_1784 ();
 sg13g2_fill_1 FILLER_73_1791 ();
 sg13g2_decap_4 FILLER_73_1801 ();
 sg13g2_fill_1 FILLER_73_1805 ();
 sg13g2_decap_4 FILLER_73_1809 ();
 sg13g2_fill_2 FILLER_73_1813 ();
 sg13g2_fill_2 FILLER_73_1823 ();
 sg13g2_decap_8 FILLER_73_1864 ();
 sg13g2_decap_4 FILLER_73_1871 ();
 sg13g2_fill_1 FILLER_73_1885 ();
 sg13g2_fill_2 FILLER_73_1920 ();
 sg13g2_fill_2 FILLER_73_1930 ();
 sg13g2_fill_1 FILLER_73_1932 ();
 sg13g2_fill_2 FILLER_73_1938 ();
 sg13g2_fill_1 FILLER_73_1940 ();
 sg13g2_decap_4 FILLER_73_1945 ();
 sg13g2_fill_2 FILLER_73_1949 ();
 sg13g2_fill_1 FILLER_73_1962 ();
 sg13g2_fill_2 FILLER_73_1967 ();
 sg13g2_fill_1 FILLER_73_2009 ();
 sg13g2_decap_8 FILLER_73_2019 ();
 sg13g2_fill_2 FILLER_73_2026 ();
 sg13g2_fill_1 FILLER_73_2028 ();
 sg13g2_fill_2 FILLER_73_2033 ();
 sg13g2_decap_4 FILLER_73_2040 ();
 sg13g2_decap_8 FILLER_73_2058 ();
 sg13g2_decap_8 FILLER_73_2065 ();
 sg13g2_fill_1 FILLER_73_2076 ();
 sg13g2_fill_1 FILLER_73_2111 ();
 sg13g2_decap_4 FILLER_73_2190 ();
 sg13g2_fill_2 FILLER_73_2194 ();
 sg13g2_fill_2 FILLER_73_2201 ();
 sg13g2_fill_1 FILLER_73_2203 ();
 sg13g2_decap_4 FILLER_73_2210 ();
 sg13g2_fill_1 FILLER_73_2214 ();
 sg13g2_fill_1 FILLER_73_2221 ();
 sg13g2_fill_2 FILLER_73_2226 ();
 sg13g2_fill_2 FILLER_73_2250 ();
 sg13g2_fill_1 FILLER_73_2252 ();
 sg13g2_fill_2 FILLER_73_2291 ();
 sg13g2_fill_1 FILLER_73_2293 ();
 sg13g2_fill_2 FILLER_73_2320 ();
 sg13g2_fill_1 FILLER_73_2322 ();
 sg13g2_fill_1 FILLER_73_2349 ();
 sg13g2_decap_4 FILLER_73_2458 ();
 sg13g2_decap_8 FILLER_73_2470 ();
 sg13g2_decap_8 FILLER_73_2477 ();
 sg13g2_fill_2 FILLER_73_2484 ();
 sg13g2_decap_4 FILLER_73_2496 ();
 sg13g2_fill_2 FILLER_73_2506 ();
 sg13g2_fill_2 FILLER_73_2529 ();
 sg13g2_decap_8 FILLER_73_2565 ();
 sg13g2_decap_4 FILLER_73_2572 ();
 sg13g2_fill_1 FILLER_73_2576 ();
 sg13g2_decap_8 FILLER_73_2612 ();
 sg13g2_decap_4 FILLER_73_2619 ();
 sg13g2_decap_8 FILLER_73_2650 ();
 sg13g2_decap_8 FILLER_73_2657 ();
 sg13g2_decap_4 FILLER_73_2664 ();
 sg13g2_fill_2 FILLER_73_2668 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_4 FILLER_74_7 ();
 sg13g2_fill_1 FILLER_74_11 ();
 sg13g2_fill_2 FILLER_74_47 ();
 sg13g2_fill_1 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_68 ();
 sg13g2_decap_8 FILLER_74_104 ();
 sg13g2_fill_1 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_142 ();
 sg13g2_decap_8 FILLER_74_154 ();
 sg13g2_decap_8 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_168 ();
 sg13g2_decap_4 FILLER_74_175 ();
 sg13g2_fill_2 FILLER_74_179 ();
 sg13g2_decap_8 FILLER_74_207 ();
 sg13g2_decap_8 FILLER_74_214 ();
 sg13g2_decap_8 FILLER_74_221 ();
 sg13g2_decap_8 FILLER_74_268 ();
 sg13g2_decap_8 FILLER_74_279 ();
 sg13g2_fill_2 FILLER_74_286 ();
 sg13g2_fill_1 FILLER_74_288 ();
 sg13g2_fill_2 FILLER_74_292 ();
 sg13g2_decap_8 FILLER_74_311 ();
 sg13g2_decap_8 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_325 ();
 sg13g2_fill_2 FILLER_74_358 ();
 sg13g2_fill_2 FILLER_74_370 ();
 sg13g2_fill_1 FILLER_74_372 ();
 sg13g2_fill_2 FILLER_74_406 ();
 sg13g2_fill_1 FILLER_74_487 ();
 sg13g2_decap_8 FILLER_74_523 ();
 sg13g2_decap_4 FILLER_74_530 ();
 sg13g2_fill_2 FILLER_74_534 ();
 sg13g2_decap_4 FILLER_74_548 ();
 sg13g2_fill_1 FILLER_74_552 ();
 sg13g2_decap_8 FILLER_74_561 ();
 sg13g2_decap_8 FILLER_74_568 ();
 sg13g2_decap_8 FILLER_74_575 ();
 sg13g2_decap_8 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_589 ();
 sg13g2_decap_8 FILLER_74_596 ();
 sg13g2_fill_2 FILLER_74_603 ();
 sg13g2_fill_1 FILLER_74_627 ();
 sg13g2_fill_2 FILLER_74_657 ();
 sg13g2_fill_2 FILLER_74_666 ();
 sg13g2_fill_1 FILLER_74_707 ();
 sg13g2_decap_4 FILLER_74_718 ();
 sg13g2_fill_2 FILLER_74_722 ();
 sg13g2_decap_8 FILLER_74_768 ();
 sg13g2_decap_8 FILLER_74_775 ();
 sg13g2_decap_4 FILLER_74_782 ();
 sg13g2_fill_1 FILLER_74_786 ();
 sg13g2_decap_8 FILLER_74_796 ();
 sg13g2_decap_4 FILLER_74_803 ();
 sg13g2_fill_1 FILLER_74_812 ();
 sg13g2_decap_8 FILLER_74_817 ();
 sg13g2_decap_4 FILLER_74_824 ();
 sg13g2_fill_1 FILLER_74_834 ();
 sg13g2_fill_2 FILLER_74_856 ();
 sg13g2_fill_2 FILLER_74_862 ();
 sg13g2_fill_2 FILLER_74_879 ();
 sg13g2_fill_1 FILLER_74_896 ();
 sg13g2_decap_8 FILLER_74_914 ();
 sg13g2_fill_1 FILLER_74_921 ();
 sg13g2_decap_8 FILLER_74_948 ();
 sg13g2_fill_1 FILLER_74_955 ();
 sg13g2_fill_2 FILLER_74_969 ();
 sg13g2_fill_1 FILLER_74_971 ();
 sg13g2_decap_8 FILLER_74_976 ();
 sg13g2_decap_8 FILLER_74_983 ();
 sg13g2_decap_8 FILLER_74_990 ();
 sg13g2_decap_8 FILLER_74_997 ();
 sg13g2_fill_2 FILLER_74_1004 ();
 sg13g2_fill_1 FILLER_74_1006 ();
 sg13g2_decap_4 FILLER_74_1028 ();
 sg13g2_decap_8 FILLER_74_1039 ();
 sg13g2_decap_8 FILLER_74_1046 ();
 sg13g2_decap_8 FILLER_74_1053 ();
 sg13g2_decap_8 FILLER_74_1060 ();
 sg13g2_decap_4 FILLER_74_1067 ();
 sg13g2_fill_1 FILLER_74_1071 ();
 sg13g2_fill_1 FILLER_74_1150 ();
 sg13g2_fill_2 FILLER_74_1156 ();
 sg13g2_decap_4 FILLER_74_1169 ();
 sg13g2_fill_1 FILLER_74_1173 ();
 sg13g2_decap_8 FILLER_74_1179 ();
 sg13g2_decap_8 FILLER_74_1186 ();
 sg13g2_decap_8 FILLER_74_1193 ();
 sg13g2_decap_8 FILLER_74_1200 ();
 sg13g2_fill_1 FILLER_74_1207 ();
 sg13g2_fill_2 FILLER_74_1212 ();
 sg13g2_fill_1 FILLER_74_1225 ();
 sg13g2_decap_4 FILLER_74_1232 ();
 sg13g2_fill_1 FILLER_74_1236 ();
 sg13g2_decap_8 FILLER_74_1243 ();
 sg13g2_decap_4 FILLER_74_1250 ();
 sg13g2_fill_2 FILLER_74_1254 ();
 sg13g2_fill_2 FILLER_74_1270 ();
 sg13g2_decap_4 FILLER_74_1298 ();
 sg13g2_decap_8 FILLER_74_1308 ();
 sg13g2_decap_8 FILLER_74_1315 ();
 sg13g2_decap_8 FILLER_74_1322 ();
 sg13g2_decap_8 FILLER_74_1329 ();
 sg13g2_decap_8 FILLER_74_1336 ();
 sg13g2_decap_8 FILLER_74_1381 ();
 sg13g2_decap_8 FILLER_74_1388 ();
 sg13g2_fill_1 FILLER_74_1395 ();
 sg13g2_decap_8 FILLER_74_1403 ();
 sg13g2_fill_2 FILLER_74_1410 ();
 sg13g2_fill_1 FILLER_74_1412 ();
 sg13g2_fill_2 FILLER_74_1417 ();
 sg13g2_fill_1 FILLER_74_1419 ();
 sg13g2_decap_8 FILLER_74_1426 ();
 sg13g2_decap_8 FILLER_74_1433 ();
 sg13g2_decap_8 FILLER_74_1440 ();
 sg13g2_decap_8 FILLER_74_1447 ();
 sg13g2_decap_8 FILLER_74_1454 ();
 sg13g2_decap_8 FILLER_74_1461 ();
 sg13g2_decap_8 FILLER_74_1468 ();
 sg13g2_fill_2 FILLER_74_1475 ();
 sg13g2_fill_1 FILLER_74_1477 ();
 sg13g2_decap_8 FILLER_74_1483 ();
 sg13g2_fill_2 FILLER_74_1490 ();
 sg13g2_decap_8 FILLER_74_1496 ();
 sg13g2_decap_8 FILLER_74_1503 ();
 sg13g2_decap_8 FILLER_74_1510 ();
 sg13g2_decap_8 FILLER_74_1517 ();
 sg13g2_decap_8 FILLER_74_1524 ();
 sg13g2_fill_1 FILLER_74_1531 ();
 sg13g2_fill_2 FILLER_74_1544 ();
 sg13g2_fill_2 FILLER_74_1553 ();
 sg13g2_decap_8 FILLER_74_1593 ();
 sg13g2_fill_1 FILLER_74_1600 ();
 sg13g2_fill_1 FILLER_74_1608 ();
 sg13g2_fill_2 FILLER_74_1638 ();
 sg13g2_fill_1 FILLER_74_1655 ();
 sg13g2_decap_8 FILLER_74_1670 ();
 sg13g2_decap_8 FILLER_74_1677 ();
 sg13g2_decap_8 FILLER_74_1684 ();
 sg13g2_decap_4 FILLER_74_1691 ();
 sg13g2_fill_1 FILLER_74_1695 ();
 sg13g2_decap_8 FILLER_74_1700 ();
 sg13g2_decap_8 FILLER_74_1707 ();
 sg13g2_fill_2 FILLER_74_1714 ();
 sg13g2_fill_1 FILLER_74_1716 ();
 sg13g2_fill_2 FILLER_74_1720 ();
 sg13g2_fill_1 FILLER_74_1722 ();
 sg13g2_fill_2 FILLER_74_1728 ();
 sg13g2_fill_1 FILLER_74_1730 ();
 sg13g2_decap_4 FILLER_74_1735 ();
 sg13g2_decap_4 FILLER_74_1769 ();
 sg13g2_fill_1 FILLER_74_1773 ();
 sg13g2_decap_8 FILLER_74_1800 ();
 sg13g2_decap_8 FILLER_74_1807 ();
 sg13g2_decap_8 FILLER_74_1814 ();
 sg13g2_decap_4 FILLER_74_1828 ();
 sg13g2_fill_1 FILLER_74_1832 ();
 sg13g2_decap_8 FILLER_74_1859 ();
 sg13g2_fill_2 FILLER_74_1866 ();
 sg13g2_decap_4 FILLER_74_1873 ();
 sg13g2_decap_4 FILLER_74_1886 ();
 sg13g2_fill_1 FILLER_74_1890 ();
 sg13g2_decap_4 FILLER_74_1921 ();
 sg13g2_fill_2 FILLER_74_1925 ();
 sg13g2_decap_4 FILLER_74_1979 ();
 sg13g2_fill_1 FILLER_74_1983 ();
 sg13g2_fill_2 FILLER_74_2036 ();
 sg13g2_decap_4 FILLER_74_2073 ();
 sg13g2_decap_4 FILLER_74_2081 ();
 sg13g2_fill_1 FILLER_74_2085 ();
 sg13g2_fill_1 FILLER_74_2107 ();
 sg13g2_fill_2 FILLER_74_2138 ();
 sg13g2_fill_1 FILLER_74_2140 ();
 sg13g2_fill_1 FILLER_74_2145 ();
 sg13g2_fill_2 FILLER_74_2151 ();
 sg13g2_fill_2 FILLER_74_2157 ();
 sg13g2_fill_2 FILLER_74_2164 ();
 sg13g2_decap_8 FILLER_74_2192 ();
 sg13g2_decap_8 FILLER_74_2199 ();
 sg13g2_decap_8 FILLER_74_2214 ();
 sg13g2_decap_8 FILLER_74_2221 ();
 sg13g2_decap_8 FILLER_74_2228 ();
 sg13g2_fill_2 FILLER_74_2235 ();
 sg13g2_decap_4 FILLER_74_2244 ();
 sg13g2_fill_2 FILLER_74_2248 ();
 sg13g2_decap_8 FILLER_74_2280 ();
 sg13g2_decap_8 FILLER_74_2287 ();
 sg13g2_decap_8 FILLER_74_2294 ();
 sg13g2_fill_1 FILLER_74_2301 ();
 sg13g2_decap_8 FILLER_74_2306 ();
 sg13g2_fill_2 FILLER_74_2313 ();
 sg13g2_fill_1 FILLER_74_2315 ();
 sg13g2_fill_1 FILLER_74_2346 ();
 sg13g2_decap_4 FILLER_74_2425 ();
 sg13g2_fill_1 FILLER_74_2429 ();
 sg13g2_decap_8 FILLER_74_2471 ();
 sg13g2_fill_2 FILLER_74_2478 ();
 sg13g2_fill_1 FILLER_74_2480 ();
 sg13g2_decap_8 FILLER_74_2557 ();
 sg13g2_decap_8 FILLER_74_2564 ();
 sg13g2_decap_8 FILLER_74_2571 ();
 sg13g2_decap_4 FILLER_74_2578 ();
 sg13g2_fill_2 FILLER_74_2595 ();
 sg13g2_decap_8 FILLER_74_2622 ();
 sg13g2_fill_2 FILLER_74_2668 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_4 FILLER_75_21 ();
 sg13g2_fill_1 FILLER_75_25 ();
 sg13g2_decap_8 FILLER_75_46 ();
 sg13g2_fill_2 FILLER_75_53 ();
 sg13g2_decap_8 FILLER_75_65 ();
 sg13g2_decap_8 FILLER_75_72 ();
 sg13g2_fill_2 FILLER_75_79 ();
 sg13g2_fill_1 FILLER_75_81 ();
 sg13g2_decap_8 FILLER_75_92 ();
 sg13g2_decap_8 FILLER_75_99 ();
 sg13g2_decap_8 FILLER_75_106 ();
 sg13g2_decap_4 FILLER_75_113 ();
 sg13g2_fill_1 FILLER_75_117 ();
 sg13g2_decap_4 FILLER_75_123 ();
 sg13g2_fill_1 FILLER_75_164 ();
 sg13g2_fill_1 FILLER_75_180 ();
 sg13g2_decap_8 FILLER_75_191 ();
 sg13g2_decap_8 FILLER_75_198 ();
 sg13g2_decap_8 FILLER_75_205 ();
 sg13g2_decap_8 FILLER_75_212 ();
 sg13g2_decap_8 FILLER_75_219 ();
 sg13g2_decap_8 FILLER_75_226 ();
 sg13g2_decap_4 FILLER_75_233 ();
 sg13g2_fill_2 FILLER_75_237 ();
 sg13g2_decap_8 FILLER_75_243 ();
 sg13g2_decap_4 FILLER_75_250 ();
 sg13g2_fill_1 FILLER_75_254 ();
 sg13g2_fill_2 FILLER_75_271 ();
 sg13g2_fill_2 FILLER_75_309 ();
 sg13g2_decap_8 FILLER_75_321 ();
 sg13g2_fill_2 FILLER_75_354 ();
 sg13g2_decap_8 FILLER_75_360 ();
 sg13g2_fill_2 FILLER_75_367 ();
 sg13g2_decap_4 FILLER_75_381 ();
 sg13g2_fill_2 FILLER_75_385 ();
 sg13g2_fill_1 FILLER_75_399 ();
 sg13g2_decap_4 FILLER_75_403 ();
 sg13g2_decap_8 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_75_418 ();
 sg13g2_decap_8 FILLER_75_425 ();
 sg13g2_decap_8 FILLER_75_432 ();
 sg13g2_decap_4 FILLER_75_439 ();
 sg13g2_fill_2 FILLER_75_443 ();
 sg13g2_fill_1 FILLER_75_450 ();
 sg13g2_decap_4 FILLER_75_455 ();
 sg13g2_fill_2 FILLER_75_459 ();
 sg13g2_decap_8 FILLER_75_471 ();
 sg13g2_decap_8 FILLER_75_478 ();
 sg13g2_fill_2 FILLER_75_485 ();
 sg13g2_decap_8 FILLER_75_491 ();
 sg13g2_fill_2 FILLER_75_498 ();
 sg13g2_fill_2 FILLER_75_515 ();
 sg13g2_fill_1 FILLER_75_517 ();
 sg13g2_decap_8 FILLER_75_523 ();
 sg13g2_decap_8 FILLER_75_530 ();
 sg13g2_decap_4 FILLER_75_537 ();
 sg13g2_fill_1 FILLER_75_541 ();
 sg13g2_fill_1 FILLER_75_555 ();
 sg13g2_fill_2 FILLER_75_572 ();
 sg13g2_decap_8 FILLER_75_600 ();
 sg13g2_decap_4 FILLER_75_607 ();
 sg13g2_fill_2 FILLER_75_611 ();
 sg13g2_decap_4 FILLER_75_657 ();
 sg13g2_fill_2 FILLER_75_661 ();
 sg13g2_decap_8 FILLER_75_671 ();
 sg13g2_decap_4 FILLER_75_678 ();
 sg13g2_fill_1 FILLER_75_682 ();
 sg13g2_fill_2 FILLER_75_713 ();
 sg13g2_decap_8 FILLER_75_741 ();
 sg13g2_decap_4 FILLER_75_748 ();
 sg13g2_fill_1 FILLER_75_752 ();
 sg13g2_decap_8 FILLER_75_762 ();
 sg13g2_fill_1 FILLER_75_769 ();
 sg13g2_decap_8 FILLER_75_775 ();
 sg13g2_fill_2 FILLER_75_782 ();
 sg13g2_fill_1 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_789 ();
 sg13g2_fill_2 FILLER_75_796 ();
 sg13g2_decap_8 FILLER_75_824 ();
 sg13g2_decap_8 FILLER_75_831 ();
 sg13g2_decap_8 FILLER_75_838 ();
 sg13g2_decap_8 FILLER_75_845 ();
 sg13g2_decap_4 FILLER_75_852 ();
 sg13g2_fill_2 FILLER_75_871 ();
 sg13g2_fill_1 FILLER_75_890 ();
 sg13g2_fill_2 FILLER_75_898 ();
 sg13g2_fill_2 FILLER_75_909 ();
 sg13g2_decap_8 FILLER_75_917 ();
 sg13g2_decap_8 FILLER_75_924 ();
 sg13g2_decap_4 FILLER_75_931 ();
 sg13g2_decap_8 FILLER_75_938 ();
 sg13g2_fill_2 FILLER_75_945 ();
 sg13g2_fill_1 FILLER_75_947 ();
 sg13g2_decap_8 FILLER_75_1006 ();
 sg13g2_decap_8 FILLER_75_1013 ();
 sg13g2_fill_1 FILLER_75_1020 ();
 sg13g2_decap_8 FILLER_75_1041 ();
 sg13g2_decap_4 FILLER_75_1048 ();
 sg13g2_decap_8 FILLER_75_1056 ();
 sg13g2_decap_8 FILLER_75_1063 ();
 sg13g2_decap_8 FILLER_75_1070 ();
 sg13g2_decap_4 FILLER_75_1077 ();
 sg13g2_fill_2 FILLER_75_1081 ();
 sg13g2_fill_2 FILLER_75_1088 ();
 sg13g2_fill_1 FILLER_75_1094 ();
 sg13g2_decap_8 FILLER_75_1104 ();
 sg13g2_fill_2 FILLER_75_1116 ();
 sg13g2_decap_8 FILLER_75_1126 ();
 sg13g2_decap_8 FILLER_75_1133 ();
 sg13g2_decap_8 FILLER_75_1140 ();
 sg13g2_decap_4 FILLER_75_1153 ();
 sg13g2_decap_8 FILLER_75_1161 ();
 sg13g2_fill_2 FILLER_75_1168 ();
 sg13g2_decap_8 FILLER_75_1202 ();
 sg13g2_decap_8 FILLER_75_1209 ();
 sg13g2_decap_8 FILLER_75_1216 ();
 sg13g2_fill_2 FILLER_75_1223 ();
 sg13g2_decap_8 FILLER_75_1235 ();
 sg13g2_decap_8 FILLER_75_1242 ();
 sg13g2_decap_4 FILLER_75_1249 ();
 sg13g2_fill_2 FILLER_75_1253 ();
 sg13g2_decap_8 FILLER_75_1286 ();
 sg13g2_decap_8 FILLER_75_1293 ();
 sg13g2_decap_8 FILLER_75_1300 ();
 sg13g2_decap_4 FILLER_75_1307 ();
 sg13g2_fill_1 FILLER_75_1324 ();
 sg13g2_fill_1 FILLER_75_1351 ();
 sg13g2_fill_2 FILLER_75_1385 ();
 sg13g2_fill_1 FILLER_75_1390 ();
 sg13g2_fill_2 FILLER_75_1394 ();
 sg13g2_fill_2 FILLER_75_1414 ();
 sg13g2_fill_1 FILLER_75_1416 ();
 sg13g2_decap_8 FILLER_75_1443 ();
 sg13g2_decap_8 FILLER_75_1450 ();
 sg13g2_decap_8 FILLER_75_1457 ();
 sg13g2_decap_8 FILLER_75_1464 ();
 sg13g2_fill_1 FILLER_75_1471 ();
 sg13g2_decap_8 FILLER_75_1501 ();
 sg13g2_decap_8 FILLER_75_1508 ();
 sg13g2_decap_8 FILLER_75_1515 ();
 sg13g2_decap_8 FILLER_75_1522 ();
 sg13g2_decap_4 FILLER_75_1529 ();
 sg13g2_decap_4 FILLER_75_1559 ();
 sg13g2_fill_1 FILLER_75_1563 ();
 sg13g2_decap_4 FILLER_75_1568 ();
 sg13g2_fill_1 FILLER_75_1575 ();
 sg13g2_fill_2 FILLER_75_1581 ();
 sg13g2_decap_4 FILLER_75_1587 ();
 sg13g2_fill_2 FILLER_75_1595 ();
 sg13g2_fill_1 FILLER_75_1602 ();
 sg13g2_fill_2 FILLER_75_1607 ();
 sg13g2_fill_1 FILLER_75_1609 ();
 sg13g2_decap_8 FILLER_75_1614 ();
 sg13g2_decap_4 FILLER_75_1621 ();
 sg13g2_fill_2 FILLER_75_1642 ();
 sg13g2_fill_1 FILLER_75_1678 ();
 sg13g2_decap_4 FILLER_75_1684 ();
 sg13g2_fill_2 FILLER_75_1688 ();
 sg13g2_fill_2 FILLER_75_1701 ();
 sg13g2_fill_1 FILLER_75_1703 ();
 sg13g2_fill_2 FILLER_75_1709 ();
 sg13g2_fill_1 FILLER_75_1711 ();
 sg13g2_fill_1 FILLER_75_1716 ();
 sg13g2_fill_2 FILLER_75_1720 ();
 sg13g2_fill_1 FILLER_75_1722 ();
 sg13g2_fill_1 FILLER_75_1728 ();
 sg13g2_decap_4 FILLER_75_1755 ();
 sg13g2_fill_2 FILLER_75_1759 ();
 sg13g2_fill_1 FILLER_75_1795 ();
 sg13g2_decap_4 FILLER_75_1800 ();
 sg13g2_fill_2 FILLER_75_1835 ();
 sg13g2_fill_1 FILLER_75_1837 ();
 sg13g2_fill_2 FILLER_75_1895 ();
 sg13g2_fill_1 FILLER_75_1897 ();
 sg13g2_decap_4 FILLER_75_1908 ();
 sg13g2_fill_1 FILLER_75_1912 ();
 sg13g2_decap_4 FILLER_75_1926 ();
 sg13g2_fill_2 FILLER_75_1930 ();
 sg13g2_decap_8 FILLER_75_1988 ();
 sg13g2_decap_8 FILLER_75_1995 ();
 sg13g2_decap_8 FILLER_75_2002 ();
 sg13g2_decap_4 FILLER_75_2009 ();
 sg13g2_decap_4 FILLER_75_2021 ();
 sg13g2_fill_1 FILLER_75_2025 ();
 sg13g2_decap_4 FILLER_75_2030 ();
 sg13g2_fill_1 FILLER_75_2034 ();
 sg13g2_fill_1 FILLER_75_2040 ();
 sg13g2_decap_8 FILLER_75_2070 ();
 sg13g2_decap_8 FILLER_75_2077 ();
 sg13g2_fill_2 FILLER_75_2084 ();
 sg13g2_decap_8 FILLER_75_2091 ();
 sg13g2_fill_1 FILLER_75_2098 ();
 sg13g2_decap_8 FILLER_75_2114 ();
 sg13g2_decap_8 FILLER_75_2121 ();
 sg13g2_decap_8 FILLER_75_2128 ();
 sg13g2_decap_8 FILLER_75_2139 ();
 sg13g2_decap_8 FILLER_75_2146 ();
 sg13g2_decap_8 FILLER_75_2153 ();
 sg13g2_decap_8 FILLER_75_2160 ();
 sg13g2_fill_2 FILLER_75_2167 ();
 sg13g2_decap_8 FILLER_75_2195 ();
 sg13g2_decap_8 FILLER_75_2202 ();
 sg13g2_decap_4 FILLER_75_2209 ();
 sg13g2_fill_2 FILLER_75_2213 ();
 sg13g2_decap_4 FILLER_75_2258 ();
 sg13g2_decap_8 FILLER_75_2266 ();
 sg13g2_decap_8 FILLER_75_2273 ();
 sg13g2_decap_8 FILLER_75_2310 ();
 sg13g2_decap_4 FILLER_75_2317 ();
 sg13g2_fill_2 FILLER_75_2321 ();
 sg13g2_fill_1 FILLER_75_2328 ();
 sg13g2_fill_1 FILLER_75_2354 ();
 sg13g2_fill_2 FILLER_75_2359 ();
 sg13g2_fill_1 FILLER_75_2408 ();
 sg13g2_decap_8 FILLER_75_2419 ();
 sg13g2_decap_8 FILLER_75_2426 ();
 sg13g2_fill_2 FILLER_75_2433 ();
 sg13g2_fill_2 FILLER_75_2447 ();
 sg13g2_fill_2 FILLER_75_2453 ();
 sg13g2_fill_2 FILLER_75_2485 ();
 sg13g2_decap_8 FILLER_75_2513 ();
 sg13g2_decap_4 FILLER_75_2520 ();
 sg13g2_fill_2 FILLER_75_2524 ();
 sg13g2_decap_8 FILLER_75_2529 ();
 sg13g2_decap_8 FILLER_75_2544 ();
 sg13g2_decap_8 FILLER_75_2551 ();
 sg13g2_decap_8 FILLER_75_2558 ();
 sg13g2_decap_8 FILLER_75_2565 ();
 sg13g2_decap_8 FILLER_75_2572 ();
 sg13g2_decap_8 FILLER_75_2579 ();
 sg13g2_decap_8 FILLER_75_2586 ();
 sg13g2_decap_4 FILLER_75_2593 ();
 sg13g2_decap_4 FILLER_75_2633 ();
 sg13g2_decap_8 FILLER_75_2653 ();
 sg13g2_decap_8 FILLER_75_2660 ();
 sg13g2_fill_2 FILLER_75_2667 ();
 sg13g2_fill_1 FILLER_75_2669 ();
 sg13g2_fill_2 FILLER_76_0 ();
 sg13g2_decap_4 FILLER_76_32 ();
 sg13g2_fill_1 FILLER_76_36 ();
 sg13g2_fill_2 FILLER_76_52 ();
 sg13g2_fill_1 FILLER_76_54 ();
 sg13g2_fill_1 FILLER_76_65 ();
 sg13g2_fill_2 FILLER_76_71 ();
 sg13g2_fill_1 FILLER_76_77 ();
 sg13g2_fill_2 FILLER_76_83 ();
 sg13g2_fill_1 FILLER_76_127 ();
 sg13g2_fill_1 FILLER_76_154 ();
 sg13g2_fill_2 FILLER_76_187 ();
 sg13g2_fill_1 FILLER_76_189 ();
 sg13g2_decap_8 FILLER_76_194 ();
 sg13g2_decap_4 FILLER_76_201 ();
 sg13g2_fill_1 FILLER_76_205 ();
 sg13g2_decap_4 FILLER_76_232 ();
 sg13g2_decap_4 FILLER_76_250 ();
 sg13g2_fill_2 FILLER_76_254 ();
 sg13g2_decap_8 FILLER_76_330 ();
 sg13g2_decap_8 FILLER_76_337 ();
 sg13g2_fill_1 FILLER_76_344 ();
 sg13g2_fill_2 FILLER_76_354 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_decap_4 FILLER_76_361 ();
 sg13g2_fill_2 FILLER_76_365 ();
 sg13g2_fill_2 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_391 ();
 sg13g2_fill_2 FILLER_76_398 ();
 sg13g2_fill_1 FILLER_76_405 ();
 sg13g2_fill_2 FILLER_76_416 ();
 sg13g2_fill_1 FILLER_76_418 ();
 sg13g2_decap_4 FILLER_76_423 ();
 sg13g2_decap_4 FILLER_76_430 ();
 sg13g2_fill_2 FILLER_76_434 ();
 sg13g2_decap_8 FILLER_76_441 ();
 sg13g2_fill_1 FILLER_76_448 ();
 sg13g2_fill_2 FILLER_76_458 ();
 sg13g2_decap_4 FILLER_76_463 ();
 sg13g2_fill_1 FILLER_76_467 ();
 sg13g2_fill_2 FILLER_76_471 ();
 sg13g2_fill_1 FILLER_76_473 ();
 sg13g2_fill_1 FILLER_76_497 ();
 sg13g2_fill_1 FILLER_76_508 ();
 sg13g2_fill_2 FILLER_76_522 ();
 sg13g2_fill_1 FILLER_76_536 ();
 sg13g2_fill_1 FILLER_76_548 ();
 sg13g2_fill_1 FILLER_76_560 ();
 sg13g2_decap_4 FILLER_76_566 ();
 sg13g2_decap_4 FILLER_76_584 ();
 sg13g2_fill_1 FILLER_76_588 ();
 sg13g2_decap_8 FILLER_76_660 ();
 sg13g2_decap_8 FILLER_76_667 ();
 sg13g2_decap_8 FILLER_76_674 ();
 sg13g2_decap_8 FILLER_76_681 ();
 sg13g2_decap_8 FILLER_76_688 ();
 sg13g2_decap_4 FILLER_76_695 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_4 FILLER_76_718 ();
 sg13g2_fill_1 FILLER_76_722 ();
 sg13g2_decap_8 FILLER_76_728 ();
 sg13g2_fill_1 FILLER_76_735 ();
 sg13g2_decap_8 FILLER_76_740 ();
 sg13g2_decap_8 FILLER_76_747 ();
 sg13g2_fill_1 FILLER_76_754 ();
 sg13g2_decap_8 FILLER_76_759 ();
 sg13g2_fill_2 FILLER_76_796 ();
 sg13g2_fill_1 FILLER_76_798 ();
 sg13g2_fill_2 FILLER_76_808 ();
 sg13g2_decap_4 FILLER_76_819 ();
 sg13g2_decap_8 FILLER_76_827 ();
 sg13g2_fill_1 FILLER_76_834 ();
 sg13g2_fill_2 FILLER_76_848 ();
 sg13g2_fill_1 FILLER_76_876 ();
 sg13g2_fill_2 FILLER_76_888 ();
 sg13g2_fill_1 FILLER_76_898 ();
 sg13g2_fill_2 FILLER_76_906 ();
 sg13g2_decap_4 FILLER_76_924 ();
 sg13g2_fill_2 FILLER_76_963 ();
 sg13g2_fill_1 FILLER_76_975 ();
 sg13g2_fill_2 FILLER_76_988 ();
 sg13g2_fill_1 FILLER_76_990 ();
 sg13g2_fill_1 FILLER_76_1029 ();
 sg13g2_decap_8 FILLER_76_1059 ();
 sg13g2_fill_2 FILLER_76_1066 ();
 sg13g2_decap_8 FILLER_76_1082 ();
 sg13g2_decap_8 FILLER_76_1089 ();
 sg13g2_decap_8 FILLER_76_1096 ();
 sg13g2_decap_8 FILLER_76_1103 ();
 sg13g2_decap_4 FILLER_76_1110 ();
 sg13g2_fill_1 FILLER_76_1114 ();
 sg13g2_decap_8 FILLER_76_1119 ();
 sg13g2_decap_8 FILLER_76_1126 ();
 sg13g2_decap_4 FILLER_76_1133 ();
 sg13g2_fill_2 FILLER_76_1137 ();
 sg13g2_decap_4 FILLER_76_1165 ();
 sg13g2_decap_8 FILLER_76_1173 ();
 sg13g2_decap_8 FILLER_76_1180 ();
 sg13g2_decap_8 FILLER_76_1187 ();
 sg13g2_decap_4 FILLER_76_1194 ();
 sg13g2_decap_8 FILLER_76_1202 ();
 sg13g2_decap_4 FILLER_76_1209 ();
 sg13g2_fill_2 FILLER_76_1213 ();
 sg13g2_fill_1 FILLER_76_1220 ();
 sg13g2_decap_8 FILLER_76_1247 ();
 sg13g2_decap_8 FILLER_76_1254 ();
 sg13g2_fill_1 FILLER_76_1261 ();
 sg13g2_fill_2 FILLER_76_1279 ();
 sg13g2_fill_1 FILLER_76_1286 ();
 sg13g2_decap_8 FILLER_76_1326 ();
 sg13g2_decap_4 FILLER_76_1333 ();
 sg13g2_fill_1 FILLER_76_1337 ();
 sg13g2_fill_2 FILLER_76_1342 ();
 sg13g2_fill_1 FILLER_76_1390 ();
 sg13g2_decap_4 FILLER_76_1430 ();
 sg13g2_fill_2 FILLER_76_1443 ();
 sg13g2_fill_1 FILLER_76_1445 ();
 sg13g2_decap_4 FILLER_76_1451 ();
 sg13g2_fill_1 FILLER_76_1455 ();
 sg13g2_decap_8 FILLER_76_1460 ();
 sg13g2_fill_2 FILLER_76_1467 ();
 sg13g2_decap_8 FILLER_76_1473 ();
 sg13g2_decap_8 FILLER_76_1480 ();
 sg13g2_decap_8 FILLER_76_1487 ();
 sg13g2_decap_4 FILLER_76_1494 ();
 sg13g2_fill_1 FILLER_76_1533 ();
 sg13g2_decap_4 FILLER_76_1550 ();
 sg13g2_fill_1 FILLER_76_1559 ();
 sg13g2_decap_8 FILLER_76_1565 ();
 sg13g2_decap_8 FILLER_76_1572 ();
 sg13g2_fill_2 FILLER_76_1584 ();
 sg13g2_fill_2 FILLER_76_1590 ();
 sg13g2_fill_1 FILLER_76_1627 ();
 sg13g2_decap_8 FILLER_76_1680 ();
 sg13g2_fill_2 FILLER_76_1687 ();
 sg13g2_fill_1 FILLER_76_1689 ();
 sg13g2_decap_8 FILLER_76_1695 ();
 sg13g2_decap_8 FILLER_76_1702 ();
 sg13g2_decap_8 FILLER_76_1709 ();
 sg13g2_fill_1 FILLER_76_1716 ();
 sg13g2_decap_8 FILLER_76_1750 ();
 sg13g2_decap_8 FILLER_76_1757 ();
 sg13g2_decap_8 FILLER_76_1764 ();
 sg13g2_decap_4 FILLER_76_1771 ();
 sg13g2_fill_2 FILLER_76_1779 ();
 sg13g2_fill_1 FILLER_76_1781 ();
 sg13g2_decap_4 FILLER_76_1786 ();
 sg13g2_decap_8 FILLER_76_1820 ();
 sg13g2_fill_2 FILLER_76_1827 ();
 sg13g2_fill_2 FILLER_76_1841 ();
 sg13g2_fill_2 FILLER_76_1874 ();
 sg13g2_fill_2 FILLER_76_1880 ();
 sg13g2_decap_8 FILLER_76_1917 ();
 sg13g2_fill_2 FILLER_76_1924 ();
 sg13g2_decap_8 FILLER_76_1974 ();
 sg13g2_decap_8 FILLER_76_1981 ();
 sg13g2_decap_8 FILLER_76_1988 ();
 sg13g2_decap_8 FILLER_76_1995 ();
 sg13g2_decap_4 FILLER_76_2002 ();
 sg13g2_fill_2 FILLER_76_2006 ();
 sg13g2_decap_8 FILLER_76_2073 ();
 sg13g2_decap_8 FILLER_76_2080 ();
 sg13g2_decap_8 FILLER_76_2087 ();
 sg13g2_decap_4 FILLER_76_2094 ();
 sg13g2_fill_1 FILLER_76_2098 ();
 sg13g2_decap_8 FILLER_76_2104 ();
 sg13g2_decap_8 FILLER_76_2111 ();
 sg13g2_decap_4 FILLER_76_2118 ();
 sg13g2_fill_2 FILLER_76_2122 ();
 sg13g2_decap_8 FILLER_76_2160 ();
 sg13g2_decap_8 FILLER_76_2167 ();
 sg13g2_decap_8 FILLER_76_2174 ();
 sg13g2_fill_1 FILLER_76_2181 ();
 sg13g2_fill_2 FILLER_76_2264 ();
 sg13g2_decap_8 FILLER_76_2304 ();
 sg13g2_decap_8 FILLER_76_2311 ();
 sg13g2_decap_4 FILLER_76_2318 ();
 sg13g2_fill_1 FILLER_76_2322 ();
 sg13g2_fill_1 FILLER_76_2365 ();
 sg13g2_fill_1 FILLER_76_2378 ();
 sg13g2_fill_2 FILLER_76_2395 ();
 sg13g2_fill_2 FILLER_76_2405 ();
 sg13g2_decap_8 FILLER_76_2420 ();
 sg13g2_decap_8 FILLER_76_2427 ();
 sg13g2_decap_8 FILLER_76_2434 ();
 sg13g2_fill_2 FILLER_76_2441 ();
 sg13g2_decap_8 FILLER_76_2449 ();
 sg13g2_fill_2 FILLER_76_2456 ();
 sg13g2_fill_1 FILLER_76_2458 ();
 sg13g2_fill_1 FILLER_76_2463 ();
 sg13g2_fill_2 FILLER_76_2490 ();
 sg13g2_fill_1 FILLER_76_2496 ();
 sg13g2_decap_8 FILLER_76_2501 ();
 sg13g2_fill_2 FILLER_76_2508 ();
 sg13g2_fill_1 FILLER_76_2510 ();
 sg13g2_fill_1 FILLER_76_2532 ();
 sg13g2_decap_4 FILLER_76_2537 ();
 sg13g2_fill_1 FILLER_76_2541 ();
 sg13g2_decap_8 FILLER_76_2546 ();
 sg13g2_decap_8 FILLER_76_2553 ();
 sg13g2_decap_8 FILLER_76_2560 ();
 sg13g2_decap_8 FILLER_76_2567 ();
 sg13g2_fill_1 FILLER_76_2574 ();
 sg13g2_fill_2 FILLER_76_2592 ();
 sg13g2_decap_8 FILLER_76_2659 ();
 sg13g2_decap_4 FILLER_76_2666 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_fill_2 FILLER_77_14 ();
 sg13g2_fill_1 FILLER_77_16 ();
 sg13g2_decap_4 FILLER_77_37 ();
 sg13g2_fill_1 FILLER_77_41 ();
 sg13g2_fill_2 FILLER_77_80 ();
 sg13g2_decap_8 FILLER_77_89 ();
 sg13g2_decap_8 FILLER_77_96 ();
 sg13g2_decap_8 FILLER_77_103 ();
 sg13g2_fill_2 FILLER_77_110 ();
 sg13g2_fill_1 FILLER_77_112 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_fill_2 FILLER_77_160 ();
 sg13g2_fill_1 FILLER_77_250 ();
 sg13g2_fill_2 FILLER_77_254 ();
 sg13g2_fill_1 FILLER_77_256 ();
 sg13g2_decap_4 FILLER_77_304 ();
 sg13g2_decap_8 FILLER_77_325 ();
 sg13g2_decap_8 FILLER_77_332 ();
 sg13g2_decap_8 FILLER_77_339 ();
 sg13g2_fill_2 FILLER_77_346 ();
 sg13g2_fill_1 FILLER_77_348 ();
 sg13g2_fill_2 FILLER_77_354 ();
 sg13g2_fill_1 FILLER_77_387 ();
 sg13g2_decap_4 FILLER_77_397 ();
 sg13g2_fill_1 FILLER_77_401 ();
 sg13g2_fill_1 FILLER_77_408 ();
 sg13g2_fill_2 FILLER_77_435 ();
 sg13g2_fill_1 FILLER_77_445 ();
 sg13g2_fill_2 FILLER_77_452 ();
 sg13g2_fill_2 FILLER_77_460 ();
 sg13g2_decap_4 FILLER_77_467 ();
 sg13g2_fill_2 FILLER_77_471 ();
 sg13g2_fill_1 FILLER_77_488 ();
 sg13g2_fill_1 FILLER_77_519 ();
 sg13g2_decap_4 FILLER_77_539 ();
 sg13g2_fill_1 FILLER_77_543 ();
 sg13g2_decap_8 FILLER_77_589 ();
 sg13g2_decap_4 FILLER_77_596 ();
 sg13g2_decap_8 FILLER_77_613 ();
 sg13g2_decap_8 FILLER_77_620 ();
 sg13g2_decap_8 FILLER_77_627 ();
 sg13g2_decap_8 FILLER_77_634 ();
 sg13g2_decap_8 FILLER_77_641 ();
 sg13g2_decap_4 FILLER_77_648 ();
 sg13g2_decap_8 FILLER_77_657 ();
 sg13g2_decap_4 FILLER_77_664 ();
 sg13g2_fill_1 FILLER_77_699 ();
 sg13g2_fill_1 FILLER_77_707 ();
 sg13g2_fill_1 FILLER_77_712 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_4 FILLER_77_759 ();
 sg13g2_fill_2 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_4 FILLER_77_784 ();
 sg13g2_fill_1 FILLER_77_788 ();
 sg13g2_fill_2 FILLER_77_824 ();
 sg13g2_fill_1 FILLER_77_826 ();
 sg13g2_fill_1 FILLER_77_858 ();
 sg13g2_fill_1 FILLER_77_910 ();
 sg13g2_fill_1 FILLER_77_915 ();
 sg13g2_decap_8 FILLER_77_924 ();
 sg13g2_fill_2 FILLER_77_931 ();
 sg13g2_fill_1 FILLER_77_933 ();
 sg13g2_fill_1 FILLER_77_965 ();
 sg13g2_fill_2 FILLER_77_971 ();
 sg13g2_decap_4 FILLER_77_1035 ();
 sg13g2_fill_2 FILLER_77_1080 ();
 sg13g2_decap_4 FILLER_77_1108 ();
 sg13g2_decap_8 FILLER_77_1138 ();
 sg13g2_fill_2 FILLER_77_1150 ();
 sg13g2_decap_8 FILLER_77_1182 ();
 sg13g2_fill_2 FILLER_77_1189 ();
 sg13g2_fill_1 FILLER_77_1231 ();
 sg13g2_fill_1 FILLER_77_1267 ();
 sg13g2_fill_2 FILLER_77_1273 ();
 sg13g2_fill_2 FILLER_77_1301 ();
 sg13g2_fill_1 FILLER_77_1303 ();
 sg13g2_decap_8 FILLER_77_1309 ();
 sg13g2_fill_1 FILLER_77_1316 ();
 sg13g2_fill_1 FILLER_77_1322 ();
 sg13g2_decap_4 FILLER_77_1328 ();
 sg13g2_fill_2 FILLER_77_1332 ();
 sg13g2_fill_2 FILLER_77_1365 ();
 sg13g2_fill_1 FILLER_77_1367 ();
 sg13g2_fill_2 FILLER_77_1381 ();
 sg13g2_fill_1 FILLER_77_1414 ();
 sg13g2_decap_4 FILLER_77_1420 ();
 sg13g2_decap_4 FILLER_77_1429 ();
 sg13g2_decap_4 FILLER_77_1473 ();
 sg13g2_decap_8 FILLER_77_1590 ();
 sg13g2_decap_8 FILLER_77_1597 ();
 sg13g2_decap_4 FILLER_77_1604 ();
 sg13g2_fill_2 FILLER_77_1621 ();
 sg13g2_decap_4 FILLER_77_1675 ();
 sg13g2_fill_1 FILLER_77_1679 ();
 sg13g2_fill_1 FILLER_77_1706 ();
 sg13g2_decap_8 FILLER_77_1760 ();
 sg13g2_decap_4 FILLER_77_1797 ();
 sg13g2_fill_2 FILLER_77_1801 ();
 sg13g2_fill_1 FILLER_77_1835 ();
 sg13g2_fill_1 FILLER_77_1844 ();
 sg13g2_decap_4 FILLER_77_1853 ();
 sg13g2_fill_2 FILLER_77_1857 ();
 sg13g2_decap_8 FILLER_77_1916 ();
 sg13g2_fill_1 FILLER_77_1949 ();
 sg13g2_decap_4 FILLER_77_2001 ();
 sg13g2_fill_1 FILLER_77_2005 ();
 sg13g2_decap_4 FILLER_77_2019 ();
 sg13g2_fill_1 FILLER_77_2023 ();
 sg13g2_fill_2 FILLER_77_2028 ();
 sg13g2_decap_8 FILLER_77_2034 ();
 sg13g2_fill_1 FILLER_77_2050 ();
 sg13g2_decap_8 FILLER_77_2087 ();
 sg13g2_decap_8 FILLER_77_2094 ();
 sg13g2_decap_4 FILLER_77_2127 ();
 sg13g2_decap_4 FILLER_77_2207 ();
 sg13g2_fill_1 FILLER_77_2211 ();
 sg13g2_fill_2 FILLER_77_2224 ();
 sg13g2_decap_8 FILLER_77_2230 ();
 sg13g2_decap_4 FILLER_77_2237 ();
 sg13g2_decap_8 FILLER_77_2245 ();
 sg13g2_fill_2 FILLER_77_2252 ();
 sg13g2_fill_2 FILLER_77_2280 ();
 sg13g2_fill_2 FILLER_77_2299 ();
 sg13g2_fill_2 FILLER_77_2357 ();
 sg13g2_fill_1 FILLER_77_2359 ();
 sg13g2_decap_8 FILLER_77_2383 ();
 sg13g2_decap_8 FILLER_77_2390 ();
 sg13g2_fill_1 FILLER_77_2397 ();
 sg13g2_fill_2 FILLER_77_2402 ();
 sg13g2_fill_1 FILLER_77_2404 ();
 sg13g2_decap_8 FILLER_77_2431 ();
 sg13g2_fill_2 FILLER_77_2438 ();
 sg13g2_fill_1 FILLER_77_2440 ();
 sg13g2_decap_8 FILLER_77_2445 ();
 sg13g2_decap_8 FILLER_77_2452 ();
 sg13g2_decap_8 FILLER_77_2459 ();
 sg13g2_fill_2 FILLER_77_2466 ();
 sg13g2_fill_2 FILLER_77_2472 ();
 sg13g2_decap_8 FILLER_77_2488 ();
 sg13g2_fill_1 FILLER_77_2495 ();
 sg13g2_decap_4 FILLER_77_2529 ();
 sg13g2_fill_1 FILLER_77_2533 ();
 sg13g2_decap_8 FILLER_77_2560 ();
 sg13g2_decap_8 FILLER_77_2567 ();
 sg13g2_decap_4 FILLER_77_2574 ();
 sg13g2_decap_8 FILLER_77_2582 ();
 sg13g2_fill_2 FILLER_77_2667 ();
 sg13g2_fill_1 FILLER_77_2669 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_7 ();
 sg13g2_fill_1 FILLER_78_34 ();
 sg13g2_fill_2 FILLER_78_39 ();
 sg13g2_fill_1 FILLER_78_41 ();
 sg13g2_fill_1 FILLER_78_71 ();
 sg13g2_fill_2 FILLER_78_94 ();
 sg13g2_decap_4 FILLER_78_100 ();
 sg13g2_decap_8 FILLER_78_130 ();
 sg13g2_fill_2 FILLER_78_137 ();
 sg13g2_fill_1 FILLER_78_139 ();
 sg13g2_fill_2 FILLER_78_165 ();
 sg13g2_fill_2 FILLER_78_172 ();
 sg13g2_decap_8 FILLER_78_204 ();
 sg13g2_fill_2 FILLER_78_254 ();
 sg13g2_decap_4 FILLER_78_282 ();
 sg13g2_fill_1 FILLER_78_286 ();
 sg13g2_fill_1 FILLER_78_292 ();
 sg13g2_decap_8 FILLER_78_329 ();
 sg13g2_decap_8 FILLER_78_336 ();
 sg13g2_decap_8 FILLER_78_343 ();
 sg13g2_decap_4 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_354 ();
 sg13g2_fill_1 FILLER_78_407 ();
 sg13g2_fill_1 FILLER_78_413 ();
 sg13g2_fill_1 FILLER_78_418 ();
 sg13g2_fill_1 FILLER_78_424 ();
 sg13g2_fill_2 FILLER_78_490 ();
 sg13g2_fill_1 FILLER_78_492 ();
 sg13g2_decap_4 FILLER_78_506 ();
 sg13g2_fill_1 FILLER_78_510 ();
 sg13g2_decap_4 FILLER_78_515 ();
 sg13g2_fill_1 FILLER_78_519 ();
 sg13g2_fill_2 FILLER_78_533 ();
 sg13g2_fill_1 FILLER_78_535 ();
 sg13g2_fill_2 FILLER_78_549 ();
 sg13g2_fill_1 FILLER_78_583 ();
 sg13g2_fill_2 FILLER_78_588 ();
 sg13g2_decap_8 FILLER_78_616 ();
 sg13g2_fill_1 FILLER_78_623 ();
 sg13g2_fill_1 FILLER_78_629 ();
 sg13g2_decap_8 FILLER_78_656 ();
 sg13g2_fill_2 FILLER_78_663 ();
 sg13g2_fill_1 FILLER_78_665 ();
 sg13g2_fill_1 FILLER_78_692 ();
 sg13g2_fill_2 FILLER_78_698 ();
 sg13g2_fill_1 FILLER_78_700 ();
 sg13g2_fill_2 FILLER_78_719 ();
 sg13g2_fill_1 FILLER_78_721 ();
 sg13g2_fill_1 FILLER_78_748 ();
 sg13g2_fill_1 FILLER_78_754 ();
 sg13g2_decap_4 FILLER_78_781 ();
 sg13g2_fill_2 FILLER_78_834 ();
 sg13g2_fill_2 FILLER_78_901 ();
 sg13g2_decap_8 FILLER_78_960 ();
 sg13g2_decap_4 FILLER_78_993 ();
 sg13g2_fill_1 FILLER_78_1031 ();
 sg13g2_fill_1 FILLER_78_1058 ();
 sg13g2_fill_1 FILLER_78_1085 ();
 sg13g2_fill_1 FILLER_78_1138 ();
 sg13g2_decap_8 FILLER_78_1170 ();
 sg13g2_decap_8 FILLER_78_1177 ();
 sg13g2_decap_8 FILLER_78_1184 ();
 sg13g2_fill_1 FILLER_78_1221 ();
 sg13g2_fill_1 FILLER_78_1244 ();
 sg13g2_fill_2 FILLER_78_1259 ();
 sg13g2_decap_8 FILLER_78_1317 ();
 sg13g2_fill_2 FILLER_78_1324 ();
 sg13g2_fill_2 FILLER_78_1356 ();
 sg13g2_fill_2 FILLER_78_1366 ();
 sg13g2_fill_2 FILLER_78_1407 ();
 sg13g2_fill_2 FILLER_78_1427 ();
 sg13g2_fill_1 FILLER_78_1512 ();
 sg13g2_fill_2 FILLER_78_1517 ();
 sg13g2_fill_2 FILLER_78_1550 ();
 sg13g2_fill_1 FILLER_78_1552 ();
 sg13g2_decap_8 FILLER_78_1561 ();
 sg13g2_decap_4 FILLER_78_1568 ();
 sg13g2_fill_1 FILLER_78_1572 ();
 sg13g2_fill_1 FILLER_78_1578 ();
 sg13g2_decap_8 FILLER_78_1605 ();
 sg13g2_decap_4 FILLER_78_1612 ();
 sg13g2_fill_1 FILLER_78_1616 ();
 sg13g2_decap_4 FILLER_78_1643 ();
 sg13g2_fill_1 FILLER_78_1647 ();
 sg13g2_decap_8 FILLER_78_1665 ();
 sg13g2_decap_4 FILLER_78_1672 ();
 sg13g2_fill_2 FILLER_78_1676 ();
 sg13g2_fill_2 FILLER_78_1827 ();
 sg13g2_decap_8 FILLER_78_1845 ();
 sg13g2_fill_2 FILLER_78_1852 ();
 sg13g2_fill_2 FILLER_78_1858 ();
 sg13g2_fill_1 FILLER_78_1860 ();
 sg13g2_fill_1 FILLER_78_1887 ();
 sg13g2_fill_1 FILLER_78_1917 ();
 sg13g2_decap_4 FILLER_78_1922 ();
 sg13g2_fill_2 FILLER_78_1926 ();
 sg13g2_decap_4 FILLER_78_1972 ();
 sg13g2_fill_1 FILLER_78_1976 ();
 sg13g2_decap_8 FILLER_78_1981 ();
 sg13g2_fill_2 FILLER_78_1988 ();
 sg13g2_fill_2 FILLER_78_2042 ();
 sg13g2_decap_8 FILLER_78_2076 ();
 sg13g2_fill_2 FILLER_78_2083 ();
 sg13g2_fill_1 FILLER_78_2085 ();
 sg13g2_fill_2 FILLER_78_2120 ();
 sg13g2_fill_2 FILLER_78_2126 ();
 sg13g2_decap_8 FILLER_78_2136 ();
 sg13g2_fill_2 FILLER_78_2143 ();
 sg13g2_decap_8 FILLER_78_2155 ();
 sg13g2_fill_2 FILLER_78_2162 ();
 sg13g2_decap_4 FILLER_78_2206 ();
 sg13g2_fill_1 FILLER_78_2210 ();
 sg13g2_decap_4 FILLER_78_2313 ();
 sg13g2_fill_1 FILLER_78_2317 ();
 sg13g2_fill_2 FILLER_78_2344 ();
 sg13g2_fill_1 FILLER_78_2346 ();
 sg13g2_fill_1 FILLER_78_2403 ();
 sg13g2_fill_2 FILLER_78_2434 ();
 sg13g2_fill_2 FILLER_78_2440 ();
 sg13g2_fill_2 FILLER_78_2468 ();
 sg13g2_fill_1 FILLER_78_2470 ();
 sg13g2_fill_1 FILLER_78_2475 ();
 sg13g2_fill_1 FILLER_78_2502 ();
 sg13g2_fill_1 FILLER_78_2533 ();
 sg13g2_fill_2 FILLER_78_2564 ();
 sg13g2_fill_1 FILLER_78_2566 ();
 sg13g2_fill_1 FILLER_78_2593 ();
 sg13g2_decap_8 FILLER_78_2663 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_fill_1 FILLER_79_14 ();
 sg13g2_fill_2 FILLER_79_41 ();
 sg13g2_fill_1 FILLER_79_43 ();
 sg13g2_decap_8 FILLER_79_48 ();
 sg13g2_decap_4 FILLER_79_55 ();
 sg13g2_fill_1 FILLER_79_67 ();
 sg13g2_decap_4 FILLER_79_102 ();
 sg13g2_fill_2 FILLER_79_106 ();
 sg13g2_decap_4 FILLER_79_118 ();
 sg13g2_decap_8 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_133 ();
 sg13g2_decap_8 FILLER_79_140 ();
 sg13g2_decap_8 FILLER_79_147 ();
 sg13g2_decap_4 FILLER_79_159 ();
 sg13g2_fill_1 FILLER_79_163 ();
 sg13g2_decap_8 FILLER_79_169 ();
 sg13g2_decap_8 FILLER_79_176 ();
 sg13g2_decap_4 FILLER_79_195 ();
 sg13g2_fill_1 FILLER_79_199 ();
 sg13g2_decap_4 FILLER_79_212 ();
 sg13g2_fill_2 FILLER_79_216 ();
 sg13g2_fill_2 FILLER_79_226 ();
 sg13g2_fill_1 FILLER_79_228 ();
 sg13g2_decap_8 FILLER_79_274 ();
 sg13g2_decap_8 FILLER_79_281 ();
 sg13g2_decap_4 FILLER_79_292 ();
 sg13g2_fill_1 FILLER_79_296 ();
 sg13g2_decap_4 FILLER_79_331 ();
 sg13g2_fill_2 FILLER_79_335 ();
 sg13g2_decap_4 FILLER_79_417 ();
 sg13g2_fill_1 FILLER_79_421 ();
 sg13g2_decap_8 FILLER_79_427 ();
 sg13g2_fill_1 FILLER_79_434 ();
 sg13g2_decap_4 FILLER_79_474 ();
 sg13g2_fill_2 FILLER_79_478 ();
 sg13g2_decap_8 FILLER_79_497 ();
 sg13g2_decap_8 FILLER_79_504 ();
 sg13g2_decap_8 FILLER_79_511 ();
 sg13g2_fill_1 FILLER_79_561 ();
 sg13g2_fill_1 FILLER_79_576 ();
 sg13g2_fill_1 FILLER_79_580 ();
 sg13g2_fill_2 FILLER_79_607 ();
 sg13g2_fill_2 FILLER_79_617 ();
 sg13g2_fill_2 FILLER_79_624 ();
 sg13g2_decap_8 FILLER_79_652 ();
 sg13g2_decap_8 FILLER_79_659 ();
 sg13g2_decap_8 FILLER_79_666 ();
 sg13g2_decap_8 FILLER_79_673 ();
 sg13g2_decap_8 FILLER_79_680 ();
 sg13g2_fill_2 FILLER_79_687 ();
 sg13g2_fill_1 FILLER_79_689 ();
 sg13g2_fill_1 FILLER_79_720 ();
 sg13g2_fill_2 FILLER_79_747 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_4 FILLER_79_760 ();
 sg13g2_fill_2 FILLER_79_764 ();
 sg13g2_fill_2 FILLER_79_792 ();
 sg13g2_decap_4 FILLER_79_820 ();
 sg13g2_decap_4 FILLER_79_850 ();
 sg13g2_fill_1 FILLER_79_862 ();
 sg13g2_fill_2 FILLER_79_889 ();
 sg13g2_decap_8 FILLER_79_935 ();
 sg13g2_fill_2 FILLER_79_942 ();
 sg13g2_fill_1 FILLER_79_944 ();
 sg13g2_decap_4 FILLER_79_953 ();
 sg13g2_decap_8 FILLER_79_962 ();
 sg13g2_decap_4 FILLER_79_969 ();
 sg13g2_fill_1 FILLER_79_973 ();
 sg13g2_fill_2 FILLER_79_1000 ();
 sg13g2_decap_4 FILLER_79_1007 ();
 sg13g2_fill_2 FILLER_79_1037 ();
 sg13g2_decap_4 FILLER_79_1065 ();
 sg13g2_fill_1 FILLER_79_1074 ();
 sg13g2_fill_2 FILLER_79_1110 ();
 sg13g2_fill_1 FILLER_79_1112 ();
 sg13g2_fill_2 FILLER_79_1135 ();
 sg13g2_fill_2 FILLER_79_1145 ();
 sg13g2_fill_1 FILLER_79_1147 ();
 sg13g2_fill_2 FILLER_79_1153 ();
 sg13g2_fill_1 FILLER_79_1155 ();
 sg13g2_fill_2 FILLER_79_1200 ();
 sg13g2_fill_1 FILLER_79_1202 ();
 sg13g2_fill_2 FILLER_79_1211 ();
 sg13g2_fill_1 FILLER_79_1213 ();
 sg13g2_fill_1 FILLER_79_1219 ();
 sg13g2_fill_2 FILLER_79_1246 ();
 sg13g2_fill_1 FILLER_79_1248 ();
 sg13g2_fill_1 FILLER_79_1275 ();
 sg13g2_decap_8 FILLER_79_1280 ();
 sg13g2_fill_2 FILLER_79_1287 ();
 sg13g2_fill_1 FILLER_79_1289 ();
 sg13g2_decap_8 FILLER_79_1298 ();
 sg13g2_decap_4 FILLER_79_1305 ();
 sg13g2_fill_1 FILLER_79_1309 ();
 sg13g2_decap_8 FILLER_79_1336 ();
 sg13g2_decap_8 FILLER_79_1343 ();
 sg13g2_decap_8 FILLER_79_1350 ();
 sg13g2_fill_2 FILLER_79_1357 ();
 sg13g2_fill_1 FILLER_79_1359 ();
 sg13g2_fill_2 FILLER_79_1376 ();
 sg13g2_decap_8 FILLER_79_1465 ();
 sg13g2_decap_8 FILLER_79_1472 ();
 sg13g2_fill_2 FILLER_79_1484 ();
 sg13g2_fill_1 FILLER_79_1486 ();
 sg13g2_fill_1 FILLER_79_1510 ();
 sg13g2_fill_2 FILLER_79_1516 ();
 sg13g2_decap_4 FILLER_79_1522 ();
 sg13g2_fill_2 FILLER_79_1526 ();
 sg13g2_fill_1 FILLER_79_1533 ();
 sg13g2_decap_4 FILLER_79_1560 ();
 sg13g2_fill_2 FILLER_79_1564 ();
 sg13g2_decap_4 FILLER_79_1574 ();
 sg13g2_decap_8 FILLER_79_1608 ();
 sg13g2_fill_1 FILLER_79_1615 ();
 sg13g2_decap_8 FILLER_79_1629 ();
 sg13g2_fill_2 FILLER_79_1636 ();
 sg13g2_fill_1 FILLER_79_1658 ();
 sg13g2_fill_1 FILLER_79_1689 ();
 sg13g2_decap_4 FILLER_79_1695 ();
 sg13g2_fill_1 FILLER_79_1699 ();
 sg13g2_fill_1 FILLER_79_1762 ();
 sg13g2_fill_2 FILLER_79_1773 ();
 sg13g2_fill_2 FILLER_79_1782 ();
 sg13g2_decap_4 FILLER_79_1788 ();
 sg13g2_fill_1 FILLER_79_1792 ();
 sg13g2_fill_1 FILLER_79_1842 ();
 sg13g2_decap_8 FILLER_79_1873 ();
 sg13g2_decap_8 FILLER_79_1880 ();
 sg13g2_fill_1 FILLER_79_1887 ();
 sg13g2_fill_2 FILLER_79_1894 ();
 sg13g2_fill_2 FILLER_79_1926 ();
 sg13g2_fill_2 FILLER_79_1932 ();
 sg13g2_fill_1 FILLER_79_1934 ();
 sg13g2_fill_2 FILLER_79_1974 ();
 sg13g2_fill_1 FILLER_79_1976 ();
 sg13g2_fill_1 FILLER_79_2011 ();
 sg13g2_fill_2 FILLER_79_2038 ();
 sg13g2_fill_1 FILLER_79_2115 ();
 sg13g2_decap_8 FILLER_79_2142 ();
 sg13g2_decap_8 FILLER_79_2149 ();
 sg13g2_decap_8 FILLER_79_2156 ();
 sg13g2_fill_1 FILLER_79_2163 ();
 sg13g2_fill_1 FILLER_79_2246 ();
 sg13g2_fill_2 FILLER_79_2251 ();
 sg13g2_fill_2 FILLER_79_2257 ();
 sg13g2_fill_2 FILLER_79_2263 ();
 sg13g2_fill_1 FILLER_79_2269 ();
 sg13g2_fill_1 FILLER_79_2274 ();
 sg13g2_fill_1 FILLER_79_2301 ();
 sg13g2_fill_2 FILLER_79_2344 ();
 sg13g2_decap_8 FILLER_79_2350 ();
 sg13g2_fill_1 FILLER_79_2357 ();
 sg13g2_decap_4 FILLER_79_2362 ();
 sg13g2_decap_8 FILLER_79_2435 ();
 sg13g2_fill_1 FILLER_79_2442 ();
 sg13g2_fill_2 FILLER_79_2499 ();
 sg13g2_fill_1 FILLER_79_2501 ();
 sg13g2_decap_4 FILLER_79_2567 ();
 sg13g2_fill_2 FILLER_79_2571 ();
 sg13g2_decap_8 FILLER_79_2648 ();
 sg13g2_decap_8 FILLER_79_2655 ();
 sg13g2_decap_8 FILLER_79_2662 ();
 sg13g2_fill_1 FILLER_79_2669 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_56 ();
 sg13g2_fill_2 FILLER_80_60 ();
 sg13g2_fill_2 FILLER_80_74 ();
 sg13g2_fill_2 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_90 ();
 sg13g2_fill_2 FILLER_80_121 ();
 sg13g2_fill_1 FILLER_80_123 ();
 sg13g2_fill_2 FILLER_80_128 ();
 sg13g2_fill_1 FILLER_80_130 ();
 sg13g2_fill_2 FILLER_80_139 ();
 sg13g2_decap_8 FILLER_80_145 ();
 sg13g2_decap_8 FILLER_80_152 ();
 sg13g2_decap_4 FILLER_80_159 ();
 sg13g2_fill_2 FILLER_80_163 ();
 sg13g2_decap_8 FILLER_80_169 ();
 sg13g2_decap_8 FILLER_80_176 ();
 sg13g2_fill_1 FILLER_80_183 ();
 sg13g2_fill_2 FILLER_80_204 ();
 sg13g2_fill_2 FILLER_80_210 ();
 sg13g2_decap_4 FILLER_80_216 ();
 sg13g2_fill_1 FILLER_80_228 ();
 sg13g2_decap_4 FILLER_80_233 ();
 sg13g2_fill_2 FILLER_80_241 ();
 sg13g2_decap_8 FILLER_80_263 ();
 sg13g2_decap_8 FILLER_80_270 ();
 sg13g2_fill_1 FILLER_80_277 ();
 sg13g2_decap_8 FILLER_80_282 ();
 sg13g2_decap_8 FILLER_80_289 ();
 sg13g2_fill_1 FILLER_80_296 ();
 sg13g2_decap_8 FILLER_80_305 ();
 sg13g2_decap_8 FILLER_80_320 ();
 sg13g2_decap_4 FILLER_80_327 ();
 sg13g2_fill_1 FILLER_80_331 ();
 sg13g2_decap_8 FILLER_80_361 ();
 sg13g2_decap_8 FILLER_80_368 ();
 sg13g2_fill_1 FILLER_80_375 ();
 sg13g2_decap_4 FILLER_80_380 ();
 sg13g2_decap_4 FILLER_80_388 ();
 sg13g2_fill_2 FILLER_80_392 ();
 sg13g2_decap_4 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_8 FILLER_80_426 ();
 sg13g2_decap_4 FILLER_80_433 ();
 sg13g2_fill_2 FILLER_80_437 ();
 sg13g2_decap_8 FILLER_80_443 ();
 sg13g2_decap_8 FILLER_80_450 ();
 sg13g2_decap_8 FILLER_80_465 ();
 sg13g2_decap_8 FILLER_80_472 ();
 sg13g2_decap_8 FILLER_80_479 ();
 sg13g2_decap_8 FILLER_80_486 ();
 sg13g2_decap_8 FILLER_80_493 ();
 sg13g2_decap_8 FILLER_80_500 ();
 sg13g2_decap_8 FILLER_80_507 ();
 sg13g2_decap_8 FILLER_80_514 ();
 sg13g2_fill_2 FILLER_80_521 ();
 sg13g2_decap_8 FILLER_80_528 ();
 sg13g2_decap_8 FILLER_80_535 ();
 sg13g2_decap_8 FILLER_80_542 ();
 sg13g2_fill_1 FILLER_80_554 ();
 sg13g2_decap_8 FILLER_80_559 ();
 sg13g2_decap_8 FILLER_80_566 ();
 sg13g2_decap_4 FILLER_80_573 ();
 sg13g2_decap_8 FILLER_80_582 ();
 sg13g2_decap_8 FILLER_80_589 ();
 sg13g2_decap_8 FILLER_80_596 ();
 sg13g2_decap_8 FILLER_80_603 ();
 sg13g2_decap_8 FILLER_80_610 ();
 sg13g2_decap_8 FILLER_80_617 ();
 sg13g2_decap_8 FILLER_80_624 ();
 sg13g2_decap_8 FILLER_80_631 ();
 sg13g2_decap_8 FILLER_80_638 ();
 sg13g2_decap_8 FILLER_80_645 ();
 sg13g2_decap_8 FILLER_80_652 ();
 sg13g2_decap_8 FILLER_80_659 ();
 sg13g2_decap_8 FILLER_80_666 ();
 sg13g2_decap_8 FILLER_80_673 ();
 sg13g2_decap_8 FILLER_80_680 ();
 sg13g2_decap_8 FILLER_80_687 ();
 sg13g2_decap_8 FILLER_80_694 ();
 sg13g2_decap_8 FILLER_80_709 ();
 sg13g2_fill_1 FILLER_80_716 ();
 sg13g2_fill_2 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_fill_2 FILLER_80_777 ();
 sg13g2_fill_1 FILLER_80_779 ();
 sg13g2_decap_8 FILLER_80_793 ();
 sg13g2_decap_8 FILLER_80_808 ();
 sg13g2_decap_8 FILLER_80_815 ();
 sg13g2_decap_8 FILLER_80_822 ();
 sg13g2_decap_8 FILLER_80_829 ();
 sg13g2_decap_8 FILLER_80_836 ();
 sg13g2_decap_8 FILLER_80_843 ();
 sg13g2_decap_8 FILLER_80_850 ();
 sg13g2_decap_8 FILLER_80_857 ();
 sg13g2_decap_8 FILLER_80_864 ();
 sg13g2_decap_8 FILLER_80_871 ();
 sg13g2_decap_8 FILLER_80_878 ();
 sg13g2_decap_8 FILLER_80_885 ();
 sg13g2_fill_2 FILLER_80_892 ();
 sg13g2_fill_1 FILLER_80_894 ();
 sg13g2_decap_8 FILLER_80_921 ();
 sg13g2_decap_8 FILLER_80_928 ();
 sg13g2_decap_8 FILLER_80_935 ();
 sg13g2_decap_8 FILLER_80_942 ();
 sg13g2_decap_8 FILLER_80_949 ();
 sg13g2_decap_8 FILLER_80_956 ();
 sg13g2_decap_8 FILLER_80_963 ();
 sg13g2_decap_8 FILLER_80_970 ();
 sg13g2_decap_8 FILLER_80_977 ();
 sg13g2_decap_8 FILLER_80_984 ();
 sg13g2_decap_8 FILLER_80_991 ();
 sg13g2_decap_8 FILLER_80_998 ();
 sg13g2_decap_4 FILLER_80_1005 ();
 sg13g2_fill_1 FILLER_80_1009 ();
 sg13g2_decap_8 FILLER_80_1018 ();
 sg13g2_decap_8 FILLER_80_1025 ();
 sg13g2_decap_8 FILLER_80_1032 ();
 sg13g2_decap_8 FILLER_80_1039 ();
 sg13g2_fill_2 FILLER_80_1046 ();
 sg13g2_decap_8 FILLER_80_1056 ();
 sg13g2_decap_8 FILLER_80_1068 ();
 sg13g2_fill_1 FILLER_80_1075 ();
 sg13g2_fill_2 FILLER_80_1080 ();
 sg13g2_decap_8 FILLER_80_1086 ();
 sg13g2_decap_8 FILLER_80_1093 ();
 sg13g2_decap_8 FILLER_80_1100 ();
 sg13g2_decap_8 FILLER_80_1107 ();
 sg13g2_decap_8 FILLER_80_1114 ();
 sg13g2_decap_8 FILLER_80_1121 ();
 sg13g2_decap_8 FILLER_80_1128 ();
 sg13g2_decap_8 FILLER_80_1135 ();
 sg13g2_decap_8 FILLER_80_1142 ();
 sg13g2_decap_8 FILLER_80_1149 ();
 sg13g2_decap_4 FILLER_80_1156 ();
 sg13g2_decap_8 FILLER_80_1164 ();
 sg13g2_decap_8 FILLER_80_1171 ();
 sg13g2_decap_8 FILLER_80_1178 ();
 sg13g2_decap_4 FILLER_80_1185 ();
 sg13g2_decap_8 FILLER_80_1215 ();
 sg13g2_decap_8 FILLER_80_1222 ();
 sg13g2_decap_8 FILLER_80_1229 ();
 sg13g2_decap_8 FILLER_80_1236 ();
 sg13g2_decap_8 FILLER_80_1243 ();
 sg13g2_decap_8 FILLER_80_1250 ();
 sg13g2_fill_2 FILLER_80_1257 ();
 sg13g2_fill_1 FILLER_80_1259 ();
 sg13g2_decap_8 FILLER_80_1268 ();
 sg13g2_decap_8 FILLER_80_1275 ();
 sg13g2_decap_8 FILLER_80_1282 ();
 sg13g2_decap_8 FILLER_80_1289 ();
 sg13g2_decap_8 FILLER_80_1296 ();
 sg13g2_decap_8 FILLER_80_1303 ();
 sg13g2_decap_8 FILLER_80_1310 ();
 sg13g2_decap_8 FILLER_80_1317 ();
 sg13g2_decap_8 FILLER_80_1324 ();
 sg13g2_decap_8 FILLER_80_1331 ();
 sg13g2_decap_8 FILLER_80_1338 ();
 sg13g2_decap_8 FILLER_80_1345 ();
 sg13g2_fill_1 FILLER_80_1352 ();
 sg13g2_decap_4 FILLER_80_1358 ();
 sg13g2_fill_1 FILLER_80_1362 ();
 sg13g2_fill_1 FILLER_80_1428 ();
 sg13g2_fill_2 FILLER_80_1443 ();
 sg13g2_decap_8 FILLER_80_1449 ();
 sg13g2_decap_4 FILLER_80_1456 ();
 sg13g2_fill_2 FILLER_80_1460 ();
 sg13g2_decap_8 FILLER_80_1470 ();
 sg13g2_decap_8 FILLER_80_1477 ();
 sg13g2_decap_8 FILLER_80_1488 ();
 sg13g2_decap_8 FILLER_80_1499 ();
 sg13g2_decap_8 FILLER_80_1506 ();
 sg13g2_decap_8 FILLER_80_1513 ();
 sg13g2_decap_8 FILLER_80_1520 ();
 sg13g2_decap_8 FILLER_80_1527 ();
 sg13g2_decap_8 FILLER_80_1534 ();
 sg13g2_decap_4 FILLER_80_1545 ();
 sg13g2_fill_1 FILLER_80_1549 ();
 sg13g2_decap_8 FILLER_80_1555 ();
 sg13g2_decap_8 FILLER_80_1562 ();
 sg13g2_decap_8 FILLER_80_1569 ();
 sg13g2_decap_8 FILLER_80_1576 ();
 sg13g2_decap_4 FILLER_80_1583 ();
 sg13g2_fill_1 FILLER_80_1587 ();
 sg13g2_decap_8 FILLER_80_1592 ();
 sg13g2_decap_8 FILLER_80_1599 ();
 sg13g2_decap_8 FILLER_80_1606 ();
 sg13g2_decap_8 FILLER_80_1613 ();
 sg13g2_decap_8 FILLER_80_1620 ();
 sg13g2_decap_8 FILLER_80_1627 ();
 sg13g2_decap_8 FILLER_80_1634 ();
 sg13g2_decap_8 FILLER_80_1641 ();
 sg13g2_fill_2 FILLER_80_1648 ();
 sg13g2_fill_1 FILLER_80_1650 ();
 sg13g2_decap_8 FILLER_80_1660 ();
 sg13g2_fill_1 FILLER_80_1667 ();
 sg13g2_decap_8 FILLER_80_1672 ();
 sg13g2_decap_8 FILLER_80_1679 ();
 sg13g2_decap_8 FILLER_80_1686 ();
 sg13g2_fill_2 FILLER_80_1693 ();
 sg13g2_fill_1 FILLER_80_1695 ();
 sg13g2_fill_2 FILLER_80_1720 ();
 sg13g2_fill_1 FILLER_80_1753 ();
 sg13g2_decap_8 FILLER_80_1784 ();
 sg13g2_decap_8 FILLER_80_1791 ();
 sg13g2_fill_1 FILLER_80_1798 ();
 sg13g2_decap_4 FILLER_80_1803 ();
 sg13g2_fill_2 FILLER_80_1807 ();
 sg13g2_fill_2 FILLER_80_1821 ();
 sg13g2_fill_1 FILLER_80_1838 ();
 sg13g2_fill_1 FILLER_80_1849 ();
 sg13g2_fill_2 FILLER_80_1857 ();
 sg13g2_decap_8 FILLER_80_1864 ();
 sg13g2_decap_8 FILLER_80_1871 ();
 sg13g2_decap_8 FILLER_80_1878 ();
 sg13g2_decap_8 FILLER_80_1885 ();
 sg13g2_decap_8 FILLER_80_1892 ();
 sg13g2_decap_4 FILLER_80_1899 ();
 sg13g2_fill_2 FILLER_80_1907 ();
 sg13g2_fill_1 FILLER_80_1909 ();
 sg13g2_decap_8 FILLER_80_1948 ();
 sg13g2_fill_1 FILLER_80_1955 ();
 sg13g2_decap_8 FILLER_80_1960 ();
 sg13g2_decap_8 FILLER_80_1967 ();
 sg13g2_decap_8 FILLER_80_1974 ();
 sg13g2_decap_8 FILLER_80_1981 ();
 sg13g2_decap_8 FILLER_80_1992 ();
 sg13g2_decap_8 FILLER_80_1999 ();
 sg13g2_decap_8 FILLER_80_2006 ();
 sg13g2_decap_4 FILLER_80_2013 ();
 sg13g2_fill_1 FILLER_80_2017 ();
 sg13g2_decap_8 FILLER_80_2022 ();
 sg13g2_decap_8 FILLER_80_2029 ();
 sg13g2_decap_4 FILLER_80_2066 ();
 sg13g2_fill_2 FILLER_80_2070 ();
 sg13g2_decap_4 FILLER_80_2085 ();
 sg13g2_fill_2 FILLER_80_2089 ();
 sg13g2_fill_1 FILLER_80_2095 ();
 sg13g2_fill_1 FILLER_80_2100 ();
 sg13g2_decap_8 FILLER_80_2105 ();
 sg13g2_decap_8 FILLER_80_2112 ();
 sg13g2_decap_8 FILLER_80_2119 ();
 sg13g2_decap_8 FILLER_80_2126 ();
 sg13g2_decap_8 FILLER_80_2133 ();
 sg13g2_decap_8 FILLER_80_2140 ();
 sg13g2_decap_8 FILLER_80_2147 ();
 sg13g2_decap_8 FILLER_80_2154 ();
 sg13g2_decap_8 FILLER_80_2161 ();
 sg13g2_decap_4 FILLER_80_2168 ();
 sg13g2_decap_4 FILLER_80_2176 ();
 sg13g2_fill_1 FILLER_80_2180 ();
 sg13g2_decap_8 FILLER_80_2185 ();
 sg13g2_decap_8 FILLER_80_2192 ();
 sg13g2_decap_8 FILLER_80_2203 ();
 sg13g2_decap_8 FILLER_80_2210 ();
 sg13g2_fill_2 FILLER_80_2217 ();
 sg13g2_fill_1 FILLER_80_2219 ();
 sg13g2_decap_8 FILLER_80_2228 ();
 sg13g2_decap_8 FILLER_80_2235 ();
 sg13g2_decap_8 FILLER_80_2242 ();
 sg13g2_decap_8 FILLER_80_2249 ();
 sg13g2_decap_8 FILLER_80_2256 ();
 sg13g2_decap_8 FILLER_80_2263 ();
 sg13g2_decap_8 FILLER_80_2270 ();
 sg13g2_decap_8 FILLER_80_2277 ();
 sg13g2_decap_8 FILLER_80_2288 ();
 sg13g2_decap_8 FILLER_80_2295 ();
 sg13g2_decap_8 FILLER_80_2302 ();
 sg13g2_decap_8 FILLER_80_2313 ();
 sg13g2_decap_8 FILLER_80_2320 ();
 sg13g2_decap_8 FILLER_80_2327 ();
 sg13g2_decap_8 FILLER_80_2334 ();
 sg13g2_decap_8 FILLER_80_2341 ();
 sg13g2_decap_8 FILLER_80_2348 ();
 sg13g2_decap_8 FILLER_80_2355 ();
 sg13g2_decap_8 FILLER_80_2362 ();
 sg13g2_fill_2 FILLER_80_2369 ();
 sg13g2_fill_1 FILLER_80_2371 ();
 sg13g2_decap_4 FILLER_80_2376 ();
 sg13g2_decap_8 FILLER_80_2384 ();
 sg13g2_decap_8 FILLER_80_2391 ();
 sg13g2_decap_4 FILLER_80_2398 ();
 sg13g2_fill_2 FILLER_80_2402 ();
 sg13g2_decap_8 FILLER_80_2434 ();
 sg13g2_decap_8 FILLER_80_2441 ();
 sg13g2_fill_1 FILLER_80_2448 ();
 sg13g2_fill_1 FILLER_80_2453 ();
 sg13g2_decap_8 FILLER_80_2458 ();
 sg13g2_decap_8 FILLER_80_2465 ();
 sg13g2_decap_8 FILLER_80_2472 ();
 sg13g2_fill_1 FILLER_80_2479 ();
 sg13g2_decap_8 FILLER_80_2488 ();
 sg13g2_decap_8 FILLER_80_2495 ();
 sg13g2_decap_8 FILLER_80_2502 ();
 sg13g2_fill_2 FILLER_80_2509 ();
 sg13g2_fill_2 FILLER_80_2519 ();
 sg13g2_fill_1 FILLER_80_2521 ();
 sg13g2_decap_8 FILLER_80_2526 ();
 sg13g2_decap_4 FILLER_80_2533 ();
 sg13g2_fill_2 FILLER_80_2537 ();
 sg13g2_fill_1 FILLER_80_2543 ();
 sg13g2_decap_8 FILLER_80_2552 ();
 sg13g2_decap_8 FILLER_80_2559 ();
 sg13g2_fill_2 FILLER_80_2566 ();
 sg13g2_fill_1 FILLER_80_2603 ();
 sg13g2_fill_2 FILLER_80_2624 ();
 sg13g2_decap_8 FILLER_80_2649 ();
 sg13g2_decap_8 FILLER_80_2656 ();
 sg13g2_decap_8 FILLER_80_2663 ();
endmodule
