module tt_um_fountaincoder_top_V2 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire clknet_leaf_0_clk;
 wire net151;
 wire \madd.count[0] ;
 wire \madd.count[10] ;
 wire \madd.count[11] ;
 wire \madd.count[1] ;
 wire \madd.count[2] ;
 wire \madd.count[3] ;
 wire \madd.count[4] ;
 wire \madd.count[5] ;
 wire \madd.count[6] ;
 wire \madd.count[7] ;
 wire \madd.count[8] ;
 wire \madd.count[9] ;
 wire \madd.delta[0] ;
 wire \madd.delta[10] ;
 wire \madd.delta[11] ;
 wire \madd.delta[1] ;
 wire \madd.delta[2] ;
 wire \madd.delta[3] ;
 wire \madd.delta[4] ;
 wire \madd.delta[5] ;
 wire \madd.delta[6] ;
 wire \madd.delta[7] ;
 wire \madd.delta[8] ;
 wire \madd.delta[9] ;
 wire \madd.i[0] ;
 wire \madd.i[1] ;
 wire \madd.i[2] ;
 wire \madd.i[3] ;
 wire \madd.i_d[0] ;
 wire \madd.i_e[0] ;
 wire \madd.mem[0][0] ;
 wire \madd.mem[0][10] ;
 wire \madd.mem[0][11] ;
 wire \madd.mem[0][1] ;
 wire \madd.mem[0][2] ;
 wire \madd.mem[0][3] ;
 wire \madd.mem[0][4] ;
 wire \madd.mem[0][5] ;
 wire \madd.mem[0][6] ;
 wire \madd.mem[0][7] ;
 wire \madd.mem[0][8] ;
 wire \madd.mem[0][9] ;
 wire \madd.mem[10][0] ;
 wire \madd.mem[10][10] ;
 wire \madd.mem[10][11] ;
 wire \madd.mem[10][1] ;
 wire \madd.mem[10][2] ;
 wire \madd.mem[10][3] ;
 wire \madd.mem[10][4] ;
 wire \madd.mem[10][5] ;
 wire \madd.mem[10][6] ;
 wire \madd.mem[10][7] ;
 wire \madd.mem[10][8] ;
 wire \madd.mem[10][9] ;
 wire \madd.mem[11][0] ;
 wire \madd.mem[11][10] ;
 wire \madd.mem[11][11] ;
 wire \madd.mem[11][1] ;
 wire \madd.mem[11][2] ;
 wire \madd.mem[11][3] ;
 wire \madd.mem[11][4] ;
 wire \madd.mem[11][5] ;
 wire \madd.mem[11][6] ;
 wire \madd.mem[11][7] ;
 wire \madd.mem[11][8] ;
 wire \madd.mem[11][9] ;
 wire \madd.mem[12][0] ;
 wire \madd.mem[12][10] ;
 wire \madd.mem[12][11] ;
 wire \madd.mem[12][1] ;
 wire \madd.mem[12][2] ;
 wire \madd.mem[12][3] ;
 wire \madd.mem[12][4] ;
 wire \madd.mem[12][5] ;
 wire \madd.mem[12][6] ;
 wire \madd.mem[12][7] ;
 wire \madd.mem[12][8] ;
 wire \madd.mem[12][9] ;
 wire \madd.mem[13][0] ;
 wire \madd.mem[13][10] ;
 wire \madd.mem[13][11] ;
 wire \madd.mem[13][1] ;
 wire \madd.mem[13][2] ;
 wire \madd.mem[13][3] ;
 wire \madd.mem[13][4] ;
 wire \madd.mem[13][5] ;
 wire \madd.mem[13][6] ;
 wire \madd.mem[13][7] ;
 wire \madd.mem[13][8] ;
 wire \madd.mem[13][9] ;
 wire \madd.mem[14][0] ;
 wire \madd.mem[14][10] ;
 wire \madd.mem[14][11] ;
 wire \madd.mem[14][1] ;
 wire \madd.mem[14][2] ;
 wire \madd.mem[14][3] ;
 wire \madd.mem[14][4] ;
 wire \madd.mem[14][5] ;
 wire \madd.mem[14][6] ;
 wire \madd.mem[14][7] ;
 wire \madd.mem[14][8] ;
 wire \madd.mem[14][9] ;
 wire \madd.mem[15][0] ;
 wire \madd.mem[15][10] ;
 wire \madd.mem[15][11] ;
 wire \madd.mem[15][1] ;
 wire \madd.mem[15][2] ;
 wire \madd.mem[15][3] ;
 wire \madd.mem[15][4] ;
 wire \madd.mem[15][5] ;
 wire \madd.mem[15][6] ;
 wire \madd.mem[15][7] ;
 wire \madd.mem[15][8] ;
 wire \madd.mem[15][9] ;
 wire \madd.mem[1][0] ;
 wire \madd.mem[1][10] ;
 wire \madd.mem[1][11] ;
 wire \madd.mem[1][1] ;
 wire \madd.mem[1][2] ;
 wire \madd.mem[1][3] ;
 wire \madd.mem[1][4] ;
 wire \madd.mem[1][5] ;
 wire \madd.mem[1][6] ;
 wire \madd.mem[1][7] ;
 wire \madd.mem[1][8] ;
 wire \madd.mem[1][9] ;
 wire \madd.mem[2][0] ;
 wire \madd.mem[2][10] ;
 wire \madd.mem[2][11] ;
 wire \madd.mem[2][1] ;
 wire \madd.mem[2][2] ;
 wire \madd.mem[2][3] ;
 wire \madd.mem[2][4] ;
 wire \madd.mem[2][5] ;
 wire \madd.mem[2][6] ;
 wire \madd.mem[2][7] ;
 wire \madd.mem[2][8] ;
 wire \madd.mem[2][9] ;
 wire \madd.mem[3][0] ;
 wire \madd.mem[3][10] ;
 wire \madd.mem[3][11] ;
 wire \madd.mem[3][1] ;
 wire \madd.mem[3][2] ;
 wire \madd.mem[3][3] ;
 wire \madd.mem[3][4] ;
 wire \madd.mem[3][5] ;
 wire \madd.mem[3][6] ;
 wire \madd.mem[3][7] ;
 wire \madd.mem[3][8] ;
 wire \madd.mem[3][9] ;
 wire \madd.mem[4][0] ;
 wire \madd.mem[4][10] ;
 wire \madd.mem[4][11] ;
 wire \madd.mem[4][1] ;
 wire \madd.mem[4][2] ;
 wire \madd.mem[4][3] ;
 wire \madd.mem[4][4] ;
 wire \madd.mem[4][5] ;
 wire \madd.mem[4][6] ;
 wire \madd.mem[4][7] ;
 wire \madd.mem[4][8] ;
 wire \madd.mem[4][9] ;
 wire \madd.mem[5][0] ;
 wire \madd.mem[5][10] ;
 wire \madd.mem[5][11] ;
 wire \madd.mem[5][1] ;
 wire \madd.mem[5][2] ;
 wire \madd.mem[5][3] ;
 wire \madd.mem[5][4] ;
 wire \madd.mem[5][5] ;
 wire \madd.mem[5][6] ;
 wire \madd.mem[5][7] ;
 wire \madd.mem[5][8] ;
 wire \madd.mem[5][9] ;
 wire \madd.mem[6][0] ;
 wire \madd.mem[6][10] ;
 wire \madd.mem[6][11] ;
 wire \madd.mem[6][1] ;
 wire \madd.mem[6][2] ;
 wire \madd.mem[6][3] ;
 wire \madd.mem[6][4] ;
 wire \madd.mem[6][5] ;
 wire \madd.mem[6][6] ;
 wire \madd.mem[6][7] ;
 wire \madd.mem[6][8] ;
 wire \madd.mem[6][9] ;
 wire \madd.mem[7][0] ;
 wire \madd.mem[7][10] ;
 wire \madd.mem[7][11] ;
 wire \madd.mem[7][1] ;
 wire \madd.mem[7][2] ;
 wire \madd.mem[7][3] ;
 wire \madd.mem[7][4] ;
 wire \madd.mem[7][5] ;
 wire \madd.mem[7][6] ;
 wire \madd.mem[7][7] ;
 wire \madd.mem[7][8] ;
 wire \madd.mem[7][9] ;
 wire \madd.mem[8][0] ;
 wire \madd.mem[8][10] ;
 wire \madd.mem[8][11] ;
 wire \madd.mem[8][1] ;
 wire \madd.mem[8][2] ;
 wire \madd.mem[8][3] ;
 wire \madd.mem[8][4] ;
 wire \madd.mem[8][5] ;
 wire \madd.mem[8][6] ;
 wire \madd.mem[8][7] ;
 wire \madd.mem[8][8] ;
 wire \madd.mem[8][9] ;
 wire \madd.mem[9][0] ;
 wire \madd.mem[9][10] ;
 wire \madd.mem[9][11] ;
 wire \madd.mem[9][1] ;
 wire \madd.mem[9][2] ;
 wire \madd.mem[9][3] ;
 wire \madd.mem[9][4] ;
 wire \madd.mem[9][5] ;
 wire \madd.mem[9][6] ;
 wire \madd.mem[9][7] ;
 wire \madd.mem[9][8] ;
 wire \madd.mem[9][9] ;
 wire \madd.set ;
 wire \madd.total[0] ;
 wire \madd.total[10] ;
 wire \madd.total[11] ;
 wire \madd.total[1] ;
 wire \madd.total[2] ;
 wire \madd.total[3] ;
 wire \madd.total[4] ;
 wire \madd.total[5] ;
 wire \madd.total[6] ;
 wire \madd.total[7] ;
 wire \madd.total[8] ;
 wire \madd.total[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sg13g2_buf_8 _2117_ (.A(uio_in[0]),
    .X(_1751_));
 sg13g2_buf_1 _2118_ (.A(uio_in[1]),
    .X(_1752_));
 sg13g2_buf_8 _2119_ (.A(uio_in[3]),
    .X(_1753_));
 sg13g2_buf_8 _2120_ (.A(uio_in[2]),
    .X(_1754_));
 sg13g2_nor3_2 _2121_ (.A(net142),
    .B(_1753_),
    .C(_1754_),
    .Y(_1755_));
 sg13g2_buf_1 _2122_ (.A(rst_n),
    .X(_1756_));
 sg13g2_inv_1 _2123_ (.Y(_1757_),
    .A(_1756_));
 sg13g2_buf_1 _2124_ (.A(_1757_),
    .X(_1758_));
 sg13g2_a21oi_2 _2125_ (.B1(net132),
    .Y(_1759_),
    .A2(_1755_),
    .A1(_1751_));
 sg13g2_buf_2 _2126_ (.A(\madd.i[0] ),
    .X(_1760_));
 sg13g2_buf_1 _2127_ (.A(_1760_),
    .X(_1761_));
 sg13g2_buf_1 _2128_ (.A(\madd.i_d[0] ),
    .X(_1762_));
 sg13g2_nand2_1 _2129_ (.Y(_1763_),
    .A(_1751_),
    .B(_1752_));
 sg13g2_nor2_1 _2130_ (.A(_1757_),
    .B(_1754_),
    .Y(_1764_));
 sg13g2_nand3_1 _2131_ (.B(_1763_),
    .C(_1764_),
    .A(_1753_),
    .Y(_1765_));
 sg13g2_buf_1 _2132_ (.A(_1765_),
    .X(_1766_));
 sg13g2_inv_1 _2133_ (.Y(_1767_),
    .A(_1751_));
 sg13g2_nand2_1 _2134_ (.Y(_1768_),
    .A(_1767_),
    .B(_1753_));
 sg13g2_a21oi_1 _2135_ (.A1(net142),
    .A2(_1768_),
    .Y(_1769_),
    .B1(_1754_));
 sg13g2_buf_1 _2136_ (.A(_1756_),
    .X(_1770_));
 sg13g2_nand2b_1 _2137_ (.Y(_1771_),
    .B(_1770_),
    .A_N(_1769_));
 sg13g2_o21ai_1 _2138_ (.B1(_1771_),
    .Y(_1772_),
    .A1(_1762_),
    .A2(_1766_));
 sg13g2_nor2b_2 _2139_ (.A(_1761_),
    .B_N(_1762_),
    .Y(_1773_));
 sg13g2_inv_1 _2140_ (.Y(_1774_),
    .A(_1766_));
 sg13g2_a22oi_1 _2141_ (.Y(_1775_),
    .B1(_1773_),
    .B2(_1774_),
    .A2(_1772_),
    .A1(_1761_));
 sg13g2_nand2_1 _2142_ (.Y(_0004_),
    .A(_1759_),
    .B(_1775_));
 sg13g2_buf_1 _2143_ (.A(\madd.i[1] ),
    .X(_1776_));
 sg13g2_xor2_1 _2144_ (.B(net142),
    .A(_1751_),
    .X(_1777_));
 sg13g2_nand3_1 _2145_ (.B(_1764_),
    .C(_1777_),
    .A(_1753_),
    .Y(_1778_));
 sg13g2_nand2_1 _2146_ (.Y(_1779_),
    .A(_1762_),
    .B(_1778_));
 sg13g2_xnor2_1 _2147_ (.Y(_1780_),
    .A(_1773_),
    .B(_1779_));
 sg13g2_o21ai_1 _2148_ (.B1(_1771_),
    .Y(_1781_),
    .A1(_1766_),
    .A2(_1780_));
 sg13g2_nor2_1 _2149_ (.A(net139),
    .B(_1766_),
    .Y(_1782_));
 sg13g2_a22oi_1 _2150_ (.Y(_1783_),
    .B1(_1782_),
    .B2(_1780_),
    .A2(_1781_),
    .A1(_1776_));
 sg13g2_nand2_1 _2151_ (.Y(_0005_),
    .A(_1759_),
    .B(_1783_));
 sg13g2_buf_2 _2152_ (.A(\madd.i[2] ),
    .X(_1784_));
 sg13g2_inv_1 _2153_ (.Y(_1785_),
    .A(_1776_));
 sg13g2_and2_1 _2154_ (.A(_1785_),
    .B(_1773_),
    .X(_1786_));
 sg13g2_nor3_1 _2155_ (.A(_1785_),
    .B(_1773_),
    .C(_1779_),
    .Y(_1787_));
 sg13g2_a21oi_1 _2156_ (.A1(_1779_),
    .A2(_1786_),
    .Y(_1788_),
    .B1(_1787_));
 sg13g2_inv_1 _2157_ (.Y(_1789_),
    .A(_1771_));
 sg13g2_a21o_1 _2158_ (.A2(_1788_),
    .A1(_1774_),
    .B1(_1789_),
    .X(_1790_));
 sg13g2_nor3_1 _2159_ (.A(_1784_),
    .B(_1766_),
    .C(_1788_),
    .Y(_1791_));
 sg13g2_a21oi_1 _2160_ (.A1(_1784_),
    .A2(_1790_),
    .Y(_1792_),
    .B1(_1791_));
 sg13g2_nand2_1 _2161_ (.Y(_0006_),
    .A(_1759_),
    .B(_1792_));
 sg13g2_buf_1 _2162_ (.A(_0162_),
    .X(_1793_));
 sg13g2_buf_2 _2163_ (.A(_0157_),
    .X(_1794_));
 sg13g2_inv_1 _2164_ (.Y(_1795_),
    .A(_1794_));
 sg13g2_a21oi_1 _2165_ (.A1(_1762_),
    .A2(_1778_),
    .Y(_1796_),
    .B1(_1795_));
 sg13g2_or2_1 _2166_ (.X(_1797_),
    .B(_1796_),
    .A(_1787_));
 sg13g2_a22oi_1 _2167_ (.Y(_1798_),
    .B1(_1797_),
    .B2(_1784_),
    .A2(_1796_),
    .A1(_1786_));
 sg13g2_xnor2_1 _2168_ (.Y(_1799_),
    .A(net138),
    .B(_1798_));
 sg13g2_inv_1 _2169_ (.Y(_1800_),
    .A(_1759_));
 sg13g2_a21oi_1 _2170_ (.A1(\madd.i[3] ),
    .A2(_1789_),
    .Y(_1801_),
    .B1(_1800_));
 sg13g2_o21ai_1 _2171_ (.B1(_1801_),
    .Y(_0007_),
    .A1(_1766_),
    .A2(_1799_));
 sg13g2_buf_1 _2172_ (.A(_1770_),
    .X(_1802_));
 sg13g2_buf_2 _2173_ (.A(\madd.count[0] ),
    .X(_1803_));
 sg13g2_nand3b_1 _2174_ (.B(net142),
    .C(_1753_),
    .Y(_1804_),
    .A_N(_1751_));
 sg13g2_buf_1 _2175_ (.A(_1804_),
    .X(_1805_));
 sg13g2_buf_8 _2176_ (.A(_1805_),
    .X(_1806_));
 sg13g2_nor2_1 _2177_ (.A(_1754_),
    .B(net118),
    .Y(_1807_));
 sg13g2_buf_1 _2178_ (.A(_1807_),
    .X(_1808_));
 sg13g2_buf_1 _2179_ (.A(net102),
    .X(_1809_));
 sg13g2_nand2_1 _2180_ (.Y(_1810_),
    .A(\madd.delta[0] ),
    .B(_1809_));
 sg13g2_xnor2_1 _2181_ (.Y(_1811_),
    .A(_1803_),
    .B(_1810_));
 sg13g2_and2_1 _2182_ (.A(net130),
    .B(_1811_),
    .X(_0187_));
 sg13g2_buf_1 _2183_ (.A(\madd.count[10] ),
    .X(_1812_));
 sg13g2_and2_1 _2184_ (.A(net140),
    .B(net137),
    .X(_1813_));
 sg13g2_buf_1 _2185_ (.A(net132),
    .X(_1814_));
 sg13g2_nor2_1 _2186_ (.A(net117),
    .B(_1812_),
    .Y(_1815_));
 sg13g2_or2_1 _2187_ (.X(_1816_),
    .B(net118),
    .A(_1754_));
 sg13g2_buf_1 _2188_ (.A(_1816_),
    .X(_1817_));
 sg13g2_buf_1 _2189_ (.A(_1817_),
    .X(_1818_));
 sg13g2_buf_2 _2190_ (.A(\madd.delta[10] ),
    .X(_1819_));
 sg13g2_buf_2 _2191_ (.A(\madd.delta[9] ),
    .X(_1820_));
 sg13g2_inv_1 _2192_ (.Y(_1821_),
    .A(_1820_));
 sg13g2_buf_2 _2193_ (.A(\madd.count[8] ),
    .X(_1822_));
 sg13g2_buf_1 _2194_ (.A(\madd.delta[8] ),
    .X(_1823_));
 sg13g2_buf_1 _2195_ (.A(\madd.delta[7] ),
    .X(_1824_));
 sg13g2_inv_1 _2196_ (.Y(_1825_),
    .A(_1824_));
 sg13g2_buf_2 _2197_ (.A(\madd.delta[6] ),
    .X(_1826_));
 sg13g2_buf_1 _2198_ (.A(\madd.count[5] ),
    .X(_1827_));
 sg13g2_inv_1 _2199_ (.Y(_1828_),
    .A(\madd.delta[5] ));
 sg13g2_buf_1 _2200_ (.A(\madd.delta[4] ),
    .X(_1829_));
 sg13g2_buf_1 _2201_ (.A(\madd.count[3] ),
    .X(_1830_));
 sg13g2_inv_1 _2202_ (.Y(_1831_),
    .A(_1830_));
 sg13g2_buf_1 _2203_ (.A(\madd.delta[3] ),
    .X(_1832_));
 sg13g2_buf_2 _2204_ (.A(\madd.count[1] ),
    .X(_1833_));
 sg13g2_buf_2 _2205_ (.A(\madd.delta[1] ),
    .X(_1834_));
 sg13g2_nor2_1 _2206_ (.A(_1833_),
    .B(_1834_),
    .Y(_1835_));
 sg13g2_a22oi_1 _2207_ (.Y(_1836_),
    .B1(\madd.delta[0] ),
    .B2(_1803_),
    .A2(_1834_),
    .A1(_1833_));
 sg13g2_buf_1 _2208_ (.A(\madd.count[2] ),
    .X(_1837_));
 sg13g2_nor2_1 _2209_ (.A(_1837_),
    .B(\madd.delta[2] ),
    .Y(_1838_));
 sg13g2_nor3_1 _2210_ (.A(_1835_),
    .B(_1836_),
    .C(_1838_),
    .Y(_1839_));
 sg13g2_inv_1 _2211_ (.Y(_1840_),
    .A(_1837_));
 sg13g2_inv_1 _2212_ (.Y(_1841_),
    .A(\madd.delta[2] ));
 sg13g2_nor2_1 _2213_ (.A(_1840_),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_nor3_1 _2214_ (.A(_1832_),
    .B(_1839_),
    .C(_1842_),
    .Y(_1843_));
 sg13g2_o21ai_1 _2215_ (.B1(_1832_),
    .Y(_1844_),
    .A1(_1839_),
    .A2(_1842_));
 sg13g2_o21ai_1 _2216_ (.B1(_1844_),
    .Y(_1845_),
    .A1(_1831_),
    .A2(_1843_));
 sg13g2_nand2_1 _2217_ (.Y(_1846_),
    .A(_1829_),
    .B(_1845_));
 sg13g2_o21ai_1 _2218_ (.B1(\madd.count[4] ),
    .Y(_1847_),
    .A1(_1829_),
    .A2(_1845_));
 sg13g2_nand3_1 _2219_ (.B(_1846_),
    .C(_1847_),
    .A(_1828_),
    .Y(_1848_));
 sg13g2_a21oi_1 _2220_ (.A1(_1846_),
    .A2(_1847_),
    .Y(_1849_),
    .B1(_1828_));
 sg13g2_a21o_1 _2221_ (.A2(_1848_),
    .A1(_1827_),
    .B1(_1849_),
    .X(_1850_));
 sg13g2_nand2_1 _2222_ (.Y(_1851_),
    .A(_1826_),
    .B(_1850_));
 sg13g2_o21ai_1 _2223_ (.B1(\madd.count[6] ),
    .Y(_1852_),
    .A1(_1826_),
    .A2(_1850_));
 sg13g2_nand3_1 _2224_ (.B(_1851_),
    .C(_1852_),
    .A(_1825_),
    .Y(_1853_));
 sg13g2_a21oi_1 _2225_ (.A1(_1851_),
    .A2(_1852_),
    .Y(_1854_),
    .B1(_1825_));
 sg13g2_a221oi_1 _2226_ (.B2(\madd.count[7] ),
    .C1(_1854_),
    .B1(_1853_),
    .A1(_1822_),
    .Y(_1855_),
    .A2(_1823_));
 sg13g2_nor2_1 _2227_ (.A(_1822_),
    .B(_1823_),
    .Y(_1856_));
 sg13g2_nor3_1 _2228_ (.A(_1821_),
    .B(_1855_),
    .C(_1856_),
    .Y(_1857_));
 sg13g2_o21ai_1 _2229_ (.B1(_1821_),
    .Y(_1858_),
    .A1(_1855_),
    .A2(_1856_));
 sg13g2_o21ai_1 _2230_ (.B1(_1858_),
    .Y(_1859_),
    .A1(\madd.count[9] ),
    .A2(_1857_));
 sg13g2_xor2_1 _2231_ (.B(_1859_),
    .A(_1819_),
    .X(_1860_));
 sg13g2_nor2_1 _2232_ (.A(net92),
    .B(_1860_),
    .Y(_1861_));
 sg13g2_mux2_1 _2233_ (.A0(_1813_),
    .A1(_1815_),
    .S(_1861_),
    .X(_0188_));
 sg13g2_buf_1 _2234_ (.A(\madd.count[11] ),
    .X(_1862_));
 sg13g2_and2_1 _2235_ (.A(net140),
    .B(_1862_),
    .X(_1863_));
 sg13g2_nor2_1 _2236_ (.A(_1758_),
    .B(_1862_),
    .Y(_1864_));
 sg13g2_and2_1 _2237_ (.A(\madd.delta[11] ),
    .B(net102),
    .X(_1865_));
 sg13g2_nor2_1 _2238_ (.A(\madd.delta[11] ),
    .B(_1817_),
    .Y(_1866_));
 sg13g2_nand2_1 _2239_ (.Y(_1867_),
    .A(net137),
    .B(_1819_));
 sg13g2_nor2_1 _2240_ (.A(net137),
    .B(_1819_),
    .Y(_1868_));
 sg13g2_a21oi_1 _2241_ (.A1(_1859_),
    .A2(_1867_),
    .Y(_1869_),
    .B1(_1868_));
 sg13g2_mux2_1 _2242_ (.A0(_1865_),
    .A1(_1866_),
    .S(_1869_),
    .X(_1870_));
 sg13g2_mux2_1 _2243_ (.A0(_1863_),
    .A1(_1864_),
    .S(_1870_),
    .X(_0189_));
 sg13g2_buf_1 _2244_ (.A(net117),
    .X(_1871_));
 sg13g2_nand2_1 _2245_ (.Y(_1872_),
    .A(_1803_),
    .B(\madd.delta[0] ));
 sg13g2_xor2_1 _2246_ (.B(_1872_),
    .A(_1834_),
    .X(_1873_));
 sg13g2_nor2_1 _2247_ (.A(net92),
    .B(_1873_),
    .Y(_1874_));
 sg13g2_xnor2_1 _2248_ (.Y(_1875_),
    .A(_1833_),
    .B(_1874_));
 sg13g2_nor2_1 _2249_ (.A(net109),
    .B(_1875_),
    .Y(_0190_));
 sg13g2_nor2_1 _2250_ (.A(_1835_),
    .B(_1836_),
    .Y(_1876_));
 sg13g2_xnor2_1 _2251_ (.Y(_1877_),
    .A(\madd.delta[2] ),
    .B(_1876_));
 sg13g2_nor2_1 _2252_ (.A(_1818_),
    .B(_1877_),
    .Y(_1878_));
 sg13g2_xnor2_1 _2253_ (.Y(_1879_),
    .A(_1837_),
    .B(_1878_));
 sg13g2_nor2_1 _2254_ (.A(_1871_),
    .B(_1879_),
    .Y(_0191_));
 sg13g2_nand3b_1 _2255_ (.B(_1844_),
    .C(net93),
    .Y(_1880_),
    .A_N(_1843_));
 sg13g2_xnor2_1 _2256_ (.Y(_1881_),
    .A(_1831_),
    .B(_1880_));
 sg13g2_nor2_1 _2257_ (.A(net109),
    .B(_1881_),
    .Y(_0192_));
 sg13g2_or2_1 _2258_ (.X(_1882_),
    .B(_1845_),
    .A(_1829_));
 sg13g2_and3_1 _2259_ (.X(_1883_),
    .A(_1808_),
    .B(_1882_),
    .C(_1846_));
 sg13g2_xnor2_1 _2260_ (.Y(_1884_),
    .A(\madd.count[4] ),
    .B(_1883_));
 sg13g2_nor2_1 _2261_ (.A(net109),
    .B(_1884_),
    .Y(_0193_));
 sg13g2_nand3b_1 _2262_ (.B(net93),
    .C(_1848_),
    .Y(_1885_),
    .A_N(_1849_));
 sg13g2_xor2_1 _2263_ (.B(_1885_),
    .A(_1827_),
    .X(_1886_));
 sg13g2_nor2_1 _2264_ (.A(_1871_),
    .B(_1886_),
    .Y(_0194_));
 sg13g2_or2_1 _2265_ (.X(_1887_),
    .B(_1850_),
    .A(_1826_));
 sg13g2_and3_1 _2266_ (.X(_1888_),
    .A(net102),
    .B(_1887_),
    .C(_1851_));
 sg13g2_xnor2_1 _2267_ (.Y(_1889_),
    .A(\madd.count[6] ),
    .B(_1888_));
 sg13g2_nor2_1 _2268_ (.A(net109),
    .B(_1889_),
    .Y(_0195_));
 sg13g2_inv_2 _2269_ (.Y(_1890_),
    .A(\madd.count[7] ));
 sg13g2_nand3b_1 _2270_ (.B(net93),
    .C(_1853_),
    .Y(_1891_),
    .A_N(_1854_));
 sg13g2_xnor2_1 _2271_ (.Y(_1892_),
    .A(_1890_),
    .B(_1891_));
 sg13g2_nor2_1 _2272_ (.A(net109),
    .B(_1892_),
    .Y(_0196_));
 sg13g2_buf_1 _2273_ (.A(_1817_),
    .X(_1893_));
 sg13g2_inv_2 _2274_ (.Y(_1894_),
    .A(_1823_));
 sg13g2_a21oi_1 _2275_ (.A1(\madd.count[7] ),
    .A2(_1853_),
    .Y(_1895_),
    .B1(_1854_));
 sg13g2_xnor2_1 _2276_ (.Y(_1896_),
    .A(_1894_),
    .B(_1895_));
 sg13g2_nor2_1 _2277_ (.A(net91),
    .B(_1896_),
    .Y(_1897_));
 sg13g2_xnor2_1 _2278_ (.Y(_1898_),
    .A(_1822_),
    .B(_1897_));
 sg13g2_nor2_1 _2279_ (.A(net109),
    .B(_1898_),
    .Y(_0197_));
 sg13g2_inv_1 _2280_ (.Y(_1899_),
    .A(\madd.count[9] ));
 sg13g2_nand3b_1 _2281_ (.B(_1858_),
    .C(net93),
    .Y(_1900_),
    .A_N(_1857_));
 sg13g2_xnor2_1 _2282_ (.Y(_1901_),
    .A(_1899_),
    .B(_1900_));
 sg13g2_nor2_1 _2283_ (.A(net109),
    .B(_1901_),
    .Y(_0198_));
 sg13g2_nand2b_1 _2284_ (.Y(_1902_),
    .B(_1756_),
    .A_N(_1754_));
 sg13g2_buf_8 _2285_ (.A(_1902_),
    .X(_1903_));
 sg13g2_or2_1 _2286_ (.X(_1904_),
    .B(net118),
    .A(net129));
 sg13g2_buf_8 _2287_ (.A(_1904_),
    .X(_1905_));
 sg13g2_buf_8 _2288_ (.A(_1905_),
    .X(_1906_));
 sg13g2_nand2b_1 _2289_ (.Y(_1907_),
    .B(net139),
    .A_N(_1760_));
 sg13g2_buf_1 _2290_ (.A(_1907_),
    .X(_1908_));
 sg13g2_nand2b_1 _2291_ (.Y(_1909_),
    .B(net131),
    .A_N(net139));
 sg13g2_buf_1 _2292_ (.A(_1909_),
    .X(_1910_));
 sg13g2_o21ai_1 _2293_ (.B1(net108),
    .Y(_1911_),
    .A1(_0168_),
    .A2(net116));
 sg13g2_buf_4 _2294_ (.X(_1912_),
    .A(ui_in[4]));
 sg13g2_buf_8 _2295_ (.A(_1912_),
    .X(_1913_));
 sg13g2_buf_1 _2296_ (.A(net136),
    .X(_1914_));
 sg13g2_buf_8 _2297_ (.A(ui_in[5]),
    .X(_1915_));
 sg13g2_buf_1 _2298_ (.A(net141),
    .X(_1916_));
 sg13g2_a21oi_1 _2299_ (.A1(_1914_),
    .A2(_0168_),
    .Y(_1917_),
    .B1(_1916_));
 sg13g2_mux2_1 _2300_ (.A0(_1911_),
    .A1(_1917_),
    .S(net101),
    .X(_1918_));
 sg13g2_or2_1 _2301_ (.X(_1919_),
    .B(\madd.i[1] ),
    .A(_1760_));
 sg13g2_buf_1 _2302_ (.A(_1919_),
    .X(_1920_));
 sg13g2_buf_1 _2303_ (.A(_1920_),
    .X(_1921_));
 sg13g2_nand2_1 _2304_ (.Y(_1922_),
    .A(net131),
    .B(net139));
 sg13g2_buf_2 _2305_ (.A(_1922_),
    .X(_1923_));
 sg13g2_o21ai_1 _2306_ (.B1(_1923_),
    .Y(_1924_),
    .A1(_0170_),
    .A2(net107));
 sg13g2_inv_2 _2307_ (.Y(_1925_),
    .A(_1915_));
 sg13g2_a21oi_1 _2308_ (.A1(net128),
    .A2(_0170_),
    .Y(_1926_),
    .B1(_1925_));
 sg13g2_mux2_1 _2309_ (.A0(_1924_),
    .A1(_1926_),
    .S(net101),
    .X(_1927_));
 sg13g2_inv_1 _2310_ (.Y(_1928_),
    .A(_1912_));
 sg13g2_o21ai_1 _2311_ (.B1(_1928_),
    .Y(_1929_),
    .A1(net129),
    .A2(_1805_));
 sg13g2_buf_2 _2312_ (.A(_1929_),
    .X(_1930_));
 sg13g2_inv_1 _2313_ (.Y(_1931_),
    .A(_1760_));
 sg13g2_or3_1 _2314_ (.A(_1931_),
    .B(net129),
    .C(_1805_),
    .X(_1932_));
 sg13g2_buf_2 _2315_ (.A(_1932_),
    .X(_1933_));
 sg13g2_and2_1 _2316_ (.A(_1930_),
    .B(_1933_),
    .X(_1934_));
 sg13g2_buf_1 _2317_ (.A(_1934_),
    .X(_1935_));
 sg13g2_o21ai_1 _2318_ (.B1(_1935_),
    .Y(_1936_),
    .A1(_1918_),
    .A2(_1927_));
 sg13g2_nand2b_1 _2319_ (.Y(_1937_),
    .B(_1927_),
    .A_N(_0169_));
 sg13g2_xnor2_1 _2320_ (.Y(_1938_),
    .A(_1784_),
    .B(net138));
 sg13g2_nor2_1 _2321_ (.A(_1920_),
    .B(_1938_),
    .Y(_1939_));
 sg13g2_nor2_2 _2322_ (.A(_1760_),
    .B(\madd.i[1] ),
    .Y(_1940_));
 sg13g2_nor3_1 _2323_ (.A(_1794_),
    .B(net138),
    .C(_1940_),
    .Y(_1941_));
 sg13g2_a21oi_1 _2324_ (.A1(_1794_),
    .A2(_1939_),
    .Y(_1942_),
    .B1(_1941_));
 sg13g2_buf_8 _2325_ (.A(net101),
    .X(_1943_));
 sg13g2_buf_2 _2326_ (.A(ui_in[6]),
    .X(_1944_));
 sg13g2_inv_2 _2327_ (.Y(_1945_),
    .A(_1944_));
 sg13g2_buf_2 _2328_ (.A(ui_in[7]),
    .X(_1946_));
 sg13g2_inv_1 _2329_ (.Y(_1947_),
    .A(_1946_));
 sg13g2_nor2_2 _2330_ (.A(_1945_),
    .B(_1947_),
    .Y(_1948_));
 sg13g2_nand2_1 _2331_ (.Y(_1949_),
    .A(net89),
    .B(_1948_));
 sg13g2_o21ai_1 _2332_ (.B1(_1949_),
    .Y(_1950_),
    .A1(net90),
    .A2(_1942_));
 sg13g2_nand2b_1 _2333_ (.Y(_1951_),
    .B(_1918_),
    .A_N(_0167_));
 sg13g2_nand4_1 _2334_ (.B(_1937_),
    .C(_1950_),
    .A(_1936_),
    .Y(_1952_),
    .D(_1951_));
 sg13g2_o21ai_1 _2335_ (.B1(_1923_),
    .Y(_1953_),
    .A1(_0156_),
    .A2(_1921_));
 sg13g2_a21oi_1 _2336_ (.A1(net136),
    .A2(_0156_),
    .Y(_1954_),
    .B1(_1925_));
 sg13g2_mux2_1 _2337_ (.A0(_1953_),
    .A1(_1954_),
    .S(net101),
    .X(_1955_));
 sg13g2_o21ai_1 _2338_ (.B1(net108),
    .Y(_1956_),
    .A1(_0154_),
    .A2(net116));
 sg13g2_a21oi_1 _2339_ (.A1(_1914_),
    .A2(_0154_),
    .Y(_1957_),
    .B1(net135));
 sg13g2_mux2_1 _2340_ (.A0(_1956_),
    .A1(_1957_),
    .S(_1905_),
    .X(_1958_));
 sg13g2_o21ai_1 _2341_ (.B1(_1935_),
    .Y(_1959_),
    .A1(_1955_),
    .A2(_1958_));
 sg13g2_nand2b_1 _2342_ (.Y(_1960_),
    .B(_1958_),
    .A_N(_0153_));
 sg13g2_nor2_1 _2343_ (.A(_1944_),
    .B(_1946_),
    .Y(_1961_));
 sg13g2_buf_1 _2344_ (.A(_1961_),
    .X(_1962_));
 sg13g2_nand3_1 _2345_ (.B(net138),
    .C(_1921_),
    .A(_1794_),
    .Y(_1963_));
 sg13g2_nand3_1 _2346_ (.B(_1940_),
    .C(_1938_),
    .A(_1795_),
    .Y(_1964_));
 sg13g2_a21oi_1 _2347_ (.A1(_1963_),
    .A2(_1964_),
    .Y(_1965_),
    .B1(_1943_));
 sg13g2_a21o_1 _2348_ (.A2(net127),
    .A1(net90),
    .B1(_1965_),
    .X(_1966_));
 sg13g2_nand2b_1 _2349_ (.Y(_1967_),
    .B(_1955_),
    .A_N(_0155_));
 sg13g2_nand4_1 _2350_ (.B(_1960_),
    .C(_1966_),
    .A(_1959_),
    .Y(_1968_),
    .D(_1967_));
 sg13g2_nor2_1 _2351_ (.A(_1903_),
    .B(net118),
    .Y(_1969_));
 sg13g2_buf_1 _2352_ (.A(_1969_),
    .X(_1970_));
 sg13g2_buf_1 _2353_ (.A(_1947_),
    .X(_1971_));
 sg13g2_nand2_2 _2354_ (.Y(_1972_),
    .A(_1944_),
    .B(net126));
 sg13g2_nand3_1 _2355_ (.B(_1940_),
    .C(_1938_),
    .A(_1794_),
    .Y(_1973_));
 sg13g2_nand3_1 _2356_ (.B(net138),
    .C(net107),
    .A(_1795_),
    .Y(_1974_));
 sg13g2_a21o_1 _2357_ (.A2(_1974_),
    .A1(_1973_),
    .B1(_1943_),
    .X(_1975_));
 sg13g2_o21ai_1 _2358_ (.B1(_1975_),
    .Y(_1976_),
    .A1(net100),
    .A2(_1972_));
 sg13g2_o21ai_1 _2359_ (.B1(net108),
    .Y(_1977_),
    .A1(_0159_),
    .A2(net116));
 sg13g2_a21oi_1 _2360_ (.A1(net128),
    .A2(_0159_),
    .Y(_1978_),
    .B1(net135));
 sg13g2_mux2_1 _2361_ (.A0(_1977_),
    .A1(_1978_),
    .S(net101),
    .X(_1979_));
 sg13g2_inv_1 _2362_ (.Y(_1980_),
    .A(_0158_));
 sg13g2_a21o_1 _2363_ (.A2(_1933_),
    .A1(_1930_),
    .B1(_1980_),
    .X(_1981_));
 sg13g2_o21ai_1 _2364_ (.B1(_1923_),
    .Y(_1982_),
    .A1(_0161_),
    .A2(net107));
 sg13g2_a21oi_1 _2365_ (.A1(net128),
    .A2(_0161_),
    .Y(_1983_),
    .B1(_1925_));
 sg13g2_mux2_1 _2366_ (.A0(_1982_),
    .A1(_1983_),
    .S(net101),
    .X(_1984_));
 sg13g2_inv_1 _2367_ (.Y(_1985_),
    .A(_0160_));
 sg13g2_a21o_1 _2368_ (.A2(_1933_),
    .A1(_1930_),
    .B1(_1985_),
    .X(_1986_));
 sg13g2_a22oi_1 _2369_ (.Y(_1987_),
    .B1(_1984_),
    .B2(_1986_),
    .A2(_1981_),
    .A1(_1979_));
 sg13g2_o21ai_1 _2370_ (.B1(_1923_),
    .Y(_1988_),
    .A1(_0166_),
    .A2(net107));
 sg13g2_and2_1 _2371_ (.A(net100),
    .B(_1988_),
    .X(_1989_));
 sg13g2_buf_1 _2372_ (.A(net128),
    .X(_1990_));
 sg13g2_buf_1 _2373_ (.A(net135),
    .X(_1991_));
 sg13g2_o21ai_1 _2374_ (.B1(net125),
    .Y(_1992_),
    .A1(net129),
    .A2(net118));
 sg13g2_a21oi_1 _2375_ (.A1(_1990_),
    .A2(_0166_),
    .Y(_1993_),
    .B1(_1992_));
 sg13g2_inv_1 _2376_ (.Y(_1994_),
    .A(_0165_));
 sg13g2_a21o_1 _2377_ (.A2(_1933_),
    .A1(_1930_),
    .B1(_1994_),
    .X(_1995_));
 sg13g2_o21ai_1 _2378_ (.B1(_1995_),
    .Y(_1996_),
    .A1(_1989_),
    .A2(_1993_));
 sg13g2_nor3_1 _2379_ (.A(_1795_),
    .B(net138),
    .C(_1940_),
    .Y(_1997_));
 sg13g2_a21oi_1 _2380_ (.A1(_1795_),
    .A2(_1939_),
    .Y(_1998_),
    .B1(_1997_));
 sg13g2_o21ai_1 _2381_ (.B1(net108),
    .Y(_1999_),
    .A1(_0164_),
    .A2(net116));
 sg13g2_a21oi_1 _2382_ (.A1(net128),
    .A2(_0164_),
    .Y(_2000_),
    .B1(net135));
 sg13g2_mux2_1 _2383_ (.A0(_1999_),
    .A1(_2000_),
    .S(net101),
    .X(_2001_));
 sg13g2_inv_1 _2384_ (.Y(_2002_),
    .A(_0163_));
 sg13g2_a21o_1 _2385_ (.A2(_1933_),
    .A1(_1930_),
    .B1(_2002_),
    .X(_2003_));
 sg13g2_nor2_2 _2386_ (.A(_1944_),
    .B(_1947_),
    .Y(_2004_));
 sg13g2_nor2_1 _2387_ (.A(net100),
    .B(_2004_),
    .Y(_2005_));
 sg13g2_a221oi_1 _2388_ (.B2(_2003_),
    .C1(_2005_),
    .B1(_2001_),
    .A1(net100),
    .Y(_2006_),
    .A2(_1998_));
 sg13g2_a22oi_1 _2389_ (.Y(_2007_),
    .B1(_1996_),
    .B2(_2006_),
    .A2(_1987_),
    .A1(_1976_));
 sg13g2_nand3_1 _2390_ (.B(_1968_),
    .C(_2007_),
    .A(_1952_),
    .Y(_2008_));
 sg13g2_xnor2_1 _2391_ (.Y(_2009_),
    .A(_0152_),
    .B(_2008_));
 sg13g2_nand3_1 _2392_ (.B(\madd.delta[0] ),
    .C(net92),
    .A(_1802_),
    .Y(_2010_));
 sg13g2_o21ai_1 _2393_ (.B1(_2010_),
    .Y(_0199_),
    .A1(_1906_),
    .A2(_2009_));
 sg13g2_nand2_1 _2394_ (.Y(_2011_),
    .A(_1930_),
    .B(_1933_));
 sg13g2_buf_2 _2395_ (.A(_2011_),
    .X(_2012_));
 sg13g2_buf_2 _2396_ (.A(_2012_),
    .X(_2013_));
 sg13g2_buf_8 _2397_ (.A(net78),
    .X(_2014_));
 sg13g2_nand2_1 _2398_ (.Y(_2015_),
    .A(net108),
    .B(_1908_));
 sg13g2_o21ai_1 _2399_ (.B1(_1992_),
    .Y(_2016_),
    .A1(net89),
    .A2(_2015_));
 sg13g2_buf_1 _2400_ (.A(_2016_),
    .X(_2017_));
 sg13g2_buf_2 _2401_ (.A(net74),
    .X(_2018_));
 sg13g2_mux4_1 _2402_ (.S0(net75),
    .A0(_0089_),
    .A1(_0088_),
    .A2(_0091_),
    .A3(_0090_),
    .S1(net68),
    .X(_2019_));
 sg13g2_mux4_1 _2403_ (.S0(net75),
    .A0(_0097_),
    .A1(_0096_),
    .A2(_0099_),
    .A3(_0098_),
    .S1(net68),
    .X(_2020_));
 sg13g2_mux4_1 _2404_ (.S0(net75),
    .A0(_0093_),
    .A1(_0092_),
    .A2(_0095_),
    .A3(_0094_),
    .S1(net74),
    .X(_2021_));
 sg13g2_mux4_1 _2405_ (.S0(net75),
    .A0(_0101_),
    .A1(_0100_),
    .A2(_0103_),
    .A3(_0102_),
    .S1(net74),
    .X(_2022_));
 sg13g2_nor3_1 _2406_ (.A(net131),
    .B(net139),
    .C(_1784_),
    .Y(_2023_));
 sg13g2_xnor2_1 _2407_ (.Y(_2024_),
    .A(_1793_),
    .B(_2023_));
 sg13g2_mux2_1 _2408_ (.A0(_1946_),
    .A1(_2024_),
    .S(net100),
    .X(_2025_));
 sg13g2_buf_2 _2409_ (.A(_2025_),
    .X(_2026_));
 sg13g2_buf_2 _2410_ (.A(_2026_),
    .X(_2027_));
 sg13g2_xnor2_1 _2411_ (.Y(_2028_),
    .A(_1794_),
    .B(_1940_));
 sg13g2_mux2_1 _2412_ (.A0(_1944_),
    .A1(_2028_),
    .S(net100),
    .X(_2029_));
 sg13g2_buf_2 _2413_ (.A(_2029_),
    .X(_2030_));
 sg13g2_buf_8 _2414_ (.A(_2030_),
    .X(_2031_));
 sg13g2_buf_2 _2415_ (.A(_2031_),
    .X(_2032_));
 sg13g2_mux4_1 _2416_ (.S0(net73),
    .A0(_2019_),
    .A1(_2020_),
    .A2(_2021_),
    .A3(_2022_),
    .S1(net67),
    .X(_2033_));
 sg13g2_inv_1 _2417_ (.Y(_2034_),
    .A(_2033_));
 sg13g2_nor2_1 _2418_ (.A(_1824_),
    .B(_2034_),
    .Y(_2035_));
 sg13g2_buf_2 _2419_ (.A(net75),
    .X(_2036_));
 sg13g2_mux4_1 _2420_ (.S0(net66),
    .A0(_0105_),
    .A1(_0104_),
    .A2(_0107_),
    .A3(_0106_),
    .S1(net68),
    .X(_2037_));
 sg13g2_mux4_1 _2421_ (.S0(net66),
    .A0(_0113_),
    .A1(_0112_),
    .A2(_0115_),
    .A3(_0114_),
    .S1(net68),
    .X(_2038_));
 sg13g2_mux4_1 _2422_ (.S0(net75),
    .A0(_0109_),
    .A1(_0108_),
    .A2(_0111_),
    .A3(_0110_),
    .S1(net68),
    .X(_2039_));
 sg13g2_mux4_1 _2423_ (.S0(net75),
    .A0(_0117_),
    .A1(_0116_),
    .A2(_0119_),
    .A3(_0118_),
    .S1(net68),
    .X(_2040_));
 sg13g2_mux4_1 _2424_ (.S0(net73),
    .A0(_2037_),
    .A1(_2038_),
    .A2(_2039_),
    .A3(_2040_),
    .S1(net67),
    .X(_2041_));
 sg13g2_mux4_1 _2425_ (.S0(net78),
    .A0(_0073_),
    .A1(_0072_),
    .A2(_0075_),
    .A3(_0074_),
    .S1(net74),
    .X(_2042_));
 sg13g2_mux4_1 _2426_ (.S0(net78),
    .A0(_0081_),
    .A1(_0080_),
    .A2(_0083_),
    .A3(_0082_),
    .S1(net74),
    .X(_0430_));
 sg13g2_mux4_1 _2427_ (.S0(net78),
    .A0(_0077_),
    .A1(_0076_),
    .A2(_0079_),
    .A3(_0078_),
    .S1(net74),
    .X(_0431_));
 sg13g2_mux4_1 _2428_ (.S0(net78),
    .A0(_0085_),
    .A1(_0084_),
    .A2(_0087_),
    .A3(_0086_),
    .S1(net74),
    .X(_0432_));
 sg13g2_mux4_1 _2429_ (.S0(net73),
    .A0(_2042_),
    .A1(_0430_),
    .A2(_0431_),
    .A3(_0432_),
    .S1(_2032_),
    .X(_0433_));
 sg13g2_buf_2 _2430_ (.A(_0433_),
    .X(_0434_));
 sg13g2_nand2b_1 _2431_ (.Y(_0435_),
    .B(_0434_),
    .A_N(_1826_));
 sg13g2_nand2b_1 _2432_ (.Y(_0436_),
    .B(_1826_),
    .A_N(_0434_));
 sg13g2_mux4_1 _2433_ (.S0(net78),
    .A0(_0057_),
    .A1(_0056_),
    .A2(_0061_),
    .A3(_0060_),
    .S1(net72),
    .X(_0437_));
 sg13g2_mux4_1 _2434_ (.S0(_2013_),
    .A0(_0059_),
    .A1(_0058_),
    .A2(_0063_),
    .A3(_0062_),
    .S1(net72),
    .X(_0438_));
 sg13g2_mux4_1 _2435_ (.S0(net78),
    .A0(_0065_),
    .A1(_0064_),
    .A2(_0069_),
    .A3(_0068_),
    .S1(net72),
    .X(_0439_));
 sg13g2_mux4_1 _2436_ (.S0(net78),
    .A0(_0067_),
    .A1(_0066_),
    .A2(_0071_),
    .A3(_0070_),
    .S1(net72),
    .X(_0440_));
 sg13g2_mux4_1 _2437_ (.S0(net74),
    .A0(_0437_),
    .A1(_0438_),
    .A2(_0439_),
    .A3(_0440_),
    .S1(net73),
    .X(_0441_));
 sg13g2_buf_2 _2438_ (.A(_0441_),
    .X(_0442_));
 sg13g2_and2_1 _2439_ (.A(_1828_),
    .B(_0442_),
    .X(_0443_));
 sg13g2_nand2_1 _2440_ (.Y(_0444_),
    .A(_0436_),
    .B(_0443_));
 sg13g2_a22oi_1 _2441_ (.Y(_0445_),
    .B1(_0435_),
    .B2(_0444_),
    .A2(_2034_),
    .A1(_1824_));
 sg13g2_or3_1 _2442_ (.A(_2035_),
    .B(_2041_),
    .C(_0445_),
    .X(_0446_));
 sg13g2_buf_1 _2443_ (.A(_0446_),
    .X(_0447_));
 sg13g2_and2_1 _2444_ (.A(_2012_),
    .B(_2017_),
    .X(_0448_));
 sg13g2_mux4_1 _2445_ (.S0(net72),
    .A0(_0026_),
    .A1(_0030_),
    .A2(_0034_),
    .A3(_0038_),
    .S1(_2027_),
    .X(_0449_));
 sg13g2_mux4_1 _2446_ (.S0(net72),
    .A0(_0027_),
    .A1(_0031_),
    .A2(_0035_),
    .A3(_0039_),
    .S1(net73),
    .X(_0450_));
 sg13g2_buf_8 _2447_ (.A(_1935_),
    .X(_0451_));
 sg13g2_and2_1 _2448_ (.A(net77),
    .B(_2017_),
    .X(_0452_));
 sg13g2_a22oi_1 _2449_ (.Y(_0453_),
    .B1(_0450_),
    .B2(_0452_),
    .A2(_0449_),
    .A1(_0448_));
 sg13g2_nand2_1 _2450_ (.Y(_0454_),
    .A(net138),
    .B(_2015_));
 sg13g2_buf_1 _2451_ (.A(_1925_),
    .X(_0455_));
 sg13g2_nand3_1 _2452_ (.B(net126),
    .C(net90),
    .A(net124),
    .Y(_0456_));
 sg13g2_o21ai_1 _2453_ (.B1(_0456_),
    .Y(_0457_),
    .A1(net90),
    .A2(_0454_));
 sg13g2_mux4_1 _2454_ (.S0(_2012_),
    .A0(_0025_),
    .A1(_0024_),
    .A2(_0029_),
    .A3(_0028_),
    .S1(net72),
    .X(_0458_));
 sg13g2_mux4_1 _2455_ (.S0(_2012_),
    .A0(_0033_),
    .A1(_0032_),
    .A2(_0037_),
    .A3(_0036_),
    .S1(net72),
    .X(_0459_));
 sg13g2_nand3b_1 _2456_ (.B(net100),
    .C(_2015_),
    .Y(_0460_),
    .A_N(net138));
 sg13g2_nand3_1 _2457_ (.B(_1946_),
    .C(net90),
    .A(net124),
    .Y(_0461_));
 sg13g2_nand2_1 _2458_ (.Y(_0462_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_a22oi_1 _2459_ (.Y(_0463_),
    .B1(_0459_),
    .B2(_0462_),
    .A2(_0458_),
    .A1(_0457_));
 sg13g2_and2_1 _2460_ (.A(_0453_),
    .B(_0463_),
    .X(_0464_));
 sg13g2_buf_2 _2461_ (.A(_0464_),
    .X(_0465_));
 sg13g2_and2_1 _2462_ (.A(_1832_),
    .B(_0465_),
    .X(_0466_));
 sg13g2_buf_1 _2463_ (.A(_0466_),
    .X(_0467_));
 sg13g2_inv_1 _2464_ (.Y(_0468_),
    .A(_1829_));
 sg13g2_nor2_1 _2465_ (.A(_1832_),
    .B(_0465_),
    .Y(_0469_));
 sg13g2_nor2_1 _2466_ (.A(_0468_),
    .B(_0469_),
    .Y(_0470_));
 sg13g2_mux4_1 _2467_ (.S0(_2030_),
    .A0(_0010_),
    .A1(_0014_),
    .A2(_0018_),
    .A3(_0022_),
    .S1(_2026_),
    .X(_0471_));
 sg13g2_mux4_1 _2468_ (.S0(_2031_),
    .A0(_0011_),
    .A1(_0015_),
    .A2(_0019_),
    .A3(_0023_),
    .S1(_2026_),
    .X(_0472_));
 sg13g2_a22oi_1 _2469_ (.Y(_0473_),
    .B1(_0452_),
    .B2(_0472_),
    .A2(_0471_),
    .A1(_0448_));
 sg13g2_buf_1 _2470_ (.A(_0473_),
    .X(_0474_));
 sg13g2_mux4_1 _2471_ (.S0(_2012_),
    .A0(_0009_),
    .A1(_0008_),
    .A2(_0013_),
    .A3(_0012_),
    .S1(_2030_),
    .X(_0475_));
 sg13g2_buf_1 _2472_ (.A(_1944_),
    .X(_0476_));
 sg13g2_nor2_1 _2473_ (.A(_1928_),
    .B(net134),
    .Y(_0477_));
 sg13g2_xor2_1 _2474_ (.B(_1794_),
    .A(net139),
    .X(_0478_));
 sg13g2_nor4_1 _2475_ (.A(net131),
    .B(net129),
    .C(net118),
    .D(_0478_),
    .Y(_0479_));
 sg13g2_a21o_1 _2476_ (.A2(_0477_),
    .A1(net90),
    .B1(_0479_),
    .X(_0480_));
 sg13g2_inv_1 _2477_ (.Y(_0481_),
    .A(_0017_));
 sg13g2_a22oi_1 _2478_ (.Y(_0482_),
    .B1(_0480_),
    .B2(_0481_),
    .A2(_0461_),
    .A1(_0460_));
 sg13g2_a21o_1 _2479_ (.A2(_1933_),
    .A1(_1930_),
    .B1(_0016_),
    .X(_0483_));
 sg13g2_buf_1 _2480_ (.A(net136),
    .X(_0484_));
 sg13g2_nor2b_1 _2481_ (.A(_0484_),
    .B_N(_0020_),
    .Y(_0485_));
 sg13g2_o21ai_1 _2482_ (.B1(_0485_),
    .Y(_0486_),
    .A1(_1903_),
    .A2(net118));
 sg13g2_and2_1 _2483_ (.A(net123),
    .B(_0021_),
    .X(_0487_));
 sg13g2_o21ai_1 _2484_ (.B1(_0487_),
    .Y(_0488_),
    .A1(net129),
    .A2(net118));
 sg13g2_nand2_1 _2485_ (.Y(_0489_),
    .A(net131),
    .B(_0020_));
 sg13g2_or3_1 _2486_ (.A(net129),
    .B(_1806_),
    .C(_0489_),
    .X(_0490_));
 sg13g2_inv_1 _2487_ (.Y(_0491_),
    .A(_0021_));
 sg13g2_or4_1 _2488_ (.A(net131),
    .B(_0491_),
    .C(net129),
    .D(_1806_),
    .X(_0492_));
 sg13g2_nand4_1 _2489_ (.B(_0488_),
    .C(_0490_),
    .A(_0486_),
    .Y(_0493_),
    .D(_0492_));
 sg13g2_mux2_1 _2490_ (.A0(_0483_),
    .A1(_0493_),
    .S(_2030_),
    .X(_0494_));
 sg13g2_a22oi_1 _2491_ (.Y(_0495_),
    .B1(_0482_),
    .B2(_0494_),
    .A2(_0475_),
    .A1(_0457_));
 sg13g2_nand2_1 _2492_ (.Y(_0496_),
    .A(_0474_),
    .B(_0495_));
 sg13g2_and2_1 _2493_ (.A(\madd.delta[2] ),
    .B(_0495_),
    .X(_0497_));
 sg13g2_nand2_1 _2494_ (.Y(_0498_),
    .A(_0474_),
    .B(_0497_));
 sg13g2_inv_1 _2495_ (.Y(_0499_),
    .A(_0152_));
 sg13g2_and4_1 _2496_ (.A(_0499_),
    .B(_1952_),
    .C(_1968_),
    .D(_2007_),
    .X(_0500_));
 sg13g2_buf_1 _2497_ (.A(_0500_),
    .X(_0501_));
 sg13g2_o21ai_1 _2498_ (.B1(net108),
    .Y(_0502_),
    .A1(_0180_),
    .A2(net116));
 sg13g2_a21oi_1 _2499_ (.A1(net123),
    .A2(_0180_),
    .Y(_0503_),
    .B1(net125));
 sg13g2_mux2_1 _2500_ (.A0(_0502_),
    .A1(_0503_),
    .S(net89),
    .X(_0504_));
 sg13g2_o21ai_1 _2501_ (.B1(_1923_),
    .Y(_0505_),
    .A1(_0182_),
    .A2(net107));
 sg13g2_a21oi_1 _2502_ (.A1(net123),
    .A2(_0182_),
    .Y(_0506_),
    .B1(_1925_));
 sg13g2_mux2_1 _2503_ (.A0(_0505_),
    .A1(_0506_),
    .S(net89),
    .X(_0507_));
 sg13g2_o21ai_1 _2504_ (.B1(net77),
    .Y(_0508_),
    .A1(_0504_),
    .A2(_0507_));
 sg13g2_nand2b_1 _2505_ (.Y(_0509_),
    .B(_0507_),
    .A_N(_0181_));
 sg13g2_inv_1 _2506_ (.Y(_0510_),
    .A(_0179_));
 sg13g2_a221oi_1 _2507_ (.B2(_0510_),
    .C1(_2005_),
    .B1(_0504_),
    .A1(net100),
    .Y(_0511_),
    .A2(_1998_));
 sg13g2_nand3_1 _2508_ (.B(_0509_),
    .C(_0511_),
    .A(_0508_),
    .Y(_0512_));
 sg13g2_o21ai_1 _2509_ (.B1(_1910_),
    .Y(_0513_),
    .A1(_0172_),
    .A2(net116));
 sg13g2_a21oi_1 _2510_ (.A1(net128),
    .A2(_0172_),
    .Y(_0514_),
    .B1(net125));
 sg13g2_mux2_1 _2511_ (.A0(_0513_),
    .A1(_0514_),
    .S(net89),
    .X(_0515_));
 sg13g2_o21ai_1 _2512_ (.B1(_1923_),
    .Y(_0516_),
    .A1(_0174_),
    .A2(net107));
 sg13g2_a21oi_1 _2513_ (.A1(_0484_),
    .A2(_0174_),
    .Y(_0517_),
    .B1(_1925_));
 sg13g2_mux2_1 _2514_ (.A0(_0516_),
    .A1(_0517_),
    .S(net89),
    .X(_0518_));
 sg13g2_o21ai_1 _2515_ (.B1(net77),
    .Y(_0519_),
    .A1(_0515_),
    .A2(_0518_));
 sg13g2_nand2b_1 _2516_ (.Y(_0520_),
    .B(_0518_),
    .A_N(_0173_));
 sg13g2_nand2b_1 _2517_ (.Y(_0521_),
    .B(_0515_),
    .A_N(_0171_));
 sg13g2_nand4_1 _2518_ (.B(_0519_),
    .C(_0520_),
    .A(_1966_),
    .Y(_0522_),
    .D(_0521_));
 sg13g2_inv_1 _2519_ (.Y(_0523_),
    .A(_0177_));
 sg13g2_o21ai_1 _2520_ (.B1(_1923_),
    .Y(_0524_),
    .A1(_0178_),
    .A2(net107));
 sg13g2_a21oi_1 _2521_ (.A1(net123),
    .A2(_0178_),
    .Y(_0525_),
    .B1(_0455_));
 sg13g2_mux2_1 _2522_ (.A0(_0524_),
    .A1(_0525_),
    .S(net90),
    .X(_0526_));
 sg13g2_o21ai_1 _2523_ (.B1(_0526_),
    .Y(_0527_),
    .A1(_0523_),
    .A2(net77));
 sg13g2_inv_1 _2524_ (.Y(_0528_),
    .A(_0175_));
 sg13g2_o21ai_1 _2525_ (.B1(net108),
    .Y(_0529_),
    .A1(_0176_),
    .A2(net116));
 sg13g2_a21oi_1 _2526_ (.A1(net123),
    .A2(_0176_),
    .Y(_0530_),
    .B1(net125));
 sg13g2_mux2_1 _2527_ (.A0(_0529_),
    .A1(_0530_),
    .S(net89),
    .X(_0531_));
 sg13g2_o21ai_1 _2528_ (.B1(_0531_),
    .Y(_0532_),
    .A1(_0528_),
    .A2(net77));
 sg13g2_nand3_1 _2529_ (.B(_0527_),
    .C(_0532_),
    .A(_1976_),
    .Y(_0533_));
 sg13g2_o21ai_1 _2530_ (.B1(_1923_),
    .Y(_0534_),
    .A1(_0186_),
    .A2(net107));
 sg13g2_a21oi_1 _2531_ (.A1(net128),
    .A2(_0186_),
    .Y(_0535_),
    .B1(_1925_));
 sg13g2_mux2_1 _2532_ (.A0(_0534_),
    .A1(_0535_),
    .S(net101),
    .X(_0536_));
 sg13g2_o21ai_1 _2533_ (.B1(net108),
    .Y(_0537_),
    .A1(_0184_),
    .A2(net116));
 sg13g2_a21oi_1 _2534_ (.A1(net128),
    .A2(_0184_),
    .Y(_0538_),
    .B1(net135));
 sg13g2_mux2_1 _2535_ (.A0(_0537_),
    .A1(_0538_),
    .S(net89),
    .X(_0539_));
 sg13g2_o21ai_1 _2536_ (.B1(_0451_),
    .Y(_0540_),
    .A1(_0536_),
    .A2(_0539_));
 sg13g2_nand2b_1 _2537_ (.Y(_0541_),
    .B(_0539_),
    .A_N(_0183_));
 sg13g2_nand2b_1 _2538_ (.Y(_0542_),
    .B(_0536_),
    .A_N(_0185_));
 sg13g2_nand4_1 _2539_ (.B(_0540_),
    .C(_0541_),
    .A(_1950_),
    .Y(_0543_),
    .D(_0542_));
 sg13g2_and4_1 _2540_ (.A(_0512_),
    .B(_0522_),
    .C(_0533_),
    .D(_0543_),
    .X(_0544_));
 sg13g2_buf_8 _2541_ (.A(_0544_),
    .X(_0545_));
 sg13g2_nor2_1 _2542_ (.A(_0501_),
    .B(_0545_),
    .Y(_0546_));
 sg13g2_a221oi_1 _2543_ (.B2(_0501_),
    .C1(_1834_),
    .B1(_0545_),
    .A1(_0474_),
    .Y(_0547_),
    .A2(_0497_));
 sg13g2_a221oi_1 _2544_ (.B2(_0546_),
    .C1(_0547_),
    .B1(_0498_),
    .A1(_1841_),
    .Y(_0548_),
    .A2(_0496_));
 sg13g2_buf_1 _2545_ (.A(_0548_),
    .X(_0549_));
 sg13g2_mux4_1 _2546_ (.S0(net75),
    .A0(_0041_),
    .A1(_0040_),
    .A2(_0045_),
    .A3(_0044_),
    .S1(net67),
    .X(_0550_));
 sg13g2_mux4_1 _2547_ (.S0(_2014_),
    .A0(_0043_),
    .A1(_0042_),
    .A2(_0047_),
    .A3(_0046_),
    .S1(net67),
    .X(_0551_));
 sg13g2_mux4_1 _2548_ (.S0(_2013_),
    .A0(_0049_),
    .A1(_0048_),
    .A2(_0053_),
    .A3(_0052_),
    .S1(net67),
    .X(_0552_));
 sg13g2_mux4_1 _2549_ (.S0(_2014_),
    .A0(_0051_),
    .A1(_0050_),
    .A2(_0055_),
    .A3(_0054_),
    .S1(_2032_),
    .X(_0553_));
 sg13g2_mux4_1 _2550_ (.S0(_2018_),
    .A0(_0550_),
    .A1(_0551_),
    .A2(_0552_),
    .A3(_0553_),
    .S1(net73),
    .X(_0554_));
 sg13g2_buf_1 _2551_ (.A(_0554_),
    .X(_0555_));
 sg13g2_nor2_1 _2552_ (.A(_0468_),
    .B(_0555_),
    .Y(_0556_));
 sg13g2_a221oi_1 _2553_ (.B2(_0549_),
    .C1(_0556_),
    .B1(_0470_),
    .A1(_1829_),
    .Y(_0557_),
    .A2(_0467_));
 sg13g2_buf_1 _2554_ (.A(_0557_),
    .X(_0558_));
 sg13g2_nor2_1 _2555_ (.A(_0555_),
    .B(_0469_),
    .Y(_0559_));
 sg13g2_o21ai_1 _2556_ (.B1(_0559_),
    .Y(_0560_),
    .A1(_0549_),
    .A2(_0467_));
 sg13g2_buf_2 _2557_ (.A(_0560_),
    .X(_0561_));
 sg13g2_nand2b_1 _2558_ (.Y(_0562_),
    .B(\madd.delta[5] ),
    .A_N(_0442_));
 sg13g2_nand2_1 _2559_ (.Y(_0563_),
    .A(_1824_),
    .B(_2034_));
 sg13g2_and3_1 _2560_ (.X(_0564_),
    .A(_0562_),
    .B(_0563_),
    .C(_0436_));
 sg13g2_nand3_1 _2561_ (.B(_0561_),
    .C(_0564_),
    .A(_0558_),
    .Y(_0565_));
 sg13g2_nand2b_1 _2562_ (.Y(_0566_),
    .B(_0565_),
    .A_N(_0447_));
 sg13g2_buf_2 _2563_ (.A(net68),
    .X(_0567_));
 sg13g2_mux4_1 _2564_ (.S0(net66),
    .A0(_0137_),
    .A1(_0136_),
    .A2(_0139_),
    .A3(_0138_),
    .S1(net63),
    .X(_0568_));
 sg13g2_mux4_1 _2565_ (.S0(_2036_),
    .A0(_0145_),
    .A1(_0144_),
    .A2(_0147_),
    .A3(_0146_),
    .S1(net63),
    .X(_0569_));
 sg13g2_mux4_1 _2566_ (.S0(net66),
    .A0(_0141_),
    .A1(_0140_),
    .A2(_0143_),
    .A3(_0142_),
    .S1(net68),
    .X(_0570_));
 sg13g2_mux4_1 _2567_ (.S0(net66),
    .A0(_0149_),
    .A1(_0148_),
    .A2(_0151_),
    .A3(_0150_),
    .S1(_2018_),
    .X(_0571_));
 sg13g2_mux4_1 _2568_ (.S0(net73),
    .A0(_0568_),
    .A1(_0569_),
    .A2(_0570_),
    .A3(_0571_),
    .S1(net67),
    .X(_0572_));
 sg13g2_buf_1 _2569_ (.A(_0572_),
    .X(_0573_));
 sg13g2_mux4_1 _2570_ (.S0(_2036_),
    .A0(_0121_),
    .A1(_0120_),
    .A2(_0123_),
    .A3(_0122_),
    .S1(_0567_),
    .X(_0574_));
 sg13g2_mux4_1 _2571_ (.S0(net66),
    .A0(_0129_),
    .A1(_0128_),
    .A2(_0131_),
    .A3(_0130_),
    .S1(net63),
    .X(_0575_));
 sg13g2_mux4_1 _2572_ (.S0(net66),
    .A0(_0125_),
    .A1(_0124_),
    .A2(_0127_),
    .A3(_0126_),
    .S1(net63),
    .X(_0576_));
 sg13g2_mux4_1 _2573_ (.S0(net66),
    .A0(_0133_),
    .A1(_0132_),
    .A2(_0135_),
    .A3(_0134_),
    .S1(net63),
    .X(_0577_));
 sg13g2_mux4_1 _2574_ (.S0(net73),
    .A0(_0574_),
    .A1(_0575_),
    .A2(_0576_),
    .A3(_0577_),
    .S1(net67),
    .X(_0578_));
 sg13g2_inv_2 _2575_ (.Y(_0579_),
    .A(_0578_));
 sg13g2_nand3_1 _2576_ (.B(net47),
    .C(_0579_),
    .A(_1807_),
    .Y(_0580_));
 sg13g2_nand3_1 _2577_ (.B(_1807_),
    .C(net47),
    .A(_1820_),
    .Y(_0581_));
 sg13g2_or2_1 _2578_ (.X(_0582_),
    .B(_0445_),
    .A(_2035_));
 sg13g2_inv_1 _2579_ (.Y(_0583_),
    .A(_0582_));
 sg13g2_inv_1 _2580_ (.Y(_0584_),
    .A(_2041_));
 sg13g2_a21oi_1 _2581_ (.A1(_0565_),
    .A2(_0583_),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a221oi_1 _2582_ (.B2(_0581_),
    .C1(_0585_),
    .B1(_0580_),
    .A1(_1894_),
    .Y(_0586_),
    .A2(_0566_));
 sg13g2_and3_1 _2583_ (.X(_0587_),
    .A(_0558_),
    .B(_0561_),
    .C(_0564_));
 sg13g2_buf_8 _2584_ (.A(_0587_),
    .X(_0588_));
 sg13g2_o21ai_1 _2585_ (.B1(_1894_),
    .Y(_0589_),
    .A1(_0588_),
    .A2(_0447_));
 sg13g2_o21ai_1 _2586_ (.B1(_2041_),
    .Y(_0590_),
    .A1(_0588_),
    .A2(_0582_));
 sg13g2_buf_1 _2587_ (.A(_0590_),
    .X(_0591_));
 sg13g2_nor2_1 _2588_ (.A(net47),
    .B(_0579_),
    .Y(_0592_));
 sg13g2_nand2_1 _2589_ (.Y(_0593_),
    .A(net102),
    .B(_0592_));
 sg13g2_or3_1 _2590_ (.A(_1820_),
    .B(_1817_),
    .C(net47),
    .X(_0594_));
 sg13g2_a22oi_1 _2591_ (.Y(_0595_),
    .B1(_0593_),
    .B2(_0594_),
    .A2(_0591_),
    .A1(_0589_));
 sg13g2_nand4_1 _2592_ (.B(net102),
    .C(net47),
    .A(_1820_),
    .Y(_0596_),
    .D(_0579_));
 sg13g2_nand3_1 _2593_ (.B(net102),
    .C(_0592_),
    .A(_1821_),
    .Y(_0597_));
 sg13g2_nand2_1 _2594_ (.Y(_0598_),
    .A(_0596_),
    .B(_0597_));
 sg13g2_nor3_1 _2595_ (.A(_0586_),
    .B(_0595_),
    .C(_0598_),
    .Y(_0599_));
 sg13g2_xor2_1 _2596_ (.B(_0599_),
    .A(_1819_),
    .X(_0600_));
 sg13g2_nor2_1 _2597_ (.A(net109),
    .B(_0600_),
    .Y(_0200_));
 sg13g2_and2_1 _2598_ (.A(net140),
    .B(\madd.delta[11] ),
    .X(_0601_));
 sg13g2_nor2_1 _2599_ (.A(_1758_),
    .B(\madd.delta[11] ),
    .Y(_0602_));
 sg13g2_mux4_1 _2600_ (.S0(net77),
    .A0(\madd.mem[0][11] ),
    .A1(\madd.mem[1][11] ),
    .A2(\madd.mem[2][11] ),
    .A3(\madd.mem[3][11] ),
    .S1(net63),
    .X(_0603_));
 sg13g2_mux4_1 _2601_ (.S0(_0451_),
    .A0(\madd.mem[8][11] ),
    .A1(\madd.mem[9][11] ),
    .A2(\madd.mem[10][11] ),
    .A3(\madd.mem[11][11] ),
    .S1(_0567_),
    .X(_0604_));
 sg13g2_mux4_1 _2602_ (.S0(net77),
    .A0(\madd.mem[4][11] ),
    .A1(\madd.mem[5][11] ),
    .A2(\madd.mem[6][11] ),
    .A3(\madd.mem[7][11] ),
    .S1(net63),
    .X(_0605_));
 sg13g2_mux4_1 _2603_ (.S0(net77),
    .A0(\madd.mem[12][11] ),
    .A1(\madd.mem[13][11] ),
    .A2(\madd.mem[14][11] ),
    .A3(\madd.mem[15][11] ),
    .S1(net63),
    .X(_0606_));
 sg13g2_mux4_1 _2604_ (.S0(_2027_),
    .A0(_0603_),
    .A1(_0604_),
    .A2(_0605_),
    .A3(_0606_),
    .S1(net67),
    .X(_0607_));
 sg13g2_and2_1 _2605_ (.A(net102),
    .B(_0607_),
    .X(_0608_));
 sg13g2_nor2_1 _2606_ (.A(_1817_),
    .B(_0607_),
    .Y(_0609_));
 sg13g2_nor2b_1 _2607_ (.A(_1819_),
    .B_N(net47),
    .Y(_0610_));
 sg13g2_nor2b_1 _2608_ (.A(_0573_),
    .B_N(_1819_),
    .Y(_0611_));
 sg13g2_nor2_1 _2609_ (.A(_0579_),
    .B(_0611_),
    .Y(_0612_));
 sg13g2_o21ai_1 _2610_ (.B1(_0612_),
    .Y(_0613_),
    .A1(_0588_),
    .A2(_0447_));
 sg13g2_nor2_1 _2611_ (.A(_1820_),
    .B(_0611_),
    .Y(_0614_));
 sg13g2_o21ai_1 _2612_ (.B1(_0614_),
    .Y(_0615_),
    .A1(_0588_),
    .A2(_0447_));
 sg13g2_nor4_1 _2613_ (.A(_1894_),
    .B(_0588_),
    .C(_2035_),
    .D(_0445_),
    .Y(_0616_));
 sg13g2_a221oi_1 _2614_ (.B2(_0615_),
    .C1(_0616_),
    .B1(_0613_),
    .A1(_1823_),
    .Y(_0617_),
    .A2(_0584_));
 sg13g2_nor3_1 _2615_ (.A(_1820_),
    .B(_0579_),
    .C(_0611_),
    .Y(_0618_));
 sg13g2_nor3_1 _2616_ (.A(_0610_),
    .B(_0617_),
    .C(_0618_),
    .Y(_0619_));
 sg13g2_mux2_1 _2617_ (.A0(_0608_),
    .A1(_0609_),
    .S(_0619_),
    .X(_0620_));
 sg13g2_mux2_1 _2618_ (.A0(_0601_),
    .A1(_0602_),
    .S(_0620_),
    .X(_0201_));
 sg13g2_buf_1 _2619_ (.A(net117),
    .X(_0621_));
 sg13g2_xnor2_1 _2620_ (.Y(_0622_),
    .A(_0501_),
    .B(_0545_));
 sg13g2_nor2_1 _2621_ (.A(_1893_),
    .B(_0622_),
    .Y(_0623_));
 sg13g2_xnor2_1 _2622_ (.Y(_0624_),
    .A(_1834_),
    .B(_0623_));
 sg13g2_nor2_1 _2623_ (.A(net106),
    .B(_0624_),
    .Y(_0202_));
 sg13g2_a21oi_1 _2624_ (.A1(_0501_),
    .A2(_0545_),
    .Y(_0625_),
    .B1(_1834_));
 sg13g2_nor2_1 _2625_ (.A(_0546_),
    .B(_0625_),
    .Y(_0626_));
 sg13g2_xnor2_1 _2626_ (.Y(_0627_),
    .A(_0496_),
    .B(_0626_));
 sg13g2_nand2_1 _2627_ (.Y(_0628_),
    .A(_1809_),
    .B(_0627_));
 sg13g2_xnor2_1 _2628_ (.Y(_0629_),
    .A(_1841_),
    .B(_0628_));
 sg13g2_nor2_1 _2629_ (.A(_0621_),
    .B(_0629_),
    .Y(_0203_));
 sg13g2_xnor2_1 _2630_ (.Y(_0630_),
    .A(_0549_),
    .B(_0465_));
 sg13g2_nor2_1 _2631_ (.A(_1893_),
    .B(_0630_),
    .Y(_0631_));
 sg13g2_xnor2_1 _2632_ (.Y(_0632_),
    .A(_1832_),
    .B(_0631_));
 sg13g2_nor2_1 _2633_ (.A(net106),
    .B(_0632_),
    .Y(_0204_));
 sg13g2_nor2_1 _2634_ (.A(_0549_),
    .B(_0467_),
    .Y(_0633_));
 sg13g2_o21ai_1 _2635_ (.B1(_0555_),
    .Y(_0634_),
    .A1(_0633_),
    .A2(_0469_));
 sg13g2_and3_1 _2636_ (.X(_0635_),
    .A(net102),
    .B(_0561_),
    .C(_0634_));
 sg13g2_xnor2_1 _2637_ (.Y(_0636_),
    .A(_1829_),
    .B(_0635_));
 sg13g2_nor2_1 _2638_ (.A(net106),
    .B(_0636_),
    .Y(_0205_));
 sg13g2_nand2_1 _2639_ (.Y(_0637_),
    .A(_0558_),
    .B(_0561_));
 sg13g2_xnor2_1 _2640_ (.Y(_0638_),
    .A(_0637_),
    .B(_0442_));
 sg13g2_nand2_1 _2641_ (.Y(_0639_),
    .A(net93),
    .B(_0638_));
 sg13g2_xnor2_1 _2642_ (.Y(_0640_),
    .A(_1828_),
    .B(_0639_));
 sg13g2_nor2_1 _2643_ (.A(_0621_),
    .B(_0640_),
    .Y(_0206_));
 sg13g2_a21o_1 _2644_ (.A2(_0561_),
    .A1(_0558_),
    .B1(_0443_),
    .X(_0641_));
 sg13g2_nand2_1 _2645_ (.Y(_0642_),
    .A(_0562_),
    .B(_0641_));
 sg13g2_xor2_1 _2646_ (.B(_0642_),
    .A(_0434_),
    .X(_0643_));
 sg13g2_nor2_1 _2647_ (.A(net91),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_xnor2_1 _2648_ (.Y(_0645_),
    .A(_1826_),
    .B(_0644_));
 sg13g2_nor2_1 _2649_ (.A(net106),
    .B(_0645_),
    .Y(_0207_));
 sg13g2_a21oi_1 _2650_ (.A1(_0562_),
    .A2(_0641_),
    .Y(_0646_),
    .B1(_0434_));
 sg13g2_nand3_1 _2651_ (.B(_0434_),
    .C(_0641_),
    .A(_0562_),
    .Y(_0647_));
 sg13g2_o21ai_1 _2652_ (.B1(_0647_),
    .Y(_0648_),
    .A1(_1826_),
    .A2(_0646_));
 sg13g2_xnor2_1 _2653_ (.Y(_0649_),
    .A(_2033_),
    .B(_0648_));
 sg13g2_o21ai_1 _2654_ (.B1(_1824_),
    .Y(_0650_),
    .A1(net92),
    .A2(_0649_));
 sg13g2_or3_1 _2655_ (.A(_1824_),
    .B(net92),
    .C(_0649_),
    .X(_0651_));
 sg13g2_a21oi_1 _2656_ (.A1(_0650_),
    .A2(_0651_),
    .Y(_0208_),
    .B1(net117));
 sg13g2_nand3_1 _2657_ (.B(_0566_),
    .C(_0591_),
    .A(net93),
    .Y(_0652_));
 sg13g2_xnor2_1 _2658_ (.Y(_0653_),
    .A(_1894_),
    .B(_0652_));
 sg13g2_nor2_1 _2659_ (.A(net106),
    .B(_0653_),
    .Y(_0209_));
 sg13g2_a21oi_1 _2660_ (.A1(_0589_),
    .A2(_0591_),
    .Y(_0654_),
    .B1(_0579_));
 sg13g2_and3_1 _2661_ (.X(_0655_),
    .A(_0589_),
    .B(_0591_),
    .C(_0579_));
 sg13g2_nor3_1 _2662_ (.A(net91),
    .B(_0654_),
    .C(_0655_),
    .Y(_0656_));
 sg13g2_xnor2_1 _2663_ (.Y(_0657_),
    .A(_1820_),
    .B(_0656_));
 sg13g2_nor2_1 _2664_ (.A(net106),
    .B(_0657_),
    .Y(_0210_));
 sg13g2_mux2_1 _2665_ (.A0(\madd.i_e[0] ),
    .A1(_1767_),
    .S(_1755_),
    .X(_0658_));
 sg13g2_and2_1 _2666_ (.A(net130),
    .B(_0658_),
    .X(_0212_));
 sg13g2_nand2_1 _2667_ (.Y(_0659_),
    .A(_1928_),
    .B(_1925_));
 sg13g2_buf_1 _2668_ (.A(_0659_),
    .X(_0660_));
 sg13g2_nand3b_1 _2669_ (.B(_1754_),
    .C(_1756_),
    .Y(_0661_),
    .A_N(_1753_));
 sg13g2_buf_1 _2670_ (.A(_0661_),
    .X(_0662_));
 sg13g2_nand2b_1 _2671_ (.Y(_0663_),
    .B(_1763_),
    .A_N(_0662_));
 sg13g2_buf_1 _2672_ (.A(_0663_),
    .X(_0664_));
 sg13g2_nor2_1 _2673_ (.A(net114),
    .B(_0664_),
    .Y(_0665_));
 sg13g2_and2_1 _2674_ (.A(net127),
    .B(_0665_),
    .X(_0666_));
 sg13g2_buf_1 _2675_ (.A(_0666_),
    .X(_0667_));
 sg13g2_buf_1 _2676_ (.A(_0667_),
    .X(_0668_));
 sg13g2_inv_1 _2677_ (.Y(_0669_),
    .A(net1));
 sg13g2_nand2_1 _2678_ (.Y(_0670_),
    .A(_0669_),
    .B(_2008_));
 sg13g2_nand4_1 _2679_ (.B(_1952_),
    .C(_1968_),
    .A(net1),
    .Y(_0671_),
    .D(_2007_));
 sg13g2_nand2_1 _2680_ (.Y(_0672_),
    .A(_1767_),
    .B(net142));
 sg13g2_or2_1 _2681_ (.X(_0673_),
    .B(_0662_),
    .A(_0672_));
 sg13g2_buf_1 _2682_ (.A(_0673_),
    .X(_0674_));
 sg13g2_buf_1 _2683_ (.A(_0674_),
    .X(_0675_));
 sg13g2_a21o_1 _2684_ (.A2(_0671_),
    .A1(_0670_),
    .B1(net99),
    .X(_0676_));
 sg13g2_buf_2 _2685_ (.A(_0676_),
    .X(_0677_));
 sg13g2_buf_1 _2686_ (.A(_1757_),
    .X(_0678_));
 sg13g2_nor2_1 _2687_ (.A(_0672_),
    .B(_0662_),
    .Y(_0679_));
 sg13g2_buf_1 _2688_ (.A(_0679_),
    .X(_0680_));
 sg13g2_nand2_2 _2689_ (.Y(_0681_),
    .A(net127),
    .B(_0680_));
 sg13g2_buf_1 _2690_ (.A(net115),
    .X(_0682_));
 sg13g2_buf_2 _2691_ (.A(net105),
    .X(_0683_));
 sg13g2_buf_1 _2692_ (.A(net98),
    .X(_0684_));
 sg13g2_nand2_1 _2693_ (.Y(_0685_),
    .A(net88),
    .B(net124));
 sg13g2_nor2_1 _2694_ (.A(_0681_),
    .B(_0685_),
    .Y(_0686_));
 sg13g2_buf_2 _2695_ (.A(_0686_),
    .X(_0687_));
 sg13g2_nor3_1 _2696_ (.A(_0678_),
    .B(_0667_),
    .C(_0687_),
    .Y(_0688_));
 sg13g2_buf_1 _2697_ (.A(_0688_),
    .X(_0689_));
 sg13g2_buf_1 _2698_ (.A(_0680_),
    .X(_0690_));
 sg13g2_buf_1 _2699_ (.A(_1928_),
    .X(_0691_));
 sg13g2_buf_1 _2700_ (.A(_1991_),
    .X(_0692_));
 sg13g2_buf_1 _2701_ (.A(net113),
    .X(_0693_));
 sg13g2_buf_1 _2702_ (.A(net104),
    .X(_0694_));
 sg13g2_buf_1 _2703_ (.A(net96),
    .X(_0695_));
 sg13g2_buf_1 _2704_ (.A(net87),
    .X(_0696_));
 sg13g2_nor2_1 _2705_ (.A(_0691_),
    .B(net76),
    .Y(_0697_));
 sg13g2_nand3_1 _2706_ (.B(_0690_),
    .C(_0697_),
    .A(_1962_),
    .Y(_0698_));
 sg13g2_buf_2 _2707_ (.A(_0698_),
    .X(_0699_));
 sg13g2_mux4_1 _2708_ (.S0(net136),
    .A0(_0170_),
    .A1(_0167_),
    .A2(_0168_),
    .A3(_0169_),
    .S1(net141),
    .X(_0700_));
 sg13g2_mux4_1 _2709_ (.S0(_1912_),
    .A0(_0161_),
    .A1(_0158_),
    .A2(_0159_),
    .A3(_0160_),
    .S1(net141),
    .X(_0701_));
 sg13g2_mux2_1 _2710_ (.A0(_0700_),
    .A1(_0701_),
    .S(_1971_),
    .X(_0702_));
 sg13g2_nand3_1 _2711_ (.B(_0660_),
    .C(_0702_),
    .A(net134),
    .Y(_0703_));
 sg13g2_nor3_1 _2712_ (.A(_1912_),
    .B(net141),
    .C(_1944_),
    .Y(_0704_));
 sg13g2_mux2_1 _2713_ (.A0(_0700_),
    .A1(_0701_),
    .S(_1946_),
    .X(_0705_));
 sg13g2_nor2_1 _2714_ (.A(_1912_),
    .B(net141),
    .Y(_0706_));
 sg13g2_buf_8 _2715_ (.A(_0706_),
    .X(_0707_));
 sg13g2_xnor2_1 _2716_ (.Y(_0708_),
    .A(_1944_),
    .B(_0707_));
 sg13g2_mux4_1 _2717_ (.S0(net136),
    .A0(_0166_),
    .A1(_0163_),
    .A2(_0164_),
    .A3(_0165_),
    .S1(net135),
    .X(_0709_));
 sg13g2_mux4_1 _2718_ (.S0(_1913_),
    .A0(_0156_),
    .A1(_0153_),
    .A2(_0154_),
    .A3(_0155_),
    .S1(net135),
    .X(_0710_));
 sg13g2_mux2_1 _2719_ (.A0(_0709_),
    .A1(_0710_),
    .S(_1971_),
    .X(_0711_));
 sg13g2_a22oi_1 _2720_ (.Y(_0712_),
    .B1(_0708_),
    .B2(_0711_),
    .A2(_0705_),
    .A1(_0704_));
 sg13g2_nand2_1 _2721_ (.Y(_0713_),
    .A(_0703_),
    .B(_0712_));
 sg13g2_xnor2_1 _2722_ (.Y(_0714_),
    .A(_0669_),
    .B(_0713_));
 sg13g2_buf_2 _2723_ (.A(_0714_),
    .X(_0715_));
 sg13g2_buf_1 _2724_ (.A(_0715_),
    .X(_0716_));
 sg13g2_nor2_1 _2725_ (.A(_0699_),
    .B(net70),
    .Y(_0717_));
 sg13g2_a221oi_1 _2726_ (.B2(\madd.mem[0][0] ),
    .C1(_0717_),
    .B1(net60),
    .A1(net71),
    .Y(_0718_),
    .A2(_0677_));
 sg13g2_inv_1 _2727_ (.Y(_0213_),
    .A(_0718_));
 sg13g2_buf_1 _2728_ (.A(_0680_),
    .X(_0719_));
 sg13g2_buf_1 _2729_ (.A(net95),
    .X(_0720_));
 sg13g2_nand2_1 _2730_ (.Y(_0721_),
    .A(net71),
    .B(net86));
 sg13g2_inv_1 _2731_ (.Y(_0722_),
    .A(net3));
 sg13g2_nand3_1 _2732_ (.B(_0474_),
    .C(_0495_),
    .A(net2),
    .Y(_0723_));
 sg13g2_buf_1 _2733_ (.A(ui_in[1]),
    .X(_0724_));
 sg13g2_nand2_1 _2734_ (.Y(_0725_),
    .A(_0724_),
    .B(_0545_));
 sg13g2_inv_1 _2735_ (.Y(_0726_),
    .A(_0724_));
 sg13g2_nand4_1 _2736_ (.B(_0522_),
    .C(_0533_),
    .A(_0512_),
    .Y(_0727_),
    .D(_0543_));
 sg13g2_a21o_1 _2737_ (.A2(_0727_),
    .A1(_0726_),
    .B1(_0671_),
    .X(_0728_));
 sg13g2_nand3_1 _2738_ (.B(_0725_),
    .C(_0728_),
    .A(_0723_),
    .Y(_0729_));
 sg13g2_inv_1 _2739_ (.Y(_0730_),
    .A(net2));
 sg13g2_nand2_1 _2740_ (.Y(_0731_),
    .A(_0730_),
    .B(_0496_));
 sg13g2_nand3_1 _2741_ (.B(_0729_),
    .C(_0731_),
    .A(_0465_),
    .Y(_0732_));
 sg13g2_a21oi_1 _2742_ (.A1(_0729_),
    .A2(_0731_),
    .Y(_0733_),
    .B1(_0465_));
 sg13g2_a21oi_2 _2743_ (.B1(_0733_),
    .Y(_0734_),
    .A2(_0732_),
    .A1(_0722_));
 sg13g2_nor3_1 _2744_ (.A(_0555_),
    .B(_0442_),
    .C(_0434_),
    .Y(_0735_));
 sg13g2_nand4_1 _2745_ (.B(_0584_),
    .C(_0734_),
    .A(_2034_),
    .Y(_0736_),
    .D(_0735_));
 sg13g2_nor2_1 _2746_ (.A(_0578_),
    .B(_0736_),
    .Y(_0737_));
 sg13g2_xor2_1 _2747_ (.B(_0737_),
    .A(net47),
    .X(_0738_));
 sg13g2_buf_2 _2748_ (.A(_0738_),
    .X(_0739_));
 sg13g2_buf_8 _2749_ (.A(_0739_),
    .X(_0740_));
 sg13g2_mux4_1 _2750_ (.S0(net87),
    .A0(\madd.mem[7][10] ),
    .A1(\madd.mem[5][10] ),
    .A2(\madd.mem[4][10] ),
    .A3(\madd.mem[6][10] ),
    .S1(net88),
    .X(_0741_));
 sg13g2_mux4_1 _2751_ (.S0(net87),
    .A0(\madd.mem[15][10] ),
    .A1(\madd.mem[13][10] ),
    .A2(\madd.mem[12][10] ),
    .A3(\madd.mem[14][10] ),
    .S1(net88),
    .X(_0742_));
 sg13g2_xnor2_1 _2752_ (.Y(_0743_),
    .A(_1947_),
    .B(_0704_));
 sg13g2_buf_1 _2753_ (.A(_0743_),
    .X(_0744_));
 sg13g2_buf_1 _2754_ (.A(net112),
    .X(_0745_));
 sg13g2_mux2_1 _2755_ (.A0(_0741_),
    .A1(_0742_),
    .S(net103),
    .X(_0746_));
 sg13g2_nor2_1 _2756_ (.A(_0708_),
    .B(_0746_),
    .Y(_0747_));
 sg13g2_nor2_1 _2757_ (.A(net124),
    .B(\madd.mem[10][10] ),
    .Y(_0748_));
 sg13g2_nor2_1 _2758_ (.A(net76),
    .B(\madd.mem[8][10] ),
    .Y(_0749_));
 sg13g2_o21ai_1 _2759_ (.B1(_0477_),
    .Y(_0750_),
    .A1(_0748_),
    .A2(_0749_));
 sg13g2_nand2b_1 _2760_ (.Y(_0751_),
    .B(net134),
    .A_N(net113));
 sg13g2_nor2_1 _2761_ (.A(\madd.mem[11][10] ),
    .B(_0751_),
    .Y(_0752_));
 sg13g2_nand2b_1 _2762_ (.Y(_0753_),
    .B(net113),
    .A_N(_0476_));
 sg13g2_nor2_1 _2763_ (.A(\madd.mem[9][10] ),
    .B(_0753_),
    .Y(_0754_));
 sg13g2_o21ai_1 _2764_ (.B1(net121),
    .Y(_0755_),
    .A1(_0752_),
    .A2(_0754_));
 sg13g2_nand2_1 _2765_ (.Y(_0756_),
    .A(_0750_),
    .B(_0755_));
 sg13g2_xnor2_1 _2766_ (.Y(_0757_),
    .A(_1945_),
    .B(_0707_));
 sg13g2_buf_2 _2767_ (.A(_0757_),
    .X(_0758_));
 sg13g2_mux4_1 _2768_ (.S0(net76),
    .A0(\madd.mem[3][10] ),
    .A1(\madd.mem[1][10] ),
    .A2(\madd.mem[0][10] ),
    .A3(\madd.mem[2][10] ),
    .S1(net88),
    .X(_0759_));
 sg13g2_nor3_1 _2769_ (.A(_0758_),
    .B(net103),
    .C(_0759_),
    .Y(_0760_));
 sg13g2_a21oi_1 _2770_ (.A1(net103),
    .A2(_0756_),
    .Y(_0761_),
    .B1(_0760_));
 sg13g2_nor2b_1 _2771_ (.A(_0747_),
    .B_N(_0761_),
    .Y(_0762_));
 sg13g2_nand2_1 _2772_ (.Y(_0763_),
    .A(net96),
    .B(net134));
 sg13g2_buf_1 _2773_ (.A(net134),
    .X(_0764_));
 sg13g2_or3_1 _2774_ (.A(net87),
    .B(net120),
    .C(_0127_),
    .X(_0765_));
 sg13g2_o21ai_1 _2775_ (.B1(_0765_),
    .Y(_0766_),
    .A1(_0133_),
    .A2(_0763_));
 sg13g2_nor2_1 _2776_ (.A(net121),
    .B(_1945_),
    .Y(_0767_));
 sg13g2_nand2b_1 _2777_ (.Y(_0768_),
    .B(net87),
    .A_N(_0134_));
 sg13g2_o21ai_1 _2778_ (.B1(_0768_),
    .Y(_0769_),
    .A1(net76),
    .A2(_0132_));
 sg13g2_a22oi_1 _2779_ (.Y(_0770_),
    .B1(_0767_),
    .B2(_0769_),
    .A2(_0766_),
    .A1(net121));
 sg13g2_buf_1 _2780_ (.A(_1946_),
    .X(_0771_));
 sg13g2_and2_1 _2781_ (.A(net87),
    .B(_0126_),
    .X(_0772_));
 sg13g2_a21oi_1 _2782_ (.A1(net124),
    .A2(_0124_),
    .Y(_0773_),
    .B1(_0772_));
 sg13g2_nor2b_1 _2783_ (.A(net136),
    .B_N(net141),
    .Y(_0774_));
 sg13g2_buf_1 _2784_ (.A(_0774_),
    .X(_0775_));
 sg13g2_inv_1 _2785_ (.Y(_0776_),
    .A(_0125_));
 sg13g2_a22oi_1 _2786_ (.Y(_0777_),
    .B1(net111),
    .B2(_0776_),
    .A2(_0773_),
    .A1(net98));
 sg13g2_mux4_1 _2787_ (.S0(net98),
    .A0(_0123_),
    .A1(_0120_),
    .A2(_0121_),
    .A3(_0122_),
    .S1(_0695_),
    .X(_0778_));
 sg13g2_mux4_1 _2788_ (.S0(net98),
    .A0(_0131_),
    .A1(_0128_),
    .A2(_0129_),
    .A3(_0130_),
    .S1(_0694_),
    .X(_0779_));
 sg13g2_and2_1 _2789_ (.A(_0771_),
    .B(_0779_),
    .X(_0780_));
 sg13g2_a21oi_1 _2790_ (.A1(net126),
    .A2(_0778_),
    .Y(_0781_),
    .B1(_0780_));
 sg13g2_nand2_1 _2791_ (.Y(_0782_),
    .A(_0707_),
    .B(_0781_));
 sg13g2_o21ai_1 _2792_ (.B1(_0782_),
    .Y(_0783_),
    .A1(net133),
    .A2(_0777_));
 sg13g2_nor3_1 _2793_ (.A(_0771_),
    .B(_0135_),
    .C(net114),
    .Y(_0784_));
 sg13g2_a21oi_1 _2794_ (.A1(_0660_),
    .A2(_0781_),
    .Y(_0785_),
    .B1(_0784_));
 sg13g2_nor2_1 _2795_ (.A(_0764_),
    .B(_0785_),
    .Y(_0786_));
 sg13g2_a21oi_1 _2796_ (.A1(_0764_),
    .A2(_0783_),
    .Y(_0787_),
    .B1(_0786_));
 sg13g2_o21ai_1 _2797_ (.B1(_0787_),
    .Y(_0788_),
    .A1(net126),
    .A2(_0770_));
 sg13g2_nand2b_1 _2798_ (.Y(_0789_),
    .B(net87),
    .A_N(_0118_));
 sg13g2_o21ai_1 _2799_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0695_),
    .A2(_0116_));
 sg13g2_or3_1 _2800_ (.A(net87),
    .B(net120),
    .C(_0111_),
    .X(_0791_));
 sg13g2_o21ai_1 _2801_ (.B1(_0791_),
    .Y(_0792_),
    .A1(_0117_),
    .A2(_0763_));
 sg13g2_a22oi_1 _2802_ (.Y(_0793_),
    .B1(_0792_),
    .B2(net121),
    .A2(_0790_),
    .A1(_0767_));
 sg13g2_inv_1 _2803_ (.Y(_0794_),
    .A(_0109_));
 sg13g2_and2_1 _2804_ (.A(net96),
    .B(_0110_),
    .X(_0795_));
 sg13g2_a21oi_1 _2805_ (.A1(net124),
    .A2(_0108_),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_a22oi_1 _2806_ (.Y(_0797_),
    .B1(_0796_),
    .B2(net98),
    .A2(net111),
    .A1(_0794_));
 sg13g2_mux4_1 _2807_ (.S0(net105),
    .A0(_0107_),
    .A1(_0104_),
    .A2(_0105_),
    .A3(_0106_),
    .S1(net104),
    .X(_0798_));
 sg13g2_mux4_1 _2808_ (.S0(net105),
    .A0(_0115_),
    .A1(_0112_),
    .A2(_0113_),
    .A3(_0114_),
    .S1(net104),
    .X(_0799_));
 sg13g2_and2_1 _2809_ (.A(_1946_),
    .B(_0799_),
    .X(_0800_));
 sg13g2_a21oi_1 _2810_ (.A1(net126),
    .A2(_0798_),
    .Y(_0801_),
    .B1(_0800_));
 sg13g2_nand2_1 _2811_ (.Y(_0802_),
    .A(_0707_),
    .B(_0801_));
 sg13g2_o21ai_1 _2812_ (.B1(_0802_),
    .Y(_0803_),
    .A1(net133),
    .A2(_0797_));
 sg13g2_nor3_1 _2813_ (.A(net133),
    .B(_0119_),
    .C(net114),
    .Y(_0804_));
 sg13g2_a21oi_1 _2814_ (.A1(net114),
    .A2(_0801_),
    .Y(_0805_),
    .B1(_0804_));
 sg13g2_nor2_1 _2815_ (.A(net120),
    .B(_0805_),
    .Y(_0806_));
 sg13g2_a21oi_1 _2816_ (.A1(net120),
    .A2(_0803_),
    .Y(_0807_),
    .B1(_0806_));
 sg13g2_o21ai_1 _2817_ (.B1(_0807_),
    .Y(_0808_),
    .A1(net126),
    .A2(_0793_));
 sg13g2_nor2_1 _2818_ (.A(_0101_),
    .B(_0763_),
    .Y(_0809_));
 sg13g2_nor3_1 _2819_ (.A(net96),
    .B(net120),
    .C(_0095_),
    .Y(_0810_));
 sg13g2_nor2_1 _2820_ (.A(_0809_),
    .B(_0810_),
    .Y(_0811_));
 sg13g2_nand2b_1 _2821_ (.Y(_0812_),
    .B(net96),
    .A_N(_0102_));
 sg13g2_o21ai_1 _2822_ (.B1(_0812_),
    .Y(_0813_),
    .A1(net96),
    .A2(_0100_));
 sg13g2_a21oi_1 _2823_ (.A1(net120),
    .A2(_0813_),
    .Y(_0814_),
    .B1(net121));
 sg13g2_a21oi_1 _2824_ (.A1(net121),
    .A2(_0811_),
    .Y(_0815_),
    .B1(_0814_));
 sg13g2_mux4_1 _2825_ (.S0(net105),
    .A0(_0091_),
    .A1(_0088_),
    .A2(_0089_),
    .A3(_0090_),
    .S1(net104),
    .X(_0816_));
 sg13g2_mux4_1 _2826_ (.S0(net115),
    .A0(_0099_),
    .A1(_0096_),
    .A2(_0097_),
    .A3(_0098_),
    .S1(_0693_),
    .X(_0817_));
 sg13g2_and2_1 _2827_ (.A(_1946_),
    .B(_0817_),
    .X(_0818_));
 sg13g2_a21oi_1 _2828_ (.A1(net126),
    .A2(_0816_),
    .Y(_0819_),
    .B1(_0818_));
 sg13g2_nor3_1 _2829_ (.A(net133),
    .B(_0103_),
    .C(net114),
    .Y(_0820_));
 sg13g2_a21oi_1 _2830_ (.A1(net114),
    .A2(_0819_),
    .Y(_0821_),
    .B1(_0820_));
 sg13g2_nand2_2 _2831_ (.Y(_0822_),
    .A(net121),
    .B(net104));
 sg13g2_nand2_1 _2832_ (.Y(_0823_),
    .A(net104),
    .B(_0094_));
 sg13g2_nand2_1 _2833_ (.Y(_0824_),
    .A(net124),
    .B(_0092_));
 sg13g2_nand3_1 _2834_ (.B(_0823_),
    .C(_0824_),
    .A(net98),
    .Y(_0825_));
 sg13g2_o21ai_1 _2835_ (.B1(_0825_),
    .Y(_0826_),
    .A1(_0093_),
    .A2(_0822_));
 sg13g2_a221oi_1 _2836_ (.B2(net126),
    .C1(_1945_),
    .B1(_0826_),
    .A1(_0707_),
    .Y(_0827_),
    .A2(_0819_));
 sg13g2_a21oi_1 _2837_ (.A1(_1945_),
    .A2(_0821_),
    .Y(_0828_),
    .B1(_0827_));
 sg13g2_a21o_1 _2838_ (.A2(_0815_),
    .A1(net133),
    .B1(_0828_),
    .X(_0829_));
 sg13g2_buf_1 _2839_ (.A(_0829_),
    .X(_0830_));
 sg13g2_mux4_1 _2840_ (.S0(net98),
    .A0(_0079_),
    .A1(_0076_),
    .A2(_0077_),
    .A3(_0078_),
    .S1(net96),
    .X(_0831_));
 sg13g2_mux4_1 _2841_ (.S0(net98),
    .A0(_0087_),
    .A1(_0084_),
    .A2(_0085_),
    .A3(_0086_),
    .S1(net96),
    .X(_0832_));
 sg13g2_mux2_1 _2842_ (.A0(_0831_),
    .A1(_0832_),
    .S(net103),
    .X(_0833_));
 sg13g2_nor2_1 _2843_ (.A(_0708_),
    .B(_0833_),
    .Y(_0834_));
 sg13g2_mux2_1 _2844_ (.A0(_0081_),
    .A1(_0082_),
    .S(_0683_),
    .X(_0835_));
 sg13g2_nor3_1 _2845_ (.A(_0682_),
    .B(_1945_),
    .C(_0083_),
    .Y(_0836_));
 sg13g2_nor3_1 _2846_ (.A(net121),
    .B(net134),
    .C(_0080_),
    .Y(_0837_));
 sg13g2_o21ai_1 _2847_ (.B1(net124),
    .Y(_0838_),
    .A1(_0836_),
    .A2(_0837_));
 sg13g2_o21ai_1 _2848_ (.B1(_0838_),
    .Y(_0839_),
    .A1(_0753_),
    .A2(_0835_));
 sg13g2_mux4_1 _2849_ (.S0(_0683_),
    .A0(_0075_),
    .A1(_0072_),
    .A2(_0073_),
    .A3(_0074_),
    .S1(_0694_),
    .X(_0840_));
 sg13g2_nor3_1 _2850_ (.A(_0758_),
    .B(net103),
    .C(_0840_),
    .Y(_0841_));
 sg13g2_a21oi_1 _2851_ (.A1(net103),
    .A2(_0839_),
    .Y(_0842_),
    .B1(_0841_));
 sg13g2_nor2b_1 _2852_ (.A(_0834_),
    .B_N(_0842_),
    .Y(_0843_));
 sg13g2_mux4_1 _2853_ (.S0(net113),
    .A0(\madd.mem[7][5] ),
    .A1(\madd.mem[5][5] ),
    .A2(\madd.mem[4][5] ),
    .A3(\madd.mem[6][5] ),
    .S1(net105),
    .X(_0844_));
 sg13g2_mux4_1 _2854_ (.S0(net113),
    .A0(\madd.mem[15][5] ),
    .A1(\madd.mem[13][5] ),
    .A2(\madd.mem[12][5] ),
    .A3(\madd.mem[14][5] ),
    .S1(net105),
    .X(_0845_));
 sg13g2_mux2_1 _2855_ (.A0(_0844_),
    .A1(_0845_),
    .S(net112),
    .X(_0846_));
 sg13g2_nor2_1 _2856_ (.A(_0708_),
    .B(_0846_),
    .Y(_0847_));
 sg13g2_nor2_1 _2857_ (.A(_0455_),
    .B(\madd.mem[10][5] ),
    .Y(_0848_));
 sg13g2_nor2_1 _2858_ (.A(_0693_),
    .B(\madd.mem[8][5] ),
    .Y(_0849_));
 sg13g2_o21ai_1 _2859_ (.B1(_0477_),
    .Y(_0850_),
    .A1(_0848_),
    .A2(_0849_));
 sg13g2_nor2_1 _2860_ (.A(\madd.mem[11][5] ),
    .B(_0751_),
    .Y(_0851_));
 sg13g2_nor2_1 _2861_ (.A(\madd.mem[9][5] ),
    .B(_0753_),
    .Y(_0852_));
 sg13g2_o21ai_1 _2862_ (.B1(_0691_),
    .Y(_0853_),
    .A1(_0851_),
    .A2(_0852_));
 sg13g2_nand2_1 _2863_ (.Y(_0854_),
    .A(_0850_),
    .B(_0853_));
 sg13g2_mux4_1 _2864_ (.S0(net113),
    .A0(\madd.mem[3][5] ),
    .A1(\madd.mem[1][5] ),
    .A2(\madd.mem[0][5] ),
    .A3(\madd.mem[2][5] ),
    .S1(net115),
    .X(_0855_));
 sg13g2_nor3_1 _2865_ (.A(_0758_),
    .B(net112),
    .C(_0855_),
    .Y(_0856_));
 sg13g2_a21oi_1 _2866_ (.A1(_0745_),
    .A2(_0854_),
    .Y(_0857_),
    .B1(_0856_));
 sg13g2_nor2b_1 _2867_ (.A(_0847_),
    .B_N(_0857_),
    .Y(_0858_));
 sg13g2_inv_1 _2868_ (.Y(_0859_),
    .A(_0858_));
 sg13g2_mux4_1 _2869_ (.S0(net104),
    .A0(\madd.mem[7][4] ),
    .A1(\madd.mem[5][4] ),
    .A2(\madd.mem[4][4] ),
    .A3(\madd.mem[6][4] ),
    .S1(net105),
    .X(_0860_));
 sg13g2_mux4_1 _2870_ (.S0(net104),
    .A0(\madd.mem[15][4] ),
    .A1(\madd.mem[13][4] ),
    .A2(\madd.mem[12][4] ),
    .A3(\madd.mem[14][4] ),
    .S1(net105),
    .X(_0861_));
 sg13g2_mux2_1 _2871_ (.A0(_0860_),
    .A1(_0861_),
    .S(_0745_),
    .X(_0862_));
 sg13g2_mux4_1 _2872_ (.S0(net113),
    .A0(\madd.mem[3][4] ),
    .A1(\madd.mem[1][4] ),
    .A2(\madd.mem[0][4] ),
    .A3(\madd.mem[2][4] ),
    .S1(_0682_),
    .X(_0863_));
 sg13g2_nand2_1 _2873_ (.Y(_0864_),
    .A(net134),
    .B(\madd.mem[11][4] ));
 sg13g2_mux2_1 _2874_ (.A0(\madd.mem[8][4] ),
    .A1(\madd.mem[10][4] ),
    .S(net113),
    .X(_0865_));
 sg13g2_a22oi_1 _2875_ (.Y(_0866_),
    .B1(_0865_),
    .B2(net115),
    .A2(net111),
    .A1(\madd.mem[9][4] ));
 sg13g2_nand3_1 _2876_ (.B(_0864_),
    .C(_0866_),
    .A(net112),
    .Y(_0867_));
 sg13g2_o21ai_1 _2877_ (.B1(_0867_),
    .Y(_0868_),
    .A1(net103),
    .A2(_0863_));
 sg13g2_nor2_1 _2878_ (.A(_0758_),
    .B(_0868_),
    .Y(_0869_));
 sg13g2_a21oi_1 _2879_ (.A1(_0758_),
    .A2(_0862_),
    .Y(_0870_),
    .B1(_0869_));
 sg13g2_mux4_1 _2880_ (.S0(_1913_),
    .A0(_0174_),
    .A1(_0171_),
    .A2(_0172_),
    .A3(_0173_),
    .S1(_1915_),
    .X(_0871_));
 sg13g2_inv_1 _2881_ (.Y(_0872_),
    .A(_0871_));
 sg13g2_mux4_1 _2882_ (.S0(net136),
    .A0(_0182_),
    .A1(_0179_),
    .A2(_0180_),
    .A3(_0181_),
    .S1(net135),
    .X(_0873_));
 sg13g2_inv_1 _2883_ (.Y(_0874_),
    .A(_0873_));
 sg13g2_mux4_1 _2884_ (.S0(_1912_),
    .A0(_0178_),
    .A1(_0175_),
    .A2(_0176_),
    .A3(_0177_),
    .S1(net141),
    .X(_0875_));
 sg13g2_inv_1 _2885_ (.Y(_0876_),
    .A(_0875_));
 sg13g2_mux4_1 _2886_ (.S0(net136),
    .A0(_0186_),
    .A1(_0183_),
    .A2(_0184_),
    .A3(_0185_),
    .S1(net141),
    .X(_0877_));
 sg13g2_inv_1 _2887_ (.Y(_0878_),
    .A(_0877_));
 sg13g2_mux4_1 _2888_ (.S0(net112),
    .A0(_0872_),
    .A1(_0874_),
    .A2(_0876_),
    .A3(_0878_),
    .S1(_0758_),
    .X(_0879_));
 sg13g2_nor2_1 _2889_ (.A(_0726_),
    .B(_0879_),
    .Y(_0880_));
 sg13g2_a221oi_1 _2890_ (.B2(_0726_),
    .C1(_0669_),
    .B1(_0879_),
    .A1(_0703_),
    .Y(_0881_),
    .A2(_0712_));
 sg13g2_mux4_1 _2891_ (.S0(net123),
    .A0(_0011_),
    .A1(_0008_),
    .A2(_0009_),
    .A3(_0010_),
    .S1(_1991_),
    .X(_0882_));
 sg13g2_nand2_1 _2892_ (.Y(_0883_),
    .A(_0476_),
    .B(_0019_));
 sg13g2_mux2_1 _2893_ (.A0(_0016_),
    .A1(_0018_),
    .S(_1916_),
    .X(_0884_));
 sg13g2_a22oi_1 _2894_ (.Y(_0885_),
    .B1(_0884_),
    .B2(_1990_),
    .A2(net111),
    .A1(_0017_));
 sg13g2_nand2_1 _2895_ (.Y(_0886_),
    .A(_0883_),
    .B(_0885_));
 sg13g2_mux4_1 _2896_ (.S0(net123),
    .A0(_0015_),
    .A1(_0012_),
    .A2(_0013_),
    .A3(_0014_),
    .S1(net125),
    .X(_0887_));
 sg13g2_mux4_1 _2897_ (.S0(net123),
    .A0(_0023_),
    .A1(_0020_),
    .A2(_0021_),
    .A3(_0022_),
    .S1(net125),
    .X(_0888_));
 sg13g2_mux4_1 _2898_ (.S0(_0744_),
    .A0(_0882_),
    .A1(_0886_),
    .A2(_0887_),
    .A3(_0888_),
    .S1(_0758_),
    .X(_0889_));
 sg13g2_o21ai_1 _2899_ (.B1(_0889_),
    .Y(_0890_),
    .A1(_0880_),
    .A2(_0881_));
 sg13g2_nor3_1 _2900_ (.A(_0889_),
    .B(_0880_),
    .C(_0881_),
    .Y(_0891_));
 sg13g2_a21oi_1 _2901_ (.A1(_0730_),
    .A2(_0890_),
    .Y(_0892_),
    .B1(_0891_));
 sg13g2_mux4_1 _2902_ (.S0(net115),
    .A0(_0027_),
    .A1(_0024_),
    .A2(_0025_),
    .A3(_0026_),
    .S1(_0692_),
    .X(_0893_));
 sg13g2_nand2_1 _2903_ (.Y(_0894_),
    .A(net134),
    .B(_0035_));
 sg13g2_mux2_1 _2904_ (.A0(_0032_),
    .A1(_0034_),
    .S(net125),
    .X(_0895_));
 sg13g2_a22oi_1 _2905_ (.Y(_0896_),
    .B1(_0895_),
    .B2(net115),
    .A2(_0775_),
    .A1(_0033_));
 sg13g2_nand3_1 _2906_ (.B(_0894_),
    .C(_0896_),
    .A(net112),
    .Y(_0897_));
 sg13g2_o21ai_1 _2907_ (.B1(_0897_),
    .Y(_0898_),
    .A1(net112),
    .A2(_0893_));
 sg13g2_mux4_1 _2908_ (.S0(net115),
    .A0(_0031_),
    .A1(_0028_),
    .A2(_0029_),
    .A3(_0030_),
    .S1(_0692_),
    .X(_0899_));
 sg13g2_mux4_1 _2909_ (.S0(net115),
    .A0(_0039_),
    .A1(_0036_),
    .A2(_0037_),
    .A3(_0038_),
    .S1(net125),
    .X(_0900_));
 sg13g2_mux2_1 _2910_ (.A0(_0899_),
    .A1(_0900_),
    .S(net112),
    .X(_0901_));
 sg13g2_nor2_1 _2911_ (.A(_0708_),
    .B(_0901_),
    .Y(_0902_));
 sg13g2_a21o_1 _2912_ (.A2(_0898_),
    .A1(_0708_),
    .B1(_0902_),
    .X(_0903_));
 sg13g2_nand2_1 _2913_ (.Y(_0904_),
    .A(_0722_),
    .B(_0903_));
 sg13g2_nor2_1 _2914_ (.A(_0722_),
    .B(_0903_),
    .Y(_0905_));
 sg13g2_a21o_1 _2915_ (.A2(_0904_),
    .A1(_0892_),
    .B1(_0905_),
    .X(_0906_));
 sg13g2_and3_1 _2916_ (.X(_0907_),
    .A(_0859_),
    .B(_0870_),
    .C(_0906_));
 sg13g2_buf_1 _2917_ (.A(_0907_),
    .X(_0908_));
 sg13g2_nand2_1 _2918_ (.Y(_0909_),
    .A(_0843_),
    .B(_0908_));
 sg13g2_nor3_1 _2919_ (.A(_0808_),
    .B(_0830_),
    .C(_0909_),
    .Y(_0910_));
 sg13g2_nor2b_1 _2920_ (.A(_0788_),
    .B_N(_0910_),
    .Y(_0911_));
 sg13g2_xnor2_1 _2921_ (.Y(_0912_),
    .A(_0762_),
    .B(_0911_));
 sg13g2_buf_2 _2922_ (.A(_0912_),
    .X(_0913_));
 sg13g2_buf_1 _2923_ (.A(_0913_),
    .X(_0914_));
 sg13g2_nor2_1 _2924_ (.A(_0699_),
    .B(net26),
    .Y(_0915_));
 sg13g2_a21oi_1 _2925_ (.A1(\madd.mem[0][10] ),
    .A2(net60),
    .Y(_0916_),
    .B1(_0915_));
 sg13g2_o21ai_1 _2926_ (.B1(_0916_),
    .Y(_0214_),
    .A1(_0721_),
    .A2(_0740_));
 sg13g2_nand2_1 _2927_ (.Y(_0917_),
    .A(\madd.mem[0][11] ),
    .B(net60));
 sg13g2_and2_1 _2928_ (.A(net71),
    .B(net86),
    .X(_0918_));
 sg13g2_nor3_1 _2929_ (.A(net47),
    .B(_0578_),
    .C(_0736_),
    .Y(_0919_));
 sg13g2_xor2_1 _2930_ (.B(_0919_),
    .A(_0607_),
    .X(_0920_));
 sg13g2_buf_2 _2931_ (.A(_0920_),
    .X(_0921_));
 sg13g2_nor2b_1 _2932_ (.A(_0762_),
    .B_N(_0911_),
    .Y(_0922_));
 sg13g2_mux4_1 _2933_ (.S0(net76),
    .A0(\madd.mem[3][11] ),
    .A1(\madd.mem[1][11] ),
    .A2(\madd.mem[0][11] ),
    .A3(\madd.mem[2][11] ),
    .S1(net88),
    .X(_0923_));
 sg13g2_nand2_1 _2934_ (.Y(_0924_),
    .A(net120),
    .B(\madd.mem[11][11] ));
 sg13g2_mux2_1 _2935_ (.A0(\madd.mem[8][11] ),
    .A1(\madd.mem[10][11] ),
    .S(_0696_),
    .X(_0925_));
 sg13g2_a22oi_1 _2936_ (.Y(_0926_),
    .B1(_0925_),
    .B2(_0684_),
    .A2(net111),
    .A1(\madd.mem[9][11] ));
 sg13g2_nand2_1 _2937_ (.Y(_0927_),
    .A(_0924_),
    .B(_0926_));
 sg13g2_mux4_1 _2938_ (.S0(net76),
    .A0(\madd.mem[7][11] ),
    .A1(\madd.mem[5][11] ),
    .A2(\madd.mem[4][11] ),
    .A3(\madd.mem[6][11] ),
    .S1(net88),
    .X(_0928_));
 sg13g2_mux4_1 _2939_ (.S0(net76),
    .A0(\madd.mem[15][11] ),
    .A1(\madd.mem[13][11] ),
    .A2(\madd.mem[12][11] ),
    .A3(\madd.mem[14][11] ),
    .S1(net88),
    .X(_0929_));
 sg13g2_mux4_1 _2940_ (.S0(net103),
    .A0(_0923_),
    .A1(_0927_),
    .A2(_0928_),
    .A3(_0929_),
    .S1(_0758_),
    .X(_0930_));
 sg13g2_xor2_1 _2941_ (.B(_0930_),
    .A(_0922_),
    .X(_0931_));
 sg13g2_buf_2 _2942_ (.A(_0931_),
    .X(_0932_));
 sg13g2_buf_8 _2943_ (.A(_0932_),
    .X(_0933_));
 sg13g2_a22oi_1 _2944_ (.Y(_0934_),
    .B1(net23),
    .B2(_0687_),
    .A2(net24),
    .A1(_0918_));
 sg13g2_nand2_1 _2945_ (.Y(_0215_),
    .A(_0917_),
    .B(_0934_));
 sg13g2_xnor2_1 _2946_ (.Y(_0935_),
    .A(_0724_),
    .B(_0545_));
 sg13g2_xnor2_1 _2947_ (.Y(_0936_),
    .A(_0671_),
    .B(_0935_));
 sg13g2_nor2_1 _2948_ (.A(net99),
    .B(_0936_),
    .Y(_0937_));
 sg13g2_buf_2 _2949_ (.A(_0937_),
    .X(_0938_));
 sg13g2_buf_1 _2950_ (.A(_0938_),
    .X(_0939_));
 sg13g2_nand2_1 _2951_ (.Y(_0940_),
    .A(net1),
    .B(_0713_));
 sg13g2_xnor2_1 _2952_ (.Y(_0941_),
    .A(_0724_),
    .B(_0879_));
 sg13g2_xnor2_1 _2953_ (.Y(_0942_),
    .A(_0940_),
    .B(_0941_));
 sg13g2_buf_2 _2954_ (.A(_0942_),
    .X(_0943_));
 sg13g2_buf_1 _2955_ (.A(_0943_),
    .X(_0944_));
 sg13g2_nor2_1 _2956_ (.A(_0699_),
    .B(net65),
    .Y(_0945_));
 sg13g2_a221oi_1 _2957_ (.B2(_0668_),
    .C1(_0945_),
    .B1(net31),
    .A1(\madd.mem[0][1] ),
    .Y(_0946_),
    .A2(net60));
 sg13g2_inv_1 _2958_ (.Y(_0216_),
    .A(_0946_));
 sg13g2_and2_1 _2959_ (.A(_0723_),
    .B(_0731_),
    .X(_0947_));
 sg13g2_a21o_1 _2960_ (.A2(_0728_),
    .A1(_0725_),
    .B1(_0947_),
    .X(_0948_));
 sg13g2_nand3_1 _2961_ (.B(_0728_),
    .C(_0947_),
    .A(_0725_),
    .Y(_0949_));
 sg13g2_a21oi_1 _2962_ (.A1(_0948_),
    .A2(_0949_),
    .Y(_0950_),
    .B1(net99));
 sg13g2_buf_2 _2963_ (.A(_0950_),
    .X(_0951_));
 sg13g2_nand2_1 _2964_ (.Y(_0952_),
    .A(_0668_),
    .B(_0951_));
 sg13g2_nor2_1 _2965_ (.A(_0880_),
    .B(_0881_),
    .Y(_0953_));
 sg13g2_xnor2_1 _2966_ (.Y(_0954_),
    .A(net2),
    .B(_0889_));
 sg13g2_xnor2_1 _2967_ (.Y(_0955_),
    .A(_0953_),
    .B(_0954_));
 sg13g2_buf_2 _2968_ (.A(_0955_),
    .X(_0956_));
 sg13g2_buf_1 _2969_ (.A(_0956_),
    .X(_0957_));
 sg13g2_a22oi_1 _2970_ (.Y(_0958_),
    .B1(net62),
    .B2(_0687_),
    .A2(net60),
    .A1(\madd.mem[0][2] ));
 sg13g2_nand2_1 _2971_ (.Y(_0217_),
    .A(_0952_),
    .B(_0958_));
 sg13g2_nand2_1 _2972_ (.Y(_0959_),
    .A(_0729_),
    .B(_0731_));
 sg13g2_xnor2_1 _2973_ (.Y(_0960_),
    .A(_0722_),
    .B(_0465_));
 sg13g2_xnor2_1 _2974_ (.Y(_0961_),
    .A(_0959_),
    .B(_0960_));
 sg13g2_buf_1 _2975_ (.A(_0961_),
    .X(_0962_));
 sg13g2_nand3_1 _2976_ (.B(net86),
    .C(net30),
    .A(net71),
    .Y(_0963_));
 sg13g2_xnor2_1 _2977_ (.Y(_0964_),
    .A(net3),
    .B(_0903_));
 sg13g2_xnor2_1 _2978_ (.Y(_0965_),
    .A(_0892_),
    .B(_0964_));
 sg13g2_buf_2 _2979_ (.A(_0965_),
    .X(_0966_));
 sg13g2_buf_1 _2980_ (.A(_0966_),
    .X(_0967_));
 sg13g2_a22oi_1 _2981_ (.Y(_0968_),
    .B1(net59),
    .B2(_0687_),
    .A2(_0689_),
    .A1(\madd.mem[0][3] ));
 sg13g2_nand2_1 _2982_ (.Y(_0218_),
    .A(_0963_),
    .B(_0968_));
 sg13g2_xor2_1 _2983_ (.B(_0734_),
    .A(_0555_),
    .X(_0969_));
 sg13g2_nor2_1 _2984_ (.A(_0675_),
    .B(_0969_),
    .Y(_0970_));
 sg13g2_buf_2 _2985_ (.A(_0970_),
    .X(_0971_));
 sg13g2_buf_1 _2986_ (.A(_0971_),
    .X(_0972_));
 sg13g2_xor2_1 _2987_ (.B(_0906_),
    .A(_0870_),
    .X(_0973_));
 sg13g2_buf_2 _2988_ (.A(_0973_),
    .X(_0974_));
 sg13g2_buf_1 _2989_ (.A(_0974_),
    .X(_0975_));
 sg13g2_nor2_1 _2990_ (.A(_0699_),
    .B(net52),
    .Y(_0976_));
 sg13g2_a221oi_1 _2991_ (.B2(net71),
    .C1(_0976_),
    .B1(net22),
    .A1(\madd.mem[0][4] ),
    .Y(_0977_),
    .A2(_0689_));
 sg13g2_inv_1 _2992_ (.Y(_0219_),
    .A(_0977_));
 sg13g2_nand2b_1 _2993_ (.Y(_0978_),
    .B(_0734_),
    .A_N(_0555_));
 sg13g2_xor2_1 _2994_ (.B(_0978_),
    .A(_0442_),
    .X(_0979_));
 sg13g2_and2_1 _2995_ (.A(_0680_),
    .B(_0979_),
    .X(_0980_));
 sg13g2_buf_2 _2996_ (.A(_0980_),
    .X(_0981_));
 sg13g2_buf_1 _2997_ (.A(_0981_),
    .X(_0982_));
 sg13g2_a21oi_1 _2998_ (.A1(_0870_),
    .A2(_0906_),
    .Y(_0983_),
    .B1(_0859_));
 sg13g2_nor2_1 _2999_ (.A(_0908_),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_buf_2 _3000_ (.A(_0984_),
    .X(_0985_));
 sg13g2_buf_1 _3001_ (.A(_0985_),
    .X(_0986_));
 sg13g2_nor2_1 _3002_ (.A(_0699_),
    .B(net33),
    .Y(_0987_));
 sg13g2_a221oi_1 _3003_ (.B2(net71),
    .C1(_0987_),
    .B1(net19),
    .A1(\madd.mem[0][5] ),
    .Y(_0988_),
    .A2(net60));
 sg13g2_inv_1 _3004_ (.Y(_0220_),
    .A(_0988_));
 sg13g2_nor2_1 _3005_ (.A(_0442_),
    .B(_0978_),
    .Y(_0989_));
 sg13g2_xor2_1 _3006_ (.B(_0989_),
    .A(_0434_),
    .X(_0990_));
 sg13g2_nor2_1 _3007_ (.A(net99),
    .B(_0990_),
    .Y(_0991_));
 sg13g2_buf_2 _3008_ (.A(_0991_),
    .X(_0992_));
 sg13g2_xor2_1 _3009_ (.B(_0908_),
    .A(_0843_),
    .X(_0993_));
 sg13g2_buf_2 _3010_ (.A(_0993_),
    .X(_0994_));
 sg13g2_buf_1 _3011_ (.A(_0994_),
    .X(_0995_));
 sg13g2_nand2_1 _3012_ (.Y(_0996_),
    .A(\madd.mem[0][6] ),
    .B(_0688_));
 sg13g2_o21ai_1 _3013_ (.B1(_0996_),
    .Y(_0997_),
    .A1(_0699_),
    .A2(net32));
 sg13g2_a21o_1 _3014_ (.A2(_0992_),
    .A1(net71),
    .B1(_0997_),
    .X(_0221_));
 sg13g2_nor4_2 _3015_ (.A(_0442_),
    .B(_2033_),
    .C(_0434_),
    .Y(_0998_),
    .D(_0978_));
 sg13g2_a21oi_1 _3016_ (.A1(_0734_),
    .A2(_0735_),
    .Y(_0999_),
    .B1(_2034_));
 sg13g2_nor3_1 _3017_ (.A(_0675_),
    .B(_0998_),
    .C(_0999_),
    .Y(_1000_));
 sg13g2_buf_2 _3018_ (.A(_1000_),
    .X(_1001_));
 sg13g2_buf_1 _3019_ (.A(_1001_),
    .X(_1002_));
 sg13g2_xor2_1 _3020_ (.B(_0909_),
    .A(_0830_),
    .X(_1003_));
 sg13g2_buf_2 _3021_ (.A(_1003_),
    .X(_1004_));
 sg13g2_buf_1 _3022_ (.A(_1004_),
    .X(_1005_));
 sg13g2_nor2_1 _3023_ (.A(_0699_),
    .B(net29),
    .Y(_1006_));
 sg13g2_a221oi_1 _3024_ (.B2(net71),
    .C1(_1006_),
    .B1(net18),
    .A1(\madd.mem[0][7] ),
    .Y(_1007_),
    .A2(_0688_));
 sg13g2_inv_1 _3025_ (.Y(_0222_),
    .A(_1007_));
 sg13g2_nand2_1 _3026_ (.Y(_1008_),
    .A(\madd.mem[0][8] ),
    .B(net60));
 sg13g2_xnor2_1 _3027_ (.Y(_1009_),
    .A(_2041_),
    .B(_0998_));
 sg13g2_buf_2 _3028_ (.A(_1009_),
    .X(_1010_));
 sg13g2_nor2_1 _3029_ (.A(_0830_),
    .B(_0909_),
    .Y(_1011_));
 sg13g2_xor2_1 _3030_ (.B(_1011_),
    .A(_0808_),
    .X(_1012_));
 sg13g2_buf_2 _3031_ (.A(_1012_),
    .X(_1013_));
 sg13g2_buf_1 _3032_ (.A(_1013_),
    .X(_1014_));
 sg13g2_a22oi_1 _3033_ (.Y(_1015_),
    .B1(_1014_),
    .B2(_0687_),
    .A2(_1010_),
    .A1(_0918_));
 sg13g2_nand2_1 _3034_ (.Y(_0223_),
    .A(_1008_),
    .B(_1015_));
 sg13g2_nand2_1 _3035_ (.Y(_1016_),
    .A(\madd.mem[0][9] ),
    .B(net60));
 sg13g2_xnor2_1 _3036_ (.Y(_1017_),
    .A(_0579_),
    .B(_0736_));
 sg13g2_buf_2 _3037_ (.A(_1017_),
    .X(_1018_));
 sg13g2_xor2_1 _3038_ (.B(_0910_),
    .A(_0788_),
    .X(_1019_));
 sg13g2_buf_2 _3039_ (.A(_1019_),
    .X(_1020_));
 sg13g2_buf_1 _3040_ (.A(_1020_),
    .X(_1021_));
 sg13g2_a22oi_1 _3041_ (.Y(_1022_),
    .B1(_1021_),
    .B2(_0687_),
    .A2(_1018_),
    .A1(_0918_));
 sg13g2_nand2_1 _3042_ (.Y(_0224_),
    .A(_1016_),
    .B(_1022_));
 sg13g2_buf_1 _3043_ (.A(_0677_),
    .X(_1023_));
 sg13g2_nand2_1 _3044_ (.Y(_1024_),
    .A(_1945_),
    .B(net133));
 sg13g2_buf_1 _3045_ (.A(_1024_),
    .X(_1025_));
 sg13g2_nor2b_2 _3046_ (.A(_0662_),
    .B_N(_1763_),
    .Y(_1026_));
 sg13g2_nand2_2 _3047_ (.Y(_1027_),
    .A(_1026_),
    .B(net111));
 sg13g2_nor2_1 _3048_ (.A(net110),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_buf_1 _3049_ (.A(_1028_),
    .X(_1029_));
 sg13g2_buf_1 _3050_ (.A(_0674_),
    .X(_1030_));
 sg13g2_nand2_2 _3051_ (.Y(_1031_),
    .A(net88),
    .B(_0696_));
 sg13g2_nor3_2 _3052_ (.A(net110),
    .B(_1030_),
    .C(_1031_),
    .Y(_1032_));
 sg13g2_nor3_1 _3053_ (.A(net132),
    .B(net85),
    .C(_1032_),
    .Y(_1033_));
 sg13g2_buf_1 _3054_ (.A(_1033_),
    .X(_1034_));
 sg13g2_nand4_1 _3055_ (.B(net76),
    .C(_2004_),
    .A(_0684_),
    .Y(_1035_),
    .D(_0680_));
 sg13g2_buf_2 _3056_ (.A(_1035_),
    .X(_1036_));
 sg13g2_nor2_1 _3057_ (.A(_0716_),
    .B(_1036_),
    .Y(_1037_));
 sg13g2_a221oi_1 _3058_ (.B2(\madd.mem[10][0] ),
    .C1(_1037_),
    .B1(net58),
    .A1(net39),
    .Y(_1038_),
    .A2(net85));
 sg13g2_inv_1 _3059_ (.Y(_0225_),
    .A(_1038_));
 sg13g2_nor3_2 _3060_ (.A(net110),
    .B(net99),
    .C(_1027_),
    .Y(_1039_));
 sg13g2_nand2b_1 _3061_ (.Y(_1040_),
    .B(_1039_),
    .A_N(_0739_));
 sg13g2_nor2_1 _3062_ (.A(net26),
    .B(_1036_),
    .Y(_1041_));
 sg13g2_a21oi_1 _3063_ (.A1(\madd.mem[10][10] ),
    .A2(net58),
    .Y(_1042_),
    .B1(_1041_));
 sg13g2_nand2_1 _3064_ (.Y(_0226_),
    .A(_1040_),
    .B(_1042_));
 sg13g2_nand2_1 _3065_ (.Y(_1043_),
    .A(\madd.mem[10][11] ),
    .B(_1034_));
 sg13g2_a22oi_1 _3066_ (.Y(_1044_),
    .B1(_1039_),
    .B2(_0921_),
    .A2(_1032_),
    .A1(net23));
 sg13g2_nand2_1 _3067_ (.Y(_0227_),
    .A(_1043_),
    .B(_1044_));
 sg13g2_nor2_1 _3068_ (.A(_0944_),
    .B(_1036_),
    .Y(_1045_));
 sg13g2_a221oi_1 _3069_ (.B2(\madd.mem[10][1] ),
    .C1(_1045_),
    .B1(net58),
    .A1(_0939_),
    .Y(_1046_),
    .A2(net85));
 sg13g2_inv_1 _3070_ (.Y(_0228_),
    .A(_1046_));
 sg13g2_buf_1 _3071_ (.A(_0951_),
    .X(_1047_));
 sg13g2_nand2_1 _3072_ (.Y(_1048_),
    .A(net25),
    .B(net85));
 sg13g2_a22oi_1 _3073_ (.Y(_1049_),
    .B1(net58),
    .B2(\madd.mem[10][2] ),
    .A2(_1032_),
    .A1(_0957_));
 sg13g2_nand2_1 _3074_ (.Y(_0229_),
    .A(_1048_),
    .B(_1049_));
 sg13g2_nand3_1 _3075_ (.B(_0962_),
    .C(_1029_),
    .A(net86),
    .Y(_1050_));
 sg13g2_a22oi_1 _3076_ (.Y(_1051_),
    .B1(_1034_),
    .B2(\madd.mem[10][3] ),
    .A2(_1032_),
    .A1(_0967_));
 sg13g2_nand2_1 _3077_ (.Y(_0230_),
    .A(_1050_),
    .B(_1051_));
 sg13g2_nor2_1 _3078_ (.A(_0975_),
    .B(_1036_),
    .Y(_1052_));
 sg13g2_a221oi_1 _3079_ (.B2(\madd.mem[10][4] ),
    .C1(_1052_),
    .B1(net58),
    .A1(_0972_),
    .Y(_1053_),
    .A2(net85));
 sg13g2_inv_1 _3080_ (.Y(_0231_),
    .A(_1053_));
 sg13g2_nor2_1 _3081_ (.A(net33),
    .B(_1036_),
    .Y(_1054_));
 sg13g2_a221oi_1 _3082_ (.B2(\madd.mem[10][5] ),
    .C1(_1054_),
    .B1(net58),
    .A1(_0982_),
    .Y(_1055_),
    .A2(net85));
 sg13g2_inv_1 _3083_ (.Y(_0232_),
    .A(_1055_));
 sg13g2_buf_1 _3084_ (.A(_0992_),
    .X(_1056_));
 sg13g2_nand2_1 _3085_ (.Y(_1057_),
    .A(\madd.mem[10][6] ),
    .B(_1033_));
 sg13g2_o21ai_1 _3086_ (.B1(_1057_),
    .Y(_1058_),
    .A1(_0995_),
    .A2(_1036_));
 sg13g2_a21o_1 _3087_ (.A2(net85),
    .A1(_1056_),
    .B1(_1058_),
    .X(_0233_));
 sg13g2_nor2_1 _3088_ (.A(_1005_),
    .B(_1036_),
    .Y(_1059_));
 sg13g2_a221oi_1 _3089_ (.B2(\madd.mem[10][7] ),
    .C1(_1059_),
    .B1(_1033_),
    .A1(_1002_),
    .Y(_1060_),
    .A2(net85));
 sg13g2_inv_1 _3090_ (.Y(_0234_),
    .A(_1060_));
 sg13g2_nand2_1 _3091_ (.Y(_1061_),
    .A(\madd.mem[10][8] ),
    .B(net58));
 sg13g2_buf_8 _3092_ (.A(_1010_),
    .X(_1062_));
 sg13g2_a22oi_1 _3093_ (.Y(_1063_),
    .B1(_1039_),
    .B2(_1062_),
    .A2(_1032_),
    .A1(_1014_));
 sg13g2_nand2_1 _3094_ (.Y(_0235_),
    .A(_1061_),
    .B(_1063_));
 sg13g2_nand2_1 _3095_ (.Y(_1064_),
    .A(\madd.mem[10][9] ),
    .B(net58));
 sg13g2_buf_1 _3096_ (.A(_1018_),
    .X(_1065_));
 sg13g2_a22oi_1 _3097_ (.Y(_1066_),
    .B1(_1039_),
    .B2(net21),
    .A2(_1032_),
    .A1(_1021_));
 sg13g2_nand2_1 _3098_ (.Y(_0236_),
    .A(_1064_),
    .B(_1066_));
 sg13g2_or2_1 _3099_ (.X(_1067_),
    .B(_1031_),
    .A(_0664_));
 sg13g2_buf_1 _3100_ (.A(_1067_),
    .X(_1068_));
 sg13g2_nor2_1 _3101_ (.A(net110),
    .B(_1068_),
    .Y(_1069_));
 sg13g2_buf_1 _3102_ (.A(_1069_),
    .X(_1070_));
 sg13g2_nand2_1 _3103_ (.Y(_1071_),
    .A(_1948_),
    .B(_0665_));
 sg13g2_nor2_1 _3104_ (.A(net94),
    .B(_1071_),
    .Y(_1072_));
 sg13g2_buf_2 _3105_ (.A(_1072_),
    .X(_1073_));
 sg13g2_nor3_1 _3106_ (.A(net132),
    .B(net51),
    .C(_1073_),
    .Y(_1074_));
 sg13g2_buf_1 _3107_ (.A(_1074_),
    .X(_1075_));
 sg13g2_nand2_1 _3108_ (.Y(_1076_),
    .A(net120),
    .B(net133));
 sg13g2_buf_2 _3109_ (.A(_1076_),
    .X(_1077_));
 sg13g2_nand2_2 _3110_ (.Y(_1078_),
    .A(_0707_),
    .B(_1026_));
 sg13g2_nor2_1 _3111_ (.A(_1077_),
    .B(_1078_),
    .Y(_1079_));
 sg13g2_buf_1 _3112_ (.A(_1079_),
    .X(_1080_));
 sg13g2_nand2_1 _3113_ (.Y(_1081_),
    .A(net95),
    .B(net84));
 sg13g2_buf_2 _3114_ (.A(_1081_),
    .X(_1082_));
 sg13g2_nor2_1 _3115_ (.A(net70),
    .B(_1082_),
    .Y(_1083_));
 sg13g2_a221oi_1 _3116_ (.B2(\madd.mem[11][0] ),
    .C1(_1083_),
    .B1(net38),
    .A1(net39),
    .Y(_1084_),
    .A2(net51));
 sg13g2_inv_1 _3117_ (.Y(_0237_),
    .A(_1084_));
 sg13g2_nor3_2 _3118_ (.A(net110),
    .B(net99),
    .C(_1068_),
    .Y(_1085_));
 sg13g2_nand2b_1 _3119_ (.Y(_1086_),
    .B(_1085_),
    .A_N(_0739_));
 sg13g2_nor2_1 _3120_ (.A(net26),
    .B(_1082_),
    .Y(_1087_));
 sg13g2_a21oi_1 _3121_ (.A1(\madd.mem[11][10] ),
    .A2(net38),
    .Y(_1088_),
    .B1(_1087_));
 sg13g2_nand2_1 _3122_ (.Y(_0238_),
    .A(_1086_),
    .B(_1088_));
 sg13g2_nand2_1 _3123_ (.Y(_1089_),
    .A(\madd.mem[11][11] ),
    .B(net38));
 sg13g2_a22oi_1 _3124_ (.Y(_1090_),
    .B1(_1085_),
    .B2(net24),
    .A2(_1073_),
    .A1(net23));
 sg13g2_nand2_1 _3125_ (.Y(_0239_),
    .A(_1089_),
    .B(_1090_));
 sg13g2_nor2_1 _3126_ (.A(net65),
    .B(_1082_),
    .Y(_1091_));
 sg13g2_a221oi_1 _3127_ (.B2(\madd.mem[11][1] ),
    .C1(_1091_),
    .B1(net38),
    .A1(net31),
    .Y(_1092_),
    .A2(net51));
 sg13g2_inv_1 _3128_ (.Y(_0240_),
    .A(_1092_));
 sg13g2_nand2_1 _3129_ (.Y(_1093_),
    .A(net25),
    .B(net51));
 sg13g2_a22oi_1 _3130_ (.Y(_1094_),
    .B1(net38),
    .B2(\madd.mem[11][2] ),
    .A2(_1073_),
    .A1(net62));
 sg13g2_nand2_1 _3131_ (.Y(_0241_),
    .A(_1093_),
    .B(_1094_));
 sg13g2_nand3_1 _3132_ (.B(net30),
    .C(net51),
    .A(net86),
    .Y(_1095_));
 sg13g2_a22oi_1 _3133_ (.Y(_1096_),
    .B1(_1075_),
    .B2(\madd.mem[11][3] ),
    .A2(_1073_),
    .A1(net59));
 sg13g2_nand2_1 _3134_ (.Y(_0242_),
    .A(_1095_),
    .B(_1096_));
 sg13g2_nor2_1 _3135_ (.A(net52),
    .B(_1082_),
    .Y(_1097_));
 sg13g2_a221oi_1 _3136_ (.B2(\madd.mem[11][4] ),
    .C1(_1097_),
    .B1(net38),
    .A1(net22),
    .Y(_1098_),
    .A2(net51));
 sg13g2_inv_1 _3137_ (.Y(_0243_),
    .A(_1098_));
 sg13g2_nor2_1 _3138_ (.A(net33),
    .B(_1082_),
    .Y(_1099_));
 sg13g2_a221oi_1 _3139_ (.B2(\madd.mem[11][5] ),
    .C1(_1099_),
    .B1(_1075_),
    .A1(net19),
    .Y(_1100_),
    .A2(_1070_));
 sg13g2_inv_1 _3140_ (.Y(_0244_),
    .A(_1100_));
 sg13g2_nand2_1 _3141_ (.Y(_1101_),
    .A(\madd.mem[11][6] ),
    .B(_1074_));
 sg13g2_o21ai_1 _3142_ (.B1(_1101_),
    .Y(_1102_),
    .A1(net32),
    .A2(_1082_));
 sg13g2_a21o_1 _3143_ (.A2(net51),
    .A1(net16),
    .B1(_1102_),
    .X(_0245_));
 sg13g2_nor2_1 _3144_ (.A(net29),
    .B(_1082_),
    .Y(_1103_));
 sg13g2_a221oi_1 _3145_ (.B2(\madd.mem[11][7] ),
    .C1(_1103_),
    .B1(_1074_),
    .A1(net18),
    .Y(_1104_),
    .A2(net51));
 sg13g2_inv_1 _3146_ (.Y(_0246_),
    .A(_1104_));
 sg13g2_nand2_1 _3147_ (.Y(_1105_),
    .A(\madd.mem[11][8] ),
    .B(net38));
 sg13g2_a22oi_1 _3148_ (.Y(_1106_),
    .B1(_1085_),
    .B2(net17),
    .A2(_1073_),
    .A1(_1013_));
 sg13g2_nand2_1 _3149_ (.Y(_0247_),
    .A(_1105_),
    .B(_1106_));
 sg13g2_nand2_1 _3150_ (.Y(_1107_),
    .A(\madd.mem[11][9] ),
    .B(net38));
 sg13g2_a22oi_1 _3151_ (.Y(_1108_),
    .B1(_1085_),
    .B2(net21),
    .A2(_1073_),
    .A1(_1020_));
 sg13g2_nand2_1 _3152_ (.Y(_0248_),
    .A(_1107_),
    .B(_1108_));
 sg13g2_nor2_2 _3153_ (.A(_0664_),
    .B(_0685_),
    .Y(_1109_));
 sg13g2_nand2_1 _3154_ (.Y(_1110_),
    .A(_1948_),
    .B(_1109_));
 sg13g2_nor2_1 _3155_ (.A(net94),
    .B(_1110_),
    .Y(_1111_));
 sg13g2_buf_2 _3156_ (.A(_1111_),
    .X(_1112_));
 sg13g2_nor3_1 _3157_ (.A(net122),
    .B(net84),
    .C(_1112_),
    .Y(_1113_));
 sg13g2_buf_1 _3158_ (.A(_1113_),
    .X(_1114_));
 sg13g2_nand2_1 _3159_ (.Y(_1115_),
    .A(_1026_),
    .B(_0697_));
 sg13g2_nor2_1 _3160_ (.A(_1077_),
    .B(_1115_),
    .Y(_1116_));
 sg13g2_buf_1 _3161_ (.A(_1116_),
    .X(_1117_));
 sg13g2_nand2_1 _3162_ (.Y(_1118_),
    .A(net95),
    .B(net57));
 sg13g2_buf_2 _3163_ (.A(_1118_),
    .X(_1119_));
 sg13g2_nor2_1 _3164_ (.A(net70),
    .B(_1119_),
    .Y(_1120_));
 sg13g2_a221oi_1 _3165_ (.B2(\madd.mem[12][0] ),
    .C1(_1120_),
    .B1(net46),
    .A1(net39),
    .Y(_1121_),
    .A2(net84));
 sg13g2_inv_1 _3166_ (.Y(_0249_),
    .A(_1121_));
 sg13g2_nor2_1 _3167_ (.A(net26),
    .B(_1119_),
    .Y(_1122_));
 sg13g2_a21oi_1 _3168_ (.A1(\madd.mem[12][10] ),
    .A2(_1113_),
    .Y(_1123_),
    .B1(_1122_));
 sg13g2_o21ai_1 _3169_ (.B1(_1123_),
    .Y(_0250_),
    .A1(net20),
    .A2(_1082_));
 sg13g2_nand2_1 _3170_ (.Y(_1124_),
    .A(net95),
    .B(net24));
 sg13g2_buf_8 _3171_ (.A(_1124_),
    .X(_1125_));
 sg13g2_a22oi_1 _3172_ (.Y(_1126_),
    .B1(_1114_),
    .B2(\madd.mem[12][11] ),
    .A2(_1112_),
    .A1(net23));
 sg13g2_o21ai_1 _3173_ (.B1(_1126_),
    .Y(_0251_),
    .A1(_1071_),
    .A2(_1125_));
 sg13g2_nor2_1 _3174_ (.A(net65),
    .B(_1119_),
    .Y(_1127_));
 sg13g2_a221oi_1 _3175_ (.B2(\madd.mem[12][1] ),
    .C1(_1127_),
    .B1(net46),
    .A1(net31),
    .Y(_1128_),
    .A2(net84));
 sg13g2_inv_1 _3176_ (.Y(_0252_),
    .A(_1128_));
 sg13g2_nand2_1 _3177_ (.Y(_1129_),
    .A(net25),
    .B(net84));
 sg13g2_a22oi_1 _3178_ (.Y(_1130_),
    .B1(net46),
    .B2(\madd.mem[12][2] ),
    .A2(_1112_),
    .A1(net62));
 sg13g2_nand2_1 _3179_ (.Y(_0253_),
    .A(_1129_),
    .B(_1130_));
 sg13g2_nand2_1 _3180_ (.Y(_1131_),
    .A(net95),
    .B(net30));
 sg13g2_buf_2 _3181_ (.A(_1131_),
    .X(_1132_));
 sg13g2_a22oi_1 _3182_ (.Y(_1133_),
    .B1(net46),
    .B2(\madd.mem[12][3] ),
    .A2(_1112_),
    .A1(net59));
 sg13g2_o21ai_1 _3183_ (.B1(_1133_),
    .Y(_0254_),
    .A1(_1132_),
    .A2(_1071_));
 sg13g2_nor2_1 _3184_ (.A(net52),
    .B(_1119_),
    .Y(_1134_));
 sg13g2_a221oi_1 _3185_ (.B2(\madd.mem[12][4] ),
    .C1(_1134_),
    .B1(net46),
    .A1(net22),
    .Y(_1135_),
    .A2(net84));
 sg13g2_inv_1 _3186_ (.Y(_0255_),
    .A(_1135_));
 sg13g2_nor2_1 _3187_ (.A(net33),
    .B(_1119_),
    .Y(_1136_));
 sg13g2_a221oi_1 _3188_ (.B2(\madd.mem[12][5] ),
    .C1(_1136_),
    .B1(_1114_),
    .A1(net19),
    .Y(_1137_),
    .A2(_1080_));
 sg13g2_inv_1 _3189_ (.Y(_0256_),
    .A(_1137_));
 sg13g2_nand2_1 _3190_ (.Y(_1138_),
    .A(\madd.mem[12][6] ),
    .B(_1113_));
 sg13g2_o21ai_1 _3191_ (.B1(_1138_),
    .Y(_1139_),
    .A1(net32),
    .A2(_1119_));
 sg13g2_a21o_1 _3192_ (.A2(net84),
    .A1(net16),
    .B1(_1139_),
    .X(_0257_));
 sg13g2_nor2_1 _3193_ (.A(net29),
    .B(_1119_),
    .Y(_1140_));
 sg13g2_a221oi_1 _3194_ (.B2(\madd.mem[12][7] ),
    .C1(_1140_),
    .B1(net46),
    .A1(net18),
    .Y(_1141_),
    .A2(net84));
 sg13g2_inv_1 _3195_ (.Y(_0258_),
    .A(_1141_));
 sg13g2_nand2_1 _3196_ (.Y(_1142_),
    .A(\madd.mem[12][8] ),
    .B(net46));
 sg13g2_a22oi_1 _3197_ (.Y(_1143_),
    .B1(_1112_),
    .B2(net28),
    .A2(_1073_),
    .A1(net17));
 sg13g2_nand2_1 _3198_ (.Y(_0259_),
    .A(_1142_),
    .B(_1143_));
 sg13g2_nand2_1 _3199_ (.Y(_1144_),
    .A(\madd.mem[12][9] ),
    .B(net46));
 sg13g2_a22oi_1 _3200_ (.Y(_1145_),
    .B1(_1112_),
    .B2(net27),
    .A2(_1073_),
    .A1(net21));
 sg13g2_nand2_1 _3201_ (.Y(_0260_),
    .A(_1144_),
    .B(_1145_));
 sg13g2_nor3_2 _3202_ (.A(_1077_),
    .B(net94),
    .C(_0822_),
    .Y(_1146_));
 sg13g2_nor3_1 _3203_ (.A(net122),
    .B(net57),
    .C(_1146_),
    .Y(_1147_));
 sg13g2_buf_1 _3204_ (.A(_1147_),
    .X(_1148_));
 sg13g2_nand3_1 _3205_ (.B(net97),
    .C(_0775_),
    .A(_1948_),
    .Y(_1149_));
 sg13g2_buf_2 _3206_ (.A(_1149_),
    .X(_1150_));
 sg13g2_nor2_1 _3207_ (.A(net70),
    .B(_1150_),
    .Y(_1151_));
 sg13g2_a221oi_1 _3208_ (.B2(\madd.mem[13][0] ),
    .C1(_1151_),
    .B1(net45),
    .A1(net39),
    .Y(_1152_),
    .A2(net57));
 sg13g2_inv_1 _3209_ (.Y(_0261_),
    .A(_1152_));
 sg13g2_nor2_1 _3210_ (.A(net26),
    .B(_1150_),
    .Y(_1153_));
 sg13g2_a21oi_1 _3211_ (.A1(\madd.mem[13][10] ),
    .A2(_1147_),
    .Y(_1154_),
    .B1(_1153_));
 sg13g2_o21ai_1 _3212_ (.B1(_1154_),
    .Y(_0262_),
    .A1(net20),
    .A2(_1119_));
 sg13g2_a22oi_1 _3213_ (.Y(_1155_),
    .B1(net45),
    .B2(\madd.mem[13][11] ),
    .A2(_1146_),
    .A1(net23));
 sg13g2_o21ai_1 _3214_ (.B1(_1155_),
    .Y(_0263_),
    .A1(_1110_),
    .A2(_1125_));
 sg13g2_nor2_1 _3215_ (.A(net65),
    .B(_1150_),
    .Y(_1156_));
 sg13g2_a221oi_1 _3216_ (.B2(\madd.mem[13][1] ),
    .C1(_1156_),
    .B1(net45),
    .A1(net31),
    .Y(_1157_),
    .A2(net57));
 sg13g2_inv_1 _3217_ (.Y(_0264_),
    .A(_1157_));
 sg13g2_nand2_1 _3218_ (.Y(_1158_),
    .A(net25),
    .B(net57));
 sg13g2_a22oi_1 _3219_ (.Y(_1159_),
    .B1(net45),
    .B2(\madd.mem[13][2] ),
    .A2(_1146_),
    .A1(net62));
 sg13g2_nand2_1 _3220_ (.Y(_0265_),
    .A(_1158_),
    .B(_1159_));
 sg13g2_a22oi_1 _3221_ (.Y(_1160_),
    .B1(_1148_),
    .B2(\madd.mem[13][3] ),
    .A2(_1146_),
    .A1(net59));
 sg13g2_o21ai_1 _3222_ (.B1(_1160_),
    .Y(_0266_),
    .A1(_1132_),
    .A2(_1110_));
 sg13g2_nor2_1 _3223_ (.A(net52),
    .B(_1150_),
    .Y(_1161_));
 sg13g2_a221oi_1 _3224_ (.B2(\madd.mem[13][4] ),
    .C1(_1161_),
    .B1(net45),
    .A1(net22),
    .Y(_1162_),
    .A2(_1117_));
 sg13g2_inv_1 _3225_ (.Y(_0267_),
    .A(_1162_));
 sg13g2_nor2_1 _3226_ (.A(net33),
    .B(_1150_),
    .Y(_1163_));
 sg13g2_a221oi_1 _3227_ (.B2(\madd.mem[13][5] ),
    .C1(_1163_),
    .B1(_1148_),
    .A1(net19),
    .Y(_1164_),
    .A2(net57));
 sg13g2_inv_1 _3228_ (.Y(_0268_),
    .A(_1164_));
 sg13g2_nand2_1 _3229_ (.Y(_1165_),
    .A(\madd.mem[13][6] ),
    .B(_1147_));
 sg13g2_o21ai_1 _3230_ (.B1(_1165_),
    .Y(_1166_),
    .A1(net32),
    .A2(_1150_));
 sg13g2_a21o_1 _3231_ (.A2(net57),
    .A1(net16),
    .B1(_1166_),
    .X(_0269_));
 sg13g2_nor2_1 _3232_ (.A(net29),
    .B(_1150_),
    .Y(_1167_));
 sg13g2_a221oi_1 _3233_ (.B2(\madd.mem[13][7] ),
    .C1(_1167_),
    .B1(net45),
    .A1(net18),
    .Y(_1168_),
    .A2(net57));
 sg13g2_inv_1 _3234_ (.Y(_0270_),
    .A(_1168_));
 sg13g2_nand2_1 _3235_ (.Y(_1169_),
    .A(\madd.mem[13][8] ),
    .B(net45));
 sg13g2_a22oi_1 _3236_ (.Y(_1170_),
    .B1(_1146_),
    .B2(net28),
    .A2(_1112_),
    .A1(net17));
 sg13g2_nand2_1 _3237_ (.Y(_0271_),
    .A(_1169_),
    .B(_1170_));
 sg13g2_nand2_1 _3238_ (.Y(_1171_),
    .A(\madd.mem[13][9] ),
    .B(net45));
 sg13g2_a22oi_1 _3239_ (.Y(_1172_),
    .B1(_1146_),
    .B2(net27),
    .A2(_1112_),
    .A1(net21));
 sg13g2_nand2_1 _3240_ (.Y(_0272_),
    .A(_1171_),
    .B(_1172_));
 sg13g2_nor2_1 _3241_ (.A(_1077_),
    .B(_1027_),
    .Y(_1173_));
 sg13g2_buf_1 _3242_ (.A(_1173_),
    .X(_1174_));
 sg13g2_nor2_1 _3243_ (.A(_0664_),
    .B(_1031_),
    .Y(_1175_));
 sg13g2_nand2_1 _3244_ (.Y(_1176_),
    .A(_1948_),
    .B(_1175_));
 sg13g2_nor2_1 _3245_ (.A(_1030_),
    .B(_1176_),
    .Y(_1177_));
 sg13g2_buf_2 _3246_ (.A(_1177_),
    .X(_1178_));
 sg13g2_nor3_1 _3247_ (.A(net132),
    .B(net83),
    .C(_1178_),
    .Y(_1179_));
 sg13g2_buf_1 _3248_ (.A(_1179_),
    .X(_1180_));
 sg13g2_nor2_1 _3249_ (.A(_1077_),
    .B(_1068_),
    .Y(_1181_));
 sg13g2_buf_1 _3250_ (.A(_1181_),
    .X(_1182_));
 sg13g2_nand2_1 _3251_ (.Y(_1183_),
    .A(net95),
    .B(net50));
 sg13g2_buf_2 _3252_ (.A(_1183_),
    .X(_1184_));
 sg13g2_nor2_1 _3253_ (.A(net70),
    .B(_1184_),
    .Y(_1185_));
 sg13g2_a221oi_1 _3254_ (.B2(\madd.mem[14][0] ),
    .C1(_1185_),
    .B1(net37),
    .A1(net39),
    .Y(_1186_),
    .A2(net83));
 sg13g2_inv_1 _3255_ (.Y(_0273_),
    .A(_1186_));
 sg13g2_nor3_2 _3256_ (.A(_1077_),
    .B(net99),
    .C(_1027_),
    .Y(_1187_));
 sg13g2_nand2b_1 _3257_ (.Y(_1188_),
    .B(_1187_),
    .A_N(_0739_));
 sg13g2_nor2_1 _3258_ (.A(net26),
    .B(_1184_),
    .Y(_1189_));
 sg13g2_a21oi_1 _3259_ (.A1(\madd.mem[14][10] ),
    .A2(net37),
    .Y(_1190_),
    .B1(_1189_));
 sg13g2_nand2_1 _3260_ (.Y(_0274_),
    .A(_1188_),
    .B(_1190_));
 sg13g2_nand2_1 _3261_ (.Y(_1191_),
    .A(\madd.mem[14][11] ),
    .B(net37));
 sg13g2_a22oi_1 _3262_ (.Y(_1192_),
    .B1(_1187_),
    .B2(net24),
    .A2(_1178_),
    .A1(net23));
 sg13g2_nand2_1 _3263_ (.Y(_0275_),
    .A(_1191_),
    .B(_1192_));
 sg13g2_nor2_1 _3264_ (.A(net65),
    .B(_1184_),
    .Y(_1193_));
 sg13g2_a221oi_1 _3265_ (.B2(\madd.mem[14][1] ),
    .C1(_1193_),
    .B1(net37),
    .A1(net31),
    .Y(_1194_),
    .A2(net83));
 sg13g2_inv_1 _3266_ (.Y(_0276_),
    .A(_1194_));
 sg13g2_nand2_1 _3267_ (.Y(_1195_),
    .A(net25),
    .B(net83));
 sg13g2_a22oi_1 _3268_ (.Y(_1196_),
    .B1(net37),
    .B2(\madd.mem[14][2] ),
    .A2(_1178_),
    .A1(net62));
 sg13g2_nand2_1 _3269_ (.Y(_0277_),
    .A(_1195_),
    .B(_1196_));
 sg13g2_nand3_1 _3270_ (.B(net30),
    .C(_1174_),
    .A(net86),
    .Y(_1197_));
 sg13g2_a22oi_1 _3271_ (.Y(_1198_),
    .B1(_1180_),
    .B2(\madd.mem[14][3] ),
    .A2(_1178_),
    .A1(net59));
 sg13g2_nand2_1 _3272_ (.Y(_0278_),
    .A(_1197_),
    .B(_1198_));
 sg13g2_nor2_1 _3273_ (.A(net52),
    .B(_1184_),
    .Y(_1199_));
 sg13g2_a221oi_1 _3274_ (.B2(\madd.mem[14][4] ),
    .C1(_1199_),
    .B1(net37),
    .A1(net22),
    .Y(_1200_),
    .A2(net83));
 sg13g2_inv_1 _3275_ (.Y(_0279_),
    .A(_1200_));
 sg13g2_nor2_1 _3276_ (.A(net33),
    .B(_1184_),
    .Y(_1201_));
 sg13g2_a221oi_1 _3277_ (.B2(\madd.mem[14][5] ),
    .C1(_1201_),
    .B1(_1180_),
    .A1(net19),
    .Y(_1202_),
    .A2(net83));
 sg13g2_inv_1 _3278_ (.Y(_0280_),
    .A(_1202_));
 sg13g2_nand2_1 _3279_ (.Y(_1203_),
    .A(\madd.mem[14][6] ),
    .B(_1179_));
 sg13g2_o21ai_1 _3280_ (.B1(_1203_),
    .Y(_1204_),
    .A1(net32),
    .A2(_1184_));
 sg13g2_a21o_1 _3281_ (.A2(net83),
    .A1(net16),
    .B1(_1204_),
    .X(_0281_));
 sg13g2_nor2_1 _3282_ (.A(net29),
    .B(_1184_),
    .Y(_1205_));
 sg13g2_a221oi_1 _3283_ (.B2(\madd.mem[14][7] ),
    .C1(_1205_),
    .B1(_1179_),
    .A1(net18),
    .Y(_1206_),
    .A2(net83));
 sg13g2_inv_1 _3284_ (.Y(_0282_),
    .A(_1206_));
 sg13g2_nand2_1 _3285_ (.Y(_1207_),
    .A(\madd.mem[14][8] ),
    .B(net37));
 sg13g2_a22oi_1 _3286_ (.Y(_1208_),
    .B1(_1187_),
    .B2(net17),
    .A2(_1178_),
    .A1(_1013_));
 sg13g2_nand2_1 _3287_ (.Y(_0283_),
    .A(_1207_),
    .B(_1208_));
 sg13g2_nand2_1 _3288_ (.Y(_1209_),
    .A(\madd.mem[14][9] ),
    .B(net37));
 sg13g2_a22oi_1 _3289_ (.Y(_1210_),
    .B1(_1187_),
    .B2(net21),
    .A2(_1178_),
    .A1(_1020_));
 sg13g2_nand2_1 _3290_ (.Y(_0284_),
    .A(_1209_),
    .B(_1210_));
 sg13g2_nor2_2 _3291_ (.A(net114),
    .B(_0681_),
    .Y(_1211_));
 sg13g2_nor3_1 _3292_ (.A(net122),
    .B(net50),
    .C(_1211_),
    .Y(_1212_));
 sg13g2_buf_1 _3293_ (.A(_1212_),
    .X(_1213_));
 sg13g2_nand3_1 _3294_ (.B(_0707_),
    .C(_0690_),
    .A(net127),
    .Y(_1214_));
 sg13g2_buf_2 _3295_ (.A(_1214_),
    .X(_1215_));
 sg13g2_nor2_1 _3296_ (.A(net70),
    .B(_1215_),
    .Y(_1216_));
 sg13g2_a221oi_1 _3297_ (.B2(\madd.mem[15][0] ),
    .C1(_1216_),
    .B1(net36),
    .A1(net39),
    .Y(_1217_),
    .A2(net50));
 sg13g2_inv_1 _3298_ (.Y(_0285_),
    .A(_1217_));
 sg13g2_nor2_1 _3299_ (.A(net26),
    .B(_1215_),
    .Y(_1218_));
 sg13g2_a21oi_1 _3300_ (.A1(\madd.mem[15][10] ),
    .A2(_1212_),
    .Y(_1219_),
    .B1(_1218_));
 sg13g2_o21ai_1 _3301_ (.B1(_1219_),
    .Y(_0286_),
    .A1(net20),
    .A2(_1184_));
 sg13g2_a22oi_1 _3302_ (.Y(_1220_),
    .B1(net36),
    .B2(\madd.mem[15][11] ),
    .A2(_1211_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3303_ (.B1(_1220_),
    .Y(_0287_),
    .A1(_1125_),
    .A2(_1176_));
 sg13g2_nor2_1 _3304_ (.A(net65),
    .B(_1215_),
    .Y(_1221_));
 sg13g2_a221oi_1 _3305_ (.B2(\madd.mem[15][1] ),
    .C1(_1221_),
    .B1(net36),
    .A1(net31),
    .Y(_1222_),
    .A2(net50));
 sg13g2_inv_1 _3306_ (.Y(_0288_),
    .A(_1222_));
 sg13g2_nand2_1 _3307_ (.Y(_1223_),
    .A(net25),
    .B(_1182_));
 sg13g2_a22oi_1 _3308_ (.Y(_1224_),
    .B1(net36),
    .B2(\madd.mem[15][2] ),
    .A2(_1211_),
    .A1(net62));
 sg13g2_nand2_1 _3309_ (.Y(_0289_),
    .A(_1223_),
    .B(_1224_));
 sg13g2_a22oi_1 _3310_ (.Y(_1225_),
    .B1(_1213_),
    .B2(\madd.mem[15][3] ),
    .A2(_1211_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3311_ (.B1(_1225_),
    .Y(_0290_),
    .A1(_1132_),
    .A2(_1176_));
 sg13g2_nor2_1 _3312_ (.A(net52),
    .B(_1215_),
    .Y(_1226_));
 sg13g2_a221oi_1 _3313_ (.B2(\madd.mem[15][4] ),
    .C1(_1226_),
    .B1(net36),
    .A1(net22),
    .Y(_1227_),
    .A2(net50));
 sg13g2_inv_1 _3314_ (.Y(_0291_),
    .A(_1227_));
 sg13g2_nor2_1 _3315_ (.A(net33),
    .B(_1215_),
    .Y(_1228_));
 sg13g2_a221oi_1 _3316_ (.B2(\madd.mem[15][5] ),
    .C1(_1228_),
    .B1(_1213_),
    .A1(net19),
    .Y(_1229_),
    .A2(net50));
 sg13g2_inv_1 _3317_ (.Y(_0292_),
    .A(_1229_));
 sg13g2_nand2_1 _3318_ (.Y(_1230_),
    .A(\madd.mem[15][6] ),
    .B(_1212_));
 sg13g2_o21ai_1 _3319_ (.B1(_1230_),
    .Y(_1231_),
    .A1(net32),
    .A2(_1215_));
 sg13g2_a21o_1 _3320_ (.A2(net50),
    .A1(net16),
    .B1(_1231_),
    .X(_0293_));
 sg13g2_nor2_1 _3321_ (.A(net29),
    .B(_1215_),
    .Y(_1232_));
 sg13g2_a221oi_1 _3322_ (.B2(\madd.mem[15][7] ),
    .C1(_1232_),
    .B1(net36),
    .A1(net18),
    .Y(_1233_),
    .A2(net50));
 sg13g2_inv_1 _3323_ (.Y(_0294_),
    .A(_1233_));
 sg13g2_nand2_1 _3324_ (.Y(_1234_),
    .A(\madd.mem[15][8] ),
    .B(net36));
 sg13g2_a22oi_1 _3325_ (.Y(_1235_),
    .B1(_1211_),
    .B2(net28),
    .A2(_1178_),
    .A1(net17));
 sg13g2_nand2_1 _3326_ (.Y(_0295_),
    .A(_1234_),
    .B(_1235_));
 sg13g2_nand2_1 _3327_ (.Y(_1236_),
    .A(\madd.mem[15][9] ),
    .B(net36));
 sg13g2_a22oi_1 _3328_ (.Y(_1237_),
    .B1(_1211_),
    .B2(net27),
    .A2(_1178_),
    .A1(net21));
 sg13g2_nand2_1 _3329_ (.Y(_0296_),
    .A(_1236_),
    .B(_1237_));
 sg13g2_and2_1 _3330_ (.A(net127),
    .B(_1109_),
    .X(_1238_));
 sg13g2_buf_1 _3331_ (.A(_1238_),
    .X(_1239_));
 sg13g2_nor2_2 _3332_ (.A(_0681_),
    .B(_0822_),
    .Y(_1240_));
 sg13g2_nor3_1 _3333_ (.A(net132),
    .B(net61),
    .C(_1240_),
    .Y(_1241_));
 sg13g2_buf_1 _3334_ (.A(_1241_),
    .X(_1242_));
 sg13g2_nand3_1 _3335_ (.B(net97),
    .C(net111),
    .A(net127),
    .Y(_1243_));
 sg13g2_buf_2 _3336_ (.A(_1243_),
    .X(_1244_));
 sg13g2_nor2_1 _3337_ (.A(net70),
    .B(_1244_),
    .Y(_1245_));
 sg13g2_a221oi_1 _3338_ (.B2(\madd.mem[1][0] ),
    .C1(_1245_),
    .B1(net49),
    .A1(net39),
    .Y(_1246_),
    .A2(net61));
 sg13g2_inv_1 _3339_ (.Y(_0297_),
    .A(_1246_));
 sg13g2_and2_1 _3340_ (.A(net95),
    .B(net61),
    .X(_1247_));
 sg13g2_buf_1 _3341_ (.A(_1247_),
    .X(_1248_));
 sg13g2_inv_1 _3342_ (.Y(_1249_),
    .A(_1248_));
 sg13g2_nor2_1 _3343_ (.A(_0914_),
    .B(_1244_),
    .Y(_1250_));
 sg13g2_a21oi_1 _3344_ (.A1(\madd.mem[1][10] ),
    .A2(_1241_),
    .Y(_1251_),
    .B1(_1250_));
 sg13g2_o21ai_1 _3345_ (.B1(_1251_),
    .Y(_0298_),
    .A1(net20),
    .A2(_1249_));
 sg13g2_nand2_1 _3346_ (.Y(_1252_),
    .A(\madd.mem[1][11] ),
    .B(net49));
 sg13g2_a22oi_1 _3347_ (.Y(_1253_),
    .B1(_1248_),
    .B2(net24),
    .A2(_1240_),
    .A1(net23));
 sg13g2_nand2_1 _3348_ (.Y(_0299_),
    .A(_1252_),
    .B(_1253_));
 sg13g2_nor2_1 _3349_ (.A(net65),
    .B(_1244_),
    .Y(_1254_));
 sg13g2_a221oi_1 _3350_ (.B2(\madd.mem[1][1] ),
    .C1(_1254_),
    .B1(net49),
    .A1(net31),
    .Y(_1255_),
    .A2(_1239_));
 sg13g2_inv_1 _3351_ (.Y(_0300_),
    .A(_1255_));
 sg13g2_nand2_1 _3352_ (.Y(_1256_),
    .A(net25),
    .B(_1239_));
 sg13g2_a22oi_1 _3353_ (.Y(_1257_),
    .B1(net49),
    .B2(\madd.mem[1][2] ),
    .A2(_1240_),
    .A1(net62));
 sg13g2_nand2_1 _3354_ (.Y(_0301_),
    .A(_1256_),
    .B(_1257_));
 sg13g2_nand3_1 _3355_ (.B(net30),
    .C(net61),
    .A(net86),
    .Y(_1258_));
 sg13g2_a22oi_1 _3356_ (.Y(_1259_),
    .B1(_1242_),
    .B2(\madd.mem[1][3] ),
    .A2(_1240_),
    .A1(net59));
 sg13g2_nand2_1 _3357_ (.Y(_0302_),
    .A(_1258_),
    .B(_1259_));
 sg13g2_nor2_1 _3358_ (.A(net52),
    .B(_1244_),
    .Y(_1260_));
 sg13g2_a221oi_1 _3359_ (.B2(\madd.mem[1][4] ),
    .C1(_1260_),
    .B1(net49),
    .A1(net22),
    .Y(_1261_),
    .A2(net61));
 sg13g2_inv_1 _3360_ (.Y(_0303_),
    .A(_1261_));
 sg13g2_nor2_1 _3361_ (.A(net33),
    .B(_1244_),
    .Y(_1262_));
 sg13g2_a221oi_1 _3362_ (.B2(\madd.mem[1][5] ),
    .C1(_1262_),
    .B1(_1242_),
    .A1(net19),
    .Y(_1263_),
    .A2(net61));
 sg13g2_inv_1 _3363_ (.Y(_0304_),
    .A(_1263_));
 sg13g2_nand2_1 _3364_ (.Y(_1264_),
    .A(\madd.mem[1][6] ),
    .B(_1241_));
 sg13g2_o21ai_1 _3365_ (.B1(_1264_),
    .Y(_1265_),
    .A1(net32),
    .A2(_1244_));
 sg13g2_a21o_1 _3366_ (.A2(net61),
    .A1(net16),
    .B1(_1265_),
    .X(_0305_));
 sg13g2_nor2_1 _3367_ (.A(net29),
    .B(_1244_),
    .Y(_1266_));
 sg13g2_a221oi_1 _3368_ (.B2(\madd.mem[1][7] ),
    .C1(_1266_),
    .B1(net49),
    .A1(net18),
    .Y(_1267_),
    .A2(net61));
 sg13g2_inv_1 _3369_ (.Y(_0306_),
    .A(_1267_));
 sg13g2_nand2_1 _3370_ (.Y(_1268_),
    .A(\madd.mem[1][8] ),
    .B(net49));
 sg13g2_a22oi_1 _3371_ (.Y(_1269_),
    .B1(_1248_),
    .B2(net17),
    .A2(_1240_),
    .A1(_1013_));
 sg13g2_nand2_1 _3372_ (.Y(_0307_),
    .A(_1268_),
    .B(_1269_));
 sg13g2_nand2_1 _3373_ (.Y(_1270_),
    .A(\madd.mem[1][9] ),
    .B(net49));
 sg13g2_a22oi_1 _3374_ (.Y(_1271_),
    .B1(_1248_),
    .B2(net21),
    .A2(_1240_),
    .A1(_1020_));
 sg13g2_nand2_1 _3375_ (.Y(_0308_),
    .A(_1270_),
    .B(_1271_));
 sg13g2_nor2_1 _3376_ (.A(_0664_),
    .B(_0822_),
    .Y(_1272_));
 sg13g2_and2_1 _3377_ (.A(net127),
    .B(_1272_),
    .X(_1273_));
 sg13g2_buf_1 _3378_ (.A(_1273_),
    .X(_1274_));
 sg13g2_nor2_2 _3379_ (.A(_0681_),
    .B(_1031_),
    .Y(_1275_));
 sg13g2_nor3_1 _3380_ (.A(net132),
    .B(net69),
    .C(_1275_),
    .Y(_1276_));
 sg13g2_buf_1 _3381_ (.A(_1276_),
    .X(_1277_));
 sg13g2_or2_1 _3382_ (.X(_1278_),
    .B(_1031_),
    .A(_0681_));
 sg13g2_buf_2 _3383_ (.A(_1278_),
    .X(_1279_));
 sg13g2_nor2_1 _3384_ (.A(net70),
    .B(_1279_),
    .Y(_1280_));
 sg13g2_a221oi_1 _3385_ (.B2(\madd.mem[2][0] ),
    .C1(_1280_),
    .B1(net56),
    .A1(_1023_),
    .Y(_1281_),
    .A2(net69));
 sg13g2_inv_1 _3386_ (.Y(_0309_),
    .A(_1281_));
 sg13g2_and2_1 _3387_ (.A(_0719_),
    .B(net69),
    .X(_1282_));
 sg13g2_buf_1 _3388_ (.A(_1282_),
    .X(_1283_));
 sg13g2_nand2b_1 _3389_ (.Y(_1284_),
    .B(_1283_),
    .A_N(_0739_));
 sg13g2_nor2_1 _3390_ (.A(_0914_),
    .B(_1279_),
    .Y(_1285_));
 sg13g2_a21oi_1 _3391_ (.A1(\madd.mem[2][10] ),
    .A2(net56),
    .Y(_1286_),
    .B1(_1285_));
 sg13g2_nand2_1 _3392_ (.Y(_0310_),
    .A(_1284_),
    .B(_1286_));
 sg13g2_nand2_1 _3393_ (.Y(_1287_),
    .A(\madd.mem[2][11] ),
    .B(net56));
 sg13g2_a22oi_1 _3394_ (.Y(_1288_),
    .B1(_1283_),
    .B2(net24),
    .A2(_1275_),
    .A1(_0933_));
 sg13g2_nand2_1 _3395_ (.Y(_0311_),
    .A(_1287_),
    .B(_1288_));
 sg13g2_nor2_1 _3396_ (.A(net65),
    .B(_1279_),
    .Y(_1289_));
 sg13g2_a221oi_1 _3397_ (.B2(\madd.mem[2][1] ),
    .C1(_1289_),
    .B1(net56),
    .A1(net31),
    .Y(_1290_),
    .A2(_1274_));
 sg13g2_inv_1 _3398_ (.Y(_0312_),
    .A(_1290_));
 sg13g2_nand2_1 _3399_ (.Y(_1291_),
    .A(_1047_),
    .B(net69));
 sg13g2_a22oi_1 _3400_ (.Y(_1292_),
    .B1(net56),
    .B2(\madd.mem[2][2] ),
    .A2(_1275_),
    .A1(_0957_));
 sg13g2_nand2_1 _3401_ (.Y(_0313_),
    .A(_1291_),
    .B(_1292_));
 sg13g2_nand3_1 _3402_ (.B(net30),
    .C(_1274_),
    .A(_0720_),
    .Y(_1293_));
 sg13g2_a22oi_1 _3403_ (.Y(_1294_),
    .B1(_1277_),
    .B2(\madd.mem[2][3] ),
    .A2(_1275_),
    .A1(net59));
 sg13g2_nand2_1 _3404_ (.Y(_0314_),
    .A(_1293_),
    .B(_1294_));
 sg13g2_nor2_1 _3405_ (.A(_0975_),
    .B(_1279_),
    .Y(_1295_));
 sg13g2_a221oi_1 _3406_ (.B2(\madd.mem[2][4] ),
    .C1(_1295_),
    .B1(net56),
    .A1(_0972_),
    .Y(_1296_),
    .A2(net69));
 sg13g2_inv_1 _3407_ (.Y(_0315_),
    .A(_1296_));
 sg13g2_nor2_1 _3408_ (.A(_0986_),
    .B(_1279_),
    .Y(_1297_));
 sg13g2_a221oi_1 _3409_ (.B2(\madd.mem[2][5] ),
    .C1(_1297_),
    .B1(_1277_),
    .A1(_0982_),
    .Y(_1298_),
    .A2(net69));
 sg13g2_inv_1 _3410_ (.Y(_0316_),
    .A(_1298_));
 sg13g2_nand2_1 _3411_ (.Y(_1299_),
    .A(\madd.mem[2][6] ),
    .B(_1276_));
 sg13g2_o21ai_1 _3412_ (.B1(_1299_),
    .Y(_1300_),
    .A1(net32),
    .A2(_1279_));
 sg13g2_a21o_1 _3413_ (.A2(net69),
    .A1(net16),
    .B1(_1300_),
    .X(_0317_));
 sg13g2_nor2_1 _3414_ (.A(net29),
    .B(_1279_),
    .Y(_1301_));
 sg13g2_a221oi_1 _3415_ (.B2(\madd.mem[2][7] ),
    .C1(_1301_),
    .B1(_1276_),
    .A1(net18),
    .Y(_1302_),
    .A2(net69));
 sg13g2_inv_1 _3416_ (.Y(_0318_),
    .A(_1302_));
 sg13g2_nand2_1 _3417_ (.Y(_1303_),
    .A(\madd.mem[2][8] ),
    .B(net56));
 sg13g2_a22oi_1 _3418_ (.Y(_1304_),
    .B1(_1283_),
    .B2(net17),
    .A2(_1275_),
    .A1(_1013_));
 sg13g2_nand2_1 _3419_ (.Y(_0319_),
    .A(_1303_),
    .B(_1304_));
 sg13g2_nand2_1 _3420_ (.Y(_1305_),
    .A(\madd.mem[2][9] ),
    .B(net56));
 sg13g2_a22oi_1 _3421_ (.Y(_1306_),
    .B1(_1283_),
    .B2(_1065_),
    .A2(_1275_),
    .A1(_1020_));
 sg13g2_nand2_1 _3422_ (.Y(_0320_),
    .A(_1305_),
    .B(_1306_));
 sg13g2_and2_1 _3423_ (.A(net127),
    .B(_1175_),
    .X(_1307_));
 sg13g2_buf_1 _3424_ (.A(_1307_),
    .X(_1308_));
 sg13g2_nor2_1 _3425_ (.A(_1945_),
    .B(net133),
    .Y(_1309_));
 sg13g2_nand2_1 _3426_ (.Y(_1310_),
    .A(_1309_),
    .B(_0665_));
 sg13g2_nor2_1 _3427_ (.A(net94),
    .B(_1310_),
    .Y(_1311_));
 sg13g2_buf_2 _3428_ (.A(_1311_),
    .X(_1312_));
 sg13g2_nor3_1 _3429_ (.A(_0678_),
    .B(net55),
    .C(_1312_),
    .Y(_1313_));
 sg13g2_buf_1 _3430_ (.A(_1313_),
    .X(_1314_));
 sg13g2_nor2_1 _3431_ (.A(_1972_),
    .B(_1078_),
    .Y(_1315_));
 sg13g2_buf_1 _3432_ (.A(_1315_),
    .X(_1316_));
 sg13g2_nand2_1 _3433_ (.Y(_1317_),
    .A(net97),
    .B(net82));
 sg13g2_buf_2 _3434_ (.A(_1317_),
    .X(_1318_));
 sg13g2_nor2_1 _3435_ (.A(_0716_),
    .B(_1318_),
    .Y(_1319_));
 sg13g2_a221oi_1 _3436_ (.B2(\madd.mem[3][0] ),
    .C1(_1319_),
    .B1(net44),
    .A1(_1023_),
    .Y(_1320_),
    .A2(net55));
 sg13g2_inv_1 _3437_ (.Y(_0321_),
    .A(_1320_));
 sg13g2_and2_1 _3438_ (.A(_0719_),
    .B(net55),
    .X(_1321_));
 sg13g2_buf_1 _3439_ (.A(_1321_),
    .X(_1322_));
 sg13g2_inv_1 _3440_ (.Y(_1323_),
    .A(_1322_));
 sg13g2_nor2_1 _3441_ (.A(_0913_),
    .B(_1318_),
    .Y(_1324_));
 sg13g2_a21oi_1 _3442_ (.A1(\madd.mem[3][10] ),
    .A2(_1313_),
    .Y(_1325_),
    .B1(_1324_));
 sg13g2_o21ai_1 _3443_ (.B1(_1325_),
    .Y(_0322_),
    .A1(_0740_),
    .A2(_1323_));
 sg13g2_nand2_1 _3444_ (.Y(_1326_),
    .A(\madd.mem[3][11] ),
    .B(net44));
 sg13g2_a22oi_1 _3445_ (.Y(_1327_),
    .B1(_1322_),
    .B2(net24),
    .A2(_1312_),
    .A1(_0933_));
 sg13g2_nand2_1 _3446_ (.Y(_0323_),
    .A(_1326_),
    .B(_1327_));
 sg13g2_nor2_1 _3447_ (.A(_0944_),
    .B(_1318_),
    .Y(_1328_));
 sg13g2_a221oi_1 _3448_ (.B2(\madd.mem[3][1] ),
    .C1(_1328_),
    .B1(net44),
    .A1(_0939_),
    .Y(_1329_),
    .A2(net55));
 sg13g2_inv_1 _3449_ (.Y(_0324_),
    .A(_1329_));
 sg13g2_nand2_1 _3450_ (.Y(_1330_),
    .A(_1047_),
    .B(_1308_));
 sg13g2_a22oi_1 _3451_ (.Y(_1331_),
    .B1(net44),
    .B2(\madd.mem[3][2] ),
    .A2(_1312_),
    .A1(net62));
 sg13g2_nand2_1 _3452_ (.Y(_0325_),
    .A(_1330_),
    .B(_1331_));
 sg13g2_nand3_1 _3453_ (.B(net30),
    .C(net55),
    .A(_0720_),
    .Y(_1332_));
 sg13g2_a22oi_1 _3454_ (.Y(_1333_),
    .B1(_1314_),
    .B2(\madd.mem[3][3] ),
    .A2(_1312_),
    .A1(_0967_));
 sg13g2_nand2_1 _3455_ (.Y(_0326_),
    .A(_1332_),
    .B(_1333_));
 sg13g2_nor2_1 _3456_ (.A(net52),
    .B(_1318_),
    .Y(_1334_));
 sg13g2_a221oi_1 _3457_ (.B2(\madd.mem[3][4] ),
    .C1(_1334_),
    .B1(net44),
    .A1(net22),
    .Y(_1335_),
    .A2(net55));
 sg13g2_inv_1 _3458_ (.Y(_0327_),
    .A(_1335_));
 sg13g2_nor2_1 _3459_ (.A(_0986_),
    .B(_1318_),
    .Y(_1336_));
 sg13g2_a221oi_1 _3460_ (.B2(\madd.mem[3][5] ),
    .C1(_1336_),
    .B1(_1314_),
    .A1(net19),
    .Y(_1337_),
    .A2(_1308_));
 sg13g2_inv_1 _3461_ (.Y(_0328_),
    .A(_1337_));
 sg13g2_nand2_1 _3462_ (.Y(_1338_),
    .A(\madd.mem[3][6] ),
    .B(_1313_));
 sg13g2_o21ai_1 _3463_ (.B1(_1338_),
    .Y(_1339_),
    .A1(_0995_),
    .A2(_1318_));
 sg13g2_a21o_1 _3464_ (.A2(net55),
    .A1(_1056_),
    .B1(_1339_),
    .X(_0329_));
 sg13g2_nor2_1 _3465_ (.A(_1005_),
    .B(_1318_),
    .Y(_1340_));
 sg13g2_a221oi_1 _3466_ (.B2(\madd.mem[3][7] ),
    .C1(_1340_),
    .B1(net44),
    .A1(_1002_),
    .Y(_1341_),
    .A2(net55));
 sg13g2_inv_1 _3467_ (.Y(_0330_),
    .A(_1341_));
 sg13g2_nand2_1 _3468_ (.Y(_1342_),
    .A(\madd.mem[3][8] ),
    .B(net44));
 sg13g2_a22oi_1 _3469_ (.Y(_1343_),
    .B1(_1322_),
    .B2(_1062_),
    .A2(_1312_),
    .A1(_1013_));
 sg13g2_nand2_1 _3470_ (.Y(_0331_),
    .A(_1342_),
    .B(_1343_));
 sg13g2_nand2_1 _3471_ (.Y(_1344_),
    .A(\madd.mem[3][9] ),
    .B(net44));
 sg13g2_a22oi_1 _3472_ (.Y(_1345_),
    .B1(_1322_),
    .B2(_1065_),
    .A2(_1312_),
    .A1(_1020_));
 sg13g2_nand2_1 _3473_ (.Y(_0332_),
    .A(_1344_),
    .B(_1345_));
 sg13g2_nand2_1 _3474_ (.Y(_1346_),
    .A(_1309_),
    .B(_1109_));
 sg13g2_nor2_1 _3475_ (.A(net94),
    .B(_1346_),
    .Y(_1347_));
 sg13g2_buf_2 _3476_ (.A(_1347_),
    .X(_1348_));
 sg13g2_nor3_1 _3477_ (.A(net122),
    .B(net82),
    .C(_1348_),
    .Y(_1349_));
 sg13g2_buf_1 _3478_ (.A(_1349_),
    .X(_1350_));
 sg13g2_nor2_1 _3479_ (.A(_1972_),
    .B(_1115_),
    .Y(_1351_));
 sg13g2_buf_1 _3480_ (.A(_1351_),
    .X(_1352_));
 sg13g2_nand2_1 _3481_ (.Y(_1353_),
    .A(net97),
    .B(net54));
 sg13g2_buf_2 _3482_ (.A(_1353_),
    .X(_1354_));
 sg13g2_nor2_1 _3483_ (.A(_0715_),
    .B(_1354_),
    .Y(_1355_));
 sg13g2_a221oi_1 _3484_ (.B2(\madd.mem[4][0] ),
    .C1(_1355_),
    .B1(net43),
    .A1(net39),
    .Y(_1356_),
    .A2(net82));
 sg13g2_inv_1 _3485_ (.Y(_0333_),
    .A(_1356_));
 sg13g2_nor2_1 _3486_ (.A(_0913_),
    .B(_1354_),
    .Y(_1357_));
 sg13g2_a21oi_1 _3487_ (.A1(\madd.mem[4][10] ),
    .A2(_1349_),
    .Y(_1358_),
    .B1(_1357_));
 sg13g2_o21ai_1 _3488_ (.B1(_1358_),
    .Y(_0334_),
    .A1(net20),
    .A2(_1318_));
 sg13g2_a22oi_1 _3489_ (.Y(_1359_),
    .B1(net43),
    .B2(\madd.mem[4][11] ),
    .A2(_1348_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3490_ (.B1(_1359_),
    .Y(_0335_),
    .A1(_1125_),
    .A2(_1310_));
 sg13g2_nor2_1 _3491_ (.A(_0943_),
    .B(_1354_),
    .Y(_1360_));
 sg13g2_a221oi_1 _3492_ (.B2(\madd.mem[4][1] ),
    .C1(_1360_),
    .B1(net43),
    .A1(_0938_),
    .Y(_1361_),
    .A2(net82));
 sg13g2_inv_1 _3493_ (.Y(_0336_),
    .A(_1361_));
 sg13g2_nand2_1 _3494_ (.Y(_1362_),
    .A(net25),
    .B(_1316_));
 sg13g2_a22oi_1 _3495_ (.Y(_1363_),
    .B1(_1350_),
    .B2(\madd.mem[4][2] ),
    .A2(_1348_),
    .A1(_0956_));
 sg13g2_nand2_1 _3496_ (.Y(_0337_),
    .A(_1362_),
    .B(_1363_));
 sg13g2_a22oi_1 _3497_ (.Y(_1364_),
    .B1(_1350_),
    .B2(\madd.mem[4][3] ),
    .A2(_1348_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3498_ (.B1(_1364_),
    .Y(_0338_),
    .A1(_1132_),
    .A2(_1310_));
 sg13g2_nor2_1 _3499_ (.A(_0974_),
    .B(_1354_),
    .Y(_1365_));
 sg13g2_a221oi_1 _3500_ (.B2(\madd.mem[4][4] ),
    .C1(_1365_),
    .B1(net43),
    .A1(_0971_),
    .Y(_1366_),
    .A2(net82));
 sg13g2_inv_1 _3501_ (.Y(_0339_),
    .A(_1366_));
 sg13g2_nor2_1 _3502_ (.A(_0985_),
    .B(_1354_),
    .Y(_1367_));
 sg13g2_a221oi_1 _3503_ (.B2(\madd.mem[4][5] ),
    .C1(_1367_),
    .B1(net43),
    .A1(_0981_),
    .Y(_1368_),
    .A2(net82));
 sg13g2_inv_1 _3504_ (.Y(_0340_),
    .A(_1368_));
 sg13g2_nand2_1 _3505_ (.Y(_1369_),
    .A(\madd.mem[4][6] ),
    .B(_1349_));
 sg13g2_o21ai_1 _3506_ (.B1(_1369_),
    .Y(_1370_),
    .A1(_0994_),
    .A2(_1354_));
 sg13g2_a21o_1 _3507_ (.A2(net82),
    .A1(net16),
    .B1(_1370_),
    .X(_0341_));
 sg13g2_nor2_1 _3508_ (.A(_1004_),
    .B(_1354_),
    .Y(_1371_));
 sg13g2_a221oi_1 _3509_ (.B2(\madd.mem[4][7] ),
    .C1(_1371_),
    .B1(net43),
    .A1(_1001_),
    .Y(_1372_),
    .A2(net82));
 sg13g2_inv_1 _3510_ (.Y(_0342_),
    .A(_1372_));
 sg13g2_nand2_1 _3511_ (.Y(_1373_),
    .A(\madd.mem[4][8] ),
    .B(net43));
 sg13g2_a22oi_1 _3512_ (.Y(_1374_),
    .B1(_1348_),
    .B2(net28),
    .A2(_1312_),
    .A1(_1010_));
 sg13g2_nand2_1 _3513_ (.Y(_0343_),
    .A(_1373_),
    .B(_1374_));
 sg13g2_nand2_1 _3514_ (.Y(_1375_),
    .A(\madd.mem[4][9] ),
    .B(net43));
 sg13g2_a22oi_1 _3515_ (.Y(_1376_),
    .B1(_1348_),
    .B2(net27),
    .A2(_1312_),
    .A1(_1018_));
 sg13g2_nand2_1 _3516_ (.Y(_0344_),
    .A(_1375_),
    .B(_1376_));
 sg13g2_nand2_1 _3517_ (.Y(_1377_),
    .A(_1309_),
    .B(_1272_));
 sg13g2_nor2_1 _3518_ (.A(_0674_),
    .B(_1377_),
    .Y(_1378_));
 sg13g2_buf_2 _3519_ (.A(_1378_),
    .X(_1379_));
 sg13g2_nor3_1 _3520_ (.A(net122),
    .B(net54),
    .C(_1379_),
    .Y(_1380_));
 sg13g2_buf_1 _3521_ (.A(_1380_),
    .X(_1381_));
 sg13g2_nor2_1 _3522_ (.A(_1972_),
    .B(_1027_),
    .Y(_1382_));
 sg13g2_buf_1 _3523_ (.A(_1382_),
    .X(_1383_));
 sg13g2_nand2_1 _3524_ (.Y(_1384_),
    .A(net97),
    .B(net81));
 sg13g2_buf_2 _3525_ (.A(_1384_),
    .X(_1385_));
 sg13g2_nor2_1 _3526_ (.A(_0715_),
    .B(_1385_),
    .Y(_1386_));
 sg13g2_a221oi_1 _3527_ (.B2(\madd.mem[5][0] ),
    .C1(_1386_),
    .B1(net42),
    .A1(_0677_),
    .Y(_1387_),
    .A2(net54));
 sg13g2_inv_1 _3528_ (.Y(_0345_),
    .A(_1387_));
 sg13g2_nor2_1 _3529_ (.A(_0913_),
    .B(_1385_),
    .Y(_1388_));
 sg13g2_a21oi_1 _3530_ (.A1(\madd.mem[5][10] ),
    .A2(_1380_),
    .Y(_1389_),
    .B1(_1388_));
 sg13g2_o21ai_1 _3531_ (.B1(_1389_),
    .Y(_0346_),
    .A1(net20),
    .A2(_1354_));
 sg13g2_a22oi_1 _3532_ (.Y(_1390_),
    .B1(_1381_),
    .B2(\madd.mem[5][11] ),
    .A2(_1379_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3533_ (.B1(_1390_),
    .Y(_0347_),
    .A1(_1125_),
    .A2(_1346_));
 sg13g2_nor2_1 _3534_ (.A(_0943_),
    .B(_1385_),
    .Y(_1391_));
 sg13g2_a221oi_1 _3535_ (.B2(\madd.mem[5][1] ),
    .C1(_1391_),
    .B1(net42),
    .A1(_0938_),
    .Y(_1392_),
    .A2(net54));
 sg13g2_inv_1 _3536_ (.Y(_0348_),
    .A(_1392_));
 sg13g2_nand2_1 _3537_ (.Y(_1393_),
    .A(_0951_),
    .B(_1352_));
 sg13g2_a22oi_1 _3538_ (.Y(_1394_),
    .B1(net42),
    .B2(\madd.mem[5][2] ),
    .A2(_1379_),
    .A1(_0956_));
 sg13g2_nand2_1 _3539_ (.Y(_0349_),
    .A(_1393_),
    .B(_1394_));
 sg13g2_a22oi_1 _3540_ (.Y(_1395_),
    .B1(net42),
    .B2(\madd.mem[5][3] ),
    .A2(_1379_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3541_ (.B1(_1395_),
    .Y(_0350_),
    .A1(_1132_),
    .A2(_1346_));
 sg13g2_nor2_1 _3542_ (.A(_0974_),
    .B(_1385_),
    .Y(_1396_));
 sg13g2_a221oi_1 _3543_ (.B2(\madd.mem[5][4] ),
    .C1(_1396_),
    .B1(_1381_),
    .A1(_0971_),
    .Y(_1397_),
    .A2(net54));
 sg13g2_inv_1 _3544_ (.Y(_0351_),
    .A(_1397_));
 sg13g2_nor2_1 _3545_ (.A(_0985_),
    .B(_1385_),
    .Y(_1398_));
 sg13g2_a221oi_1 _3546_ (.B2(\madd.mem[5][5] ),
    .C1(_1398_),
    .B1(net42),
    .A1(_0981_),
    .Y(_1399_),
    .A2(net54));
 sg13g2_inv_1 _3547_ (.Y(_0352_),
    .A(_1399_));
 sg13g2_nand2_1 _3548_ (.Y(_1400_),
    .A(\madd.mem[5][6] ),
    .B(_1380_));
 sg13g2_o21ai_1 _3549_ (.B1(_1400_),
    .Y(_1401_),
    .A1(_0994_),
    .A2(_1385_));
 sg13g2_a21o_1 _3550_ (.A2(net54),
    .A1(_0992_),
    .B1(_1401_),
    .X(_0353_));
 sg13g2_nor2_1 _3551_ (.A(_1004_),
    .B(_1385_),
    .Y(_1402_));
 sg13g2_a221oi_1 _3552_ (.B2(\madd.mem[5][7] ),
    .C1(_1402_),
    .B1(net42),
    .A1(_1001_),
    .Y(_1403_),
    .A2(net54));
 sg13g2_inv_1 _3553_ (.Y(_0354_),
    .A(_1403_));
 sg13g2_nand2_1 _3554_ (.Y(_1404_),
    .A(\madd.mem[5][8] ),
    .B(net42));
 sg13g2_a22oi_1 _3555_ (.Y(_1405_),
    .B1(_1379_),
    .B2(net28),
    .A2(_1348_),
    .A1(_1010_));
 sg13g2_nand2_1 _3556_ (.Y(_0355_),
    .A(_1404_),
    .B(_1405_));
 sg13g2_nand2_1 _3557_ (.Y(_1406_),
    .A(\madd.mem[5][9] ),
    .B(net42));
 sg13g2_a22oi_1 _3558_ (.Y(_1407_),
    .B1(_1379_),
    .B2(net27),
    .A2(_1348_),
    .A1(_1018_));
 sg13g2_nand2_1 _3559_ (.Y(_0356_),
    .A(_1406_),
    .B(_1407_));
 sg13g2_nand2_1 _3560_ (.Y(_1408_),
    .A(_1309_),
    .B(_1175_));
 sg13g2_nor2_1 _3561_ (.A(_0674_),
    .B(_1408_),
    .Y(_1409_));
 sg13g2_buf_2 _3562_ (.A(_1409_),
    .X(_1410_));
 sg13g2_nor3_1 _3563_ (.A(net122),
    .B(net81),
    .C(_1410_),
    .Y(_1411_));
 sg13g2_buf_1 _3564_ (.A(_1411_),
    .X(_1412_));
 sg13g2_nor2_1 _3565_ (.A(_1972_),
    .B(_1068_),
    .Y(_1413_));
 sg13g2_buf_1 _3566_ (.A(_1413_),
    .X(_1414_));
 sg13g2_nand2_1 _3567_ (.Y(_1415_),
    .A(net97),
    .B(net48));
 sg13g2_buf_2 _3568_ (.A(_1415_),
    .X(_1416_));
 sg13g2_nor2_1 _3569_ (.A(_0715_),
    .B(_1416_),
    .Y(_1417_));
 sg13g2_a221oi_1 _3570_ (.B2(\madd.mem[6][0] ),
    .C1(_1417_),
    .B1(net35),
    .A1(_0677_),
    .Y(_1418_),
    .A2(net81));
 sg13g2_inv_1 _3571_ (.Y(_0357_),
    .A(_1418_));
 sg13g2_nor2_1 _3572_ (.A(_0913_),
    .B(_1416_),
    .Y(_1419_));
 sg13g2_a21oi_1 _3573_ (.A1(\madd.mem[6][10] ),
    .A2(_1411_),
    .Y(_1420_),
    .B1(_1419_));
 sg13g2_o21ai_1 _3574_ (.B1(_1420_),
    .Y(_0358_),
    .A1(net20),
    .A2(_1385_));
 sg13g2_a22oi_1 _3575_ (.Y(_1421_),
    .B1(net35),
    .B2(\madd.mem[6][11] ),
    .A2(_1410_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3576_ (.B1(_1421_),
    .Y(_0359_),
    .A1(_1125_),
    .A2(_1377_));
 sg13g2_nor2_1 _3577_ (.A(_0943_),
    .B(_1416_),
    .Y(_1422_));
 sg13g2_a221oi_1 _3578_ (.B2(\madd.mem[6][1] ),
    .C1(_1422_),
    .B1(net35),
    .A1(_0938_),
    .Y(_1423_),
    .A2(net81));
 sg13g2_inv_1 _3579_ (.Y(_0360_),
    .A(_1423_));
 sg13g2_nand2_1 _3580_ (.Y(_1424_),
    .A(_0951_),
    .B(_1383_));
 sg13g2_a22oi_1 _3581_ (.Y(_1425_),
    .B1(net35),
    .B2(\madd.mem[6][2] ),
    .A2(_1410_),
    .A1(_0956_));
 sg13g2_nand2_1 _3582_ (.Y(_0361_),
    .A(_1424_),
    .B(_1425_));
 sg13g2_a22oi_1 _3583_ (.Y(_1426_),
    .B1(_1412_),
    .B2(\madd.mem[6][3] ),
    .A2(_1410_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3584_ (.B1(_1426_),
    .Y(_0362_),
    .A1(_1132_),
    .A2(_1377_));
 sg13g2_nor2_1 _3585_ (.A(_0974_),
    .B(_1416_),
    .Y(_1427_));
 sg13g2_a221oi_1 _3586_ (.B2(\madd.mem[6][4] ),
    .C1(_1427_),
    .B1(net35),
    .A1(_0971_),
    .Y(_1428_),
    .A2(net81));
 sg13g2_inv_1 _3587_ (.Y(_0363_),
    .A(_1428_));
 sg13g2_nor2_1 _3588_ (.A(_0985_),
    .B(_1416_),
    .Y(_1429_));
 sg13g2_a221oi_1 _3589_ (.B2(\madd.mem[6][5] ),
    .C1(_1429_),
    .B1(_1412_),
    .A1(_0981_),
    .Y(_1430_),
    .A2(net81));
 sg13g2_inv_1 _3590_ (.Y(_0364_),
    .A(_1430_));
 sg13g2_nand2_1 _3591_ (.Y(_1431_),
    .A(\madd.mem[6][6] ),
    .B(_1411_));
 sg13g2_o21ai_1 _3592_ (.B1(_1431_),
    .Y(_1432_),
    .A1(_0994_),
    .A2(_1416_));
 sg13g2_a21o_1 _3593_ (.A2(net81),
    .A1(_0992_),
    .B1(_1432_),
    .X(_0365_));
 sg13g2_nor2_1 _3594_ (.A(_1004_),
    .B(_1416_),
    .Y(_1433_));
 sg13g2_a221oi_1 _3595_ (.B2(\madd.mem[6][7] ),
    .C1(_1433_),
    .B1(net35),
    .A1(_1001_),
    .Y(_1434_),
    .A2(net81));
 sg13g2_inv_1 _3596_ (.Y(_0366_),
    .A(_1434_));
 sg13g2_nand2_1 _3597_ (.Y(_1435_),
    .A(\madd.mem[6][8] ),
    .B(net35));
 sg13g2_a22oi_1 _3598_ (.Y(_1436_),
    .B1(_1410_),
    .B2(net28),
    .A2(_1379_),
    .A1(_1010_));
 sg13g2_nand2_1 _3599_ (.Y(_0367_),
    .A(_1435_),
    .B(_1436_));
 sg13g2_nand2_1 _3600_ (.Y(_1437_),
    .A(\madd.mem[6][9] ),
    .B(net35));
 sg13g2_a22oi_1 _3601_ (.Y(_1438_),
    .B1(_1410_),
    .B2(net27),
    .A2(_1379_),
    .A1(_1018_));
 sg13g2_nand2_1 _3602_ (.Y(_0368_),
    .A(_1437_),
    .B(_1438_));
 sg13g2_nor3_2 _3603_ (.A(net110),
    .B(net114),
    .C(net94),
    .Y(_1439_));
 sg13g2_nor3_1 _3604_ (.A(net122),
    .B(net48),
    .C(_1439_),
    .Y(_1440_));
 sg13g2_buf_1 _3605_ (.A(_1440_),
    .X(_1441_));
 sg13g2_nand3_1 _3606_ (.B(_0707_),
    .C(net97),
    .A(_2004_),
    .Y(_1442_));
 sg13g2_buf_2 _3607_ (.A(_1442_),
    .X(_1443_));
 sg13g2_nor2_1 _3608_ (.A(_0715_),
    .B(_1443_),
    .Y(_1444_));
 sg13g2_a221oi_1 _3609_ (.B2(\madd.mem[7][0] ),
    .C1(_1444_),
    .B1(net34),
    .A1(_0677_),
    .Y(_1445_),
    .A2(net48));
 sg13g2_inv_1 _3610_ (.Y(_0369_),
    .A(_1445_));
 sg13g2_nor2_1 _3611_ (.A(_0913_),
    .B(_1443_),
    .Y(_1446_));
 sg13g2_a21oi_1 _3612_ (.A1(\madd.mem[7][10] ),
    .A2(_1440_),
    .Y(_1447_),
    .B1(_1446_));
 sg13g2_o21ai_1 _3613_ (.B1(_1447_),
    .Y(_0370_),
    .A1(net20),
    .A2(_1416_));
 sg13g2_a22oi_1 _3614_ (.Y(_1448_),
    .B1(net34),
    .B2(\madd.mem[7][11] ),
    .A2(_1439_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3615_ (.B1(_1448_),
    .Y(_0371_),
    .A1(_1125_),
    .A2(_1408_));
 sg13g2_nor2_1 _3616_ (.A(_0943_),
    .B(_1443_),
    .Y(_1449_));
 sg13g2_a221oi_1 _3617_ (.B2(\madd.mem[7][1] ),
    .C1(_1449_),
    .B1(net34),
    .A1(_0938_),
    .Y(_1450_),
    .A2(net48));
 sg13g2_inv_1 _3618_ (.Y(_0372_),
    .A(_1450_));
 sg13g2_nand2_1 _3619_ (.Y(_1451_),
    .A(_0951_),
    .B(_1414_));
 sg13g2_a22oi_1 _3620_ (.Y(_1452_),
    .B1(net34),
    .B2(\madd.mem[7][2] ),
    .A2(_1439_),
    .A1(_0956_));
 sg13g2_nand2_1 _3621_ (.Y(_0373_),
    .A(_1451_),
    .B(_1452_));
 sg13g2_a22oi_1 _3622_ (.Y(_1453_),
    .B1(net34),
    .B2(\madd.mem[7][3] ),
    .A2(_1439_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3623_ (.B1(_1453_),
    .Y(_0374_),
    .A1(_1132_),
    .A2(_1408_));
 sg13g2_nor2_1 _3624_ (.A(_0974_),
    .B(_1443_),
    .Y(_1454_));
 sg13g2_a221oi_1 _3625_ (.B2(\madd.mem[7][4] ),
    .C1(_1454_),
    .B1(_1441_),
    .A1(_0971_),
    .Y(_1455_),
    .A2(net48));
 sg13g2_inv_1 _3626_ (.Y(_0375_),
    .A(_1455_));
 sg13g2_nor2_1 _3627_ (.A(_0985_),
    .B(_1443_),
    .Y(_1456_));
 sg13g2_a221oi_1 _3628_ (.B2(\madd.mem[7][5] ),
    .C1(_1456_),
    .B1(_1441_),
    .A1(_0981_),
    .Y(_1457_),
    .A2(net48));
 sg13g2_inv_1 _3629_ (.Y(_0376_),
    .A(_1457_));
 sg13g2_nand2_1 _3630_ (.Y(_1458_),
    .A(\madd.mem[7][6] ),
    .B(_1440_));
 sg13g2_o21ai_1 _3631_ (.B1(_1458_),
    .Y(_1459_),
    .A1(_0994_),
    .A2(_1443_));
 sg13g2_a21o_1 _3632_ (.A2(net48),
    .A1(_0992_),
    .B1(_1459_),
    .X(_0377_));
 sg13g2_nor2_1 _3633_ (.A(_1004_),
    .B(_1443_),
    .Y(_1460_));
 sg13g2_a221oi_1 _3634_ (.B2(\madd.mem[7][7] ),
    .C1(_1460_),
    .B1(net34),
    .A1(_1001_),
    .Y(_1461_),
    .A2(net48));
 sg13g2_inv_1 _3635_ (.Y(_0378_),
    .A(_1461_));
 sg13g2_nand2_1 _3636_ (.Y(_1462_),
    .A(\madd.mem[7][8] ),
    .B(net34));
 sg13g2_a22oi_1 _3637_ (.Y(_1463_),
    .B1(_1439_),
    .B2(net28),
    .A2(_1410_),
    .A1(_1010_));
 sg13g2_nand2_1 _3638_ (.Y(_0379_),
    .A(_1462_),
    .B(_1463_));
 sg13g2_nand2_1 _3639_ (.Y(_1464_),
    .A(\madd.mem[7][9] ),
    .B(net34));
 sg13g2_a22oi_1 _3640_ (.Y(_1465_),
    .B1(_1439_),
    .B2(net27),
    .A2(_1410_),
    .A1(_1018_));
 sg13g2_nand2_1 _3641_ (.Y(_0380_),
    .A(_1464_),
    .B(_1465_));
 sg13g2_nor2_1 _3642_ (.A(_1025_),
    .B(_1078_),
    .Y(_1466_));
 sg13g2_buf_1 _3643_ (.A(_1466_),
    .X(_1467_));
 sg13g2_nand2_1 _3644_ (.Y(_1468_),
    .A(_2004_),
    .B(_1109_));
 sg13g2_nor2_1 _3645_ (.A(net94),
    .B(_1468_),
    .Y(_1469_));
 sg13g2_buf_2 _3646_ (.A(_1469_),
    .X(_1470_));
 sg13g2_nor3_1 _3647_ (.A(net132),
    .B(net80),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_buf_1 _3648_ (.A(_1471_),
    .X(_1472_));
 sg13g2_nor2_1 _3649_ (.A(net110),
    .B(_1115_),
    .Y(_1473_));
 sg13g2_buf_1 _3650_ (.A(_1473_),
    .X(_1474_));
 sg13g2_nand2_1 _3651_ (.Y(_1475_),
    .A(net95),
    .B(net53));
 sg13g2_buf_2 _3652_ (.A(_1475_),
    .X(_1476_));
 sg13g2_nor2_1 _3653_ (.A(_0715_),
    .B(_1476_),
    .Y(_1477_));
 sg13g2_a221oi_1 _3654_ (.B2(\madd.mem[8][0] ),
    .C1(_1477_),
    .B1(net41),
    .A1(_0677_),
    .Y(_1478_),
    .A2(net80));
 sg13g2_inv_1 _3655_ (.Y(_0381_),
    .A(_1478_));
 sg13g2_nor3_2 _3656_ (.A(_1025_),
    .B(_1078_),
    .C(net99),
    .Y(_1479_));
 sg13g2_nand2b_1 _3657_ (.Y(_1480_),
    .B(_1479_),
    .A_N(_0739_));
 sg13g2_nor2_1 _3658_ (.A(net26),
    .B(_1476_),
    .Y(_1481_));
 sg13g2_a21oi_1 _3659_ (.A1(\madd.mem[8][10] ),
    .A2(net41),
    .Y(_1482_),
    .B1(_1481_));
 sg13g2_nand2_1 _3660_ (.Y(_0382_),
    .A(_1480_),
    .B(_1482_));
 sg13g2_nand2_1 _3661_ (.Y(_1483_),
    .A(\madd.mem[8][11] ),
    .B(net41));
 sg13g2_a22oi_1 _3662_ (.Y(_1484_),
    .B1(_1479_),
    .B2(net24),
    .A2(_1470_),
    .A1(net23));
 sg13g2_nand2_1 _3663_ (.Y(_0383_),
    .A(_1483_),
    .B(_1484_));
 sg13g2_nor2_1 _3664_ (.A(_0943_),
    .B(_1476_),
    .Y(_1485_));
 sg13g2_a221oi_1 _3665_ (.B2(\madd.mem[8][1] ),
    .C1(_1485_),
    .B1(net41),
    .A1(_0938_),
    .Y(_1486_),
    .A2(net80));
 sg13g2_inv_1 _3666_ (.Y(_0384_),
    .A(_1486_));
 sg13g2_nand2_1 _3667_ (.Y(_1487_),
    .A(_0951_),
    .B(net80));
 sg13g2_a22oi_1 _3668_ (.Y(_1488_),
    .B1(net41),
    .B2(\madd.mem[8][2] ),
    .A2(_1470_),
    .A1(_0956_));
 sg13g2_nand2_1 _3669_ (.Y(_0385_),
    .A(_1487_),
    .B(_1488_));
 sg13g2_nand3_1 _3670_ (.B(net30),
    .C(net80),
    .A(net86),
    .Y(_1489_));
 sg13g2_a22oi_1 _3671_ (.Y(_1490_),
    .B1(_1472_),
    .B2(\madd.mem[8][3] ),
    .A2(_1470_),
    .A1(net59));
 sg13g2_nand2_1 _3672_ (.Y(_0386_),
    .A(_1489_),
    .B(_1490_));
 sg13g2_nor2_1 _3673_ (.A(_0974_),
    .B(_1476_),
    .Y(_1491_));
 sg13g2_a221oi_1 _3674_ (.B2(\madd.mem[8][4] ),
    .C1(_1491_),
    .B1(net41),
    .A1(_0971_),
    .Y(_1492_),
    .A2(net80));
 sg13g2_inv_1 _3675_ (.Y(_0387_),
    .A(_1492_));
 sg13g2_nor2_1 _3676_ (.A(_0985_),
    .B(_1476_),
    .Y(_1493_));
 sg13g2_a221oi_1 _3677_ (.B2(\madd.mem[8][5] ),
    .C1(_1493_),
    .B1(_1472_),
    .A1(_0981_),
    .Y(_1494_),
    .A2(_1467_));
 sg13g2_inv_1 _3678_ (.Y(_0388_),
    .A(_1494_));
 sg13g2_nand2_1 _3679_ (.Y(_1495_),
    .A(\madd.mem[8][6] ),
    .B(_1471_));
 sg13g2_o21ai_1 _3680_ (.B1(_1495_),
    .Y(_1496_),
    .A1(_0994_),
    .A2(_1476_));
 sg13g2_a21o_1 _3681_ (.A2(net80),
    .A1(_0992_),
    .B1(_1496_),
    .X(_0389_));
 sg13g2_nor2_1 _3682_ (.A(_1004_),
    .B(_1476_),
    .Y(_1497_));
 sg13g2_a221oi_1 _3683_ (.B2(\madd.mem[8][7] ),
    .C1(_1497_),
    .B1(_1471_),
    .A1(_1001_),
    .Y(_1498_),
    .A2(net80));
 sg13g2_inv_1 _3684_ (.Y(_0390_),
    .A(_1498_));
 sg13g2_nand2_1 _3685_ (.Y(_1499_),
    .A(\madd.mem[8][8] ),
    .B(net41));
 sg13g2_a22oi_1 _3686_ (.Y(_1500_),
    .B1(_1479_),
    .B2(net17),
    .A2(_1470_),
    .A1(_1013_));
 sg13g2_nand2_1 _3687_ (.Y(_0391_),
    .A(_1499_),
    .B(_1500_));
 sg13g2_nand2_1 _3688_ (.Y(_1501_),
    .A(\madd.mem[8][9] ),
    .B(net41));
 sg13g2_a22oi_1 _3689_ (.Y(_1502_),
    .B1(_1479_),
    .B2(net21),
    .A2(_1470_),
    .A1(_1020_));
 sg13g2_nand2_1 _3690_ (.Y(_0392_),
    .A(_1501_),
    .B(_1502_));
 sg13g2_nor3_2 _3691_ (.A(net110),
    .B(net94),
    .C(_0822_),
    .Y(_1503_));
 sg13g2_nor3_1 _3692_ (.A(net122),
    .B(net53),
    .C(_1503_),
    .Y(_1504_));
 sg13g2_buf_1 _3693_ (.A(_1504_),
    .X(_1505_));
 sg13g2_nand3_1 _3694_ (.B(net97),
    .C(net111),
    .A(_2004_),
    .Y(_1506_));
 sg13g2_buf_2 _3695_ (.A(_1506_),
    .X(_1507_));
 sg13g2_nor2_1 _3696_ (.A(_0715_),
    .B(_1507_),
    .Y(_1508_));
 sg13g2_a221oi_1 _3697_ (.B2(\madd.mem[9][0] ),
    .C1(_1508_),
    .B1(net40),
    .A1(_0677_),
    .Y(_1509_),
    .A2(net53));
 sg13g2_inv_1 _3698_ (.Y(_0393_),
    .A(_1509_));
 sg13g2_nor2_1 _3699_ (.A(_0913_),
    .B(_1507_),
    .Y(_1510_));
 sg13g2_a21oi_1 _3700_ (.A1(\madd.mem[9][10] ),
    .A2(_1504_),
    .Y(_1511_),
    .B1(_1510_));
 sg13g2_o21ai_1 _3701_ (.B1(_1511_),
    .Y(_0394_),
    .A1(_0739_),
    .A2(_1476_));
 sg13g2_a22oi_1 _3702_ (.Y(_1512_),
    .B1(net40),
    .B2(\madd.mem[9][11] ),
    .A2(_1503_),
    .A1(_0932_));
 sg13g2_o21ai_1 _3703_ (.B1(_1512_),
    .Y(_0395_),
    .A1(_1125_),
    .A2(_1468_));
 sg13g2_nor2_1 _3704_ (.A(_0943_),
    .B(_1507_),
    .Y(_1513_));
 sg13g2_a221oi_1 _3705_ (.B2(\madd.mem[9][1] ),
    .C1(_1513_),
    .B1(net40),
    .A1(_0938_),
    .Y(_1514_),
    .A2(net53));
 sg13g2_inv_1 _3706_ (.Y(_0396_),
    .A(_1514_));
 sg13g2_nand2_1 _3707_ (.Y(_1515_),
    .A(_0951_),
    .B(net53));
 sg13g2_a22oi_1 _3708_ (.Y(_1516_),
    .B1(net40),
    .B2(\madd.mem[9][2] ),
    .A2(_1503_),
    .A1(_0956_));
 sg13g2_nand2_1 _3709_ (.Y(_0397_),
    .A(_1515_),
    .B(_1516_));
 sg13g2_a22oi_1 _3710_ (.Y(_1517_),
    .B1(_1505_),
    .B2(\madd.mem[9][3] ),
    .A2(_1503_),
    .A1(_0966_));
 sg13g2_o21ai_1 _3711_ (.B1(_1517_),
    .Y(_0398_),
    .A1(_1132_),
    .A2(_1468_));
 sg13g2_nor2_1 _3712_ (.A(_0974_),
    .B(_1507_),
    .Y(_1518_));
 sg13g2_a221oi_1 _3713_ (.B2(\madd.mem[9][4] ),
    .C1(_1518_),
    .B1(net40),
    .A1(_0971_),
    .Y(_1519_),
    .A2(net53));
 sg13g2_inv_1 _3714_ (.Y(_0399_),
    .A(_1519_));
 sg13g2_nor2_1 _3715_ (.A(_0985_),
    .B(_1507_),
    .Y(_1520_));
 sg13g2_a221oi_1 _3716_ (.B2(\madd.mem[9][5] ),
    .C1(_1520_),
    .B1(_1505_),
    .A1(_0981_),
    .Y(_1521_),
    .A2(_1474_));
 sg13g2_inv_1 _3717_ (.Y(_0400_),
    .A(_1521_));
 sg13g2_nand2_1 _3718_ (.Y(_1522_),
    .A(\madd.mem[9][6] ),
    .B(_1504_));
 sg13g2_o21ai_1 _3719_ (.B1(_1522_),
    .Y(_1523_),
    .A1(_0994_),
    .A2(_1507_));
 sg13g2_a21o_1 _3720_ (.A2(net53),
    .A1(_0992_),
    .B1(_1523_),
    .X(_0401_));
 sg13g2_nor2_1 _3721_ (.A(_1004_),
    .B(_1507_),
    .Y(_1524_));
 sg13g2_a221oi_1 _3722_ (.B2(\madd.mem[9][7] ),
    .C1(_1524_),
    .B1(net40),
    .A1(_1001_),
    .Y(_1525_),
    .A2(net53));
 sg13g2_inv_1 _3723_ (.Y(_0402_),
    .A(_1525_));
 sg13g2_nand2_1 _3724_ (.Y(_1526_),
    .A(\madd.mem[9][8] ),
    .B(net40));
 sg13g2_a22oi_1 _3725_ (.Y(_1527_),
    .B1(_1503_),
    .B2(net28),
    .A2(_1470_),
    .A1(_1010_));
 sg13g2_nand2_1 _3726_ (.Y(_0403_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_nand2_1 _3727_ (.Y(_1528_),
    .A(\madd.mem[9][9] ),
    .B(net40));
 sg13g2_a22oi_1 _3728_ (.Y(_1529_),
    .B1(_1503_),
    .B2(net27),
    .A2(_1470_),
    .A1(_1018_));
 sg13g2_nand2_1 _3729_ (.Y(_0404_),
    .A(_1528_),
    .B(_1529_));
 sg13g2_inv_1 _3730_ (.Y(_1530_),
    .A(net8));
 sg13g2_buf_2 _3731_ (.A(_0002_),
    .X(_1531_));
 sg13g2_nor2_1 _3732_ (.A(\madd.mem[0][3] ),
    .B(\madd.mem[0][4] ),
    .Y(_1532_));
 sg13g2_buf_1 _3733_ (.A(_0000_),
    .X(_1533_));
 sg13g2_buf_1 _3734_ (.A(_1533_),
    .X(_1534_));
 sg13g2_nor4_1 _3735_ (.A(\madd.mem[0][0] ),
    .B(net119),
    .C(\madd.mem[0][1] ),
    .D(\madd.mem[0][2] ),
    .Y(_1535_));
 sg13g2_nor4_1 _3736_ (.A(\madd.mem[0][5] ),
    .B(\madd.mem[0][6] ),
    .C(\madd.mem[0][7] ),
    .D(\madd.mem[0][11] ),
    .Y(_1536_));
 sg13g2_nor3_1 _3737_ (.A(\madd.mem[0][8] ),
    .B(\madd.mem[0][9] ),
    .C(\madd.mem[0][10] ),
    .Y(_1537_));
 sg13g2_nand4_1 _3738_ (.B(_1535_),
    .C(_1536_),
    .A(_1532_),
    .Y(_1538_),
    .D(_1537_));
 sg13g2_nor2b_1 _3739_ (.A(\madd.mem[1][0] ),
    .B_N(net119),
    .Y(_1539_));
 sg13g2_nor4_1 _3740_ (.A(\madd.mem[1][1] ),
    .B(\madd.mem[1][2] ),
    .C(\madd.mem[1][3] ),
    .D(\madd.mem[1][4] ),
    .Y(_1540_));
 sg13g2_nor4_1 _3741_ (.A(\madd.mem[1][5] ),
    .B(\madd.mem[1][6] ),
    .C(\madd.mem[1][7] ),
    .D(\madd.mem[1][11] ),
    .Y(_1541_));
 sg13g2_nor3_1 _3742_ (.A(\madd.mem[1][8] ),
    .B(\madd.mem[1][9] ),
    .C(\madd.mem[1][10] ),
    .Y(_1542_));
 sg13g2_nand4_1 _3743_ (.B(_1540_),
    .C(_1541_),
    .A(_1539_),
    .Y(_1543_),
    .D(_1542_));
 sg13g2_nand2_1 _3744_ (.Y(_1544_),
    .A(_1538_),
    .B(_1543_));
 sg13g2_nor2b_1 _3745_ (.A(\madd.mem[5][0] ),
    .B_N(net119),
    .Y(_1545_));
 sg13g2_nor4_1 _3746_ (.A(\madd.mem[5][1] ),
    .B(\madd.mem[5][2] ),
    .C(\madd.mem[5][3] ),
    .D(\madd.mem[5][4] ),
    .Y(_1546_));
 sg13g2_nor4_1 _3747_ (.A(\madd.mem[5][5] ),
    .B(\madd.mem[5][6] ),
    .C(\madd.mem[5][7] ),
    .D(\madd.mem[5][11] ),
    .Y(_1547_));
 sg13g2_nor3_1 _3748_ (.A(\madd.mem[5][8] ),
    .B(\madd.mem[5][9] ),
    .C(\madd.mem[5][10] ),
    .Y(_1548_));
 sg13g2_nand4_1 _3749_ (.B(_1546_),
    .C(_1547_),
    .A(_1545_),
    .Y(_1549_),
    .D(_1548_));
 sg13g2_nor2_1 _3750_ (.A(\madd.mem[4][3] ),
    .B(\madd.mem[4][4] ),
    .Y(_1550_));
 sg13g2_nor4_1 _3751_ (.A(_1533_),
    .B(\madd.mem[4][0] ),
    .C(\madd.mem[4][1] ),
    .D(\madd.mem[4][2] ),
    .Y(_1551_));
 sg13g2_nor4_1 _3752_ (.A(\madd.mem[4][5] ),
    .B(\madd.mem[4][6] ),
    .C(\madd.mem[4][7] ),
    .D(\madd.mem[4][11] ),
    .Y(_1552_));
 sg13g2_nor3_1 _3753_ (.A(\madd.mem[4][8] ),
    .B(\madd.mem[4][9] ),
    .C(\madd.mem[4][10] ),
    .Y(_1553_));
 sg13g2_nand4_1 _3754_ (.B(_1551_),
    .C(_1552_),
    .A(_1550_),
    .Y(_1554_),
    .D(_1553_));
 sg13g2_nand3_1 _3755_ (.B(_1549_),
    .C(_1554_),
    .A(_1531_),
    .Y(_1555_));
 sg13g2_o21ai_1 _3756_ (.B1(_1555_),
    .Y(_1556_),
    .A1(_1531_),
    .A2(_1544_));
 sg13g2_nor2_1 _3757_ (.A(\madd.mem[6][3] ),
    .B(\madd.mem[6][4] ),
    .Y(_1557_));
 sg13g2_nor4_1 _3758_ (.A(net119),
    .B(\madd.mem[6][0] ),
    .C(\madd.mem[6][1] ),
    .D(\madd.mem[6][2] ),
    .Y(_1558_));
 sg13g2_nor4_1 _3759_ (.A(\madd.mem[6][5] ),
    .B(\madd.mem[6][6] ),
    .C(\madd.mem[6][7] ),
    .D(\madd.mem[6][11] ),
    .Y(_1559_));
 sg13g2_nor3_1 _3760_ (.A(\madd.mem[6][8] ),
    .B(\madd.mem[6][9] ),
    .C(\madd.mem[6][10] ),
    .Y(_1560_));
 sg13g2_nand4_1 _3761_ (.B(_1558_),
    .C(_1559_),
    .A(_1557_),
    .Y(_1561_),
    .D(_1560_));
 sg13g2_nor2b_1 _3762_ (.A(\madd.mem[7][0] ),
    .B_N(net119),
    .Y(_1562_));
 sg13g2_nor4_1 _3763_ (.A(\madd.mem[7][1] ),
    .B(\madd.mem[7][2] ),
    .C(\madd.mem[7][3] ),
    .D(\madd.mem[7][4] ),
    .Y(_1563_));
 sg13g2_nor4_1 _3764_ (.A(\madd.mem[7][5] ),
    .B(\madd.mem[7][6] ),
    .C(\madd.mem[7][7] ),
    .D(\madd.mem[7][11] ),
    .Y(_1564_));
 sg13g2_nor3_1 _3765_ (.A(\madd.mem[7][8] ),
    .B(\madd.mem[7][9] ),
    .C(\madd.mem[7][10] ),
    .Y(_1565_));
 sg13g2_nand4_1 _3766_ (.B(_1563_),
    .C(_1564_),
    .A(_1562_),
    .Y(_1566_),
    .D(_1565_));
 sg13g2_nand2_1 _3767_ (.Y(_1567_),
    .A(_1561_),
    .B(_1566_));
 sg13g2_nor2b_1 _3768_ (.A(\madd.mem[3][0] ),
    .B_N(net119),
    .Y(_1568_));
 sg13g2_nor4_1 _3769_ (.A(\madd.mem[3][1] ),
    .B(\madd.mem[3][2] ),
    .C(\madd.mem[3][3] ),
    .D(\madd.mem[3][4] ),
    .Y(_1569_));
 sg13g2_nor4_1 _3770_ (.A(\madd.mem[3][5] ),
    .B(\madd.mem[3][6] ),
    .C(\madd.mem[3][7] ),
    .D(\madd.mem[3][11] ),
    .Y(_1570_));
 sg13g2_nor3_1 _3771_ (.A(\madd.mem[3][8] ),
    .B(\madd.mem[3][9] ),
    .C(\madd.mem[3][10] ),
    .Y(_1571_));
 sg13g2_nand4_1 _3772_ (.B(_1569_),
    .C(_1570_),
    .A(_1568_),
    .Y(_1572_),
    .D(_1571_));
 sg13g2_nor2_1 _3773_ (.A(\madd.mem[2][3] ),
    .B(\madd.mem[2][4] ),
    .Y(_1573_));
 sg13g2_nor4_1 _3774_ (.A(_1533_),
    .B(\madd.mem[2][0] ),
    .C(\madd.mem[2][1] ),
    .D(\madd.mem[2][2] ),
    .Y(_1574_));
 sg13g2_nor4_1 _3775_ (.A(\madd.mem[2][5] ),
    .B(\madd.mem[2][6] ),
    .C(\madd.mem[2][7] ),
    .D(\madd.mem[2][11] ),
    .Y(_1575_));
 sg13g2_nor3_1 _3776_ (.A(\madd.mem[2][8] ),
    .B(\madd.mem[2][9] ),
    .C(\madd.mem[2][10] ),
    .Y(_1576_));
 sg13g2_nand4_1 _3777_ (.B(_1574_),
    .C(_1575_),
    .A(_1573_),
    .Y(_1577_),
    .D(_1576_));
 sg13g2_a21oi_1 _3778_ (.A1(_1572_),
    .A2(_1577_),
    .Y(_1578_),
    .B1(_1531_));
 sg13g2_a21oi_1 _3779_ (.A1(_1531_),
    .A2(_1567_),
    .Y(_1579_),
    .B1(_1578_));
 sg13g2_nor4_1 _3780_ (.A(\madd.mem[8][0] ),
    .B(\madd.mem[8][1] ),
    .C(\madd.mem[8][2] ),
    .D(\madd.mem[8][5] ),
    .Y(_1580_));
 sg13g2_nor4_1 _3781_ (.A(\madd.mem[8][3] ),
    .B(\madd.mem[8][4] ),
    .C(\madd.mem[8][6] ),
    .D(\madd.mem[8][11] ),
    .Y(_1581_));
 sg13g2_nor4_1 _3782_ (.A(\madd.mem[8][7] ),
    .B(\madd.mem[8][8] ),
    .C(\madd.mem[8][9] ),
    .D(\madd.mem[8][10] ),
    .Y(_1582_));
 sg13g2_nand3_1 _3783_ (.B(_1581_),
    .C(_1582_),
    .A(_1580_),
    .Y(_1583_));
 sg13g2_nor4_1 _3784_ (.A(\madd.mem[9][0] ),
    .B(\madd.mem[9][1] ),
    .C(\madd.mem[9][2] ),
    .D(\madd.mem[9][5] ),
    .Y(_1584_));
 sg13g2_nor4_1 _3785_ (.A(\madd.mem[9][3] ),
    .B(\madd.mem[9][4] ),
    .C(\madd.mem[9][6] ),
    .D(\madd.mem[9][11] ),
    .Y(_1585_));
 sg13g2_nor4_1 _3786_ (.A(\madd.mem[9][7] ),
    .B(\madd.mem[9][8] ),
    .C(\madd.mem[9][9] ),
    .D(\madd.mem[9][10] ),
    .Y(_1586_));
 sg13g2_nand3_1 _3787_ (.B(_1585_),
    .C(_1586_),
    .A(_1584_),
    .Y(_1587_));
 sg13g2_nor4_1 _3788_ (.A(\madd.mem[12][0] ),
    .B(\madd.mem[12][1] ),
    .C(\madd.mem[12][2] ),
    .D(\madd.mem[12][5] ),
    .Y(_1588_));
 sg13g2_nor4_1 _3789_ (.A(\madd.mem[12][3] ),
    .B(\madd.mem[12][4] ),
    .C(\madd.mem[12][6] ),
    .D(\madd.mem[12][11] ),
    .Y(_1589_));
 sg13g2_nor4_1 _3790_ (.A(\madd.mem[12][7] ),
    .B(\madd.mem[12][8] ),
    .C(\madd.mem[12][9] ),
    .D(\madd.mem[12][10] ),
    .Y(_1590_));
 sg13g2_nand3_1 _3791_ (.B(_1589_),
    .C(_1590_),
    .A(_1588_),
    .Y(_1591_));
 sg13g2_nor4_1 _3792_ (.A(\madd.mem[13][0] ),
    .B(\madd.mem[13][1] ),
    .C(\madd.mem[13][2] ),
    .D(\madd.mem[13][5] ),
    .Y(_1592_));
 sg13g2_nor4_1 _3793_ (.A(\madd.mem[13][3] ),
    .B(\madd.mem[13][4] ),
    .C(\madd.mem[13][6] ),
    .D(\madd.mem[13][11] ),
    .Y(_1593_));
 sg13g2_nor4_1 _3794_ (.A(\madd.mem[13][7] ),
    .B(\madd.mem[13][8] ),
    .C(\madd.mem[13][9] ),
    .D(\madd.mem[13][10] ),
    .Y(_1594_));
 sg13g2_nand3_1 _3795_ (.B(_1593_),
    .C(_1594_),
    .A(_1592_),
    .Y(_1595_));
 sg13g2_mux4_1 _3796_ (.S0(net119),
    .A0(_1583_),
    .A1(_1587_),
    .A2(_1591_),
    .A3(_1595_),
    .S1(_1531_),
    .X(_1596_));
 sg13g2_nor4_1 _3797_ (.A(\madd.mem[10][0] ),
    .B(\madd.mem[10][1] ),
    .C(\madd.mem[10][2] ),
    .D(\madd.mem[10][5] ),
    .Y(_1597_));
 sg13g2_nor4_1 _3798_ (.A(\madd.mem[10][3] ),
    .B(\madd.mem[10][4] ),
    .C(\madd.mem[10][6] ),
    .D(\madd.mem[10][11] ),
    .Y(_1598_));
 sg13g2_nor4_1 _3799_ (.A(\madd.mem[10][7] ),
    .B(\madd.mem[10][8] ),
    .C(\madd.mem[10][9] ),
    .D(\madd.mem[10][10] ),
    .Y(_1599_));
 sg13g2_nand3_1 _3800_ (.B(_1598_),
    .C(_1599_),
    .A(_1597_),
    .Y(_1600_));
 sg13g2_nor4_1 _3801_ (.A(\madd.mem[11][0] ),
    .B(\madd.mem[11][1] ),
    .C(\madd.mem[11][2] ),
    .D(\madd.mem[11][5] ),
    .Y(_1601_));
 sg13g2_nor4_1 _3802_ (.A(\madd.mem[11][3] ),
    .B(\madd.mem[11][4] ),
    .C(\madd.mem[11][6] ),
    .D(\madd.mem[11][11] ),
    .Y(_1602_));
 sg13g2_nor4_1 _3803_ (.A(\madd.mem[11][7] ),
    .B(\madd.mem[11][8] ),
    .C(\madd.mem[11][9] ),
    .D(\madd.mem[11][10] ),
    .Y(_1603_));
 sg13g2_nand4_1 _3804_ (.B(_1601_),
    .C(_1602_),
    .A(_1534_),
    .Y(_1604_),
    .D(_1603_));
 sg13g2_o21ai_1 _3805_ (.B1(_1604_),
    .Y(_1605_),
    .A1(_1534_),
    .A2(_1600_));
 sg13g2_nor2_1 _3806_ (.A(\madd.mem[14][3] ),
    .B(\madd.mem[14][4] ),
    .Y(_1606_));
 sg13g2_nor4_1 _3807_ (.A(_1533_),
    .B(\madd.mem[14][0] ),
    .C(\madd.mem[14][1] ),
    .D(\madd.mem[14][2] ),
    .Y(_1607_));
 sg13g2_nor4_1 _3808_ (.A(\madd.mem[14][5] ),
    .B(\madd.mem[14][6] ),
    .C(\madd.mem[14][7] ),
    .D(\madd.mem[14][11] ),
    .Y(_1608_));
 sg13g2_nor3_1 _3809_ (.A(\madd.mem[14][8] ),
    .B(\madd.mem[14][9] ),
    .C(\madd.mem[14][10] ),
    .Y(_1609_));
 sg13g2_nand4_1 _3810_ (.B(_1607_),
    .C(_1608_),
    .A(_1606_),
    .Y(_1610_),
    .D(_1609_));
 sg13g2_nor2b_1 _3811_ (.A(\madd.mem[15][0] ),
    .B_N(net119),
    .Y(_1611_));
 sg13g2_nor4_1 _3812_ (.A(\madd.mem[15][1] ),
    .B(\madd.mem[15][2] ),
    .C(\madd.mem[15][3] ),
    .D(\madd.mem[15][4] ),
    .Y(_1612_));
 sg13g2_nor4_1 _3813_ (.A(\madd.mem[15][5] ),
    .B(\madd.mem[15][6] ),
    .C(\madd.mem[15][7] ),
    .D(\madd.mem[15][11] ),
    .Y(_1613_));
 sg13g2_nor3_1 _3814_ (.A(\madd.mem[15][8] ),
    .B(\madd.mem[15][9] ),
    .C(\madd.mem[15][10] ),
    .Y(_1614_));
 sg13g2_nand4_1 _3815_ (.B(_1612_),
    .C(_1613_),
    .A(_1611_),
    .Y(_1615_),
    .D(_1614_));
 sg13g2_nand3_1 _3816_ (.B(_1610_),
    .C(_1615_),
    .A(_1531_),
    .Y(_1616_));
 sg13g2_o21ai_1 _3817_ (.B1(_1616_),
    .Y(_1617_),
    .A1(_1531_),
    .A2(_1605_));
 sg13g2_mux4_1 _3818_ (.S0(_0001_),
    .A0(_1556_),
    .A1(_1579_),
    .A2(_1596_),
    .A3(_1617_),
    .S1(_0003_),
    .X(_1618_));
 sg13g2_nor2_1 _3819_ (.A(net142),
    .B(\madd.set ),
    .Y(_1619_));
 sg13g2_nand2_1 _3820_ (.Y(_1620_),
    .A(_1618_),
    .B(_1619_));
 sg13g2_and4_1 _3821_ (.A(\madd.i_e[0] ),
    .B(net131),
    .C(net139),
    .D(_1784_),
    .X(_1621_));
 sg13g2_nor2_1 _3822_ (.A(\madd.i_e[0] ),
    .B(\madd.i[3] ),
    .Y(_1622_));
 sg13g2_a22oi_1 _3823_ (.Y(_1623_),
    .B1(_1622_),
    .B2(_2023_),
    .A2(_1621_),
    .A1(\madd.i[3] ));
 sg13g2_nand2b_1 _3824_ (.Y(_1624_),
    .B(net142),
    .A_N(_1623_));
 sg13g2_nand3_1 _3825_ (.B(_1620_),
    .C(_1624_),
    .A(net140),
    .Y(_1625_));
 sg13g2_buf_1 _3826_ (.A(_1625_),
    .X(_1626_));
 sg13g2_inv_1 _3827_ (.Y(_1627_),
    .A(_1620_));
 sg13g2_nor2b_1 _3828_ (.A(_1623_),
    .B_N(net142),
    .Y(_1628_));
 sg13g2_buf_2 _3829_ (.A(_1628_),
    .X(_1629_));
 sg13g2_buf_1 _3830_ (.A(\madd.total[0] ),
    .X(_1630_));
 sg13g2_xor2_1 _3831_ (.B(_1803_),
    .A(_1630_),
    .X(_1631_));
 sg13g2_a22oi_1 _3832_ (.Y(_1632_),
    .B1(_1629_),
    .B2(_1631_),
    .A2(net64),
    .A1(net131));
 sg13g2_o21ai_1 _3833_ (.B1(_1632_),
    .Y(_0405_),
    .A1(_1530_),
    .A2(_1626_));
 sg13g2_inv_1 _3834_ (.Y(_1633_),
    .A(net9));
 sg13g2_nand2_1 _3835_ (.Y(_1634_),
    .A(_1630_),
    .B(_1803_));
 sg13g2_buf_2 _3836_ (.A(\madd.total[1] ),
    .X(_1635_));
 sg13g2_xor2_1 _3837_ (.B(_1833_),
    .A(_1635_),
    .X(_1636_));
 sg13g2_xnor2_1 _3838_ (.Y(_1637_),
    .A(_1634_),
    .B(_1636_));
 sg13g2_a22oi_1 _3839_ (.Y(_1638_),
    .B1(_1629_),
    .B2(_1637_),
    .A2(net64),
    .A1(net139));
 sg13g2_o21ai_1 _3840_ (.B1(_1638_),
    .Y(_0408_),
    .A1(_1633_),
    .A2(_1626_));
 sg13g2_inv_1 _3841_ (.Y(_1639_),
    .A(net10));
 sg13g2_nor2_1 _3842_ (.A(_1635_),
    .B(_1833_),
    .Y(_1640_));
 sg13g2_a22oi_1 _3843_ (.Y(_1641_),
    .B1(_1635_),
    .B2(_1833_),
    .A2(_1803_),
    .A1(_1630_));
 sg13g2_nor2_1 _3844_ (.A(_1640_),
    .B(_1641_),
    .Y(_1642_));
 sg13g2_xnor2_1 _3845_ (.Y(_1643_),
    .A(\madd.total[2] ),
    .B(_1837_));
 sg13g2_xnor2_1 _3846_ (.Y(_1644_),
    .A(_1642_),
    .B(_1643_));
 sg13g2_a22oi_1 _3847_ (.Y(_1645_),
    .B1(_1629_),
    .B2(_1644_),
    .A2(net64),
    .A1(_1784_));
 sg13g2_o21ai_1 _3848_ (.B1(_1645_),
    .Y(_0409_),
    .A1(_1639_),
    .A2(_1626_));
 sg13g2_inv_1 _3849_ (.Y(_1646_),
    .A(net11));
 sg13g2_o21ai_1 _3850_ (.B1(_1840_),
    .Y(_1647_),
    .A1(_1640_),
    .A2(_1641_));
 sg13g2_nor3_1 _3851_ (.A(_1840_),
    .B(_1640_),
    .C(_1641_),
    .Y(_1648_));
 sg13g2_a21o_1 _3852_ (.A2(_1647_),
    .A1(\madd.total[2] ),
    .B1(_1648_),
    .X(_1649_));
 sg13g2_buf_1 _3853_ (.A(_1649_),
    .X(_1650_));
 sg13g2_xnor2_1 _3854_ (.Y(_1651_),
    .A(_1830_),
    .B(_1650_));
 sg13g2_xnor2_1 _3855_ (.Y(_1652_),
    .A(\madd.total[3] ),
    .B(_1651_));
 sg13g2_a22oi_1 _3856_ (.Y(_1653_),
    .B1(_1629_),
    .B2(_1652_),
    .A2(net64),
    .A1(\madd.i[3] ));
 sg13g2_o21ai_1 _3857_ (.B1(_1653_),
    .Y(_0410_),
    .A1(_1646_),
    .A2(_1626_));
 sg13g2_nand2_1 _3858_ (.Y(_1654_),
    .A(_1803_),
    .B(_1808_));
 sg13g2_xnor2_1 _3859_ (.Y(_1655_),
    .A(_1630_),
    .B(_1654_));
 sg13g2_and2_1 _3860_ (.A(_1802_),
    .B(_1655_),
    .X(_0418_));
 sg13g2_buf_2 _3861_ (.A(\madd.total[10] ),
    .X(_1656_));
 sg13g2_buf_1 _3862_ (.A(\madd.total[6] ),
    .X(_1657_));
 sg13g2_buf_1 _3863_ (.A(\madd.total[5] ),
    .X(_1658_));
 sg13g2_nor2_1 _3864_ (.A(_1658_),
    .B(_1827_),
    .Y(_1659_));
 sg13g2_inv_1 _3865_ (.Y(_1660_),
    .A(\madd.count[4] ));
 sg13g2_nand2_1 _3866_ (.Y(_1661_),
    .A(_1830_),
    .B(_1650_));
 sg13g2_o21ai_1 _3867_ (.B1(\madd.total[3] ),
    .Y(_1662_),
    .A1(_1830_),
    .A2(_1650_));
 sg13g2_nand3_1 _3868_ (.B(_1661_),
    .C(_1662_),
    .A(_1660_),
    .Y(_1663_));
 sg13g2_buf_1 _3869_ (.A(\madd.total[4] ),
    .X(_1664_));
 sg13g2_a21oi_1 _3870_ (.A1(_1661_),
    .A2(_1662_),
    .Y(_1665_),
    .B1(_1660_));
 sg13g2_a221oi_1 _3871_ (.B2(_1664_),
    .C1(_1665_),
    .B1(_1663_),
    .A1(_1658_),
    .Y(_1666_),
    .A2(_1827_));
 sg13g2_inv_1 _3872_ (.Y(_1667_),
    .A(\madd.count[6] ));
 sg13g2_o21ai_1 _3873_ (.B1(_1667_),
    .Y(_1668_),
    .A1(_1659_),
    .A2(_1666_));
 sg13g2_buf_1 _3874_ (.A(\madd.total[8] ),
    .X(_1669_));
 sg13g2_nand2_1 _3875_ (.Y(_1670_),
    .A(_1669_),
    .B(_1822_));
 sg13g2_nand2_1 _3876_ (.Y(_1671_),
    .A(_1890_),
    .B(_1670_));
 sg13g2_inv_1 _3877_ (.Y(_1672_),
    .A(\madd.total[7] ));
 sg13g2_nand2_1 _3878_ (.Y(_1673_),
    .A(_1672_),
    .B(_1670_));
 sg13g2_nor3_1 _3879_ (.A(_1667_),
    .B(_1659_),
    .C(_1666_),
    .Y(_1674_));
 sg13g2_a221oi_1 _3880_ (.B2(_1673_),
    .C1(_1674_),
    .B1(_1671_),
    .A1(_1657_),
    .Y(_1675_),
    .A2(_1668_));
 sg13g2_nand3_1 _3881_ (.B(_1890_),
    .C(_1670_),
    .A(_1672_),
    .Y(_1676_));
 sg13g2_o21ai_1 _3882_ (.B1(_1676_),
    .Y(_1677_),
    .A1(_1669_),
    .A2(_1822_));
 sg13g2_o21ai_1 _3883_ (.B1(_1899_),
    .Y(_1678_),
    .A1(_1675_),
    .A2(_1677_));
 sg13g2_nor3_1 _3884_ (.A(_1899_),
    .B(_1675_),
    .C(_1677_),
    .Y(_1679_));
 sg13g2_a21oi_1 _3885_ (.A1(\madd.total[9] ),
    .A2(_1678_),
    .Y(_1680_),
    .B1(_1679_));
 sg13g2_xor2_1 _3886_ (.B(_1680_),
    .A(net137),
    .X(_1681_));
 sg13g2_nor2_1 _3887_ (.A(net91),
    .B(_1681_),
    .Y(_1682_));
 sg13g2_xnor2_1 _3888_ (.Y(_1683_),
    .A(_1656_),
    .B(_1682_));
 sg13g2_nor2_1 _3889_ (.A(net106),
    .B(_1683_),
    .Y(_0419_));
 sg13g2_nand2b_1 _3890_ (.Y(_1684_),
    .B(net137),
    .A_N(_1862_));
 sg13g2_nand2b_1 _3891_ (.Y(_1685_),
    .B(_1656_),
    .A_N(_1862_));
 sg13g2_a21o_1 _3892_ (.A2(_1685_),
    .A1(_1684_),
    .B1(_1680_),
    .X(_1686_));
 sg13g2_nor2b_1 _3893_ (.A(net137),
    .B_N(_1862_),
    .Y(_1687_));
 sg13g2_nor2b_1 _3894_ (.A(_1656_),
    .B_N(_1862_),
    .Y(_1688_));
 sg13g2_o21ai_1 _3895_ (.B1(_1680_),
    .Y(_1689_),
    .A1(_1687_),
    .A2(_1688_));
 sg13g2_nand3b_1 _3896_ (.B(net137),
    .C(_1656_),
    .Y(_1690_),
    .A_N(_1862_));
 sg13g2_nor2_1 _3897_ (.A(_1656_),
    .B(net137),
    .Y(_1691_));
 sg13g2_nand2_1 _3898_ (.Y(_1692_),
    .A(_1862_),
    .B(_1691_));
 sg13g2_nand4_1 _3899_ (.B(_1689_),
    .C(_1690_),
    .A(_1686_),
    .Y(_1693_),
    .D(_1692_));
 sg13g2_nand2_1 _3900_ (.Y(_1694_),
    .A(net93),
    .B(_1693_));
 sg13g2_xor2_1 _3901_ (.B(_1694_),
    .A(\madd.total[11] ),
    .X(_1695_));
 sg13g2_nor2_1 _3902_ (.A(net106),
    .B(_1695_),
    .Y(_0420_));
 sg13g2_nand2_1 _3903_ (.Y(_1696_),
    .A(_1970_),
    .B(_1637_));
 sg13g2_nand3_1 _3904_ (.B(_1635_),
    .C(net92),
    .A(net130),
    .Y(_1697_));
 sg13g2_nand2_1 _3905_ (.Y(_0421_),
    .A(_1696_),
    .B(_1697_));
 sg13g2_nand2_1 _3906_ (.Y(_1698_),
    .A(_1970_),
    .B(_1644_));
 sg13g2_nand3_1 _3907_ (.B(\madd.total[2] ),
    .C(_1818_),
    .A(net130),
    .Y(_1699_));
 sg13g2_nand2_1 _3908_ (.Y(_0422_),
    .A(_1698_),
    .B(_1699_));
 sg13g2_nor2_1 _3909_ (.A(net91),
    .B(_1651_),
    .Y(_1700_));
 sg13g2_xnor2_1 _3910_ (.Y(_1701_),
    .A(\madd.total[3] ),
    .B(_1700_));
 sg13g2_nor2_1 _3911_ (.A(net117),
    .B(_1701_),
    .Y(_0423_));
 sg13g2_a21o_1 _3912_ (.A2(_1662_),
    .A1(_1661_),
    .B1(_1660_),
    .X(_1702_));
 sg13g2_nand2_1 _3913_ (.Y(_1703_),
    .A(_1663_),
    .B(_1702_));
 sg13g2_nor2_1 _3914_ (.A(net91),
    .B(_1703_),
    .Y(_1704_));
 sg13g2_xnor2_1 _3915_ (.Y(_1705_),
    .A(_1664_),
    .B(_1704_));
 sg13g2_nor2_1 _3916_ (.A(_1814_),
    .B(_1705_),
    .Y(_0424_));
 sg13g2_a21oi_1 _3917_ (.A1(_1664_),
    .A2(_1663_),
    .Y(_1706_),
    .B1(_1665_));
 sg13g2_xor2_1 _3918_ (.B(_1706_),
    .A(_1827_),
    .X(_1707_));
 sg13g2_nor2_1 _3919_ (.A(net91),
    .B(_1707_),
    .Y(_1708_));
 sg13g2_xnor2_1 _3920_ (.Y(_1709_),
    .A(_1658_),
    .B(_1708_));
 sg13g2_nor2_1 _3921_ (.A(_1814_),
    .B(_1709_),
    .Y(_0425_));
 sg13g2_or3_1 _3922_ (.A(_1667_),
    .B(_1659_),
    .C(_1666_),
    .X(_1710_));
 sg13g2_and2_1 _3923_ (.A(_1668_),
    .B(_1710_),
    .X(_1711_));
 sg13g2_nand2_1 _3924_ (.Y(_1712_),
    .A(net93),
    .B(_1711_));
 sg13g2_xor2_1 _3925_ (.B(_1712_),
    .A(_1657_),
    .X(_1713_));
 sg13g2_nor2_1 _3926_ (.A(net117),
    .B(_1713_),
    .Y(_0426_));
 sg13g2_a21oi_1 _3927_ (.A1(_1657_),
    .A2(_1668_),
    .Y(_1714_),
    .B1(_1674_));
 sg13g2_xnor2_1 _3928_ (.Y(_1715_),
    .A(_1890_),
    .B(_1714_));
 sg13g2_nor2_1 _3929_ (.A(net91),
    .B(_1715_),
    .Y(_1716_));
 sg13g2_xnor2_1 _3930_ (.Y(_1717_),
    .A(\madd.total[7] ),
    .B(_1716_));
 sg13g2_nor2_1 _3931_ (.A(net117),
    .B(_1717_),
    .Y(_0427_));
 sg13g2_o21ai_1 _3932_ (.B1(_1672_),
    .Y(_1718_),
    .A1(_1890_),
    .A2(_1714_));
 sg13g2_nand2_1 _3933_ (.Y(_1719_),
    .A(_1890_),
    .B(_1714_));
 sg13g2_nand2_1 _3934_ (.Y(_1720_),
    .A(_1718_),
    .B(_1719_));
 sg13g2_xor2_1 _3935_ (.B(_1822_),
    .A(_1669_),
    .X(_1721_));
 sg13g2_xnor2_1 _3936_ (.Y(_1722_),
    .A(_1720_),
    .B(_1721_));
 sg13g2_inv_1 _3937_ (.Y(_1723_),
    .A(_1722_));
 sg13g2_nand3_1 _3938_ (.B(_1669_),
    .C(net92),
    .A(net130),
    .Y(_1724_));
 sg13g2_o21ai_1 _3939_ (.B1(_1724_),
    .Y(_0428_),
    .A1(net90),
    .A2(_1723_));
 sg13g2_nor2_1 _3940_ (.A(_1675_),
    .B(_1677_),
    .Y(_1725_));
 sg13g2_xor2_1 _3941_ (.B(\madd.count[9] ),
    .A(\madd.total[9] ),
    .X(_1726_));
 sg13g2_xnor2_1 _3942_ (.Y(_1727_),
    .A(_1725_),
    .B(_1726_));
 sg13g2_nand3_1 _3943_ (.B(\madd.total[9] ),
    .C(net92),
    .A(net130),
    .Y(_1728_));
 sg13g2_o21ai_1 _3944_ (.B1(_1728_),
    .Y(_0429_),
    .A1(_1906_),
    .A2(_1727_));
 sg13g2_nor2_1 _3945_ (.A(net117),
    .B(_1762_),
    .Y(_1729_));
 sg13g2_nor3_1 _3946_ (.A(net64),
    .B(_1629_),
    .C(_1729_),
    .Y(_0211_));
 sg13g2_buf_1 _3947_ (.A(_1624_),
    .X(_1730_));
 sg13g2_xor2_1 _3948_ (.B(_1681_),
    .A(_1656_),
    .X(_1731_));
 sg13g2_inv_1 _3949_ (.Y(_1732_),
    .A(_1626_));
 sg13g2_nand2_1 _3950_ (.Y(_1733_),
    .A(net6),
    .B(_1732_));
 sg13g2_o21ai_1 _3951_ (.B1(_1733_),
    .Y(_0406_),
    .A1(net79),
    .A2(_1731_));
 sg13g2_xnor2_1 _3952_ (.Y(_1734_),
    .A(\madd.total[11] ),
    .B(_1693_));
 sg13g2_nand2_1 _3953_ (.Y(_1735_),
    .A(net7),
    .B(_1732_));
 sg13g2_o21ai_1 _3954_ (.B1(_1735_),
    .Y(_0407_),
    .A1(net79),
    .A2(_1734_));
 sg13g2_xor2_1 _3955_ (.B(_1703_),
    .A(_1664_),
    .X(_1736_));
 sg13g2_nand2_1 _3956_ (.Y(_1737_),
    .A(net12),
    .B(_1732_));
 sg13g2_o21ai_1 _3957_ (.B1(_1737_),
    .Y(_0411_),
    .A1(net79),
    .A2(_1736_));
 sg13g2_nand3_1 _3958_ (.B(net13),
    .C(net79),
    .A(net130),
    .Y(_1738_));
 sg13g2_xnor2_1 _3959_ (.Y(_1739_),
    .A(_1658_),
    .B(_1707_));
 sg13g2_nand2_1 _3960_ (.Y(_1740_),
    .A(_1629_),
    .B(_1739_));
 sg13g2_a21oi_1 _3961_ (.A1(_1738_),
    .A2(_1740_),
    .Y(_0412_),
    .B1(net64));
 sg13g2_xnor2_1 _3962_ (.Y(_1741_),
    .A(_1657_),
    .B(_1711_));
 sg13g2_nand3_1 _3963_ (.B(net14),
    .C(_1730_),
    .A(net140),
    .Y(_1742_));
 sg13g2_o21ai_1 _3964_ (.B1(_1742_),
    .Y(_1743_),
    .A1(_1730_),
    .A2(_1741_));
 sg13g2_and2_1 _3965_ (.A(_1620_),
    .B(_1743_),
    .X(_0413_));
 sg13g2_nand3_1 _3966_ (.B(net15),
    .C(net79),
    .A(net140),
    .Y(_1744_));
 sg13g2_xnor2_1 _3967_ (.Y(_1745_),
    .A(\madd.total[7] ),
    .B(_1715_));
 sg13g2_nand2_1 _3968_ (.Y(_1746_),
    .A(_1629_),
    .B(_1745_));
 sg13g2_a21oi_1 _3969_ (.A1(_1744_),
    .A2(_1746_),
    .Y(_0414_),
    .B1(net64));
 sg13g2_nand2_1 _3970_ (.Y(_1747_),
    .A(_1629_),
    .B(_1722_));
 sg13g2_nand3_1 _3971_ (.B(net4),
    .C(net79),
    .A(net140),
    .Y(_1748_));
 sg13g2_a21oi_1 _3972_ (.A1(_1747_),
    .A2(_1748_),
    .Y(_0415_),
    .B1(net64));
 sg13g2_nand3_1 _3973_ (.B(net5),
    .C(net79),
    .A(net140),
    .Y(_1749_));
 sg13g2_o21ai_1 _3974_ (.B1(_1749_),
    .Y(_1750_),
    .A1(net79),
    .A2(_1727_));
 sg13g2_and2_1 _3975_ (.A(_1620_),
    .B(_1750_),
    .X(_0416_));
 sg13g2_a21o_1 _3976_ (.A2(\madd.set ),
    .A1(net130),
    .B1(_1627_),
    .X(_0417_));
 sg13g2_dfrbp_1 _3977_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net151),
    .D(_0004_),
    .Q_N(_2112_),
    .Q(_0000_));
 sg13g2_dfrbp_1 _3978_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net152),
    .D(_0005_),
    .Q_N(_2113_),
    .Q(_0001_));
 sg13g2_dfrbp_1 _3979_ (.CLK(clknet_leaf_19_clk),
    .RESET_B(net153),
    .D(_0006_),
    .Q_N(_2114_),
    .Q(_0002_));
 sg13g2_dfrbp_1 _3980_ (.CLK(clknet_leaf_18_clk),
    .RESET_B(net154),
    .D(_0007_),
    .Q_N(_2111_),
    .Q(_0003_));
 sg13g2_buf_2 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sg13g2_tiehi _3977__151 (.L_HI(net151));
 sg13g2_buf_1 _3983_ (.A(net143),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3984_ (.A(net144),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3985_ (.A(net145),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3986_ (.A(net146),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3987_ (.A(net155),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3988_ (.A(net156),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3989_ (.A(net157),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3990_ (.A(net158),
    .X(uio_oe[7]));
 sg13g2_buf_1 _3991_ (.A(net147),
    .X(uio_out[0]));
 sg13g2_buf_1 _3992_ (.A(net148),
    .X(uio_out[1]));
 sg13g2_buf_1 _3993_ (.A(net149),
    .X(uio_out[2]));
 sg13g2_buf_1 _3994_ (.A(net150),
    .X(uio_out[3]));
 sg13g2_dfrbp_1 \madd.count[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net159),
    .D(_0187_),
    .Q_N(_2110_),
    .Q(\madd.count[0] ));
 sg13g2_dfrbp_1 \madd.count[10]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net160),
    .D(_0188_),
    .Q_N(_2109_),
    .Q(\madd.count[10] ));
 sg13g2_dfrbp_1 \madd.count[11]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net161),
    .D(_0189_),
    .Q_N(_2108_),
    .Q(\madd.count[11] ));
 sg13g2_dfrbp_1 \madd.count[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net162),
    .D(_0190_),
    .Q_N(_2107_),
    .Q(\madd.count[1] ));
 sg13g2_dfrbp_1 \madd.count[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net163),
    .D(_0191_),
    .Q_N(_2106_),
    .Q(\madd.count[2] ));
 sg13g2_dfrbp_1 \madd.count[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net164),
    .D(_0192_),
    .Q_N(_2105_),
    .Q(\madd.count[3] ));
 sg13g2_dfrbp_1 \madd.count[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net165),
    .D(_0193_),
    .Q_N(_2104_),
    .Q(\madd.count[4] ));
 sg13g2_dfrbp_1 \madd.count[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net166),
    .D(_0194_),
    .Q_N(_2103_),
    .Q(\madd.count[5] ));
 sg13g2_dfrbp_1 \madd.count[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net167),
    .D(_0195_),
    .Q_N(_2102_),
    .Q(\madd.count[6] ));
 sg13g2_dfrbp_1 \madd.count[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net168),
    .D(_0196_),
    .Q_N(_2101_),
    .Q(\madd.count[7] ));
 sg13g2_dfrbp_1 \madd.count[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net169),
    .D(_0197_),
    .Q_N(_2100_),
    .Q(\madd.count[8] ));
 sg13g2_dfrbp_1 \madd.count[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net170),
    .D(_0198_),
    .Q_N(_2099_),
    .Q(\madd.count[9] ));
 sg13g2_dfrbp_1 \madd.delta[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net171),
    .D(_0199_),
    .Q_N(_0152_),
    .Q(\madd.delta[0] ));
 sg13g2_dfrbp_1 \madd.delta[10]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net172),
    .D(_0200_),
    .Q_N(_2098_),
    .Q(\madd.delta[10] ));
 sg13g2_dfrbp_1 \madd.delta[11]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net173),
    .D(_0201_),
    .Q_N(_2097_),
    .Q(\madd.delta[11] ));
 sg13g2_dfrbp_1 \madd.delta[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net174),
    .D(_0202_),
    .Q_N(_2096_),
    .Q(\madd.delta[1] ));
 sg13g2_dfrbp_1 \madd.delta[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net175),
    .D(_0203_),
    .Q_N(_2095_),
    .Q(\madd.delta[2] ));
 sg13g2_dfrbp_1 \madd.delta[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net176),
    .D(_0204_),
    .Q_N(_2094_),
    .Q(\madd.delta[3] ));
 sg13g2_dfrbp_1 \madd.delta[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net177),
    .D(_0205_),
    .Q_N(_2093_),
    .Q(\madd.delta[4] ));
 sg13g2_dfrbp_1 \madd.delta[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net178),
    .D(_0206_),
    .Q_N(_2092_),
    .Q(\madd.delta[5] ));
 sg13g2_dfrbp_1 \madd.delta[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net179),
    .D(_0207_),
    .Q_N(_2091_),
    .Q(\madd.delta[6] ));
 sg13g2_dfrbp_1 \madd.delta[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net180),
    .D(_0208_),
    .Q_N(_2090_),
    .Q(\madd.delta[7] ));
 sg13g2_dfrbp_1 \madd.delta[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net181),
    .D(_0209_),
    .Q_N(_2089_),
    .Q(\madd.delta[8] ));
 sg13g2_dfrbp_1 \madd.delta[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net182),
    .D(_0210_),
    .Q_N(_2088_),
    .Q(\madd.delta[9] ));
 sg13g2_dfrbp_1 \madd.i[0]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net183),
    .D(_0004_),
    .Q_N(_2087_),
    .Q(\madd.i[0] ));
 sg13g2_dfrbp_1 \madd.i[1]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net184),
    .D(_0005_),
    .Q_N(_2086_),
    .Q(\madd.i[1] ));
 sg13g2_dfrbp_1 \madd.i[2]$_DFFE_PN_  (.CLK(clknet_leaf_19_clk),
    .RESET_B(net185),
    .D(_0006_),
    .Q_N(_0157_),
    .Q(\madd.i[2] ));
 sg13g2_dfrbp_1 \madd.i[3]$_DFFE_PN_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net186),
    .D(_0007_),
    .Q_N(_0162_),
    .Q(\madd.i[3] ));
 sg13g2_dfrbp_1 \madd.i_d[0]$_SDFFE_PP0N_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net187),
    .D(_0211_),
    .Q_N(_2085_),
    .Q(\madd.i_d[0] ));
 sg13g2_dfrbp_1 \madd.i_e[2]$_DFFE_PP_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net188),
    .D(_0212_),
    .Q_N(_2084_),
    .Q(\madd.i_e[0] ));
 sg13g2_dfrbp_1 \madd.mem[0][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net189),
    .D(_0213_),
    .Q_N(_0153_),
    .Q(\madd.mem[0][0] ));
 sg13g2_dfrbp_1 \madd.mem[0][10]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net190),
    .D(_0214_),
    .Q_N(_0136_),
    .Q(\madd.mem[0][10] ));
 sg13g2_dfrbp_1 \madd.mem[0][11]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net191),
    .D(_0215_),
    .Q_N(_2083_),
    .Q(\madd.mem[0][11] ));
 sg13g2_dfrbp_1 \madd.mem[0][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net192),
    .D(_0216_),
    .Q_N(_0171_),
    .Q(\madd.mem[0][1] ));
 sg13g2_dfrbp_1 \madd.mem[0][2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net193),
    .D(_0217_),
    .Q_N(_0008_),
    .Q(\madd.mem[0][2] ));
 sg13g2_dfrbp_1 \madd.mem[0][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net194),
    .D(_0218_),
    .Q_N(_0024_),
    .Q(\madd.mem[0][3] ));
 sg13g2_dfrbp_1 \madd.mem[0][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net195),
    .D(_0219_),
    .Q_N(_0040_),
    .Q(\madd.mem[0][4] ));
 sg13g2_dfrbp_1 \madd.mem[0][5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net196),
    .D(_0220_),
    .Q_N(_0056_),
    .Q(\madd.mem[0][5] ));
 sg13g2_dfrbp_1 \madd.mem[0][6]$_DFFE_PP_  (.CLK(clknet_leaf_12_clk),
    .RESET_B(net197),
    .D(_0221_),
    .Q_N(_0072_),
    .Q(\madd.mem[0][6] ));
 sg13g2_dfrbp_1 \madd.mem[0][7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net198),
    .D(_0222_),
    .Q_N(_0088_),
    .Q(\madd.mem[0][7] ));
 sg13g2_dfrbp_1 \madd.mem[0][8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net199),
    .D(_0223_),
    .Q_N(_0104_),
    .Q(\madd.mem[0][8] ));
 sg13g2_dfrbp_1 \madd.mem[0][9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net200),
    .D(_0224_),
    .Q_N(_0120_),
    .Q(\madd.mem[0][9] ));
 sg13g2_dfrbp_1 \madd.mem[10][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net201),
    .D(_0225_),
    .Q_N(_0165_),
    .Q(\madd.mem[10][0] ));
 sg13g2_dfrbp_1 \madd.mem[10][10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net202),
    .D(_0226_),
    .Q_N(_0146_),
    .Q(\madd.mem[10][10] ));
 sg13g2_dfrbp_1 \madd.mem[10][11]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net203),
    .D(_0227_),
    .Q_N(_2082_),
    .Q(\madd.mem[10][11] ));
 sg13g2_dfrbp_1 \madd.mem[10][1]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net204),
    .D(_0228_),
    .Q_N(_0181_),
    .Q(\madd.mem[10][1] ));
 sg13g2_dfrbp_1 \madd.mem[10][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net205),
    .D(_0229_),
    .Q_N(_0018_),
    .Q(\madd.mem[10][2] ));
 sg13g2_dfrbp_1 \madd.mem[10][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net206),
    .D(_0230_),
    .Q_N(_0034_),
    .Q(\madd.mem[10][3] ));
 sg13g2_dfrbp_1 \madd.mem[10][4]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net207),
    .D(_0231_),
    .Q_N(_0050_),
    .Q(\madd.mem[10][4] ));
 sg13g2_dfrbp_1 \madd.mem[10][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net208),
    .D(_0232_),
    .Q_N(_0066_),
    .Q(\madd.mem[10][5] ));
 sg13g2_dfrbp_1 \madd.mem[10][6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net209),
    .D(_0233_),
    .Q_N(_0082_),
    .Q(\madd.mem[10][6] ));
 sg13g2_dfrbp_1 \madd.mem[10][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net210),
    .D(_0234_),
    .Q_N(_0098_),
    .Q(\madd.mem[10][7] ));
 sg13g2_dfrbp_1 \madd.mem[10][8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net211),
    .D(_0235_),
    .Q_N(_0114_),
    .Q(\madd.mem[10][8] ));
 sg13g2_dfrbp_1 \madd.mem[10][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net212),
    .D(_0236_),
    .Q_N(_0130_),
    .Q(\madd.mem[10][9] ));
 sg13g2_dfrbp_1 \madd.mem[11][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net213),
    .D(_0237_),
    .Q_N(_0166_),
    .Q(\madd.mem[11][0] ));
 sg13g2_dfrbp_1 \madd.mem[11][10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net214),
    .D(_0238_),
    .Q_N(_0147_),
    .Q(\madd.mem[11][10] ));
 sg13g2_dfrbp_1 \madd.mem[11][11]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net215),
    .D(_0239_),
    .Q_N(_2081_),
    .Q(\madd.mem[11][11] ));
 sg13g2_dfrbp_1 \madd.mem[11][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net216),
    .D(_0240_),
    .Q_N(_0182_),
    .Q(\madd.mem[11][1] ));
 sg13g2_dfrbp_1 \madd.mem[11][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net217),
    .D(_0241_),
    .Q_N(_0019_),
    .Q(\madd.mem[11][2] ));
 sg13g2_dfrbp_1 \madd.mem[11][3]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net218),
    .D(_0242_),
    .Q_N(_0035_),
    .Q(\madd.mem[11][3] ));
 sg13g2_dfrbp_1 \madd.mem[11][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net219),
    .D(_0243_),
    .Q_N(_0051_),
    .Q(\madd.mem[11][4] ));
 sg13g2_dfrbp_1 \madd.mem[11][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net220),
    .D(_0244_),
    .Q_N(_0067_),
    .Q(\madd.mem[11][5] ));
 sg13g2_dfrbp_1 \madd.mem[11][6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net221),
    .D(_0245_),
    .Q_N(_0083_),
    .Q(\madd.mem[11][6] ));
 sg13g2_dfrbp_1 \madd.mem[11][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net222),
    .D(_0246_),
    .Q_N(_0099_),
    .Q(\madd.mem[11][7] ));
 sg13g2_dfrbp_1 \madd.mem[11][8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net223),
    .D(_0247_),
    .Q_N(_0115_),
    .Q(\madd.mem[11][8] ));
 sg13g2_dfrbp_1 \madd.mem[11][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net224),
    .D(_0248_),
    .Q_N(_0131_),
    .Q(\madd.mem[11][9] ));
 sg13g2_dfrbp_1 \madd.mem[12][0]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net225),
    .D(_0249_),
    .Q_N(_0167_),
    .Q(\madd.mem[12][0] ));
 sg13g2_dfrbp_1 \madd.mem[12][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net226),
    .D(_0250_),
    .Q_N(_0148_),
    .Q(\madd.mem[12][10] ));
 sg13g2_dfrbp_1 \madd.mem[12][11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net227),
    .D(_0251_),
    .Q_N(_2080_),
    .Q(\madd.mem[12][11] ));
 sg13g2_dfrbp_1 \madd.mem[12][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net228),
    .D(_0252_),
    .Q_N(_0183_),
    .Q(\madd.mem[12][1] ));
 sg13g2_dfrbp_1 \madd.mem[12][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net229),
    .D(_0253_),
    .Q_N(_0020_),
    .Q(\madd.mem[12][2] ));
 sg13g2_dfrbp_1 \madd.mem[12][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net230),
    .D(_0254_),
    .Q_N(_0036_),
    .Q(\madd.mem[12][3] ));
 sg13g2_dfrbp_1 \madd.mem[12][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net231),
    .D(_0255_),
    .Q_N(_0052_),
    .Q(\madd.mem[12][4] ));
 sg13g2_dfrbp_1 \madd.mem[12][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net232),
    .D(_0256_),
    .Q_N(_0068_),
    .Q(\madd.mem[12][5] ));
 sg13g2_dfrbp_1 \madd.mem[12][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net233),
    .D(_0257_),
    .Q_N(_0084_),
    .Q(\madd.mem[12][6] ));
 sg13g2_dfrbp_1 \madd.mem[12][7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net234),
    .D(_0258_),
    .Q_N(_0100_),
    .Q(\madd.mem[12][7] ));
 sg13g2_dfrbp_1 \madd.mem[12][8]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net235),
    .D(_0259_),
    .Q_N(_0116_),
    .Q(\madd.mem[12][8] ));
 sg13g2_dfrbp_1 \madd.mem[12][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net236),
    .D(_0260_),
    .Q_N(_0132_),
    .Q(\madd.mem[12][9] ));
 sg13g2_dfrbp_1 \madd.mem[13][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net237),
    .D(_0261_),
    .Q_N(_0168_),
    .Q(\madd.mem[13][0] ));
 sg13g2_dfrbp_1 \madd.mem[13][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net238),
    .D(_0262_),
    .Q_N(_0149_),
    .Q(\madd.mem[13][10] ));
 sg13g2_dfrbp_1 \madd.mem[13][11]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net239),
    .D(_0263_),
    .Q_N(_2079_),
    .Q(\madd.mem[13][11] ));
 sg13g2_dfrbp_1 \madd.mem[13][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net240),
    .D(_0264_),
    .Q_N(_0184_),
    .Q(\madd.mem[13][1] ));
 sg13g2_dfrbp_1 \madd.mem[13][2]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net241),
    .D(_0265_),
    .Q_N(_0021_),
    .Q(\madd.mem[13][2] ));
 sg13g2_dfrbp_1 \madd.mem[13][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net242),
    .D(_0266_),
    .Q_N(_0037_),
    .Q(\madd.mem[13][3] ));
 sg13g2_dfrbp_1 \madd.mem[13][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net243),
    .D(_0267_),
    .Q_N(_0053_),
    .Q(\madd.mem[13][4] ));
 sg13g2_dfrbp_1 \madd.mem[13][5]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net244),
    .D(_0268_),
    .Q_N(_0069_),
    .Q(\madd.mem[13][5] ));
 sg13g2_dfrbp_1 \madd.mem[13][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net245),
    .D(_0269_),
    .Q_N(_0085_),
    .Q(\madd.mem[13][6] ));
 sg13g2_dfrbp_1 \madd.mem[13][7]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net246),
    .D(_0270_),
    .Q_N(_0101_),
    .Q(\madd.mem[13][7] ));
 sg13g2_dfrbp_1 \madd.mem[13][8]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net247),
    .D(_0271_),
    .Q_N(_0117_),
    .Q(\madd.mem[13][8] ));
 sg13g2_dfrbp_1 \madd.mem[13][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net248),
    .D(_0272_),
    .Q_N(_0133_),
    .Q(\madd.mem[13][9] ));
 sg13g2_dfrbp_1 \madd.mem[14][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net249),
    .D(_0273_),
    .Q_N(_0169_),
    .Q(\madd.mem[14][0] ));
 sg13g2_dfrbp_1 \madd.mem[14][10]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net250),
    .D(_0274_),
    .Q_N(_0150_),
    .Q(\madd.mem[14][10] ));
 sg13g2_dfrbp_1 \madd.mem[14][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net251),
    .D(_0275_),
    .Q_N(_2078_),
    .Q(\madd.mem[14][11] ));
 sg13g2_dfrbp_1 \madd.mem[14][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net252),
    .D(_0276_),
    .Q_N(_0185_),
    .Q(\madd.mem[14][1] ));
 sg13g2_dfrbp_1 \madd.mem[14][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net253),
    .D(_0277_),
    .Q_N(_0022_),
    .Q(\madd.mem[14][2] ));
 sg13g2_dfrbp_1 \madd.mem[14][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net254),
    .D(_0278_),
    .Q_N(_0038_),
    .Q(\madd.mem[14][3] ));
 sg13g2_dfrbp_1 \madd.mem[14][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net255),
    .D(_0279_),
    .Q_N(_0054_),
    .Q(\madd.mem[14][4] ));
 sg13g2_dfrbp_1 \madd.mem[14][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net256),
    .D(_0280_),
    .Q_N(_0070_),
    .Q(\madd.mem[14][5] ));
 sg13g2_dfrbp_1 \madd.mem[14][6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net257),
    .D(_0281_),
    .Q_N(_0086_),
    .Q(\madd.mem[14][6] ));
 sg13g2_dfrbp_1 \madd.mem[14][7]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net258),
    .D(_0282_),
    .Q_N(_0102_),
    .Q(\madd.mem[14][7] ));
 sg13g2_dfrbp_1 \madd.mem[14][8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net259),
    .D(_0283_),
    .Q_N(_0118_),
    .Q(\madd.mem[14][8] ));
 sg13g2_dfrbp_1 \madd.mem[14][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net260),
    .D(_0284_),
    .Q_N(_0134_),
    .Q(\madd.mem[14][9] ));
 sg13g2_dfrbp_1 \madd.mem[15][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net261),
    .D(_0285_),
    .Q_N(_0170_),
    .Q(\madd.mem[15][0] ));
 sg13g2_dfrbp_1 \madd.mem[15][10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net262),
    .D(_0286_),
    .Q_N(_0151_),
    .Q(\madd.mem[15][10] ));
 sg13g2_dfrbp_1 \madd.mem[15][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net263),
    .D(_0287_),
    .Q_N(_2077_),
    .Q(\madd.mem[15][11] ));
 sg13g2_dfrbp_1 \madd.mem[15][1]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net264),
    .D(_0288_),
    .Q_N(_0186_),
    .Q(\madd.mem[15][1] ));
 sg13g2_dfrbp_1 \madd.mem[15][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net265),
    .D(_0289_),
    .Q_N(_0023_),
    .Q(\madd.mem[15][2] ));
 sg13g2_dfrbp_1 \madd.mem[15][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net266),
    .D(_0290_),
    .Q_N(_0039_),
    .Q(\madd.mem[15][3] ));
 sg13g2_dfrbp_1 \madd.mem[15][4]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net267),
    .D(_0291_),
    .Q_N(_0055_),
    .Q(\madd.mem[15][4] ));
 sg13g2_dfrbp_1 \madd.mem[15][5]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net268),
    .D(_0292_),
    .Q_N(_0071_),
    .Q(\madd.mem[15][5] ));
 sg13g2_dfrbp_1 \madd.mem[15][6]$_DFFE_PP_  (.CLK(clknet_leaf_32_clk),
    .RESET_B(net269),
    .D(_0293_),
    .Q_N(_0087_),
    .Q(\madd.mem[15][6] ));
 sg13g2_dfrbp_1 \madd.mem[15][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net270),
    .D(_0294_),
    .Q_N(_0103_),
    .Q(\madd.mem[15][7] ));
 sg13g2_dfrbp_1 \madd.mem[15][8]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net271),
    .D(_0295_),
    .Q_N(_0119_),
    .Q(\madd.mem[15][8] ));
 sg13g2_dfrbp_1 \madd.mem[15][9]$_DFFE_PP_  (.CLK(clknet_leaf_1_clk),
    .RESET_B(net272),
    .D(_0296_),
    .Q_N(_0135_),
    .Q(\madd.mem[15][9] ));
 sg13g2_dfrbp_1 \madd.mem[1][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net273),
    .D(_0297_),
    .Q_N(_0154_),
    .Q(\madd.mem[1][0] ));
 sg13g2_dfrbp_1 \madd.mem[1][10]$_DFFE_PP_  (.CLK(clknet_leaf_8_clk),
    .RESET_B(net274),
    .D(_0298_),
    .Q_N(_0137_),
    .Q(\madd.mem[1][10] ));
 sg13g2_dfrbp_1 \madd.mem[1][11]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net275),
    .D(_0299_),
    .Q_N(_2076_),
    .Q(\madd.mem[1][11] ));
 sg13g2_dfrbp_1 \madd.mem[1][1]$_DFFE_PP_  (.CLK(clknet_leaf_15_clk),
    .RESET_B(net276),
    .D(_0300_),
    .Q_N(_0172_),
    .Q(\madd.mem[1][1] ));
 sg13g2_dfrbp_1 \madd.mem[1][2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net277),
    .D(_0301_),
    .Q_N(_0009_),
    .Q(\madd.mem[1][2] ));
 sg13g2_dfrbp_1 \madd.mem[1][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net278),
    .D(_0302_),
    .Q_N(_0025_),
    .Q(\madd.mem[1][3] ));
 sg13g2_dfrbp_1 \madd.mem[1][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net279),
    .D(_0303_),
    .Q_N(_0041_),
    .Q(\madd.mem[1][4] ));
 sg13g2_dfrbp_1 \madd.mem[1][5]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net280),
    .D(_0304_),
    .Q_N(_0057_),
    .Q(\madd.mem[1][5] ));
 sg13g2_dfrbp_1 \madd.mem[1][6]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net281),
    .D(_0305_),
    .Q_N(_0073_),
    .Q(\madd.mem[1][6] ));
 sg13g2_dfrbp_1 \madd.mem[1][7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net282),
    .D(_0306_),
    .Q_N(_0089_),
    .Q(\madd.mem[1][7] ));
 sg13g2_dfrbp_1 \madd.mem[1][8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net283),
    .D(_0307_),
    .Q_N(_0105_),
    .Q(\madd.mem[1][8] ));
 sg13g2_dfrbp_1 \madd.mem[1][9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net284),
    .D(_0308_),
    .Q_N(_0121_),
    .Q(\madd.mem[1][9] ));
 sg13g2_dfrbp_1 \madd.mem[2][0]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net285),
    .D(_0309_),
    .Q_N(_0155_),
    .Q(\madd.mem[2][0] ));
 sg13g2_dfrbp_1 \madd.mem[2][10]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net286),
    .D(_0310_),
    .Q_N(_0138_),
    .Q(\madd.mem[2][10] ));
 sg13g2_dfrbp_1 \madd.mem[2][11]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net287),
    .D(_0311_),
    .Q_N(_2075_),
    .Q(\madd.mem[2][11] ));
 sg13g2_dfrbp_1 \madd.mem[2][1]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net288),
    .D(_0312_),
    .Q_N(_0173_),
    .Q(\madd.mem[2][1] ));
 sg13g2_dfrbp_1 \madd.mem[2][2]$_DFFE_PP_  (.CLK(clknet_leaf_20_clk),
    .RESET_B(net289),
    .D(_0313_),
    .Q_N(_0010_),
    .Q(\madd.mem[2][2] ));
 sg13g2_dfrbp_1 \madd.mem[2][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net290),
    .D(_0314_),
    .Q_N(_0026_),
    .Q(\madd.mem[2][3] ));
 sg13g2_dfrbp_1 \madd.mem[2][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net291),
    .D(_0315_),
    .Q_N(_0042_),
    .Q(\madd.mem[2][4] ));
 sg13g2_dfrbp_1 \madd.mem[2][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net292),
    .D(_0316_),
    .Q_N(_0058_),
    .Q(\madd.mem[2][5] ));
 sg13g2_dfrbp_1 \madd.mem[2][6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net293),
    .D(_0317_),
    .Q_N(_0074_),
    .Q(\madd.mem[2][6] ));
 sg13g2_dfrbp_1 \madd.mem[2][7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net294),
    .D(_0318_),
    .Q_N(_0090_),
    .Q(\madd.mem[2][7] ));
 sg13g2_dfrbp_1 \madd.mem[2][8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net295),
    .D(_0319_),
    .Q_N(_0106_),
    .Q(\madd.mem[2][8] ));
 sg13g2_dfrbp_1 \madd.mem[2][9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net296),
    .D(_0320_),
    .Q_N(_0122_),
    .Q(\madd.mem[2][9] ));
 sg13g2_dfrbp_1 \madd.mem[3][0]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net297),
    .D(_0321_),
    .Q_N(_0156_),
    .Q(\madd.mem[3][0] ));
 sg13g2_dfrbp_1 \madd.mem[3][10]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net298),
    .D(_0322_),
    .Q_N(_0139_),
    .Q(\madd.mem[3][10] ));
 sg13g2_dfrbp_1 \madd.mem[3][11]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net299),
    .D(_0323_),
    .Q_N(_2074_),
    .Q(\madd.mem[3][11] ));
 sg13g2_dfrbp_1 \madd.mem[3][1]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net300),
    .D(_0324_),
    .Q_N(_0174_),
    .Q(\madd.mem[3][1] ));
 sg13g2_dfrbp_1 \madd.mem[3][2]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net301),
    .D(_0325_),
    .Q_N(_0011_),
    .Q(\madd.mem[3][2] ));
 sg13g2_dfrbp_1 \madd.mem[3][3]$_DFFE_PP_  (.CLK(clknet_leaf_14_clk),
    .RESET_B(net302),
    .D(_0326_),
    .Q_N(_0027_),
    .Q(\madd.mem[3][3] ));
 sg13g2_dfrbp_1 \madd.mem[3][4]$_DFFE_PP_  (.CLK(clknet_leaf_13_clk),
    .RESET_B(net303),
    .D(_0327_),
    .Q_N(_0043_),
    .Q(\madd.mem[3][4] ));
 sg13g2_dfrbp_1 \madd.mem[3][5]$_DFFE_PP_  (.CLK(clknet_leaf_21_clk),
    .RESET_B(net304),
    .D(_0328_),
    .Q_N(_0059_),
    .Q(\madd.mem[3][5] ));
 sg13g2_dfrbp_1 \madd.mem[3][6]$_DFFE_PP_  (.CLK(clknet_leaf_5_clk),
    .RESET_B(net305),
    .D(_0329_),
    .Q_N(_0075_),
    .Q(\madd.mem[3][6] ));
 sg13g2_dfrbp_1 \madd.mem[3][7]$_DFFE_PP_  (.CLK(clknet_leaf_6_clk),
    .RESET_B(net306),
    .D(_0330_),
    .Q_N(_0091_),
    .Q(\madd.mem[3][7] ));
 sg13g2_dfrbp_1 \madd.mem[3][8]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net307),
    .D(_0331_),
    .Q_N(_0107_),
    .Q(\madd.mem[3][8] ));
 sg13g2_dfrbp_1 \madd.mem[3][9]$_DFFE_PP_  (.CLK(clknet_leaf_7_clk),
    .RESET_B(net308),
    .D(_0332_),
    .Q_N(_0123_),
    .Q(\madd.mem[3][9] ));
 sg13g2_dfrbp_1 \madd.mem[4][0]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net309),
    .D(_0333_),
    .Q_N(_0158_),
    .Q(\madd.mem[4][0] ));
 sg13g2_dfrbp_1 \madd.mem[4][10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net310),
    .D(_0334_),
    .Q_N(_0140_),
    .Q(\madd.mem[4][10] ));
 sg13g2_dfrbp_1 \madd.mem[4][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net311),
    .D(_0335_),
    .Q_N(_2073_),
    .Q(\madd.mem[4][11] ));
 sg13g2_dfrbp_1 \madd.mem[4][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net312),
    .D(_0336_),
    .Q_N(_0175_),
    .Q(\madd.mem[4][1] ));
 sg13g2_dfrbp_1 \madd.mem[4][2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net313),
    .D(_0337_),
    .Q_N(_0012_),
    .Q(\madd.mem[4][2] ));
 sg13g2_dfrbp_1 \madd.mem[4][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net314),
    .D(_0338_),
    .Q_N(_0028_),
    .Q(\madd.mem[4][3] ));
 sg13g2_dfrbp_1 \madd.mem[4][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net315),
    .D(_0339_),
    .Q_N(_0044_),
    .Q(\madd.mem[4][4] ));
 sg13g2_dfrbp_1 \madd.mem[4][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net316),
    .D(_0340_),
    .Q_N(_0060_),
    .Q(\madd.mem[4][5] ));
 sg13g2_dfrbp_1 \madd.mem[4][6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net317),
    .D(_0341_),
    .Q_N(_0076_),
    .Q(\madd.mem[4][6] ));
 sg13g2_dfrbp_1 \madd.mem[4][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net318),
    .D(_0342_),
    .Q_N(_0092_),
    .Q(\madd.mem[4][7] ));
 sg13g2_dfrbp_1 \madd.mem[4][8]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net319),
    .D(_0343_),
    .Q_N(_0108_),
    .Q(\madd.mem[4][8] ));
 sg13g2_dfrbp_1 \madd.mem[4][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net320),
    .D(_0344_),
    .Q_N(_0124_),
    .Q(\madd.mem[4][9] ));
 sg13g2_dfrbp_1 \madd.mem[5][0]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net321),
    .D(_0345_),
    .Q_N(_0159_),
    .Q(\madd.mem[5][0] ));
 sg13g2_dfrbp_1 \madd.mem[5][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net322),
    .D(_0346_),
    .Q_N(_0141_),
    .Q(\madd.mem[5][10] ));
 sg13g2_dfrbp_1 \madd.mem[5][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net323),
    .D(_0347_),
    .Q_N(_2072_),
    .Q(\madd.mem[5][11] ));
 sg13g2_dfrbp_1 \madd.mem[5][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net324),
    .D(_0348_),
    .Q_N(_0176_),
    .Q(\madd.mem[5][1] ));
 sg13g2_dfrbp_1 \madd.mem[5][2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net325),
    .D(_0349_),
    .Q_N(_0013_),
    .Q(\madd.mem[5][2] ));
 sg13g2_dfrbp_1 \madd.mem[5][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net326),
    .D(_0350_),
    .Q_N(_0029_),
    .Q(\madd.mem[5][3] ));
 sg13g2_dfrbp_1 \madd.mem[5][4]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net327),
    .D(_0351_),
    .Q_N(_0045_),
    .Q(\madd.mem[5][4] ));
 sg13g2_dfrbp_1 \madd.mem[5][5]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net328),
    .D(_0352_),
    .Q_N(_0061_),
    .Q(\madd.mem[5][5] ));
 sg13g2_dfrbp_1 \madd.mem[5][6]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net329),
    .D(_0353_),
    .Q_N(_0077_),
    .Q(\madd.mem[5][6] ));
 sg13g2_dfrbp_1 \madd.mem[5][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net330),
    .D(_0354_),
    .Q_N(_0093_),
    .Q(\madd.mem[5][7] ));
 sg13g2_dfrbp_1 \madd.mem[5][8]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net331),
    .D(_0355_),
    .Q_N(_0109_),
    .Q(\madd.mem[5][8] ));
 sg13g2_dfrbp_1 \madd.mem[5][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net332),
    .D(_0356_),
    .Q_N(_0125_),
    .Q(\madd.mem[5][9] ));
 sg13g2_dfrbp_1 \madd.mem[6][0]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net333),
    .D(_0357_),
    .Q_N(_0160_),
    .Q(\madd.mem[6][0] ));
 sg13g2_dfrbp_1 \madd.mem[6][10]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net334),
    .D(_0358_),
    .Q_N(_0142_),
    .Q(\madd.mem[6][10] ));
 sg13g2_dfrbp_1 \madd.mem[6][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net335),
    .D(_0359_),
    .Q_N(_2071_),
    .Q(\madd.mem[6][11] ));
 sg13g2_dfrbp_1 \madd.mem[6][1]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net336),
    .D(_0360_),
    .Q_N(_0177_),
    .Q(\madd.mem[6][1] ));
 sg13g2_dfrbp_1 \madd.mem[6][2]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net337),
    .D(_0361_),
    .Q_N(_0014_),
    .Q(\madd.mem[6][2] ));
 sg13g2_dfrbp_1 \madd.mem[6][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net338),
    .D(_0362_),
    .Q_N(_0030_),
    .Q(\madd.mem[6][3] ));
 sg13g2_dfrbp_1 \madd.mem[6][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net339),
    .D(_0363_),
    .Q_N(_0046_),
    .Q(\madd.mem[6][4] ));
 sg13g2_dfrbp_1 \madd.mem[6][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net340),
    .D(_0364_),
    .Q_N(_0062_),
    .Q(\madd.mem[6][5] ));
 sg13g2_dfrbp_1 \madd.mem[6][6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net341),
    .D(_0365_),
    .Q_N(_0078_),
    .Q(\madd.mem[6][6] ));
 sg13g2_dfrbp_1 \madd.mem[6][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net342),
    .D(_0366_),
    .Q_N(_0094_),
    .Q(\madd.mem[6][7] ));
 sg13g2_dfrbp_1 \madd.mem[6][8]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net343),
    .D(_0367_),
    .Q_N(_0110_),
    .Q(\madd.mem[6][8] ));
 sg13g2_dfrbp_1 \madd.mem[6][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net344),
    .D(_0368_),
    .Q_N(_0126_),
    .Q(\madd.mem[6][9] ));
 sg13g2_dfrbp_1 \madd.mem[7][0]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net345),
    .D(_0369_),
    .Q_N(_0161_),
    .Q(\madd.mem[7][0] ));
 sg13g2_dfrbp_1 \madd.mem[7][10]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net346),
    .D(_0370_),
    .Q_N(_0143_),
    .Q(\madd.mem[7][10] ));
 sg13g2_dfrbp_1 \madd.mem[7][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net347),
    .D(_0371_),
    .Q_N(_2070_),
    .Q(\madd.mem[7][11] ));
 sg13g2_dfrbp_1 \madd.mem[7][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net348),
    .D(_0372_),
    .Q_N(_0178_),
    .Q(\madd.mem[7][1] ));
 sg13g2_dfrbp_1 \madd.mem[7][2]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net349),
    .D(_0373_),
    .Q_N(_0015_),
    .Q(\madd.mem[7][2] ));
 sg13g2_dfrbp_1 \madd.mem[7][3]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net350),
    .D(_0374_),
    .Q_N(_0031_),
    .Q(\madd.mem[7][3] ));
 sg13g2_dfrbp_1 \madd.mem[7][4]$_DFFE_PP_  (.CLK(clknet_leaf_28_clk),
    .RESET_B(net351),
    .D(_0375_),
    .Q_N(_0047_),
    .Q(\madd.mem[7][4] ));
 sg13g2_dfrbp_1 \madd.mem[7][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net352),
    .D(_0376_),
    .Q_N(_0063_),
    .Q(\madd.mem[7][5] ));
 sg13g2_dfrbp_1 \madd.mem[7][6]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net353),
    .D(_0377_),
    .Q_N(_0079_),
    .Q(\madd.mem[7][6] ));
 sg13g2_dfrbp_1 \madd.mem[7][7]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net354),
    .D(_0378_),
    .Q_N(_0095_),
    .Q(\madd.mem[7][7] ));
 sg13g2_dfrbp_1 \madd.mem[7][8]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net355),
    .D(_0379_),
    .Q_N(_0111_),
    .Q(\madd.mem[7][8] ));
 sg13g2_dfrbp_1 \madd.mem[7][9]$_DFFE_PP_  (.CLK(clknet_leaf_36_clk),
    .RESET_B(net356),
    .D(_0380_),
    .Q_N(_0127_),
    .Q(\madd.mem[7][9] ));
 sg13g2_dfrbp_1 \madd.mem[8][0]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net357),
    .D(_0381_),
    .Q_N(_0163_),
    .Q(\madd.mem[8][0] ));
 sg13g2_dfrbp_1 \madd.mem[8][10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net358),
    .D(_0382_),
    .Q_N(_0144_),
    .Q(\madd.mem[8][10] ));
 sg13g2_dfrbp_1 \madd.mem[8][11]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net359),
    .D(_0383_),
    .Q_N(_2069_),
    .Q(\madd.mem[8][11] ));
 sg13g2_dfrbp_1 \madd.mem[8][1]$_DFFE_PP_  (.CLK(clknet_leaf_23_clk),
    .RESET_B(net360),
    .D(_0384_),
    .Q_N(_0179_),
    .Q(\madd.mem[8][1] ));
 sg13g2_dfrbp_1 \madd.mem[8][2]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net361),
    .D(_0385_),
    .Q_N(_0016_),
    .Q(\madd.mem[8][2] ));
 sg13g2_dfrbp_1 \madd.mem[8][3]$_DFFE_PP_  (.CLK(clknet_leaf_30_clk),
    .RESET_B(net362),
    .D(_0386_),
    .Q_N(_0032_),
    .Q(\madd.mem[8][3] ));
 sg13g2_dfrbp_1 \madd.mem[8][4]$_DFFE_PP_  (.CLK(clknet_leaf_31_clk),
    .RESET_B(net363),
    .D(_0387_),
    .Q_N(_0048_),
    .Q(\madd.mem[8][4] ));
 sg13g2_dfrbp_1 \madd.mem[8][5]$_DFFE_PP_  (.CLK(clknet_leaf_22_clk),
    .RESET_B(net364),
    .D(_0388_),
    .Q_N(_0064_),
    .Q(\madd.mem[8][5] ));
 sg13g2_dfrbp_1 \madd.mem[8][6]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net365),
    .D(_0389_),
    .Q_N(_0080_),
    .Q(\madd.mem[8][6] ));
 sg13g2_dfrbp_1 \madd.mem[8][7]$_DFFE_PP_  (.CLK(clknet_leaf_4_clk),
    .RESET_B(net366),
    .D(_0390_),
    .Q_N(_0096_),
    .Q(\madd.mem[8][7] ));
 sg13g2_dfrbp_1 \madd.mem[8][8]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net367),
    .D(_0391_),
    .Q_N(_0112_),
    .Q(\madd.mem[8][8] ));
 sg13g2_dfrbp_1 \madd.mem[8][9]$_DFFE_PP_  (.CLK(clknet_leaf_2_clk),
    .RESET_B(net368),
    .D(_0392_),
    .Q_N(_0128_),
    .Q(\madd.mem[8][9] ));
 sg13g2_dfrbp_1 \madd.mem[9][0]$_DFFE_PP_  (.CLK(clknet_leaf_24_clk),
    .RESET_B(net369),
    .D(_0393_),
    .Q_N(_0164_),
    .Q(\madd.mem[9][0] ));
 sg13g2_dfrbp_1 \madd.mem[9][10]$_DFFE_PP_  (.CLK(clknet_leaf_3_clk),
    .RESET_B(net370),
    .D(_0394_),
    .Q_N(_0145_),
    .Q(\madd.mem[9][10] ));
 sg13g2_dfrbp_1 \madd.mem[9][11]$_DFFE_PP_  (.CLK(clknet_leaf_33_clk),
    .RESET_B(net371),
    .D(_0395_),
    .Q_N(_2068_),
    .Q(\madd.mem[9][11] ));
 sg13g2_dfrbp_1 \madd.mem[9][1]$_DFFE_PP_  (.CLK(clknet_leaf_25_clk),
    .RESET_B(net372),
    .D(_0396_),
    .Q_N(_0180_),
    .Q(\madd.mem[9][1] ));
 sg13g2_dfrbp_1 \madd.mem[9][2]$_DFFE_PP_  (.CLK(clknet_leaf_26_clk),
    .RESET_B(net373),
    .D(_0397_),
    .Q_N(_0017_),
    .Q(\madd.mem[9][2] ));
 sg13g2_dfrbp_1 \madd.mem[9][3]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net374),
    .D(_0398_),
    .Q_N(_0033_),
    .Q(\madd.mem[9][3] ));
 sg13g2_dfrbp_1 \madd.mem[9][4]$_DFFE_PP_  (.CLK(clknet_leaf_29_clk),
    .RESET_B(net375),
    .D(_0399_),
    .Q_N(_0049_),
    .Q(\madd.mem[9][4] ));
 sg13g2_dfrbp_1 \madd.mem[9][5]$_DFFE_PP_  (.CLK(clknet_leaf_27_clk),
    .RESET_B(net376),
    .D(_0400_),
    .Q_N(_0065_),
    .Q(\madd.mem[9][5] ));
 sg13g2_dfrbp_1 \madd.mem[9][6]$_DFFE_PP_  (.CLK(clknet_leaf_34_clk),
    .RESET_B(net377),
    .D(_0401_),
    .Q_N(_0081_),
    .Q(\madd.mem[9][6] ));
 sg13g2_dfrbp_1 \madd.mem[9][7]$_DFFE_PP_  (.CLK(clknet_leaf_35_clk),
    .RESET_B(net378),
    .D(_0402_),
    .Q_N(_0097_),
    .Q(\madd.mem[9][7] ));
 sg13g2_dfrbp_1 \madd.mem[9][8]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net379),
    .D(_0403_),
    .Q_N(_0113_),
    .Q(\madd.mem[9][8] ));
 sg13g2_dfrbp_1 \madd.mem[9][9]$_DFFE_PP_  (.CLK(clknet_leaf_0_clk),
    .RESET_B(net380),
    .D(_0404_),
    .Q_N(_0129_),
    .Q(\madd.mem[9][9] ));
 sg13g2_dfrbp_1 \madd.out_reg[0]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net381),
    .D(_0405_),
    .Q_N(_2067_),
    .Q(net8));
 sg13g2_dfrbp_1 \madd.out_reg[10]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net382),
    .D(_0406_),
    .Q_N(_2066_),
    .Q(net6));
 sg13g2_dfrbp_1 \madd.out_reg[11]$_SDFFE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net383),
    .D(_0407_),
    .Q_N(_2065_),
    .Q(net7));
 sg13g2_dfrbp_1 \madd.out_reg[1]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net384),
    .D(_0408_),
    .Q_N(_2064_),
    .Q(net9));
 sg13g2_dfrbp_1 \madd.out_reg[2]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net385),
    .D(_0409_),
    .Q_N(_2063_),
    .Q(net10));
 sg13g2_dfrbp_1 \madd.out_reg[3]$_DFFE_PP_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net386),
    .D(_0410_),
    .Q_N(_2062_),
    .Q(net11));
 sg13g2_dfrbp_1 \madd.out_reg[4]$_SDFFE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net387),
    .D(_0411_),
    .Q_N(_2061_),
    .Q(net12));
 sg13g2_dfrbp_1 \madd.out_reg[5]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net388),
    .D(_0412_),
    .Q_N(_2060_),
    .Q(net13));
 sg13g2_dfrbp_1 \madd.out_reg[6]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net389),
    .D(_0413_),
    .Q_N(_2059_),
    .Q(net14));
 sg13g2_dfrbp_1 \madd.out_reg[7]$_SDFFE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net390),
    .D(_0414_),
    .Q_N(_2058_),
    .Q(net15));
 sg13g2_dfrbp_1 \madd.out_reg[8]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net391),
    .D(_0415_),
    .Q_N(_2057_),
    .Q(net4));
 sg13g2_dfrbp_1 \madd.out_reg[9]$_SDFFE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net392),
    .D(_0416_),
    .Q_N(_2056_),
    .Q(net5));
 sg13g2_dfrbp_1 \madd.set$_SDFFE_PP1N_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net393),
    .D(_0417_),
    .Q_N(_2055_),
    .Q(\madd.set ));
 sg13g2_dfrbp_1 \madd.total[0]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_17_clk),
    .RESET_B(net394),
    .D(_0418_),
    .Q_N(_2054_),
    .Q(\madd.total[0] ));
 sg13g2_dfrbp_1 \madd.total[10]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net395),
    .D(_0419_),
    .Q_N(_2053_),
    .Q(\madd.total[10] ));
 sg13g2_dfrbp_1 \madd.total[11]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net396),
    .D(_0420_),
    .Q_N(_2052_),
    .Q(\madd.total[11] ));
 sg13g2_dfrbp_1 \madd.total[1]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net397),
    .D(_0421_),
    .Q_N(_2051_),
    .Q(\madd.total[1] ));
 sg13g2_dfrbp_1 \madd.total[2]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_18_clk),
    .RESET_B(net398),
    .D(_0422_),
    .Q_N(_2050_),
    .Q(\madd.total[2] ));
 sg13g2_dfrbp_1 \madd.total[3]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net399),
    .D(_0423_),
    .Q_N(_2049_),
    .Q(\madd.total[3] ));
 sg13g2_dfrbp_1 \madd.total[4]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_16_clk),
    .RESET_B(net400),
    .D(_0424_),
    .Q_N(_2048_),
    .Q(\madd.total[4] ));
 sg13g2_dfrbp_1 \madd.total[5]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net401),
    .D(_0425_),
    .Q_N(_2047_),
    .Q(\madd.total[5] ));
 sg13g2_dfrbp_1 \madd.total[6]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_10_clk),
    .RESET_B(net402),
    .D(_0426_),
    .Q_N(_2046_),
    .Q(\madd.total[6] ));
 sg13g2_dfrbp_1 \madd.total[7]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_9_clk),
    .RESET_B(net403),
    .D(_0427_),
    .Q_N(_2045_),
    .Q(\madd.total[7] ));
 sg13g2_dfrbp_1 \madd.total[8]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net404),
    .D(_0428_),
    .Q_N(_2044_),
    .Q(\madd.total[8] ));
 sg13g2_dfrbp_1 \madd.total[9]$_SDFFCE_PP0P_  (.CLK(clknet_leaf_11_clk),
    .RESET_B(net405),
    .D(_0429_),
    .Q_N(_2043_),
    .Q(\madd.total[9] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[2]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[4]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[5]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[6]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[7]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout16 (.A(_1056_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_1062_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_1002_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_0982_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_0740_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1065_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0972_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0933_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0921_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_1047_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0914_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_1021_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_1014_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_1005_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0962_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0939_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0995_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0986_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_1441_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_1412_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1213_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1180_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1075_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_1023_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_1505_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_1472_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_1381_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_1350_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_1314_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_1148_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_1114_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_0573_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1414_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1242_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1182_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_1070_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0975_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1474_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1352_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_1308_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1277_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1117_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1034_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_0967_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_0689_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1239_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_0957_),
    .X(net62));
 sg13g2_buf_4 fanout63 (.X(net63),
    .A(_0567_));
 sg13g2_buf_2 fanout64 (.A(_1627_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_0944_),
    .X(net65));
 sg13g2_buf_8 fanout66 (.A(_2036_),
    .X(net66));
 sg13g2_buf_4 fanout67 (.X(net67),
    .A(_2032_));
 sg13g2_buf_4 fanout68 (.X(net68),
    .A(_2018_));
 sg13g2_buf_2 fanout69 (.A(_1274_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0716_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0668_),
    .X(net71));
 sg13g2_buf_4 fanout72 (.X(net72),
    .A(_2031_));
 sg13g2_buf_4 fanout73 (.X(net73),
    .A(_2027_));
 sg13g2_buf_4 fanout74 (.X(net74),
    .A(_2017_));
 sg13g2_buf_4 fanout75 (.X(net75),
    .A(_2014_));
 sg13g2_buf_4 fanout76 (.X(net76),
    .A(_0696_));
 sg13g2_buf_4 fanout77 (.X(net77),
    .A(_0451_));
 sg13g2_buf_4 fanout78 (.X(net78),
    .A(_2013_));
 sg13g2_buf_2 fanout79 (.A(_1730_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_1467_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_1383_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_1316_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_1174_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_1080_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1029_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0720_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0695_),
    .X(net87));
 sg13g2_buf_4 fanout88 (.X(net88),
    .A(_0684_));
 sg13g2_buf_2 fanout89 (.A(_1943_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_1906_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_1893_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_1818_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_1809_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_1030_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_0719_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_0694_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_0690_),
    .X(net97));
 sg13g2_buf_4 fanout98 (.X(net98),
    .A(_0683_));
 sg13g2_buf_2 fanout99 (.A(_0675_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_1970_),
    .X(net100));
 sg13g2_buf_4 fanout101 (.X(net101),
    .A(_1905_));
 sg13g2_buf_2 fanout102 (.A(_1808_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_0745_),
    .X(net103));
 sg13g2_buf_4 fanout104 (.X(net104),
    .A(_0693_));
 sg13g2_buf_4 fanout105 (.X(net105),
    .A(_0682_));
 sg13g2_buf_2 fanout106 (.A(_0621_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_1921_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_1910_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_1871_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_1025_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_0775_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_0744_),
    .X(net112));
 sg13g2_buf_4 fanout113 (.X(net113),
    .A(_0692_));
 sg13g2_buf_2 fanout114 (.A(_0660_),
    .X(net114));
 sg13g2_buf_4 fanout115 (.X(net115),
    .A(_1990_));
 sg13g2_buf_2 fanout116 (.A(_1908_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_1814_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_1806_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_1534_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_0764_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_0691_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_0678_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(_0484_));
 sg13g2_buf_2 fanout124 (.A(_0455_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_1991_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_1971_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_1962_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_1914_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_1903_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_1802_),
    .X(net130));
 sg13g2_buf_2 fanout131 (.A(_1761_),
    .X(net131));
 sg13g2_buf_2 fanout132 (.A(_1758_),
    .X(net132));
 sg13g2_buf_2 fanout133 (.A(_0771_),
    .X(net133));
 sg13g2_buf_2 fanout134 (.A(_0476_),
    .X(net134));
 sg13g2_buf_2 fanout135 (.A(_1916_),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(_1913_));
 sg13g2_buf_2 fanout137 (.A(_1812_),
    .X(net137));
 sg13g2_buf_2 fanout138 (.A(_1793_),
    .X(net138));
 sg13g2_buf_2 fanout139 (.A(_1776_),
    .X(net139));
 sg13g2_buf_2 fanout140 (.A(_1770_),
    .X(net140));
 sg13g2_buf_2 fanout141 (.A(_1915_),
    .X(net141));
 sg13g2_buf_2 fanout142 (.A(_1752_),
    .X(net142));
 sg13g2_tielo _3983__143 (.L_LO(net143));
 sg13g2_tielo _3984__144 (.L_LO(net144));
 sg13g2_tielo _3985__145 (.L_LO(net145));
 sg13g2_tielo _3986__146 (.L_LO(net146));
 sg13g2_tielo _3991__147 (.L_LO(net147));
 sg13g2_tielo _3992__148 (.L_LO(net148));
 sg13g2_tielo _3993__149 (.L_LO(net149));
 sg13g2_tielo _3994__150 (.L_LO(net150));
 sg13g2_tiehi _3978__152 (.L_HI(net152));
 sg13g2_tiehi _3979__153 (.L_HI(net153));
 sg13g2_tiehi _3980__154 (.L_HI(net154));
 sg13g2_tiehi _3987__155 (.L_HI(net155));
 sg13g2_tiehi _3988__156 (.L_HI(net156));
 sg13g2_tiehi _3989__157 (.L_HI(net157));
 sg13g2_tiehi _3990__158 (.L_HI(net158));
 sg13g2_tiehi \madd.count[0]$_SDFFCE_PP0P__159  (.L_HI(net159));
 sg13g2_tiehi \madd.count[10]$_SDFFCE_PP0P__160  (.L_HI(net160));
 sg13g2_tiehi \madd.count[11]$_SDFFCE_PP0P__161  (.L_HI(net161));
 sg13g2_tiehi \madd.count[1]$_SDFFCE_PP0P__162  (.L_HI(net162));
 sg13g2_tiehi \madd.count[2]$_SDFFCE_PP0P__163  (.L_HI(net163));
 sg13g2_tiehi \madd.count[3]$_SDFFCE_PP0P__164  (.L_HI(net164));
 sg13g2_tiehi \madd.count[4]$_SDFFCE_PP0P__165  (.L_HI(net165));
 sg13g2_tiehi \madd.count[5]$_SDFFCE_PP0P__166  (.L_HI(net166));
 sg13g2_tiehi \madd.count[6]$_SDFFCE_PP0P__167  (.L_HI(net167));
 sg13g2_tiehi \madd.count[7]$_SDFFCE_PP0P__168  (.L_HI(net168));
 sg13g2_tiehi \madd.count[8]$_SDFFCE_PP0P__169  (.L_HI(net169));
 sg13g2_tiehi \madd.count[9]$_SDFFCE_PP0P__170  (.L_HI(net170));
 sg13g2_tiehi \madd.delta[0]$_SDFFCE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \madd.delta[10]$_SDFFCE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \madd.delta[11]$_SDFFCE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \madd.delta[1]$_SDFFCE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \madd.delta[2]$_SDFFCE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \madd.delta[3]$_SDFFCE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \madd.delta[4]$_SDFFCE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \madd.delta[5]$_SDFFCE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \madd.delta[6]$_SDFFCE_PP0P__179  (.L_HI(net179));
 sg13g2_tiehi \madd.delta[7]$_SDFFCE_PP0P__180  (.L_HI(net180));
 sg13g2_tiehi \madd.delta[8]$_SDFFCE_PP0P__181  (.L_HI(net181));
 sg13g2_tiehi \madd.delta[9]$_SDFFCE_PP0P__182  (.L_HI(net182));
 sg13g2_tiehi \madd.i[0]$_DFFE_PN__183  (.L_HI(net183));
 sg13g2_tiehi \madd.i[1]$_DFFE_PN__184  (.L_HI(net184));
 sg13g2_tiehi \madd.i[2]$_DFFE_PN__185  (.L_HI(net185));
 sg13g2_tiehi \madd.i[3]$_DFFE_PN__186  (.L_HI(net186));
 sg13g2_tiehi \madd.i_d[0]$_SDFFE_PP0N__187  (.L_HI(net187));
 sg13g2_tiehi \madd.i_e[2]$_DFFE_PP__188  (.L_HI(net188));
 sg13g2_tiehi \madd.mem[0][0]$_DFFE_PP__189  (.L_HI(net189));
 sg13g2_tiehi \madd.mem[0][10]$_DFFE_PP__190  (.L_HI(net190));
 sg13g2_tiehi \madd.mem[0][11]$_DFFE_PP__191  (.L_HI(net191));
 sg13g2_tiehi \madd.mem[0][1]$_DFFE_PP__192  (.L_HI(net192));
 sg13g2_tiehi \madd.mem[0][2]$_DFFE_PP__193  (.L_HI(net193));
 sg13g2_tiehi \madd.mem[0][3]$_DFFE_PP__194  (.L_HI(net194));
 sg13g2_tiehi \madd.mem[0][4]$_DFFE_PP__195  (.L_HI(net195));
 sg13g2_tiehi \madd.mem[0][5]$_DFFE_PP__196  (.L_HI(net196));
 sg13g2_tiehi \madd.mem[0][6]$_DFFE_PP__197  (.L_HI(net197));
 sg13g2_tiehi \madd.mem[0][7]$_DFFE_PP__198  (.L_HI(net198));
 sg13g2_tiehi \madd.mem[0][8]$_DFFE_PP__199  (.L_HI(net199));
 sg13g2_tiehi \madd.mem[0][9]$_DFFE_PP__200  (.L_HI(net200));
 sg13g2_tiehi \madd.mem[10][0]$_DFFE_PP__201  (.L_HI(net201));
 sg13g2_tiehi \madd.mem[10][10]$_DFFE_PP__202  (.L_HI(net202));
 sg13g2_tiehi \madd.mem[10][11]$_DFFE_PP__203  (.L_HI(net203));
 sg13g2_tiehi \madd.mem[10][1]$_DFFE_PP__204  (.L_HI(net204));
 sg13g2_tiehi \madd.mem[10][2]$_DFFE_PP__205  (.L_HI(net205));
 sg13g2_tiehi \madd.mem[10][3]$_DFFE_PP__206  (.L_HI(net206));
 sg13g2_tiehi \madd.mem[10][4]$_DFFE_PP__207  (.L_HI(net207));
 sg13g2_tiehi \madd.mem[10][5]$_DFFE_PP__208  (.L_HI(net208));
 sg13g2_tiehi \madd.mem[10][6]$_DFFE_PP__209  (.L_HI(net209));
 sg13g2_tiehi \madd.mem[10][7]$_DFFE_PP__210  (.L_HI(net210));
 sg13g2_tiehi \madd.mem[10][8]$_DFFE_PP__211  (.L_HI(net211));
 sg13g2_tiehi \madd.mem[10][9]$_DFFE_PP__212  (.L_HI(net212));
 sg13g2_tiehi \madd.mem[11][0]$_DFFE_PP__213  (.L_HI(net213));
 sg13g2_tiehi \madd.mem[11][10]$_DFFE_PP__214  (.L_HI(net214));
 sg13g2_tiehi \madd.mem[11][11]$_DFFE_PP__215  (.L_HI(net215));
 sg13g2_tiehi \madd.mem[11][1]$_DFFE_PP__216  (.L_HI(net216));
 sg13g2_tiehi \madd.mem[11][2]$_DFFE_PP__217  (.L_HI(net217));
 sg13g2_tiehi \madd.mem[11][3]$_DFFE_PP__218  (.L_HI(net218));
 sg13g2_tiehi \madd.mem[11][4]$_DFFE_PP__219  (.L_HI(net219));
 sg13g2_tiehi \madd.mem[11][5]$_DFFE_PP__220  (.L_HI(net220));
 sg13g2_tiehi \madd.mem[11][6]$_DFFE_PP__221  (.L_HI(net221));
 sg13g2_tiehi \madd.mem[11][7]$_DFFE_PP__222  (.L_HI(net222));
 sg13g2_tiehi \madd.mem[11][8]$_DFFE_PP__223  (.L_HI(net223));
 sg13g2_tiehi \madd.mem[11][9]$_DFFE_PP__224  (.L_HI(net224));
 sg13g2_tiehi \madd.mem[12][0]$_DFFE_PP__225  (.L_HI(net225));
 sg13g2_tiehi \madd.mem[12][10]$_DFFE_PP__226  (.L_HI(net226));
 sg13g2_tiehi \madd.mem[12][11]$_DFFE_PP__227  (.L_HI(net227));
 sg13g2_tiehi \madd.mem[12][1]$_DFFE_PP__228  (.L_HI(net228));
 sg13g2_tiehi \madd.mem[12][2]$_DFFE_PP__229  (.L_HI(net229));
 sg13g2_tiehi \madd.mem[12][3]$_DFFE_PP__230  (.L_HI(net230));
 sg13g2_tiehi \madd.mem[12][4]$_DFFE_PP__231  (.L_HI(net231));
 sg13g2_tiehi \madd.mem[12][5]$_DFFE_PP__232  (.L_HI(net232));
 sg13g2_tiehi \madd.mem[12][6]$_DFFE_PP__233  (.L_HI(net233));
 sg13g2_tiehi \madd.mem[12][7]$_DFFE_PP__234  (.L_HI(net234));
 sg13g2_tiehi \madd.mem[12][8]$_DFFE_PP__235  (.L_HI(net235));
 sg13g2_tiehi \madd.mem[12][9]$_DFFE_PP__236  (.L_HI(net236));
 sg13g2_tiehi \madd.mem[13][0]$_DFFE_PP__237  (.L_HI(net237));
 sg13g2_tiehi \madd.mem[13][10]$_DFFE_PP__238  (.L_HI(net238));
 sg13g2_tiehi \madd.mem[13][11]$_DFFE_PP__239  (.L_HI(net239));
 sg13g2_tiehi \madd.mem[13][1]$_DFFE_PP__240  (.L_HI(net240));
 sg13g2_tiehi \madd.mem[13][2]$_DFFE_PP__241  (.L_HI(net241));
 sg13g2_tiehi \madd.mem[13][3]$_DFFE_PP__242  (.L_HI(net242));
 sg13g2_tiehi \madd.mem[13][4]$_DFFE_PP__243  (.L_HI(net243));
 sg13g2_tiehi \madd.mem[13][5]$_DFFE_PP__244  (.L_HI(net244));
 sg13g2_tiehi \madd.mem[13][6]$_DFFE_PP__245  (.L_HI(net245));
 sg13g2_tiehi \madd.mem[13][7]$_DFFE_PP__246  (.L_HI(net246));
 sg13g2_tiehi \madd.mem[13][8]$_DFFE_PP__247  (.L_HI(net247));
 sg13g2_tiehi \madd.mem[13][9]$_DFFE_PP__248  (.L_HI(net248));
 sg13g2_tiehi \madd.mem[14][0]$_DFFE_PP__249  (.L_HI(net249));
 sg13g2_tiehi \madd.mem[14][10]$_DFFE_PP__250  (.L_HI(net250));
 sg13g2_tiehi \madd.mem[14][11]$_DFFE_PP__251  (.L_HI(net251));
 sg13g2_tiehi \madd.mem[14][1]$_DFFE_PP__252  (.L_HI(net252));
 sg13g2_tiehi \madd.mem[14][2]$_DFFE_PP__253  (.L_HI(net253));
 sg13g2_tiehi \madd.mem[14][3]$_DFFE_PP__254  (.L_HI(net254));
 sg13g2_tiehi \madd.mem[14][4]$_DFFE_PP__255  (.L_HI(net255));
 sg13g2_tiehi \madd.mem[14][5]$_DFFE_PP__256  (.L_HI(net256));
 sg13g2_tiehi \madd.mem[14][6]$_DFFE_PP__257  (.L_HI(net257));
 sg13g2_tiehi \madd.mem[14][7]$_DFFE_PP__258  (.L_HI(net258));
 sg13g2_tiehi \madd.mem[14][8]$_DFFE_PP__259  (.L_HI(net259));
 sg13g2_tiehi \madd.mem[14][9]$_DFFE_PP__260  (.L_HI(net260));
 sg13g2_tiehi \madd.mem[15][0]$_DFFE_PP__261  (.L_HI(net261));
 sg13g2_tiehi \madd.mem[15][10]$_DFFE_PP__262  (.L_HI(net262));
 sg13g2_tiehi \madd.mem[15][11]$_DFFE_PP__263  (.L_HI(net263));
 sg13g2_tiehi \madd.mem[15][1]$_DFFE_PP__264  (.L_HI(net264));
 sg13g2_tiehi \madd.mem[15][2]$_DFFE_PP__265  (.L_HI(net265));
 sg13g2_tiehi \madd.mem[15][3]$_DFFE_PP__266  (.L_HI(net266));
 sg13g2_tiehi \madd.mem[15][4]$_DFFE_PP__267  (.L_HI(net267));
 sg13g2_tiehi \madd.mem[15][5]$_DFFE_PP__268  (.L_HI(net268));
 sg13g2_tiehi \madd.mem[15][6]$_DFFE_PP__269  (.L_HI(net269));
 sg13g2_tiehi \madd.mem[15][7]$_DFFE_PP__270  (.L_HI(net270));
 sg13g2_tiehi \madd.mem[15][8]$_DFFE_PP__271  (.L_HI(net271));
 sg13g2_tiehi \madd.mem[15][9]$_DFFE_PP__272  (.L_HI(net272));
 sg13g2_tiehi \madd.mem[1][0]$_DFFE_PP__273  (.L_HI(net273));
 sg13g2_tiehi \madd.mem[1][10]$_DFFE_PP__274  (.L_HI(net274));
 sg13g2_tiehi \madd.mem[1][11]$_DFFE_PP__275  (.L_HI(net275));
 sg13g2_tiehi \madd.mem[1][1]$_DFFE_PP__276  (.L_HI(net276));
 sg13g2_tiehi \madd.mem[1][2]$_DFFE_PP__277  (.L_HI(net277));
 sg13g2_tiehi \madd.mem[1][3]$_DFFE_PP__278  (.L_HI(net278));
 sg13g2_tiehi \madd.mem[1][4]$_DFFE_PP__279  (.L_HI(net279));
 sg13g2_tiehi \madd.mem[1][5]$_DFFE_PP__280  (.L_HI(net280));
 sg13g2_tiehi \madd.mem[1][6]$_DFFE_PP__281  (.L_HI(net281));
 sg13g2_tiehi \madd.mem[1][7]$_DFFE_PP__282  (.L_HI(net282));
 sg13g2_tiehi \madd.mem[1][8]$_DFFE_PP__283  (.L_HI(net283));
 sg13g2_tiehi \madd.mem[1][9]$_DFFE_PP__284  (.L_HI(net284));
 sg13g2_tiehi \madd.mem[2][0]$_DFFE_PP__285  (.L_HI(net285));
 sg13g2_tiehi \madd.mem[2][10]$_DFFE_PP__286  (.L_HI(net286));
 sg13g2_tiehi \madd.mem[2][11]$_DFFE_PP__287  (.L_HI(net287));
 sg13g2_tiehi \madd.mem[2][1]$_DFFE_PP__288  (.L_HI(net288));
 sg13g2_tiehi \madd.mem[2][2]$_DFFE_PP__289  (.L_HI(net289));
 sg13g2_tiehi \madd.mem[2][3]$_DFFE_PP__290  (.L_HI(net290));
 sg13g2_tiehi \madd.mem[2][4]$_DFFE_PP__291  (.L_HI(net291));
 sg13g2_tiehi \madd.mem[2][5]$_DFFE_PP__292  (.L_HI(net292));
 sg13g2_tiehi \madd.mem[2][6]$_DFFE_PP__293  (.L_HI(net293));
 sg13g2_tiehi \madd.mem[2][7]$_DFFE_PP__294  (.L_HI(net294));
 sg13g2_tiehi \madd.mem[2][8]$_DFFE_PP__295  (.L_HI(net295));
 sg13g2_tiehi \madd.mem[2][9]$_DFFE_PP__296  (.L_HI(net296));
 sg13g2_tiehi \madd.mem[3][0]$_DFFE_PP__297  (.L_HI(net297));
 sg13g2_tiehi \madd.mem[3][10]$_DFFE_PP__298  (.L_HI(net298));
 sg13g2_tiehi \madd.mem[3][11]$_DFFE_PP__299  (.L_HI(net299));
 sg13g2_tiehi \madd.mem[3][1]$_DFFE_PP__300  (.L_HI(net300));
 sg13g2_tiehi \madd.mem[3][2]$_DFFE_PP__301  (.L_HI(net301));
 sg13g2_tiehi \madd.mem[3][3]$_DFFE_PP__302  (.L_HI(net302));
 sg13g2_tiehi \madd.mem[3][4]$_DFFE_PP__303  (.L_HI(net303));
 sg13g2_tiehi \madd.mem[3][5]$_DFFE_PP__304  (.L_HI(net304));
 sg13g2_tiehi \madd.mem[3][6]$_DFFE_PP__305  (.L_HI(net305));
 sg13g2_tiehi \madd.mem[3][7]$_DFFE_PP__306  (.L_HI(net306));
 sg13g2_tiehi \madd.mem[3][8]$_DFFE_PP__307  (.L_HI(net307));
 sg13g2_tiehi \madd.mem[3][9]$_DFFE_PP__308  (.L_HI(net308));
 sg13g2_tiehi \madd.mem[4][0]$_DFFE_PP__309  (.L_HI(net309));
 sg13g2_tiehi \madd.mem[4][10]$_DFFE_PP__310  (.L_HI(net310));
 sg13g2_tiehi \madd.mem[4][11]$_DFFE_PP__311  (.L_HI(net311));
 sg13g2_tiehi \madd.mem[4][1]$_DFFE_PP__312  (.L_HI(net312));
 sg13g2_tiehi \madd.mem[4][2]$_DFFE_PP__313  (.L_HI(net313));
 sg13g2_tiehi \madd.mem[4][3]$_DFFE_PP__314  (.L_HI(net314));
 sg13g2_tiehi \madd.mem[4][4]$_DFFE_PP__315  (.L_HI(net315));
 sg13g2_tiehi \madd.mem[4][5]$_DFFE_PP__316  (.L_HI(net316));
 sg13g2_tiehi \madd.mem[4][6]$_DFFE_PP__317  (.L_HI(net317));
 sg13g2_tiehi \madd.mem[4][7]$_DFFE_PP__318  (.L_HI(net318));
 sg13g2_tiehi \madd.mem[4][8]$_DFFE_PP__319  (.L_HI(net319));
 sg13g2_tiehi \madd.mem[4][9]$_DFFE_PP__320  (.L_HI(net320));
 sg13g2_tiehi \madd.mem[5][0]$_DFFE_PP__321  (.L_HI(net321));
 sg13g2_tiehi \madd.mem[5][10]$_DFFE_PP__322  (.L_HI(net322));
 sg13g2_tiehi \madd.mem[5][11]$_DFFE_PP__323  (.L_HI(net323));
 sg13g2_tiehi \madd.mem[5][1]$_DFFE_PP__324  (.L_HI(net324));
 sg13g2_tiehi \madd.mem[5][2]$_DFFE_PP__325  (.L_HI(net325));
 sg13g2_tiehi \madd.mem[5][3]$_DFFE_PP__326  (.L_HI(net326));
 sg13g2_tiehi \madd.mem[5][4]$_DFFE_PP__327  (.L_HI(net327));
 sg13g2_tiehi \madd.mem[5][5]$_DFFE_PP__328  (.L_HI(net328));
 sg13g2_tiehi \madd.mem[5][6]$_DFFE_PP__329  (.L_HI(net329));
 sg13g2_tiehi \madd.mem[5][7]$_DFFE_PP__330  (.L_HI(net330));
 sg13g2_tiehi \madd.mem[5][8]$_DFFE_PP__331  (.L_HI(net331));
 sg13g2_tiehi \madd.mem[5][9]$_DFFE_PP__332  (.L_HI(net332));
 sg13g2_tiehi \madd.mem[6][0]$_DFFE_PP__333  (.L_HI(net333));
 sg13g2_tiehi \madd.mem[6][10]$_DFFE_PP__334  (.L_HI(net334));
 sg13g2_tiehi \madd.mem[6][11]$_DFFE_PP__335  (.L_HI(net335));
 sg13g2_tiehi \madd.mem[6][1]$_DFFE_PP__336  (.L_HI(net336));
 sg13g2_tiehi \madd.mem[6][2]$_DFFE_PP__337  (.L_HI(net337));
 sg13g2_tiehi \madd.mem[6][3]$_DFFE_PP__338  (.L_HI(net338));
 sg13g2_tiehi \madd.mem[6][4]$_DFFE_PP__339  (.L_HI(net339));
 sg13g2_tiehi \madd.mem[6][5]$_DFFE_PP__340  (.L_HI(net340));
 sg13g2_tiehi \madd.mem[6][6]$_DFFE_PP__341  (.L_HI(net341));
 sg13g2_tiehi \madd.mem[6][7]$_DFFE_PP__342  (.L_HI(net342));
 sg13g2_tiehi \madd.mem[6][8]$_DFFE_PP__343  (.L_HI(net343));
 sg13g2_tiehi \madd.mem[6][9]$_DFFE_PP__344  (.L_HI(net344));
 sg13g2_tiehi \madd.mem[7][0]$_DFFE_PP__345  (.L_HI(net345));
 sg13g2_tiehi \madd.mem[7][10]$_DFFE_PP__346  (.L_HI(net346));
 sg13g2_tiehi \madd.mem[7][11]$_DFFE_PP__347  (.L_HI(net347));
 sg13g2_tiehi \madd.mem[7][1]$_DFFE_PP__348  (.L_HI(net348));
 sg13g2_tiehi \madd.mem[7][2]$_DFFE_PP__349  (.L_HI(net349));
 sg13g2_tiehi \madd.mem[7][3]$_DFFE_PP__350  (.L_HI(net350));
 sg13g2_tiehi \madd.mem[7][4]$_DFFE_PP__351  (.L_HI(net351));
 sg13g2_tiehi \madd.mem[7][5]$_DFFE_PP__352  (.L_HI(net352));
 sg13g2_tiehi \madd.mem[7][6]$_DFFE_PP__353  (.L_HI(net353));
 sg13g2_tiehi \madd.mem[7][7]$_DFFE_PP__354  (.L_HI(net354));
 sg13g2_tiehi \madd.mem[7][8]$_DFFE_PP__355  (.L_HI(net355));
 sg13g2_tiehi \madd.mem[7][9]$_DFFE_PP__356  (.L_HI(net356));
 sg13g2_tiehi \madd.mem[8][0]$_DFFE_PP__357  (.L_HI(net357));
 sg13g2_tiehi \madd.mem[8][10]$_DFFE_PP__358  (.L_HI(net358));
 sg13g2_tiehi \madd.mem[8][11]$_DFFE_PP__359  (.L_HI(net359));
 sg13g2_tiehi \madd.mem[8][1]$_DFFE_PP__360  (.L_HI(net360));
 sg13g2_tiehi \madd.mem[8][2]$_DFFE_PP__361  (.L_HI(net361));
 sg13g2_tiehi \madd.mem[8][3]$_DFFE_PP__362  (.L_HI(net362));
 sg13g2_tiehi \madd.mem[8][4]$_DFFE_PP__363  (.L_HI(net363));
 sg13g2_tiehi \madd.mem[8][5]$_DFFE_PP__364  (.L_HI(net364));
 sg13g2_tiehi \madd.mem[8][6]$_DFFE_PP__365  (.L_HI(net365));
 sg13g2_tiehi \madd.mem[8][7]$_DFFE_PP__366  (.L_HI(net366));
 sg13g2_tiehi \madd.mem[8][8]$_DFFE_PP__367  (.L_HI(net367));
 sg13g2_tiehi \madd.mem[8][9]$_DFFE_PP__368  (.L_HI(net368));
 sg13g2_tiehi \madd.mem[9][0]$_DFFE_PP__369  (.L_HI(net369));
 sg13g2_tiehi \madd.mem[9][10]$_DFFE_PP__370  (.L_HI(net370));
 sg13g2_tiehi \madd.mem[9][11]$_DFFE_PP__371  (.L_HI(net371));
 sg13g2_tiehi \madd.mem[9][1]$_DFFE_PP__372  (.L_HI(net372));
 sg13g2_tiehi \madd.mem[9][2]$_DFFE_PP__373  (.L_HI(net373));
 sg13g2_tiehi \madd.mem[9][3]$_DFFE_PP__374  (.L_HI(net374));
 sg13g2_tiehi \madd.mem[9][4]$_DFFE_PP__375  (.L_HI(net375));
 sg13g2_tiehi \madd.mem[9][5]$_DFFE_PP__376  (.L_HI(net376));
 sg13g2_tiehi \madd.mem[9][6]$_DFFE_PP__377  (.L_HI(net377));
 sg13g2_tiehi \madd.mem[9][7]$_DFFE_PP__378  (.L_HI(net378));
 sg13g2_tiehi \madd.mem[9][8]$_DFFE_PP__379  (.L_HI(net379));
 sg13g2_tiehi \madd.mem[9][9]$_DFFE_PP__380  (.L_HI(net380));
 sg13g2_tiehi \madd.out_reg[0]$_DFFE_PP__381  (.L_HI(net381));
 sg13g2_tiehi \madd.out_reg[10]$_SDFFE_PP0P__382  (.L_HI(net382));
 sg13g2_tiehi \madd.out_reg[11]$_SDFFE_PP0P__383  (.L_HI(net383));
 sg13g2_tiehi \madd.out_reg[1]$_DFFE_PP__384  (.L_HI(net384));
 sg13g2_tiehi \madd.out_reg[2]$_DFFE_PP__385  (.L_HI(net385));
 sg13g2_tiehi \madd.out_reg[3]$_DFFE_PP__386  (.L_HI(net386));
 sg13g2_tiehi \madd.out_reg[4]$_SDFFE_PP0P__387  (.L_HI(net387));
 sg13g2_tiehi \madd.out_reg[5]$_SDFFE_PP0P__388  (.L_HI(net388));
 sg13g2_tiehi \madd.out_reg[6]$_SDFFE_PP0P__389  (.L_HI(net389));
 sg13g2_tiehi \madd.out_reg[7]$_SDFFE_PP0P__390  (.L_HI(net390));
 sg13g2_tiehi \madd.out_reg[8]$_SDFFE_PP0P__391  (.L_HI(net391));
 sg13g2_tiehi \madd.out_reg[9]$_SDFFE_PP0P__392  (.L_HI(net392));
 sg13g2_tiehi \madd.set$_SDFFE_PP1N__393  (.L_HI(net393));
 sg13g2_tiehi \madd.total[0]$_SDFFCE_PP0P__394  (.L_HI(net394));
 sg13g2_tiehi \madd.total[10]$_SDFFCE_PP0P__395  (.L_HI(net395));
 sg13g2_tiehi \madd.total[11]$_SDFFCE_PP0P__396  (.L_HI(net396));
 sg13g2_tiehi \madd.total[1]$_SDFFCE_PP0P__397  (.L_HI(net397));
 sg13g2_tiehi \madd.total[2]$_SDFFCE_PP0P__398  (.L_HI(net398));
 sg13g2_tiehi \madd.total[3]$_SDFFCE_PP0P__399  (.L_HI(net399));
 sg13g2_tiehi \madd.total[4]$_SDFFCE_PP0P__400  (.L_HI(net400));
 sg13g2_tiehi \madd.total[5]$_SDFFCE_PP0P__401  (.L_HI(net401));
 sg13g2_tiehi \madd.total[6]$_SDFFCE_PP0P__402  (.L_HI(net402));
 sg13g2_tiehi \madd.total[7]$_SDFFCE_PP0P__403  (.L_HI(net403));
 sg13g2_tiehi \madd.total[8]$_SDFFCE_PP0P__404  (.L_HI(net404));
 sg13g2_tiehi \madd.total[9]$_SDFFCE_PP0P__405  (.L_HI(net405));
 sg13g2_buf_2 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sg13g2_buf_2 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sg13g2_buf_2 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sg13g2_buf_2 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sg13g2_buf_2 clkbuf_leaf_5_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sg13g2_buf_2 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_6_clk));
 sg13g2_buf_2 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_7_clk));
 sg13g2_buf_2 clkbuf_leaf_8_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_8_clk));
 sg13g2_buf_2 clkbuf_leaf_9_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_9_clk));
 sg13g2_buf_2 clkbuf_leaf_10_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_10_clk));
 sg13g2_buf_2 clkbuf_leaf_11_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_11_clk));
 sg13g2_buf_2 clkbuf_leaf_12_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_12_clk));
 sg13g2_buf_2 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_13_clk));
 sg13g2_buf_2 clkbuf_leaf_14_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_14_clk));
 sg13g2_buf_2 clkbuf_leaf_15_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_15_clk));
 sg13g2_buf_2 clkbuf_leaf_16_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_16_clk));
 sg13g2_buf_2 clkbuf_leaf_17_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_17_clk));
 sg13g2_buf_2 clkbuf_leaf_18_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_18_clk));
 sg13g2_buf_2 clkbuf_leaf_19_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_19_clk));
 sg13g2_buf_2 clkbuf_leaf_20_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_20_clk));
 sg13g2_buf_2 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk));
 sg13g2_buf_2 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sg13g2_buf_2 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sg13g2_buf_2 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sg13g2_buf_2 clkbuf_leaf_25_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_25_clk));
 sg13g2_buf_2 clkbuf_leaf_26_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_26_clk));
 sg13g2_buf_2 clkbuf_leaf_27_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_27_clk));
 sg13g2_buf_2 clkbuf_leaf_28_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_28_clk));
 sg13g2_buf_2 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_29_clk));
 sg13g2_buf_2 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sg13g2_buf_2 clkbuf_leaf_31_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_31_clk));
 sg13g2_buf_2 clkbuf_leaf_32_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_32_clk));
 sg13g2_buf_2 clkbuf_leaf_33_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_33_clk));
 sg13g2_buf_2 clkbuf_leaf_34_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_34_clk));
 sg13g2_buf_2 clkbuf_leaf_35_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_35_clk));
 sg13g2_buf_2 clkbuf_leaf_36_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_36_clk));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_2 clkload0 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_2 clkload1 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_2 clkload2 (.A(clknet_3_7__leaf_clk));
 sg13g2_inv_2 clkload3 (.A(clknet_leaf_34_clk));
 sg13g2_buf_8 clkload4 (.A(clknet_leaf_35_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_leaf_1_clk));
 sg13g2_inv_2 clkload6 (.A(clknet_leaf_4_clk));
 sg13g2_buf_8 clkload7 (.A(clknet_leaf_32_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_leaf_25_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_leaf_26_clk));
 sg13g2_inv_2 clkload10 (.A(clknet_leaf_29_clk));
 sg13g2_buf_8 clkload11 (.A(clknet_leaf_23_clk));
 sg13g2_buf_8 clkload12 (.A(clknet_leaf_5_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_leaf_6_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_leaf_13_clk));
 sg13g2_buf_8 clkload15 (.A(clknet_leaf_31_clk));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_12_clk));
 sg13g2_inv_2 clkload17 (.A(clknet_leaf_14_clk));
 sg13g2_inv_2 clkload18 (.A(clknet_leaf_15_clk));
 sg13g2_buf_8 clkload19 (.A(clknet_leaf_19_clk));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_17_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_fill_2 FILLER_0_203 ();
 sg13g2_fill_1 FILLER_0_205 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_fill_1 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_228 ();
 sg13g2_decap_8 FILLER_0_235 ();
 sg13g2_decap_8 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_249 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_decap_8 FILLER_0_263 ();
 sg13g2_decap_8 FILLER_0_270 ();
 sg13g2_decap_8 FILLER_0_277 ();
 sg13g2_decap_8 FILLER_0_284 ();
 sg13g2_decap_8 FILLER_0_291 ();
 sg13g2_decap_8 FILLER_0_298 ();
 sg13g2_decap_8 FILLER_0_305 ();
 sg13g2_decap_8 FILLER_0_312 ();
 sg13g2_decap_8 FILLER_0_319 ();
 sg13g2_decap_8 FILLER_0_326 ();
 sg13g2_fill_2 FILLER_0_333 ();
 sg13g2_fill_1 FILLER_0_335 ();
 sg13g2_decap_8 FILLER_0_340 ();
 sg13g2_decap_8 FILLER_0_347 ();
 sg13g2_decap_8 FILLER_0_354 ();
 sg13g2_decap_8 FILLER_0_361 ();
 sg13g2_decap_8 FILLER_0_368 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_403 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_4 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_83 ();
 sg13g2_fill_2 FILLER_1_90 ();
 sg13g2_decap_4 FILLER_1_96 ();
 sg13g2_fill_2 FILLER_1_100 ();
 sg13g2_decap_8 FILLER_1_106 ();
 sg13g2_decap_8 FILLER_1_113 ();
 sg13g2_decap_4 FILLER_1_120 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_fill_2 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_fill_2 FILLER_1_196 ();
 sg13g2_fill_1 FILLER_1_198 ();
 sg13g2_decap_4 FILLER_1_251 ();
 sg13g2_fill_2 FILLER_1_255 ();
 sg13g2_fill_1 FILLER_1_283 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_4 FILLER_1_301 ();
 sg13g2_fill_2 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_311 ();
 sg13g2_fill_1 FILLER_1_318 ();
 sg13g2_fill_2 FILLER_1_323 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_4 FILLER_2_42 ();
 sg13g2_fill_2 FILLER_2_46 ();
 sg13g2_fill_1 FILLER_2_161 ();
 sg13g2_fill_1 FILLER_2_166 ();
 sg13g2_fill_2 FILLER_2_219 ();
 sg13g2_fill_1 FILLER_2_225 ();
 sg13g2_fill_2 FILLER_2_252 ();
 sg13g2_fill_2 FILLER_2_358 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_decap_8 FILLER_2_406 ();
 sg13g2_decap_8 FILLER_2_413 ();
 sg13g2_decap_8 FILLER_2_420 ();
 sg13g2_fill_2 FILLER_2_427 ();
 sg13g2_fill_1 FILLER_2_429 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_4 FILLER_3_49 ();
 sg13g2_fill_1 FILLER_3_53 ();
 sg13g2_fill_2 FILLER_3_132 ();
 sg13g2_fill_1 FILLER_3_141 ();
 sg13g2_fill_1 FILLER_3_150 ();
 sg13g2_fill_1 FILLER_3_156 ();
 sg13g2_fill_1 FILLER_3_161 ();
 sg13g2_fill_2 FILLER_3_169 ();
 sg13g2_fill_1 FILLER_3_171 ();
 sg13g2_decap_4 FILLER_3_183 ();
 sg13g2_fill_2 FILLER_3_187 ();
 sg13g2_fill_2 FILLER_3_200 ();
 sg13g2_fill_2 FILLER_3_206 ();
 sg13g2_fill_1 FILLER_3_208 ();
 sg13g2_fill_2 FILLER_3_215 ();
 sg13g2_fill_1 FILLER_3_217 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_fill_1 FILLER_3_228 ();
 sg13g2_fill_1 FILLER_3_233 ();
 sg13g2_fill_1 FILLER_3_242 ();
 sg13g2_fill_2 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_271 ();
 sg13g2_fill_1 FILLER_3_329 ();
 sg13g2_fill_1 FILLER_3_349 ();
 sg13g2_decap_8 FILLER_3_376 ();
 sg13g2_decap_8 FILLER_3_383 ();
 sg13g2_decap_8 FILLER_3_390 ();
 sg13g2_decap_8 FILLER_3_397 ();
 sg13g2_decap_8 FILLER_3_404 ();
 sg13g2_decap_8 FILLER_3_411 ();
 sg13g2_decap_8 FILLER_3_418 ();
 sg13g2_decap_4 FILLER_3_425 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_4 FILLER_4_49 ();
 sg13g2_fill_2 FILLER_4_53 ();
 sg13g2_fill_1 FILLER_4_61 ();
 sg13g2_fill_2 FILLER_4_72 ();
 sg13g2_fill_1 FILLER_4_105 ();
 sg13g2_fill_1 FILLER_4_110 ();
 sg13g2_fill_1 FILLER_4_116 ();
 sg13g2_fill_1 FILLER_4_122 ();
 sg13g2_fill_1 FILLER_4_127 ();
 sg13g2_decap_4 FILLER_4_144 ();
 sg13g2_fill_1 FILLER_4_148 ();
 sg13g2_fill_1 FILLER_4_159 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_fill_1 FILLER_4_184 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_4_211 ();
 sg13g2_fill_2 FILLER_4_218 ();
 sg13g2_decap_8 FILLER_4_225 ();
 sg13g2_decap_4 FILLER_4_236 ();
 sg13g2_fill_1 FILLER_4_240 ();
 sg13g2_decap_4 FILLER_4_245 ();
 sg13g2_fill_1 FILLER_4_249 ();
 sg13g2_fill_1 FILLER_4_255 ();
 sg13g2_fill_1 FILLER_4_298 ();
 sg13g2_fill_1 FILLER_4_312 ();
 sg13g2_fill_1 FILLER_4_317 ();
 sg13g2_fill_1 FILLER_4_322 ();
 sg13g2_fill_2 FILLER_4_348 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_decap_8 FILLER_4_381 ();
 sg13g2_decap_8 FILLER_4_388 ();
 sg13g2_decap_8 FILLER_4_395 ();
 sg13g2_decap_8 FILLER_4_402 ();
 sg13g2_decap_8 FILLER_4_409 ();
 sg13g2_decap_8 FILLER_4_416 ();
 sg13g2_decap_8 FILLER_4_423 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_fill_2 FILLER_5_49 ();
 sg13g2_fill_1 FILLER_5_51 ();
 sg13g2_fill_2 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_83 ();
 sg13g2_decap_8 FILLER_5_90 ();
 sg13g2_decap_8 FILLER_5_97 ();
 sg13g2_decap_8 FILLER_5_104 ();
 sg13g2_decap_4 FILLER_5_111 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_decap_8 FILLER_5_120 ();
 sg13g2_decap_8 FILLER_5_127 ();
 sg13g2_fill_2 FILLER_5_134 ();
 sg13g2_fill_1 FILLER_5_136 ();
 sg13g2_fill_1 FILLER_5_161 ();
 sg13g2_decap_4 FILLER_5_169 ();
 sg13g2_decap_4 FILLER_5_178 ();
 sg13g2_fill_2 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_188 ();
 sg13g2_decap_8 FILLER_5_195 ();
 sg13g2_fill_2 FILLER_5_202 ();
 sg13g2_fill_1 FILLER_5_204 ();
 sg13g2_fill_2 FILLER_5_210 ();
 sg13g2_fill_1 FILLER_5_212 ();
 sg13g2_fill_2 FILLER_5_217 ();
 sg13g2_fill_1 FILLER_5_219 ();
 sg13g2_decap_8 FILLER_5_233 ();
 sg13g2_decap_8 FILLER_5_240 ();
 sg13g2_decap_8 FILLER_5_247 ();
 sg13g2_fill_2 FILLER_5_254 ();
 sg13g2_fill_1 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_261 ();
 sg13g2_decap_8 FILLER_5_267 ();
 sg13g2_fill_2 FILLER_5_274 ();
 sg13g2_decap_4 FILLER_5_280 ();
 sg13g2_fill_2 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_290 ();
 sg13g2_decap_8 FILLER_5_297 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_4 FILLER_5_311 ();
 sg13g2_fill_2 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_fill_2 FILLER_5_337 ();
 sg13g2_fill_2 FILLER_5_343 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_decap_4 FILLER_5_352 ();
 sg13g2_fill_1 FILLER_5_356 ();
 sg13g2_fill_1 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_decap_8 FILLER_5_406 ();
 sg13g2_decap_8 FILLER_5_413 ();
 sg13g2_decap_8 FILLER_5_420 ();
 sg13g2_fill_2 FILLER_5_427 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_65 ();
 sg13g2_decap_8 FILLER_6_72 ();
 sg13g2_decap_8 FILLER_6_79 ();
 sg13g2_decap_8 FILLER_6_86 ();
 sg13g2_fill_1 FILLER_6_123 ();
 sg13g2_fill_2 FILLER_6_159 ();
 sg13g2_fill_1 FILLER_6_161 ();
 sg13g2_fill_2 FILLER_6_188 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_decap_4 FILLER_6_263 ();
 sg13g2_fill_2 FILLER_6_279 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_296 ();
 sg13g2_fill_2 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_333 ();
 sg13g2_decap_8 FILLER_6_340 ();
 sg13g2_fill_2 FILLER_6_347 ();
 sg13g2_fill_1 FILLER_6_349 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_decap_8 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_6_414 ();
 sg13g2_decap_8 FILLER_6_421 ();
 sg13g2_fill_2 FILLER_6_428 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_fill_2 FILLER_7_28 ();
 sg13g2_fill_1 FILLER_7_30 ();
 sg13g2_decap_8 FILLER_7_65 ();
 sg13g2_decap_8 FILLER_7_72 ();
 sg13g2_fill_2 FILLER_7_84 ();
 sg13g2_decap_4 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_121 ();
 sg13g2_fill_2 FILLER_7_128 ();
 sg13g2_fill_1 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_134 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_fill_2 FILLER_7_156 ();
 sg13g2_fill_1 FILLER_7_162 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_decap_4 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_183 ();
 sg13g2_decap_8 FILLER_7_210 ();
 sg13g2_decap_4 FILLER_7_217 ();
 sg13g2_fill_2 FILLER_7_221 ();
 sg13g2_fill_1 FILLER_7_230 ();
 sg13g2_decap_8 FILLER_7_243 ();
 sg13g2_fill_1 FILLER_7_250 ();
 sg13g2_fill_1 FILLER_7_313 ();
 sg13g2_fill_1 FILLER_7_323 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_4 FILLER_8_35 ();
 sg13g2_fill_1 FILLER_8_43 ();
 sg13g2_fill_1 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_59 ();
 sg13g2_fill_2 FILLER_8_64 ();
 sg13g2_decap_4 FILLER_8_112 ();
 sg13g2_decap_4 FILLER_8_154 ();
 sg13g2_decap_4 FILLER_8_170 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_decap_4 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_184 ();
 sg13g2_fill_1 FILLER_8_190 ();
 sg13g2_fill_2 FILLER_8_197 ();
 sg13g2_fill_2 FILLER_8_220 ();
 sg13g2_fill_2 FILLER_8_248 ();
 sg13g2_fill_1 FILLER_8_250 ();
 sg13g2_fill_2 FILLER_8_272 ();
 sg13g2_fill_1 FILLER_8_274 ();
 sg13g2_fill_2 FILLER_8_279 ();
 sg13g2_fill_2 FILLER_8_309 ();
 sg13g2_decap_8 FILLER_8_337 ();
 sg13g2_fill_1 FILLER_8_344 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_decap_8 FILLER_8_381 ();
 sg13g2_decap_8 FILLER_8_388 ();
 sg13g2_decap_8 FILLER_8_395 ();
 sg13g2_decap_8 FILLER_8_402 ();
 sg13g2_decap_8 FILLER_8_409 ();
 sg13g2_decap_8 FILLER_8_416 ();
 sg13g2_decap_8 FILLER_8_423 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_fill_2 FILLER_9_100 ();
 sg13g2_fill_1 FILLER_9_102 ();
 sg13g2_fill_1 FILLER_9_128 ();
 sg13g2_decap_4 FILLER_9_133 ();
 sg13g2_decap_4 FILLER_9_150 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_221 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_decap_8 FILLER_9_258 ();
 sg13g2_decap_8 FILLER_9_265 ();
 sg13g2_decap_8 FILLER_9_272 ();
 sg13g2_decap_4 FILLER_9_279 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_4 FILLER_9_306 ();
 sg13g2_fill_1 FILLER_9_310 ();
 sg13g2_fill_2 FILLER_9_316 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_4 FILLER_9_350 ();
 sg13g2_fill_1 FILLER_9_354 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_8 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_9_412 ();
 sg13g2_decap_8 FILLER_9_419 ();
 sg13g2_decap_4 FILLER_9_426 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_fill_1 FILLER_10_49 ();
 sg13g2_fill_1 FILLER_10_56 ();
 sg13g2_decap_4 FILLER_10_63 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_73 ();
 sg13g2_fill_2 FILLER_10_80 ();
 sg13g2_fill_1 FILLER_10_82 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_fill_1 FILLER_10_95 ();
 sg13g2_fill_2 FILLER_10_101 ();
 sg13g2_fill_1 FILLER_10_103 ();
 sg13g2_fill_1 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_fill_1 FILLER_10_144 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_decap_8 FILLER_10_192 ();
 sg13g2_decap_8 FILLER_10_203 ();
 sg13g2_fill_2 FILLER_10_210 ();
 sg13g2_fill_1 FILLER_10_212 ();
 sg13g2_decap_8 FILLER_10_218 ();
 sg13g2_fill_2 FILLER_10_225 ();
 sg13g2_decap_4 FILLER_10_246 ();
 sg13g2_fill_1 FILLER_10_250 ();
 sg13g2_decap_4 FILLER_10_261 ();
 sg13g2_fill_1 FILLER_10_265 ();
 sg13g2_decap_8 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_279 ();
 sg13g2_fill_1 FILLER_10_284 ();
 sg13g2_fill_2 FILLER_10_306 ();
 sg13g2_fill_1 FILLER_10_308 ();
 sg13g2_decap_4 FILLER_10_315 ();
 sg13g2_fill_1 FILLER_10_319 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_fill_1 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_fill_1 FILLER_10_355 ();
 sg13g2_fill_2 FILLER_10_359 ();
 sg13g2_decap_8 FILLER_10_391 ();
 sg13g2_decap_8 FILLER_10_398 ();
 sg13g2_decap_8 FILLER_10_405 ();
 sg13g2_decap_8 FILLER_10_412 ();
 sg13g2_decap_8 FILLER_10_419 ();
 sg13g2_decap_4 FILLER_10_426 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_4 FILLER_11_79 ();
 sg13g2_fill_1 FILLER_11_83 ();
 sg13g2_fill_2 FILLER_11_90 ();
 sg13g2_fill_2 FILLER_11_100 ();
 sg13g2_fill_1 FILLER_11_102 ();
 sg13g2_fill_2 FILLER_11_111 ();
 sg13g2_decap_8 FILLER_11_118 ();
 sg13g2_fill_2 FILLER_11_125 ();
 sg13g2_fill_1 FILLER_11_127 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_4 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_193 ();
 sg13g2_decap_8 FILLER_11_200 ();
 sg13g2_decap_8 FILLER_11_207 ();
 sg13g2_fill_2 FILLER_11_214 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_decap_4 FILLER_11_221 ();
 sg13g2_decap_8 FILLER_11_230 ();
 sg13g2_decap_8 FILLER_11_237 ();
 sg13g2_decap_8 FILLER_11_244 ();
 sg13g2_fill_2 FILLER_11_251 ();
 sg13g2_fill_1 FILLER_11_310 ();
 sg13g2_fill_1 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_fill_2 FILLER_12_56 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_decap_8 FILLER_12_63 ();
 sg13g2_decap_4 FILLER_12_70 ();
 sg13g2_fill_1 FILLER_12_100 ();
 sg13g2_decap_8 FILLER_12_135 ();
 sg13g2_decap_8 FILLER_12_142 ();
 sg13g2_fill_1 FILLER_12_149 ();
 sg13g2_decap_8 FILLER_12_155 ();
 sg13g2_fill_2 FILLER_12_175 ();
 sg13g2_fill_2 FILLER_12_185 ();
 sg13g2_fill_1 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_192 ();
 sg13g2_fill_1 FILLER_12_203 ();
 sg13g2_fill_1 FILLER_12_208 ();
 sg13g2_fill_1 FILLER_12_239 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_fill_2 FILLER_12_251 ();
 sg13g2_decap_8 FILLER_12_258 ();
 sg13g2_decap_4 FILLER_12_265 ();
 sg13g2_decap_4 FILLER_12_273 ();
 sg13g2_fill_2 FILLER_12_277 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_290 ();
 sg13g2_decap_4 FILLER_12_301 ();
 sg13g2_fill_1 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_310 ();
 sg13g2_fill_2 FILLER_12_317 ();
 sg13g2_fill_1 FILLER_12_319 ();
 sg13g2_decap_4 FILLER_12_325 ();
 sg13g2_decap_8 FILLER_12_337 ();
 sg13g2_fill_2 FILLER_12_344 ();
 sg13g2_decap_4 FILLER_12_349 ();
 sg13g2_fill_2 FILLER_12_353 ();
 sg13g2_decap_8 FILLER_12_381 ();
 sg13g2_decap_8 FILLER_12_388 ();
 sg13g2_decap_8 FILLER_12_395 ();
 sg13g2_decap_8 FILLER_12_402 ();
 sg13g2_decap_8 FILLER_12_409 ();
 sg13g2_decap_8 FILLER_12_416 ();
 sg13g2_decap_8 FILLER_12_423 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_76 ();
 sg13g2_decap_4 FILLER_13_81 ();
 sg13g2_fill_1 FILLER_13_85 ();
 sg13g2_fill_1 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_96 ();
 sg13g2_decap_8 FILLER_13_103 ();
 sg13g2_fill_2 FILLER_13_110 ();
 sg13g2_fill_1 FILLER_13_112 ();
 sg13g2_fill_2 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_165 ();
 sg13g2_fill_1 FILLER_13_167 ();
 sg13g2_fill_2 FILLER_13_172 ();
 sg13g2_fill_1 FILLER_13_174 ();
 sg13g2_fill_2 FILLER_13_180 ();
 sg13g2_fill_1 FILLER_13_182 ();
 sg13g2_fill_2 FILLER_13_195 ();
 sg13g2_fill_2 FILLER_13_207 ();
 sg13g2_fill_1 FILLER_13_209 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_225 ();
 sg13g2_fill_2 FILLER_13_258 ();
 sg13g2_decap_8 FILLER_13_270 ();
 sg13g2_decap_4 FILLER_13_277 ();
 sg13g2_fill_2 FILLER_13_289 ();
 sg13g2_fill_2 FILLER_13_317 ();
 sg13g2_fill_2 FILLER_13_324 ();
 sg13g2_decap_8 FILLER_13_353 ();
 sg13g2_decap_4 FILLER_13_360 ();
 sg13g2_fill_2 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_fill_2 FILLER_13_427 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_decap_8 FILLER_14_71 ();
 sg13g2_decap_4 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_82 ();
 sg13g2_fill_2 FILLER_14_89 ();
 sg13g2_decap_8 FILLER_14_96 ();
 sg13g2_fill_1 FILLER_14_103 ();
 sg13g2_decap_8 FILLER_14_109 ();
 sg13g2_fill_2 FILLER_14_116 ();
 sg13g2_fill_1 FILLER_14_118 ();
 sg13g2_decap_4 FILLER_14_130 ();
 sg13g2_decap_8 FILLER_14_143 ();
 sg13g2_fill_1 FILLER_14_150 ();
 sg13g2_fill_2 FILLER_14_181 ();
 sg13g2_fill_1 FILLER_14_183 ();
 sg13g2_decap_4 FILLER_14_201 ();
 sg13g2_fill_1 FILLER_14_209 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_228 ();
 sg13g2_fill_1 FILLER_14_232 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_decap_4 FILLER_14_251 ();
 sg13g2_decap_8 FILLER_14_286 ();
 sg13g2_decap_8 FILLER_14_293 ();
 sg13g2_decap_8 FILLER_14_304 ();
 sg13g2_decap_8 FILLER_14_311 ();
 sg13g2_fill_1 FILLER_14_318 ();
 sg13g2_fill_2 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_fill_2 FILLER_14_371 ();
 sg13g2_fill_1 FILLER_14_373 ();
 sg13g2_decap_8 FILLER_14_386 ();
 sg13g2_decap_8 FILLER_14_393 ();
 sg13g2_decap_8 FILLER_14_400 ();
 sg13g2_decap_8 FILLER_14_407 ();
 sg13g2_decap_8 FILLER_14_414 ();
 sg13g2_decap_8 FILLER_14_421 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_decap_8 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_35 ();
 sg13g2_fill_2 FILLER_15_42 ();
 sg13g2_decap_4 FILLER_15_48 ();
 sg13g2_decap_8 FILLER_15_69 ();
 sg13g2_decap_4 FILLER_15_76 ();
 sg13g2_fill_2 FILLER_15_80 ();
 sg13g2_decap_8 FILLER_15_89 ();
 sg13g2_decap_8 FILLER_15_145 ();
 sg13g2_decap_8 FILLER_15_152 ();
 sg13g2_decap_4 FILLER_15_163 ();
 sg13g2_fill_2 FILLER_15_167 ();
 sg13g2_decap_8 FILLER_15_175 ();
 sg13g2_decap_4 FILLER_15_182 ();
 sg13g2_fill_2 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_197 ();
 sg13g2_decap_4 FILLER_15_204 ();
 sg13g2_fill_2 FILLER_15_208 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_8 FILLER_15_239 ();
 sg13g2_decap_8 FILLER_15_246 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_4 FILLER_15_294 ();
 sg13g2_fill_1 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_325 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_15_384 ();
 sg13g2_decap_8 FILLER_15_391 ();
 sg13g2_decap_8 FILLER_15_398 ();
 sg13g2_decap_8 FILLER_15_405 ();
 sg13g2_decap_8 FILLER_15_412 ();
 sg13g2_decap_8 FILLER_15_419 ();
 sg13g2_decap_4 FILLER_15_426 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_4 FILLER_16_77 ();
 sg13g2_decap_4 FILLER_16_88 ();
 sg13g2_decap_4 FILLER_16_122 ();
 sg13g2_fill_2 FILLER_16_133 ();
 sg13g2_fill_2 FILLER_16_140 ();
 sg13g2_fill_2 FILLER_16_147 ();
 sg13g2_fill_1 FILLER_16_149 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_163 ();
 sg13g2_fill_1 FILLER_16_165 ();
 sg13g2_decap_4 FILLER_16_170 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_1 FILLER_16_198 ();
 sg13g2_decap_4 FILLER_16_238 ();
 sg13g2_decap_4 FILLER_16_247 ();
 sg13g2_fill_1 FILLER_16_290 ();
 sg13g2_decap_8 FILLER_16_320 ();
 sg13g2_decap_8 FILLER_16_327 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_decap_8 FILLER_16_341 ();
 sg13g2_decap_8 FILLER_16_348 ();
 sg13g2_decap_4 FILLER_16_355 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_8 FILLER_17_35 ();
 sg13g2_decap_8 FILLER_17_42 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_2 FILLER_17_59 ();
 sg13g2_fill_1 FILLER_17_61 ();
 sg13g2_fill_2 FILLER_17_66 ();
 sg13g2_fill_2 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_108 ();
 sg13g2_fill_1 FILLER_17_115 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_129 ();
 sg13g2_fill_2 FILLER_17_156 ();
 sg13g2_fill_1 FILLER_17_158 ();
 sg13g2_fill_2 FILLER_17_185 ();
 sg13g2_fill_1 FILLER_17_187 ();
 sg13g2_decap_4 FILLER_17_287 ();
 sg13g2_fill_1 FILLER_17_291 ();
 sg13g2_fill_2 FILLER_17_300 ();
 sg13g2_decap_4 FILLER_17_341 ();
 sg13g2_fill_1 FILLER_17_345 ();
 sg13g2_decap_4 FILLER_17_353 ();
 sg13g2_fill_2 FILLER_17_357 ();
 sg13g2_decap_8 FILLER_17_385 ();
 sg13g2_decap_8 FILLER_17_392 ();
 sg13g2_decap_8 FILLER_17_399 ();
 sg13g2_decap_8 FILLER_17_406 ();
 sg13g2_decap_8 FILLER_17_413 ();
 sg13g2_decap_8 FILLER_17_420 ();
 sg13g2_fill_2 FILLER_17_427 ();
 sg13g2_fill_1 FILLER_17_429 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_28 ();
 sg13g2_fill_1 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_94 ();
 sg13g2_decap_8 FILLER_18_99 ();
 sg13g2_fill_2 FILLER_18_106 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_2 FILLER_18_218 ();
 sg13g2_decap_4 FILLER_18_224 ();
 sg13g2_fill_2 FILLER_18_231 ();
 sg13g2_fill_1 FILLER_18_233 ();
 sg13g2_fill_1 FILLER_18_240 ();
 sg13g2_fill_1 FILLER_18_247 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_fill_1 FILLER_18_260 ();
 sg13g2_fill_2 FILLER_18_271 ();
 sg13g2_fill_2 FILLER_18_277 ();
 sg13g2_fill_2 FILLER_18_296 ();
 sg13g2_fill_1 FILLER_18_298 ();
 sg13g2_fill_1 FILLER_18_309 ();
 sg13g2_fill_1 FILLER_18_314 ();
 sg13g2_fill_1 FILLER_18_327 ();
 sg13g2_fill_1 FILLER_18_342 ();
 sg13g2_fill_2 FILLER_18_373 ();
 sg13g2_fill_2 FILLER_18_379 ();
 sg13g2_fill_1 FILLER_18_381 ();
 sg13g2_decap_8 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_18_415 ();
 sg13g2_decap_8 FILLER_18_422 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_4 FILLER_19_28 ();
 sg13g2_fill_1 FILLER_19_36 ();
 sg13g2_fill_1 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_74 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_2 FILLER_19_91 ();
 sg13g2_fill_1 FILLER_19_93 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_fill_2 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_112 ();
 sg13g2_decap_4 FILLER_19_123 ();
 sg13g2_decap_4 FILLER_19_132 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_1 FILLER_19_147 ();
 sg13g2_fill_1 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_161 ();
 sg13g2_fill_2 FILLER_19_167 ();
 sg13g2_fill_1 FILLER_19_169 ();
 sg13g2_fill_1 FILLER_19_211 ();
 sg13g2_fill_1 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_221 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_decap_8 FILLER_19_264 ();
 sg13g2_fill_2 FILLER_19_275 ();
 sg13g2_fill_1 FILLER_19_282 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_4 FILLER_19_319 ();
 sg13g2_fill_1 FILLER_19_393 ();
 sg13g2_decap_8 FILLER_19_398 ();
 sg13g2_decap_8 FILLER_19_405 ();
 sg13g2_decap_8 FILLER_19_412 ();
 sg13g2_decap_8 FILLER_19_419 ();
 sg13g2_decap_4 FILLER_19_426 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_8 FILLER_20_28 ();
 sg13g2_decap_8 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_58 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_decap_8 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_80 ();
 sg13g2_decap_4 FILLER_20_121 ();
 sg13g2_fill_1 FILLER_20_155 ();
 sg13g2_fill_1 FILLER_20_160 ();
 sg13g2_fill_2 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_175 ();
 sg13g2_fill_2 FILLER_20_182 ();
 sg13g2_fill_1 FILLER_20_184 ();
 sg13g2_fill_2 FILLER_20_190 ();
 sg13g2_decap_8 FILLER_20_197 ();
 sg13g2_decap_8 FILLER_20_204 ();
 sg13g2_decap_8 FILLER_20_211 ();
 sg13g2_decap_4 FILLER_20_218 ();
 sg13g2_fill_1 FILLER_20_222 ();
 sg13g2_fill_2 FILLER_20_239 ();
 sg13g2_fill_1 FILLER_20_241 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_decap_8 FILLER_20_260 ();
 sg13g2_decap_8 FILLER_20_267 ();
 sg13g2_decap_4 FILLER_20_274 ();
 sg13g2_fill_1 FILLER_20_278 ();
 sg13g2_decap_8 FILLER_20_282 ();
 sg13g2_decap_8 FILLER_20_289 ();
 sg13g2_decap_4 FILLER_20_296 ();
 sg13g2_decap_8 FILLER_20_310 ();
 sg13g2_decap_4 FILLER_20_317 ();
 sg13g2_fill_2 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_349 ();
 sg13g2_fill_1 FILLER_20_351 ();
 sg13g2_decap_4 FILLER_20_359 ();
 sg13g2_fill_1 FILLER_20_363 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_fill_2 FILLER_20_374 ();
 sg13g2_fill_1 FILLER_20_376 ();
 sg13g2_fill_2 FILLER_20_380 ();
 sg13g2_fill_1 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_fill_2 FILLER_21_70 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_fill_2 FILLER_21_122 ();
 sg13g2_fill_1 FILLER_21_124 ();
 sg13g2_decap_4 FILLER_21_128 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_decap_8 FILLER_21_163 ();
 sg13g2_decap_8 FILLER_21_170 ();
 sg13g2_decap_8 FILLER_21_190 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_decap_8 FILLER_21_219 ();
 sg13g2_fill_1 FILLER_21_226 ();
 sg13g2_decap_8 FILLER_21_230 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_fill_1 FILLER_21_244 ();
 sg13g2_fill_1 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_273 ();
 sg13g2_decap_4 FILLER_21_309 ();
 sg13g2_fill_1 FILLER_21_313 ();
 sg13g2_decap_8 FILLER_21_318 ();
 sg13g2_decap_8 FILLER_21_325 ();
 sg13g2_decap_8 FILLER_21_332 ();
 sg13g2_decap_8 FILLER_21_339 ();
 sg13g2_decap_8 FILLER_21_346 ();
 sg13g2_decap_8 FILLER_21_353 ();
 sg13g2_fill_1 FILLER_21_360 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_4 FILLER_21_380 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_decap_8 FILLER_21_390 ();
 sg13g2_decap_8 FILLER_21_397 ();
 sg13g2_decap_8 FILLER_21_404 ();
 sg13g2_decap_8 FILLER_21_411 ();
 sg13g2_decap_8 FILLER_21_418 ();
 sg13g2_decap_4 FILLER_21_425 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_34 ();
 sg13g2_fill_1 FILLER_22_61 ();
 sg13g2_fill_1 FILLER_22_71 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_1 FILLER_22_97 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_fill_2 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_127 ();
 sg13g2_decap_8 FILLER_22_134 ();
 sg13g2_fill_2 FILLER_22_141 ();
 sg13g2_fill_1 FILLER_22_143 ();
 sg13g2_decap_8 FILLER_22_160 ();
 sg13g2_fill_1 FILLER_22_167 ();
 sg13g2_decap_4 FILLER_22_189 ();
 sg13g2_fill_1 FILLER_22_193 ();
 sg13g2_fill_1 FILLER_22_224 ();
 sg13g2_fill_2 FILLER_22_282 ();
 sg13g2_fill_1 FILLER_22_284 ();
 sg13g2_fill_2 FILLER_22_289 ();
 sg13g2_decap_8 FILLER_22_295 ();
 sg13g2_fill_2 FILLER_22_302 ();
 sg13g2_fill_1 FILLER_22_304 ();
 sg13g2_fill_2 FILLER_22_333 ();
 sg13g2_fill_1 FILLER_22_335 ();
 sg13g2_fill_2 FILLER_22_362 ();
 sg13g2_fill_1 FILLER_22_364 ();
 sg13g2_fill_2 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_fill_1 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_409 ();
 sg13g2_decap_8 FILLER_22_416 ();
 sg13g2_decap_8 FILLER_22_423 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_fill_1 FILLER_23_103 ();
 sg13g2_decap_8 FILLER_23_130 ();
 sg13g2_decap_4 FILLER_23_137 ();
 sg13g2_fill_2 FILLER_23_141 ();
 sg13g2_fill_1 FILLER_23_199 ();
 sg13g2_decap_8 FILLER_23_204 ();
 sg13g2_decap_8 FILLER_23_211 ();
 sg13g2_fill_1 FILLER_23_218 ();
 sg13g2_fill_2 FILLER_23_258 ();
 sg13g2_fill_2 FILLER_23_274 ();
 sg13g2_decap_8 FILLER_23_282 ();
 sg13g2_fill_2 FILLER_23_289 ();
 sg13g2_fill_1 FILLER_23_291 ();
 sg13g2_decap_8 FILLER_23_298 ();
 sg13g2_decap_4 FILLER_23_313 ();
 sg13g2_fill_2 FILLER_23_317 ();
 sg13g2_decap_8 FILLER_23_345 ();
 sg13g2_decap_4 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_356 ();
 sg13g2_decap_8 FILLER_23_362 ();
 sg13g2_fill_2 FILLER_23_369 ();
 sg13g2_decap_8 FILLER_23_377 ();
 sg13g2_decap_4 FILLER_23_384 ();
 sg13g2_fill_2 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_decap_8 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_23_415 ();
 sg13g2_decap_8 FILLER_23_422 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_decap_8 FILLER_24_21 ();
 sg13g2_decap_8 FILLER_24_28 ();
 sg13g2_decap_4 FILLER_24_35 ();
 sg13g2_decap_8 FILLER_24_63 ();
 sg13g2_fill_1 FILLER_24_70 ();
 sg13g2_decap_4 FILLER_24_76 ();
 sg13g2_fill_1 FILLER_24_84 ();
 sg13g2_fill_2 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_98 ();
 sg13g2_decap_8 FILLER_24_104 ();
 sg13g2_fill_2 FILLER_24_111 ();
 sg13g2_fill_2 FILLER_24_118 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_fill_2 FILLER_24_137 ();
 sg13g2_fill_1 FILLER_24_139 ();
 sg13g2_fill_2 FILLER_24_149 ();
 sg13g2_fill_1 FILLER_24_151 ();
 sg13g2_fill_1 FILLER_24_157 ();
 sg13g2_decap_8 FILLER_24_162 ();
 sg13g2_decap_4 FILLER_24_169 ();
 sg13g2_decap_4 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_192 ();
 sg13g2_fill_2 FILLER_24_204 ();
 sg13g2_fill_1 FILLER_24_206 ();
 sg13g2_decap_8 FILLER_24_212 ();
 sg13g2_decap_4 FILLER_24_219 ();
 sg13g2_fill_1 FILLER_24_223 ();
 sg13g2_decap_8 FILLER_24_250 ();
 sg13g2_decap_4 FILLER_24_257 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_276 ();
 sg13g2_decap_4 FILLER_24_283 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_decap_8 FILLER_24_292 ();
 sg13g2_fill_1 FILLER_24_299 ();
 sg13g2_fill_2 FILLER_24_304 ();
 sg13g2_decap_8 FILLER_24_315 ();
 sg13g2_fill_2 FILLER_24_322 ();
 sg13g2_fill_1 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_379 ();
 sg13g2_fill_2 FILLER_24_384 ();
 sg13g2_fill_1 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_decap_8 FILLER_25_71 ();
 sg13g2_fill_1 FILLER_25_78 ();
 sg13g2_decap_4 FILLER_25_89 ();
 sg13g2_decap_4 FILLER_25_119 ();
 sg13g2_fill_2 FILLER_25_123 ();
 sg13g2_decap_4 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_141 ();
 sg13g2_fill_1 FILLER_25_150 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_fill_2 FILLER_25_175 ();
 sg13g2_decap_4 FILLER_25_181 ();
 sg13g2_decap_4 FILLER_25_189 ();
 sg13g2_fill_2 FILLER_25_193 ();
 sg13g2_decap_8 FILLER_25_222 ();
 sg13g2_fill_2 FILLER_25_229 ();
 sg13g2_decap_8 FILLER_25_235 ();
 sg13g2_decap_8 FILLER_25_242 ();
 sg13g2_decap_8 FILLER_25_249 ();
 sg13g2_fill_1 FILLER_25_256 ();
 sg13g2_decap_8 FILLER_25_267 ();
 sg13g2_decap_4 FILLER_25_274 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_fill_2 FILLER_25_342 ();
 sg13g2_decap_8 FILLER_25_348 ();
 sg13g2_fill_2 FILLER_25_355 ();
 sg13g2_fill_1 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_362 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_fill_2 FILLER_25_382 ();
 sg13g2_fill_1 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_401 ();
 sg13g2_decap_8 FILLER_25_408 ();
 sg13g2_decap_8 FILLER_25_415 ();
 sg13g2_decap_8 FILLER_25_422 ();
 sg13g2_fill_1 FILLER_25_429 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_4 FILLER_26_28 ();
 sg13g2_fill_1 FILLER_26_32 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_decap_8 FILLER_26_74 ();
 sg13g2_fill_1 FILLER_26_81 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_119 ();
 sg13g2_fill_2 FILLER_26_176 ();
 sg13g2_fill_1 FILLER_26_178 ();
 sg13g2_decap_8 FILLER_26_195 ();
 sg13g2_decap_4 FILLER_26_223 ();
 sg13g2_fill_2 FILLER_26_227 ();
 sg13g2_decap_8 FILLER_26_241 ();
 sg13g2_fill_2 FILLER_26_248 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_269 ();
 sg13g2_decap_8 FILLER_26_274 ();
 sg13g2_decap_8 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_288 ();
 sg13g2_fill_2 FILLER_26_292 ();
 sg13g2_fill_1 FILLER_26_324 ();
 sg13g2_decap_4 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_337 ();
 sg13g2_fill_1 FILLER_26_364 ();
 sg13g2_fill_1 FILLER_26_386 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_8 FILLER_27_7 ();
 sg13g2_decap_8 FILLER_27_14 ();
 sg13g2_decap_8 FILLER_27_21 ();
 sg13g2_decap_4 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_68 ();
 sg13g2_fill_2 FILLER_27_75 ();
 sg13g2_fill_1 FILLER_27_77 ();
 sg13g2_fill_2 FILLER_27_90 ();
 sg13g2_fill_1 FILLER_27_92 ();
 sg13g2_decap_8 FILLER_27_119 ();
 sg13g2_fill_1 FILLER_27_126 ();
 sg13g2_decap_4 FILLER_27_144 ();
 sg13g2_fill_1 FILLER_27_148 ();
 sg13g2_fill_1 FILLER_27_158 ();
 sg13g2_decap_4 FILLER_27_164 ();
 sg13g2_fill_2 FILLER_27_168 ();
 sg13g2_decap_8 FILLER_27_212 ();
 sg13g2_fill_2 FILLER_27_224 ();
 sg13g2_decap_8 FILLER_27_289 ();
 sg13g2_fill_2 FILLER_27_303 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_4 FILLER_27_354 ();
 sg13g2_fill_1 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_378 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_decap_4 FILLER_27_424 ();
 sg13g2_fill_2 FILLER_27_428 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_35 ();
 sg13g2_fill_1 FILLER_28_39 ();
 sg13g2_decap_8 FILLER_28_60 ();
 sg13g2_decap_8 FILLER_28_67 ();
 sg13g2_decap_4 FILLER_28_79 ();
 sg13g2_fill_1 FILLER_28_83 ();
 sg13g2_fill_1 FILLER_28_94 ();
 sg13g2_fill_1 FILLER_28_103 ();
 sg13g2_fill_2 FILLER_28_125 ();
 sg13g2_fill_1 FILLER_28_127 ();
 sg13g2_decap_4 FILLER_28_137 ();
 sg13g2_decap_8 FILLER_28_145 ();
 sg13g2_decap_8 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_169 ();
 sg13g2_fill_2 FILLER_28_191 ();
 sg13g2_decap_4 FILLER_28_197 ();
 sg13g2_decap_4 FILLER_28_222 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_4 FILLER_28_242 ();
 sg13g2_decap_8 FILLER_28_251 ();
 sg13g2_decap_8 FILLER_28_258 ();
 sg13g2_fill_1 FILLER_28_274 ();
 sg13g2_fill_1 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_310 ();
 sg13g2_decap_8 FILLER_28_317 ();
 sg13g2_decap_4 FILLER_28_324 ();
 sg13g2_decap_8 FILLER_28_332 ();
 sg13g2_decap_8 FILLER_28_339 ();
 sg13g2_decap_8 FILLER_28_346 ();
 sg13g2_decap_4 FILLER_28_353 ();
 sg13g2_decap_4 FILLER_28_361 ();
 sg13g2_fill_1 FILLER_28_404 ();
 sg13g2_decap_8 FILLER_28_411 ();
 sg13g2_decap_8 FILLER_28_418 ();
 sg13g2_decap_4 FILLER_28_425 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_decap_8 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_14 ();
 sg13g2_decap_8 FILLER_29_21 ();
 sg13g2_decap_8 FILLER_29_28 ();
 sg13g2_decap_8 FILLER_29_35 ();
 sg13g2_decap_8 FILLER_29_42 ();
 sg13g2_decap_8 FILLER_29_49 ();
 sg13g2_decap_8 FILLER_29_56 ();
 sg13g2_fill_2 FILLER_29_63 ();
 sg13g2_fill_1 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_103 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_decap_4 FILLER_29_117 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_4 FILLER_29_151 ();
 sg13g2_fill_2 FILLER_29_155 ();
 sg13g2_decap_4 FILLER_29_165 ();
 sg13g2_fill_2 FILLER_29_169 ();
 sg13g2_fill_2 FILLER_29_181 ();
 sg13g2_fill_1 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_213 ();
 sg13g2_decap_8 FILLER_29_220 ();
 sg13g2_fill_2 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_4 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_decap_4 FILLER_29_259 ();
 sg13g2_fill_1 FILLER_29_263 ();
 sg13g2_fill_2 FILLER_29_345 ();
 sg13g2_fill_1 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_377 ();
 sg13g2_decap_4 FILLER_29_394 ();
 sg13g2_decap_8 FILLER_29_401 ();
 sg13g2_decap_8 FILLER_29_408 ();
 sg13g2_decap_8 FILLER_29_415 ();
 sg13g2_decap_8 FILLER_29_422 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_4 FILLER_30_42 ();
 sg13g2_fill_2 FILLER_30_50 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_fill_2 FILLER_30_59 ();
 sg13g2_fill_1 FILLER_30_61 ();
 sg13g2_decap_8 FILLER_30_68 ();
 sg13g2_decap_4 FILLER_30_75 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_109 ();
 sg13g2_decap_8 FILLER_30_116 ();
 sg13g2_decap_8 FILLER_30_123 ();
 sg13g2_decap_8 FILLER_30_130 ();
 sg13g2_fill_2 FILLER_30_137 ();
 sg13g2_fill_1 FILLER_30_142 ();
 sg13g2_decap_4 FILLER_30_161 ();
 sg13g2_fill_2 FILLER_30_170 ();
 sg13g2_fill_1 FILLER_30_172 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_fill_1 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_221 ();
 sg13g2_decap_8 FILLER_30_260 ();
 sg13g2_decap_8 FILLER_30_267 ();
 sg13g2_decap_4 FILLER_30_274 ();
 sg13g2_fill_2 FILLER_30_278 ();
 sg13g2_decap_8 FILLER_30_288 ();
 sg13g2_decap_8 FILLER_30_295 ();
 sg13g2_decap_8 FILLER_30_302 ();
 sg13g2_decap_8 FILLER_30_309 ();
 sg13g2_decap_4 FILLER_30_316 ();
 sg13g2_fill_1 FILLER_30_383 ();
 sg13g2_decap_4 FILLER_30_394 ();
 sg13g2_fill_1 FILLER_30_398 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_fill_2 FILLER_31_35 ();
 sg13g2_fill_2 FILLER_31_67 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_decap_4 FILLER_31_90 ();
 sg13g2_fill_1 FILLER_31_94 ();
 sg13g2_fill_1 FILLER_31_100 ();
 sg13g2_fill_2 FILLER_31_105 ();
 sg13g2_fill_2 FILLER_31_112 ();
 sg13g2_fill_2 FILLER_31_120 ();
 sg13g2_fill_2 FILLER_31_164 ();
 sg13g2_decap_8 FILLER_31_170 ();
 sg13g2_decap_4 FILLER_31_177 ();
 sg13g2_fill_2 FILLER_31_187 ();
 sg13g2_decap_8 FILLER_31_215 ();
 sg13g2_fill_1 FILLER_31_222 ();
 sg13g2_decap_4 FILLER_31_264 ();
 sg13g2_fill_2 FILLER_31_268 ();
 sg13g2_decap_4 FILLER_31_278 ();
 sg13g2_decap_8 FILLER_31_291 ();
 sg13g2_decap_8 FILLER_31_298 ();
 sg13g2_decap_4 FILLER_31_305 ();
 sg13g2_fill_2 FILLER_31_309 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_341 ();
 sg13g2_fill_1 FILLER_31_343 ();
 sg13g2_fill_2 FILLER_31_347 ();
 sg13g2_decap_4 FILLER_31_375 ();
 sg13g2_fill_2 FILLER_31_389 ();
 sg13g2_fill_1 FILLER_31_412 ();
 sg13g2_decap_8 FILLER_31_419 ();
 sg13g2_decap_4 FILLER_31_426 ();
 sg13g2_decap_8 FILLER_32_0 ();
 sg13g2_decap_8 FILLER_32_7 ();
 sg13g2_decap_8 FILLER_32_14 ();
 sg13g2_decap_8 FILLER_32_21 ();
 sg13g2_decap_8 FILLER_32_28 ();
 sg13g2_decap_8 FILLER_32_35 ();
 sg13g2_fill_2 FILLER_32_46 ();
 sg13g2_decap_4 FILLER_32_74 ();
 sg13g2_decap_4 FILLER_32_83 ();
 sg13g2_fill_2 FILLER_32_92 ();
 sg13g2_fill_1 FILLER_32_94 ();
 sg13g2_fill_1 FILLER_32_134 ();
 sg13g2_decap_4 FILLER_32_139 ();
 sg13g2_fill_1 FILLER_32_143 ();
 sg13g2_fill_1 FILLER_32_179 ();
 sg13g2_fill_2 FILLER_32_185 ();
 sg13g2_fill_1 FILLER_32_187 ();
 sg13g2_fill_2 FILLER_32_192 ();
 sg13g2_fill_2 FILLER_32_198 ();
 sg13g2_fill_1 FILLER_32_200 ();
 sg13g2_decap_4 FILLER_32_222 ();
 sg13g2_fill_2 FILLER_32_226 ();
 sg13g2_fill_2 FILLER_32_232 ();
 sg13g2_decap_8 FILLER_32_240 ();
 sg13g2_fill_2 FILLER_32_247 ();
 sg13g2_fill_1 FILLER_32_249 ();
 sg13g2_fill_2 FILLER_32_285 ();
 sg13g2_fill_1 FILLER_32_287 ();
 sg13g2_decap_4 FILLER_32_321 ();
 sg13g2_decap_8 FILLER_32_329 ();
 sg13g2_decap_4 FILLER_32_336 ();
 sg13g2_decap_8 FILLER_32_358 ();
 sg13g2_decap_8 FILLER_32_365 ();
 sg13g2_fill_2 FILLER_32_372 ();
 sg13g2_decap_8 FILLER_32_379 ();
 sg13g2_decap_8 FILLER_32_386 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_fill_1 FILLER_32_398 ();
 sg13g2_decap_8 FILLER_32_420 ();
 sg13g2_fill_2 FILLER_32_427 ();
 sg13g2_fill_1 FILLER_32_429 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_fill_1 FILLER_33_56 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_83 ();
 sg13g2_fill_1 FILLER_33_114 ();
 sg13g2_fill_2 FILLER_33_119 ();
 sg13g2_fill_1 FILLER_33_121 ();
 sg13g2_decap_8 FILLER_33_136 ();
 sg13g2_decap_8 FILLER_33_143 ();
 sg13g2_decap_8 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_209 ();
 sg13g2_fill_1 FILLER_33_211 ();
 sg13g2_decap_8 FILLER_33_233 ();
 sg13g2_decap_4 FILLER_33_240 ();
 sg13g2_decap_8 FILLER_33_249 ();
 sg13g2_fill_2 FILLER_33_256 ();
 sg13g2_decap_8 FILLER_33_262 ();
 sg13g2_decap_4 FILLER_33_269 ();
 sg13g2_fill_2 FILLER_33_273 ();
 sg13g2_fill_2 FILLER_33_284 ();
 sg13g2_decap_4 FILLER_33_291 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_fill_1 FILLER_33_304 ();
 sg13g2_fill_2 FILLER_33_311 ();
 sg13g2_fill_2 FILLER_33_317 ();
 sg13g2_fill_1 FILLER_33_331 ();
 sg13g2_fill_2 FILLER_33_335 ();
 sg13g2_fill_1 FILLER_33_363 ();
 sg13g2_fill_2 FILLER_33_385 ();
 sg13g2_fill_1 FILLER_33_392 ();
 sg13g2_fill_2 FILLER_33_398 ();
 sg13g2_decap_8 FILLER_33_403 ();
 sg13g2_fill_2 FILLER_33_410 ();
 sg13g2_decap_8 FILLER_33_417 ();
 sg13g2_decap_4 FILLER_33_424 ();
 sg13g2_fill_2 FILLER_33_428 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_14 ();
 sg13g2_decap_8 FILLER_34_21 ();
 sg13g2_decap_8 FILLER_34_28 ();
 sg13g2_decap_8 FILLER_34_35 ();
 sg13g2_fill_1 FILLER_34_51 ();
 sg13g2_fill_1 FILLER_34_56 ();
 sg13g2_decap_4 FILLER_34_61 ();
 sg13g2_decap_4 FILLER_34_86 ();
 sg13g2_decap_4 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_133 ();
 sg13g2_decap_8 FILLER_34_140 ();
 sg13g2_fill_2 FILLER_34_147 ();
 sg13g2_fill_1 FILLER_34_149 ();
 sg13g2_decap_8 FILLER_34_202 ();
 sg13g2_decap_8 FILLER_34_209 ();
 sg13g2_decap_4 FILLER_34_216 ();
 sg13g2_fill_1 FILLER_34_220 ();
 sg13g2_decap_8 FILLER_34_229 ();
 sg13g2_decap_8 FILLER_34_236 ();
 sg13g2_decap_8 FILLER_34_243 ();
 sg13g2_decap_8 FILLER_34_250 ();
 sg13g2_decap_4 FILLER_34_257 ();
 sg13g2_decap_8 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_272 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_2 FILLER_34_368 ();
 sg13g2_fill_1 FILLER_34_370 ();
 sg13g2_fill_1 FILLER_34_424 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_fill_1 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_62 ();
 sg13g2_decap_8 FILLER_35_69 ();
 sg13g2_decap_8 FILLER_35_76 ();
 sg13g2_decap_8 FILLER_35_83 ();
 sg13g2_decap_8 FILLER_35_90 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_1 FILLER_35_159 ();
 sg13g2_decap_4 FILLER_35_164 ();
 sg13g2_fill_1 FILLER_35_176 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_1 FILLER_35_218 ();
 sg13g2_decap_8 FILLER_35_223 ();
 sg13g2_fill_1 FILLER_35_230 ();
 sg13g2_fill_1 FILLER_35_237 ();
 sg13g2_decap_8 FILLER_35_264 ();
 sg13g2_decap_8 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_278 ();
 sg13g2_decap_4 FILLER_35_284 ();
 sg13g2_fill_2 FILLER_35_288 ();
 sg13g2_decap_4 FILLER_35_293 ();
 sg13g2_fill_1 FILLER_35_297 ();
 sg13g2_decap_8 FILLER_35_302 ();
 sg13g2_decap_8 FILLER_35_327 ();
 sg13g2_decap_4 FILLER_35_334 ();
 sg13g2_fill_2 FILLER_35_338 ();
 sg13g2_decap_4 FILLER_35_347 ();
 sg13g2_decap_8 FILLER_35_355 ();
 sg13g2_decap_8 FILLER_35_362 ();
 sg13g2_decap_4 FILLER_35_369 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_419 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_4 FILLER_36_42 ();
 sg13g2_fill_2 FILLER_36_46 ();
 sg13g2_decap_8 FILLER_36_64 ();
 sg13g2_decap_8 FILLER_36_71 ();
 sg13g2_decap_8 FILLER_36_78 ();
 sg13g2_decap_4 FILLER_36_85 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_1 FILLER_36_104 ();
 sg13g2_fill_1 FILLER_36_109 ();
 sg13g2_fill_1 FILLER_36_113 ();
 sg13g2_fill_1 FILLER_36_148 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_1 FILLER_36_195 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_4 FILLER_36_212 ();
 sg13g2_fill_2 FILLER_36_216 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_269 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_fill_2 FILLER_36_315 ();
 sg13g2_fill_1 FILLER_36_317 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_4 FILLER_36_371 ();
 sg13g2_fill_2 FILLER_36_382 ();
 sg13g2_decap_8 FILLER_36_397 ();
 sg13g2_fill_2 FILLER_36_409 ();
 sg13g2_fill_1 FILLER_36_411 ();
 sg13g2_fill_2 FILLER_36_427 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_decap_8 FILLER_37_7 ();
 sg13g2_decap_8 FILLER_37_14 ();
 sg13g2_decap_8 FILLER_37_21 ();
 sg13g2_decap_4 FILLER_37_28 ();
 sg13g2_fill_2 FILLER_37_32 ();
 sg13g2_fill_2 FILLER_37_38 ();
 sg13g2_fill_2 FILLER_37_66 ();
 sg13g2_fill_1 FILLER_37_68 ();
 sg13g2_fill_2 FILLER_37_90 ();
 sg13g2_fill_1 FILLER_37_92 ();
 sg13g2_fill_2 FILLER_37_119 ();
 sg13g2_fill_1 FILLER_37_121 ();
 sg13g2_decap_4 FILLER_37_126 ();
 sg13g2_fill_1 FILLER_37_130 ();
 sg13g2_fill_1 FILLER_37_157 ();
 sg13g2_decap_8 FILLER_37_167 ();
 sg13g2_decap_8 FILLER_37_174 ();
 sg13g2_fill_2 FILLER_37_181 ();
 sg13g2_fill_2 FILLER_37_272 ();
 sg13g2_decap_8 FILLER_37_299 ();
 sg13g2_decap_8 FILLER_37_306 ();
 sg13g2_decap_8 FILLER_37_313 ();
 sg13g2_decap_4 FILLER_37_320 ();
 sg13g2_fill_1 FILLER_37_350 ();
 sg13g2_fill_2 FILLER_37_372 ();
 sg13g2_fill_2 FILLER_37_381 ();
 sg13g2_fill_1 FILLER_37_383 ();
 sg13g2_decap_4 FILLER_37_391 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_416 ();
 sg13g2_fill_1 FILLER_37_418 ();
 sg13g2_decap_4 FILLER_37_424 ();
 sg13g2_fill_2 FILLER_37_428 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_fill_2 FILLER_38_42 ();
 sg13g2_fill_1 FILLER_38_44 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_4 FILLER_38_63 ();
 sg13g2_fill_1 FILLER_38_67 ();
 sg13g2_fill_2 FILLER_38_94 ();
 sg13g2_fill_1 FILLER_38_96 ();
 sg13g2_decap_8 FILLER_38_122 ();
 sg13g2_decap_8 FILLER_38_129 ();
 sg13g2_decap_8 FILLER_38_136 ();
 sg13g2_decap_4 FILLER_38_143 ();
 sg13g2_fill_2 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_170 ();
 sg13g2_fill_2 FILLER_38_177 ();
 sg13g2_fill_1 FILLER_38_179 ();
 sg13g2_fill_2 FILLER_38_190 ();
 sg13g2_fill_1 FILLER_38_192 ();
 sg13g2_decap_4 FILLER_38_197 ();
 sg13g2_decap_4 FILLER_38_210 ();
 sg13g2_fill_1 FILLER_38_221 ();
 sg13g2_fill_2 FILLER_38_228 ();
 sg13g2_fill_1 FILLER_38_230 ();
 sg13g2_fill_2 FILLER_38_236 ();
 sg13g2_fill_1 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_2 FILLER_38_304 ();
 sg13g2_fill_2 FILLER_38_317 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_decap_4 FILLER_38_324 ();
 sg13g2_fill_1 FILLER_38_400 ();
 sg13g2_fill_2 FILLER_38_409 ();
 sg13g2_fill_1 FILLER_38_411 ();
 sg13g2_decap_4 FILLER_38_425 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_decap_8 FILLER_39_14 ();
 sg13g2_decap_8 FILLER_39_21 ();
 sg13g2_decap_8 FILLER_39_28 ();
 sg13g2_decap_8 FILLER_39_35 ();
 sg13g2_decap_4 FILLER_39_42 ();
 sg13g2_fill_1 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_81 ();
 sg13g2_fill_2 FILLER_39_88 ();
 sg13g2_fill_2 FILLER_39_95 ();
 sg13g2_decap_4 FILLER_39_106 ();
 sg13g2_fill_2 FILLER_39_110 ();
 sg13g2_fill_1 FILLER_39_123 ();
 sg13g2_decap_4 FILLER_39_128 ();
 sg13g2_decap_8 FILLER_39_136 ();
 sg13g2_decap_8 FILLER_39_143 ();
 sg13g2_decap_8 FILLER_39_150 ();
 sg13g2_decap_8 FILLER_39_157 ();
 sg13g2_decap_8 FILLER_39_164 ();
 sg13g2_decap_8 FILLER_39_171 ();
 sg13g2_fill_2 FILLER_39_178 ();
 sg13g2_fill_1 FILLER_39_180 ();
 sg13g2_fill_1 FILLER_39_194 ();
 sg13g2_fill_1 FILLER_39_209 ();
 sg13g2_decap_4 FILLER_39_214 ();
 sg13g2_fill_1 FILLER_39_218 ();
 sg13g2_decap_4 FILLER_39_231 ();
 sg13g2_decap_8 FILLER_39_245 ();
 sg13g2_fill_2 FILLER_39_256 ();
 sg13g2_fill_1 FILLER_39_258 ();
 sg13g2_fill_1 FILLER_39_263 ();
 sg13g2_fill_1 FILLER_39_294 ();
 sg13g2_fill_2 FILLER_39_299 ();
 sg13g2_fill_2 FILLER_39_309 ();
 sg13g2_decap_8 FILLER_39_337 ();
 sg13g2_fill_1 FILLER_39_356 ();
 sg13g2_decap_8 FILLER_39_361 ();
 sg13g2_decap_4 FILLER_39_376 ();
 sg13g2_fill_1 FILLER_39_380 ();
 sg13g2_decap_8 FILLER_39_391 ();
 sg13g2_decap_8 FILLER_39_398 ();
 sg13g2_fill_1 FILLER_39_405 ();
 sg13g2_fill_1 FILLER_39_416 ();
 sg13g2_decap_8 FILLER_39_422 ();
 sg13g2_fill_1 FILLER_39_429 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_fill_1 FILLER_40_74 ();
 sg13g2_fill_1 FILLER_40_79 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_fill_1 FILLER_40_91 ();
 sg13g2_fill_2 FILLER_40_118 ();
 sg13g2_decap_4 FILLER_40_146 ();
 sg13g2_fill_2 FILLER_40_155 ();
 sg13g2_fill_1 FILLER_40_157 ();
 sg13g2_fill_2 FILLER_40_184 ();
 sg13g2_fill_2 FILLER_40_191 ();
 sg13g2_fill_2 FILLER_40_202 ();
 sg13g2_fill_1 FILLER_40_204 ();
 sg13g2_decap_8 FILLER_40_235 ();
 sg13g2_decap_8 FILLER_40_242 ();
 sg13g2_decap_8 FILLER_40_249 ();
 sg13g2_fill_1 FILLER_40_256 ();
 sg13g2_decap_8 FILLER_40_262 ();
 sg13g2_decap_4 FILLER_40_269 ();
 sg13g2_fill_2 FILLER_40_273 ();
 sg13g2_decap_4 FILLER_40_286 ();
 sg13g2_decap_8 FILLER_40_317 ();
 sg13g2_decap_4 FILLER_40_324 ();
 sg13g2_fill_2 FILLER_40_328 ();
 sg13g2_decap_8 FILLER_40_335 ();
 sg13g2_decap_8 FILLER_40_342 ();
 sg13g2_decap_8 FILLER_40_349 ();
 sg13g2_decap_8 FILLER_40_362 ();
 sg13g2_decap_8 FILLER_40_369 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_fill_1 FILLER_40_378 ();
 sg13g2_decap_4 FILLER_40_394 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_fill_2 FILLER_40_403 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_fill_2 FILLER_40_427 ();
 sg13g2_fill_1 FILLER_40_429 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_fill_2 FILLER_41_49 ();
 sg13g2_decap_4 FILLER_41_55 ();
 sg13g2_fill_2 FILLER_41_59 ();
 sg13g2_decap_4 FILLER_41_92 ();
 sg13g2_fill_2 FILLER_41_96 ();
 sg13g2_decap_8 FILLER_41_102 ();
 sg13g2_decap_8 FILLER_41_109 ();
 sg13g2_fill_1 FILLER_41_126 ();
 sg13g2_fill_2 FILLER_41_131 ();
 sg13g2_fill_2 FILLER_41_136 ();
 sg13g2_fill_1 FILLER_41_150 ();
 sg13g2_fill_1 FILLER_41_167 ();
 sg13g2_decap_8 FILLER_41_172 ();
 sg13g2_fill_1 FILLER_41_185 ();
 sg13g2_fill_2 FILLER_41_190 ();
 sg13g2_fill_1 FILLER_41_196 ();
 sg13g2_fill_2 FILLER_41_202 ();
 sg13g2_fill_2 FILLER_41_209 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_4 FILLER_41_259 ();
 sg13g2_fill_2 FILLER_41_263 ();
 sg13g2_fill_2 FILLER_41_301 ();
 sg13g2_fill_1 FILLER_41_303 ();
 sg13g2_fill_2 FILLER_41_351 ();
 sg13g2_fill_1 FILLER_41_353 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_4 FILLER_41_378 ();
 sg13g2_fill_2 FILLER_41_382 ();
 sg13g2_fill_1 FILLER_41_399 ();
 sg13g2_fill_1 FILLER_41_404 ();
 sg13g2_decap_4 FILLER_41_425 ();
 sg13g2_fill_1 FILLER_41_429 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_decap_8 FILLER_42_7 ();
 sg13g2_decap_8 FILLER_42_14 ();
 sg13g2_decap_8 FILLER_42_21 ();
 sg13g2_decap_8 FILLER_42_28 ();
 sg13g2_decap_8 FILLER_42_35 ();
 sg13g2_decap_8 FILLER_42_42 ();
 sg13g2_decap_8 FILLER_42_49 ();
 sg13g2_decap_8 FILLER_42_56 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_108 ();
 sg13g2_fill_1 FILLER_42_110 ();
 sg13g2_decap_8 FILLER_42_153 ();
 sg13g2_decap_4 FILLER_42_160 ();
 sg13g2_fill_1 FILLER_42_164 ();
 sg13g2_fill_1 FILLER_42_186 ();
 sg13g2_fill_2 FILLER_42_213 ();
 sg13g2_fill_1 FILLER_42_228 ();
 sg13g2_decap_8 FILLER_42_265 ();
 sg13g2_fill_2 FILLER_42_293 ();
 sg13g2_fill_2 FILLER_42_301 ();
 sg13g2_fill_1 FILLER_42_303 ();
 sg13g2_fill_2 FILLER_42_308 ();
 sg13g2_fill_1 FILLER_42_310 ();
 sg13g2_fill_2 FILLER_42_325 ();
 sg13g2_fill_2 FILLER_42_338 ();
 sg13g2_decap_8 FILLER_42_361 ();
 sg13g2_decap_4 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_372 ();
 sg13g2_decap_4 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_382 ();
 sg13g2_fill_1 FILLER_42_388 ();
 sg13g2_decap_8 FILLER_42_404 ();
 sg13g2_fill_2 FILLER_42_411 ();
 sg13g2_decap_4 FILLER_42_424 ();
 sg13g2_fill_2 FILLER_42_428 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_fill_2 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_100 ();
 sg13g2_decap_8 FILLER_43_107 ();
 sg13g2_decap_8 FILLER_43_114 ();
 sg13g2_decap_8 FILLER_43_121 ();
 sg13g2_fill_2 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_130 ();
 sg13g2_decap_8 FILLER_43_152 ();
 sg13g2_decap_8 FILLER_43_188 ();
 sg13g2_fill_2 FILLER_43_199 ();
 sg13g2_fill_1 FILLER_43_201 ();
 sg13g2_fill_1 FILLER_43_208 ();
 sg13g2_decap_8 FILLER_43_213 ();
 sg13g2_decap_8 FILLER_43_220 ();
 sg13g2_decap_8 FILLER_43_227 ();
 sg13g2_decap_8 FILLER_43_234 ();
 sg13g2_decap_4 FILLER_43_241 ();
 sg13g2_fill_2 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_251 ();
 sg13g2_decap_8 FILLER_43_258 ();
 sg13g2_decap_8 FILLER_43_286 ();
 sg13g2_decap_8 FILLER_43_293 ();
 sg13g2_decap_4 FILLER_43_300 ();
 sg13g2_decap_8 FILLER_43_312 ();
 sg13g2_decap_8 FILLER_43_319 ();
 sg13g2_fill_1 FILLER_43_326 ();
 sg13g2_decap_8 FILLER_43_340 ();
 sg13g2_decap_4 FILLER_43_347 ();
 sg13g2_fill_2 FILLER_43_351 ();
 sg13g2_decap_4 FILLER_43_361 ();
 sg13g2_decap_4 FILLER_43_372 ();
 sg13g2_fill_1 FILLER_43_376 ();
 sg13g2_fill_1 FILLER_43_403 ();
 sg13g2_decap_8 FILLER_43_418 ();
 sg13g2_decap_4 FILLER_43_425 ();
 sg13g2_fill_1 FILLER_43_429 ();
 sg13g2_decap_8 FILLER_44_0 ();
 sg13g2_decap_8 FILLER_44_7 ();
 sg13g2_decap_8 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_21 ();
 sg13g2_decap_8 FILLER_44_28 ();
 sg13g2_decap_8 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_42 ();
 sg13g2_fill_1 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_61 ();
 sg13g2_decap_4 FILLER_44_68 ();
 sg13g2_decap_8 FILLER_44_93 ();
 sg13g2_decap_8 FILLER_44_100 ();
 sg13g2_decap_8 FILLER_44_107 ();
 sg13g2_decap_8 FILLER_44_118 ();
 sg13g2_decap_8 FILLER_44_125 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_1 FILLER_44_134 ();
 sg13g2_decap_8 FILLER_44_139 ();
 sg13g2_decap_8 FILLER_44_146 ();
 sg13g2_fill_2 FILLER_44_153 ();
 sg13g2_fill_1 FILLER_44_155 ();
 sg13g2_decap_8 FILLER_44_191 ();
 sg13g2_decap_4 FILLER_44_198 ();
 sg13g2_fill_2 FILLER_44_202 ();
 sg13g2_decap_8 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_217 ();
 sg13g2_decap_8 FILLER_44_223 ();
 sg13g2_decap_4 FILLER_44_230 ();
 sg13g2_decap_8 FILLER_44_239 ();
 sg13g2_fill_1 FILLER_44_246 ();
 sg13g2_decap_8 FILLER_44_253 ();
 sg13g2_decap_4 FILLER_44_260 ();
 sg13g2_decap_8 FILLER_44_285 ();
 sg13g2_fill_2 FILLER_44_292 ();
 sg13g2_fill_1 FILLER_44_294 ();
 sg13g2_decap_8 FILLER_44_306 ();
 sg13g2_decap_8 FILLER_44_313 ();
 sg13g2_decap_8 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_327 ();
 sg13g2_fill_1 FILLER_44_329 ();
 sg13g2_fill_1 FILLER_44_367 ();
 sg13g2_fill_2 FILLER_44_372 ();
 sg13g2_fill_1 FILLER_44_378 ();
 sg13g2_fill_2 FILLER_44_384 ();
 sg13g2_fill_1 FILLER_44_390 ();
 sg13g2_decap_8 FILLER_44_404 ();
 sg13g2_decap_8 FILLER_44_411 ();
 sg13g2_decap_8 FILLER_44_418 ();
 sg13g2_decap_4 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_72 ();
 sg13g2_decap_8 FILLER_45_79 ();
 sg13g2_decap_8 FILLER_45_86 ();
 sg13g2_fill_2 FILLER_45_93 ();
 sg13g2_fill_1 FILLER_45_124 ();
 sg13g2_decap_4 FILLER_45_130 ();
 sg13g2_fill_2 FILLER_45_134 ();
 sg13g2_decap_4 FILLER_45_144 ();
 sg13g2_fill_2 FILLER_45_148 ();
 sg13g2_fill_2 FILLER_45_166 ();
 sg13g2_fill_1 FILLER_45_168 ();
 sg13g2_fill_2 FILLER_45_175 ();
 sg13g2_fill_1 FILLER_45_177 ();
 sg13g2_decap_8 FILLER_45_212 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_decap_8 FILLER_45_263 ();
 sg13g2_decap_8 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_277 ();
 sg13g2_fill_1 FILLER_45_284 ();
 sg13g2_fill_2 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_306 ();
 sg13g2_decap_8 FILLER_45_312 ();
 sg13g2_decap_4 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_323 ();
 sg13g2_fill_1 FILLER_45_350 ();
 sg13g2_fill_1 FILLER_45_355 ();
 sg13g2_fill_1 FILLER_45_362 ();
 sg13g2_fill_1 FILLER_45_373 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_387 ();
 sg13g2_fill_1 FILLER_45_396 ();
 sg13g2_decap_8 FILLER_45_410 ();
 sg13g2_decap_8 FILLER_45_417 ();
 sg13g2_decap_4 FILLER_45_424 ();
 sg13g2_fill_2 FILLER_45_428 ();
 sg13g2_decap_8 FILLER_46_0 ();
 sg13g2_decap_8 FILLER_46_7 ();
 sg13g2_decap_8 FILLER_46_14 ();
 sg13g2_decap_8 FILLER_46_21 ();
 sg13g2_decap_8 FILLER_46_28 ();
 sg13g2_decap_8 FILLER_46_35 ();
 sg13g2_fill_1 FILLER_46_72 ();
 sg13g2_decap_8 FILLER_46_78 ();
 sg13g2_fill_2 FILLER_46_85 ();
 sg13g2_fill_1 FILLER_46_87 ();
 sg13g2_fill_1 FILLER_46_117 ();
 sg13g2_fill_1 FILLER_46_153 ();
 sg13g2_fill_1 FILLER_46_159 ();
 sg13g2_fill_1 FILLER_46_164 ();
 sg13g2_decap_4 FILLER_46_201 ();
 sg13g2_fill_2 FILLER_46_212 ();
 sg13g2_decap_4 FILLER_46_240 ();
 sg13g2_fill_2 FILLER_46_244 ();
 sg13g2_decap_8 FILLER_46_256 ();
 sg13g2_fill_1 FILLER_46_263 ();
 sg13g2_decap_8 FILLER_46_280 ();
 sg13g2_decap_4 FILLER_46_287 ();
 sg13g2_fill_2 FILLER_46_291 ();
 sg13g2_decap_8 FILLER_46_327 ();
 sg13g2_decap_8 FILLER_46_334 ();
 sg13g2_decap_8 FILLER_46_341 ();
 sg13g2_decap_4 FILLER_46_348 ();
 sg13g2_decap_4 FILLER_46_364 ();
 sg13g2_fill_1 FILLER_46_368 ();
 sg13g2_fill_2 FILLER_46_373 ();
 sg13g2_decap_8 FILLER_46_379 ();
 sg13g2_decap_8 FILLER_46_386 ();
 sg13g2_decap_4 FILLER_46_393 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_decap_8 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_4 FILLER_46_424 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_4 FILLER_47_42 ();
 sg13g2_fill_1 FILLER_47_46 ();
 sg13g2_decap_8 FILLER_47_61 ();
 sg13g2_fill_1 FILLER_47_68 ();
 sg13g2_decap_8 FILLER_47_73 ();
 sg13g2_decap_8 FILLER_47_80 ();
 sg13g2_decap_8 FILLER_47_87 ();
 sg13g2_fill_1 FILLER_47_94 ();
 sg13g2_fill_1 FILLER_47_103 ();
 sg13g2_fill_2 FILLER_47_125 ();
 sg13g2_decap_8 FILLER_47_131 ();
 sg13g2_decap_8 FILLER_47_138 ();
 sg13g2_fill_2 FILLER_47_145 ();
 sg13g2_fill_1 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_157 ();
 sg13g2_decap_8 FILLER_47_164 ();
 sg13g2_decap_4 FILLER_47_171 ();
 sg13g2_fill_1 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_180 ();
 sg13g2_decap_8 FILLER_47_212 ();
 sg13g2_fill_1 FILLER_47_219 ();
 sg13g2_decap_8 FILLER_47_228 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_fill_2 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_244 ();
 sg13g2_fill_2 FILLER_47_251 ();
 sg13g2_fill_1 FILLER_47_253 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_fill_1 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_333 ();
 sg13g2_decap_8 FILLER_47_340 ();
 sg13g2_decap_8 FILLER_47_347 ();
 sg13g2_decap_8 FILLER_47_354 ();
 sg13g2_decap_8 FILLER_47_361 ();
 sg13g2_decap_8 FILLER_47_368 ();
 sg13g2_decap_8 FILLER_47_375 ();
 sg13g2_decap_4 FILLER_47_382 ();
 sg13g2_fill_1 FILLER_47_386 ();
 sg13g2_decap_4 FILLER_47_392 ();
 sg13g2_fill_1 FILLER_47_396 ();
 sg13g2_fill_2 FILLER_47_411 ();
 sg13g2_fill_1 FILLER_47_413 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_56 ();
 sg13g2_fill_1 FILLER_48_58 ();
 sg13g2_decap_8 FILLER_48_95 ();
 sg13g2_decap_8 FILLER_48_102 ();
 sg13g2_decap_8 FILLER_48_109 ();
 sg13g2_decap_8 FILLER_48_116 ();
 sg13g2_decap_8 FILLER_48_123 ();
 sg13g2_decap_8 FILLER_48_130 ();
 sg13g2_decap_8 FILLER_48_137 ();
 sg13g2_decap_4 FILLER_48_144 ();
 sg13g2_fill_1 FILLER_48_148 ();
 sg13g2_fill_2 FILLER_48_162 ();
 sg13g2_fill_1 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_180 ();
 sg13g2_decap_8 FILLER_48_187 ();
 sg13g2_decap_8 FILLER_48_194 ();
 sg13g2_fill_2 FILLER_48_201 ();
 sg13g2_fill_2 FILLER_48_208 ();
 sg13g2_decap_8 FILLER_48_221 ();
 sg13g2_decap_4 FILLER_48_228 ();
 sg13g2_fill_2 FILLER_48_232 ();
 sg13g2_decap_8 FILLER_48_240 ();
 sg13g2_fill_1 FILLER_48_247 ();
 sg13g2_fill_1 FILLER_48_253 ();
 sg13g2_decap_8 FILLER_48_263 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_2 FILLER_48_276 ();
 sg13g2_decap_4 FILLER_48_282 ();
 sg13g2_fill_1 FILLER_48_286 ();
 sg13g2_fill_1 FILLER_48_299 ();
 sg13g2_decap_4 FILLER_48_330 ();
 sg13g2_decap_4 FILLER_48_340 ();
 sg13g2_fill_2 FILLER_48_344 ();
 sg13g2_decap_8 FILLER_48_349 ();
 sg13g2_decap_4 FILLER_48_356 ();
 sg13g2_fill_2 FILLER_48_360 ();
 sg13g2_fill_2 FILLER_48_419 ();
 sg13g2_decap_4 FILLER_48_426 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_8 FILLER_49_7 ();
 sg13g2_decap_8 FILLER_49_14 ();
 sg13g2_decap_8 FILLER_49_21 ();
 sg13g2_decap_8 FILLER_49_28 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_decap_4 FILLER_49_42 ();
 sg13g2_fill_1 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_98 ();
 sg13g2_decap_4 FILLER_49_105 ();
 sg13g2_fill_2 FILLER_49_109 ();
 sg13g2_fill_2 FILLER_49_123 ();
 sg13g2_fill_1 FILLER_49_156 ();
 sg13g2_fill_2 FILLER_49_183 ();
 sg13g2_decap_8 FILLER_49_195 ();
 sg13g2_decap_4 FILLER_49_213 ();
 sg13g2_fill_1 FILLER_49_217 ();
 sg13g2_fill_1 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_259 ();
 sg13g2_fill_1 FILLER_49_266 ();
 sg13g2_decap_8 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_307 ();
 sg13g2_fill_1 FILLER_49_312 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_fill_2 FILLER_49_347 ();
 sg13g2_fill_2 FILLER_49_375 ();
 sg13g2_fill_1 FILLER_49_377 ();
 sg13g2_fill_1 FILLER_49_410 ();
 sg13g2_fill_2 FILLER_49_420 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_4 FILLER_50_61 ();
 sg13g2_fill_1 FILLER_50_70 ();
 sg13g2_fill_2 FILLER_50_75 ();
 sg13g2_fill_2 FILLER_50_85 ();
 sg13g2_fill_1 FILLER_50_87 ();
 sg13g2_decap_8 FILLER_50_123 ();
 sg13g2_fill_2 FILLER_50_138 ();
 sg13g2_fill_2 FILLER_50_148 ();
 sg13g2_fill_1 FILLER_50_170 ();
 sg13g2_fill_1 FILLER_50_211 ();
 sg13g2_fill_1 FILLER_50_217 ();
 sg13g2_fill_1 FILLER_50_244 ();
 sg13g2_fill_1 FILLER_50_271 ();
 sg13g2_decap_8 FILLER_50_302 ();
 sg13g2_decap_4 FILLER_50_309 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_fill_1 FILLER_50_322 ();
 sg13g2_fill_1 FILLER_50_342 ();
 sg13g2_fill_1 FILLER_50_374 ();
 sg13g2_fill_2 FILLER_50_406 ();
 sg13g2_fill_1 FILLER_50_413 ();
 sg13g2_fill_1 FILLER_50_424 ();
 sg13g2_decap_8 FILLER_51_0 ();
 sg13g2_decap_8 FILLER_51_7 ();
 sg13g2_decap_8 FILLER_51_14 ();
 sg13g2_decap_8 FILLER_51_21 ();
 sg13g2_decap_8 FILLER_51_28 ();
 sg13g2_decap_8 FILLER_51_35 ();
 sg13g2_decap_8 FILLER_51_42 ();
 sg13g2_decap_4 FILLER_51_49 ();
 sg13g2_fill_1 FILLER_51_53 ();
 sg13g2_decap_8 FILLER_51_77 ();
 sg13g2_decap_8 FILLER_51_84 ();
 sg13g2_fill_2 FILLER_51_91 ();
 sg13g2_fill_1 FILLER_51_93 ();
 sg13g2_decap_8 FILLER_51_107 ();
 sg13g2_decap_8 FILLER_51_114 ();
 sg13g2_decap_8 FILLER_51_129 ();
 sg13g2_fill_2 FILLER_51_136 ();
 sg13g2_fill_1 FILLER_51_151 ();
 sg13g2_fill_2 FILLER_51_159 ();
 sg13g2_fill_1 FILLER_51_161 ();
 sg13g2_decap_8 FILLER_51_166 ();
 sg13g2_decap_8 FILLER_51_173 ();
 sg13g2_fill_1 FILLER_51_180 ();
 sg13g2_fill_1 FILLER_51_185 ();
 sg13g2_fill_2 FILLER_51_191 ();
 sg13g2_fill_1 FILLER_51_193 ();
 sg13g2_decap_4 FILLER_51_198 ();
 sg13g2_fill_1 FILLER_51_202 ();
 sg13g2_decap_4 FILLER_51_213 ();
 sg13g2_fill_1 FILLER_51_227 ();
 sg13g2_fill_1 FILLER_51_232 ();
 sg13g2_fill_2 FILLER_51_250 ();
 sg13g2_decap_8 FILLER_51_258 ();
 sg13g2_decap_8 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_272 ();
 sg13g2_fill_1 FILLER_51_292 ();
 sg13g2_decap_8 FILLER_51_296 ();
 sg13g2_decap_8 FILLER_51_303 ();
 sg13g2_decap_8 FILLER_51_310 ();
 sg13g2_fill_1 FILLER_51_317 ();
 sg13g2_fill_2 FILLER_51_322 ();
 sg13g2_fill_1 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_337 ();
 sg13g2_decap_8 FILLER_51_344 ();
 sg13g2_fill_2 FILLER_51_355 ();
 sg13g2_fill_2 FILLER_51_361 ();
 sg13g2_fill_1 FILLER_51_363 ();
 sg13g2_fill_1 FILLER_51_367 ();
 sg13g2_decap_4 FILLER_51_373 ();
 sg13g2_fill_1 FILLER_51_377 ();
 sg13g2_decap_4 FILLER_51_397 ();
 sg13g2_fill_2 FILLER_51_401 ();
 sg13g2_fill_2 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_51_410 ();
 sg13g2_decap_8 FILLER_51_421 ();
 sg13g2_fill_2 FILLER_51_428 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_fill_1 FILLER_52_49 ();
 sg13g2_fill_1 FILLER_52_115 ();
 sg13g2_fill_2 FILLER_52_127 ();
 sg13g2_fill_1 FILLER_52_129 ();
 sg13g2_decap_4 FILLER_52_138 ();
 sg13g2_fill_2 FILLER_52_187 ();
 sg13g2_fill_2 FILLER_52_193 ();
 sg13g2_fill_1 FILLER_52_195 ();
 sg13g2_fill_2 FILLER_52_202 ();
 sg13g2_decap_4 FILLER_52_207 ();
 sg13g2_decap_8 FILLER_52_216 ();
 sg13g2_decap_4 FILLER_52_223 ();
 sg13g2_decap_4 FILLER_52_231 ();
 sg13g2_decap_4 FILLER_52_239 ();
 sg13g2_decap_4 FILLER_52_252 ();
 sg13g2_fill_2 FILLER_52_256 ();
 sg13g2_fill_1 FILLER_52_262 ();
 sg13g2_decap_8 FILLER_52_268 ();
 sg13g2_decap_8 FILLER_52_275 ();
 sg13g2_fill_2 FILLER_52_282 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_fill_1 FILLER_52_374 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_4 FILLER_52_399 ();
 sg13g2_fill_1 FILLER_52_403 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_fill_1 FILLER_52_415 ();
 sg13g2_decap_4 FILLER_52_425 ();
 sg13g2_fill_1 FILLER_52_429 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_4 FILLER_53_49 ();
 sg13g2_fill_1 FILLER_53_79 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_fill_2 FILLER_53_91 ();
 sg13g2_fill_1 FILLER_53_115 ();
 sg13g2_fill_2 FILLER_53_146 ();
 sg13g2_fill_1 FILLER_53_148 ();
 sg13g2_fill_1 FILLER_53_154 ();
 sg13g2_fill_1 FILLER_53_164 ();
 sg13g2_decap_8 FILLER_53_170 ();
 sg13g2_decap_4 FILLER_53_177 ();
 sg13g2_fill_1 FILLER_53_181 ();
 sg13g2_decap_4 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_221 ();
 sg13g2_fill_1 FILLER_53_226 ();
 sg13g2_decap_8 FILLER_53_232 ();
 sg13g2_decap_4 FILLER_53_239 ();
 sg13g2_fill_1 FILLER_53_243 ();
 sg13g2_fill_2 FILLER_53_270 ();
 sg13g2_decap_8 FILLER_53_284 ();
 sg13g2_fill_1 FILLER_53_311 ();
 sg13g2_decap_8 FILLER_53_316 ();
 sg13g2_fill_2 FILLER_53_323 ();
 sg13g2_fill_1 FILLER_53_342 ();
 sg13g2_fill_2 FILLER_53_374 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_decap_4 FILLER_53_390 ();
 sg13g2_fill_2 FILLER_53_394 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_fill_1 FILLER_53_406 ();
 sg13g2_decap_4 FILLER_53_412 ();
 sg13g2_decap_4 FILLER_53_425 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_8 FILLER_54_14 ();
 sg13g2_decap_8 FILLER_54_21 ();
 sg13g2_decap_8 FILLER_54_28 ();
 sg13g2_decap_8 FILLER_54_35 ();
 sg13g2_decap_8 FILLER_54_42 ();
 sg13g2_decap_8 FILLER_54_49 ();
 sg13g2_fill_1 FILLER_54_56 ();
 sg13g2_decap_4 FILLER_54_65 ();
 sg13g2_decap_8 FILLER_54_79 ();
 sg13g2_decap_8 FILLER_54_86 ();
 sg13g2_decap_4 FILLER_54_93 ();
 sg13g2_fill_1 FILLER_54_110 ();
 sg13g2_decap_8 FILLER_54_120 ();
 sg13g2_fill_1 FILLER_54_127 ();
 sg13g2_decap_4 FILLER_54_132 ();
 sg13g2_fill_2 FILLER_54_157 ();
 sg13g2_fill_1 FILLER_54_159 ();
 sg13g2_decap_4 FILLER_54_167 ();
 sg13g2_decap_8 FILLER_54_181 ();
 sg13g2_fill_1 FILLER_54_188 ();
 sg13g2_fill_2 FILLER_54_193 ();
 sg13g2_fill_2 FILLER_54_204 ();
 sg13g2_fill_1 FILLER_54_206 ();
 sg13g2_fill_1 FILLER_54_212 ();
 sg13g2_fill_1 FILLER_54_217 ();
 sg13g2_fill_2 FILLER_54_222 ();
 sg13g2_fill_1 FILLER_54_232 ();
 sg13g2_fill_2 FILLER_54_237 ();
 sg13g2_fill_1 FILLER_54_244 ();
 sg13g2_fill_2 FILLER_54_331 ();
 sg13g2_fill_1 FILLER_54_333 ();
 sg13g2_fill_2 FILLER_54_392 ();
 sg13g2_fill_1 FILLER_54_394 ();
 sg13g2_decap_8 FILLER_54_408 ();
 sg13g2_decap_8 FILLER_54_415 ();
 sg13g2_decap_8 FILLER_54_422 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_4 FILLER_55_63 ();
 sg13g2_fill_2 FILLER_55_67 ();
 sg13g2_decap_4 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_83 ();
 sg13g2_fill_1 FILLER_55_119 ();
 sg13g2_fill_2 FILLER_55_154 ();
 sg13g2_fill_1 FILLER_55_156 ();
 sg13g2_decap_4 FILLER_55_188 ();
 sg13g2_fill_2 FILLER_55_192 ();
 sg13g2_fill_2 FILLER_55_199 ();
 sg13g2_fill_1 FILLER_55_259 ();
 sg13g2_decap_4 FILLER_55_289 ();
 sg13g2_fill_1 FILLER_55_304 ();
 sg13g2_fill_1 FILLER_55_310 ();
 sg13g2_fill_2 FILLER_55_319 ();
 sg13g2_fill_1 FILLER_55_338 ();
 sg13g2_fill_1 FILLER_55_344 ();
 sg13g2_fill_1 FILLER_55_353 ();
 sg13g2_decap_4 FILLER_55_358 ();
 sg13g2_fill_2 FILLER_55_386 ();
 sg13g2_fill_1 FILLER_55_388 ();
 sg13g2_fill_1 FILLER_55_402 ();
 sg13g2_decap_8 FILLER_55_408 ();
 sg13g2_decap_8 FILLER_55_415 ();
 sg13g2_decap_8 FILLER_55_422 ();
 sg13g2_fill_1 FILLER_55_429 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_8 FILLER_56_35 ();
 sg13g2_decap_8 FILLER_56_42 ();
 sg13g2_decap_8 FILLER_56_49 ();
 sg13g2_fill_2 FILLER_56_56 ();
 sg13g2_fill_1 FILLER_56_58 ();
 sg13g2_fill_2 FILLER_56_93 ();
 sg13g2_decap_8 FILLER_56_104 ();
 sg13g2_decap_8 FILLER_56_116 ();
 sg13g2_fill_2 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_129 ();
 sg13g2_decap_8 FILLER_56_136 ();
 sg13g2_decap_8 FILLER_56_143 ();
 sg13g2_decap_8 FILLER_56_150 ();
 sg13g2_decap_8 FILLER_56_157 ();
 sg13g2_decap_4 FILLER_56_182 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_2 FILLER_56_192 ();
 sg13g2_fill_1 FILLER_56_194 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_fill_2 FILLER_56_207 ();
 sg13g2_fill_2 FILLER_56_247 ();
 sg13g2_decap_8 FILLER_56_263 ();
 sg13g2_decap_4 FILLER_56_299 ();
 sg13g2_fill_2 FILLER_56_303 ();
 sg13g2_decap_8 FILLER_56_315 ();
 sg13g2_decap_8 FILLER_56_322 ();
 sg13g2_decap_8 FILLER_56_329 ();
 sg13g2_decap_8 FILLER_56_336 ();
 sg13g2_decap_8 FILLER_56_343 ();
 sg13g2_decap_8 FILLER_56_350 ();
 sg13g2_decap_8 FILLER_56_357 ();
 sg13g2_decap_8 FILLER_56_364 ();
 sg13g2_decap_8 FILLER_56_371 ();
 sg13g2_fill_2 FILLER_56_378 ();
 sg13g2_fill_1 FILLER_56_380 ();
 sg13g2_fill_2 FILLER_56_391 ();
 sg13g2_fill_1 FILLER_56_393 ();
 sg13g2_fill_2 FILLER_56_407 ();
 sg13g2_decap_4 FILLER_56_424 ();
 sg13g2_fill_2 FILLER_56_428 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_103 ();
 sg13g2_fill_2 FILLER_57_110 ();
 sg13g2_fill_1 FILLER_57_112 ();
 sg13g2_decap_4 FILLER_57_125 ();
 sg13g2_decap_8 FILLER_57_142 ();
 sg13g2_decap_8 FILLER_57_149 ();
 sg13g2_fill_1 FILLER_57_156 ();
 sg13g2_fill_2 FILLER_57_165 ();
 sg13g2_decap_4 FILLER_57_172 ();
 sg13g2_fill_1 FILLER_57_176 ();
 sg13g2_decap_4 FILLER_57_207 ();
 sg13g2_decap_4 FILLER_57_216 ();
 sg13g2_fill_1 FILLER_57_220 ();
 sg13g2_decap_8 FILLER_57_225 ();
 sg13g2_fill_1 FILLER_57_232 ();
 sg13g2_fill_2 FILLER_57_244 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_fill_1 FILLER_57_279 ();
 sg13g2_decap_8 FILLER_57_284 ();
 sg13g2_decap_4 FILLER_57_291 ();
 sg13g2_fill_2 FILLER_57_295 ();
 sg13g2_decap_4 FILLER_57_300 ();
 sg13g2_fill_1 FILLER_57_304 ();
 sg13g2_fill_2 FILLER_57_344 ();
 sg13g2_fill_1 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_352 ();
 sg13g2_fill_2 FILLER_57_358 ();
 sg13g2_fill_1 FILLER_57_360 ();
 sg13g2_decap_8 FILLER_57_381 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_4 FILLER_57_395 ();
 sg13g2_fill_1 FILLER_57_421 ();
 sg13g2_decap_4 FILLER_57_426 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_fill_2 FILLER_58_70 ();
 sg13g2_fill_1 FILLER_58_72 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_4 FILLER_58_105 ();
 sg13g2_fill_1 FILLER_58_117 ();
 sg13g2_decap_4 FILLER_58_126 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_decap_8 FILLER_58_136 ();
 sg13g2_decap_8 FILLER_58_143 ();
 sg13g2_decap_8 FILLER_58_150 ();
 sg13g2_decap_8 FILLER_58_157 ();
 sg13g2_decap_8 FILLER_58_164 ();
 sg13g2_decap_4 FILLER_58_171 ();
 sg13g2_fill_2 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_201 ();
 sg13g2_decap_4 FILLER_58_212 ();
 sg13g2_decap_8 FILLER_58_220 ();
 sg13g2_fill_2 FILLER_58_227 ();
 sg13g2_fill_1 FILLER_58_233 ();
 sg13g2_decap_8 FILLER_58_239 ();
 sg13g2_fill_1 FILLER_58_246 ();
 sg13g2_fill_2 FILLER_58_251 ();
 sg13g2_decap_4 FILLER_58_257 ();
 sg13g2_fill_2 FILLER_58_261 ();
 sg13g2_fill_2 FILLER_58_267 ();
 sg13g2_decap_4 FILLER_58_274 ();
 sg13g2_fill_1 FILLER_58_278 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_fill_2 FILLER_58_294 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_1 FILLER_58_323 ();
 sg13g2_fill_2 FILLER_58_328 ();
 sg13g2_fill_2 FILLER_58_340 ();
 sg13g2_fill_1 FILLER_58_364 ();
 sg13g2_fill_2 FILLER_58_372 ();
 sg13g2_decap_4 FILLER_58_390 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_fill_2 FILLER_58_400 ();
 sg13g2_fill_1 FILLER_58_413 ();
 sg13g2_fill_2 FILLER_58_418 ();
 sg13g2_fill_1 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_decap_8 FILLER_59_7 ();
 sg13g2_decap_8 FILLER_59_14 ();
 sg13g2_decap_8 FILLER_59_21 ();
 sg13g2_decap_8 FILLER_59_28 ();
 sg13g2_decap_8 FILLER_59_35 ();
 sg13g2_decap_8 FILLER_59_42 ();
 sg13g2_decap_8 FILLER_59_49 ();
 sg13g2_decap_8 FILLER_59_56 ();
 sg13g2_decap_8 FILLER_59_63 ();
 sg13g2_decap_8 FILLER_59_70 ();
 sg13g2_decap_8 FILLER_59_77 ();
 sg13g2_fill_2 FILLER_59_84 ();
 sg13g2_fill_1 FILLER_59_86 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_decap_8 FILLER_59_134 ();
 sg13g2_decap_8 FILLER_59_141 ();
 sg13g2_decap_8 FILLER_59_148 ();
 sg13g2_decap_8 FILLER_59_155 ();
 sg13g2_decap_8 FILLER_59_162 ();
 sg13g2_fill_2 FILLER_59_169 ();
 sg13g2_fill_1 FILLER_59_171 ();
 sg13g2_decap_4 FILLER_59_189 ();
 sg13g2_decap_8 FILLER_59_198 ();
 sg13g2_decap_4 FILLER_59_205 ();
 sg13g2_fill_2 FILLER_59_209 ();
 sg13g2_fill_2 FILLER_59_215 ();
 sg13g2_decap_4 FILLER_59_221 ();
 sg13g2_decap_8 FILLER_59_237 ();
 sg13g2_decap_8 FILLER_59_244 ();
 sg13g2_fill_2 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_253 ();
 sg13g2_decap_8 FILLER_59_286 ();
 sg13g2_fill_2 FILLER_59_298 ();
 sg13g2_fill_1 FILLER_59_300 ();
 sg13g2_decap_8 FILLER_59_305 ();
 sg13g2_decap_8 FILLER_59_312 ();
 sg13g2_decap_8 FILLER_59_319 ();
 sg13g2_decap_4 FILLER_59_326 ();
 sg13g2_decap_8 FILLER_59_334 ();
 sg13g2_fill_1 FILLER_59_341 ();
 sg13g2_fill_2 FILLER_59_345 ();
 sg13g2_fill_1 FILLER_59_347 ();
 sg13g2_decap_4 FILLER_59_361 ();
 sg13g2_fill_2 FILLER_59_365 ();
 sg13g2_fill_1 FILLER_59_388 ();
 sg13g2_decap_8 FILLER_59_394 ();
 sg13g2_decap_4 FILLER_59_401 ();
 sg13g2_fill_1 FILLER_59_405 ();
 sg13g2_decap_8 FILLER_59_410 ();
 sg13g2_decap_8 FILLER_59_417 ();
 sg13g2_decap_4 FILLER_59_424 ();
 sg13g2_fill_2 FILLER_59_428 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_8 FILLER_60_14 ();
 sg13g2_decap_8 FILLER_60_21 ();
 sg13g2_decap_8 FILLER_60_28 ();
 sg13g2_decap_8 FILLER_60_35 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_8 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_77 ();
 sg13g2_fill_2 FILLER_60_84 ();
 sg13g2_decap_8 FILLER_60_99 ();
 sg13g2_decap_8 FILLER_60_106 ();
 sg13g2_fill_1 FILLER_60_113 ();
 sg13g2_decap_8 FILLER_60_118 ();
 sg13g2_decap_8 FILLER_60_129 ();
 sg13g2_decap_4 FILLER_60_141 ();
 sg13g2_fill_2 FILLER_60_145 ();
 sg13g2_fill_2 FILLER_60_153 ();
 sg13g2_fill_1 FILLER_60_155 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_decap_8 FILLER_60_187 ();
 sg13g2_decap_8 FILLER_60_194 ();
 sg13g2_fill_2 FILLER_60_201 ();
 sg13g2_fill_2 FILLER_60_215 ();
 sg13g2_fill_1 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_227 ();
 sg13g2_decap_8 FILLER_60_234 ();
 sg13g2_decap_8 FILLER_60_241 ();
 sg13g2_decap_8 FILLER_60_248 ();
 sg13g2_decap_8 FILLER_60_255 ();
 sg13g2_decap_8 FILLER_60_262 ();
 sg13g2_decap_8 FILLER_60_269 ();
 sg13g2_fill_2 FILLER_60_276 ();
 sg13g2_decap_8 FILLER_60_293 ();
 sg13g2_decap_8 FILLER_60_300 ();
 sg13g2_decap_8 FILLER_60_307 ();
 sg13g2_decap_8 FILLER_60_314 ();
 sg13g2_decap_8 FILLER_60_321 ();
 sg13g2_fill_2 FILLER_60_328 ();
 sg13g2_fill_1 FILLER_60_334 ();
 sg13g2_decap_4 FILLER_60_345 ();
 sg13g2_fill_1 FILLER_60_349 ();
 sg13g2_fill_1 FILLER_60_354 ();
 sg13g2_decap_8 FILLER_60_390 ();
 sg13g2_fill_2 FILLER_60_397 ();
 sg13g2_decap_4 FILLER_60_425 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_decap_8 FILLER_61_0 ();
 sg13g2_decap_8 FILLER_61_7 ();
 sg13g2_decap_8 FILLER_61_14 ();
 sg13g2_decap_8 FILLER_61_21 ();
 sg13g2_decap_8 FILLER_61_28 ();
 sg13g2_decap_8 FILLER_61_35 ();
 sg13g2_decap_8 FILLER_61_42 ();
 sg13g2_decap_8 FILLER_61_49 ();
 sg13g2_decap_8 FILLER_61_56 ();
 sg13g2_decap_8 FILLER_61_63 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_109 ();
 sg13g2_fill_1 FILLER_61_128 ();
 sg13g2_fill_1 FILLER_61_135 ();
 sg13g2_fill_1 FILLER_61_150 ();
 sg13g2_fill_2 FILLER_61_169 ();
 sg13g2_fill_1 FILLER_61_171 ();
 sg13g2_fill_1 FILLER_61_196 ();
 sg13g2_decap_8 FILLER_61_201 ();
 sg13g2_decap_8 FILLER_61_208 ();
 sg13g2_decap_8 FILLER_61_215 ();
 sg13g2_decap_4 FILLER_61_222 ();
 sg13g2_fill_2 FILLER_61_226 ();
 sg13g2_decap_4 FILLER_61_232 ();
 sg13g2_fill_2 FILLER_61_244 ();
 sg13g2_decap_8 FILLER_61_250 ();
 sg13g2_decap_8 FILLER_61_257 ();
 sg13g2_decap_8 FILLER_61_264 ();
 sg13g2_fill_2 FILLER_61_271 ();
 sg13g2_fill_1 FILLER_61_289 ();
 sg13g2_fill_1 FILLER_61_321 ();
 sg13g2_fill_2 FILLER_61_334 ();
 sg13g2_decap_4 FILLER_61_350 ();
 sg13g2_fill_2 FILLER_61_354 ();
 sg13g2_fill_2 FILLER_61_364 ();
 sg13g2_fill_1 FILLER_61_366 ();
 sg13g2_fill_2 FILLER_61_371 ();
 sg13g2_fill_1 FILLER_61_373 ();
 sg13g2_fill_2 FILLER_61_382 ();
 sg13g2_fill_1 FILLER_61_384 ();
 sg13g2_decap_8 FILLER_61_421 ();
 sg13g2_fill_2 FILLER_61_428 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_decap_8 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_63 ();
 sg13g2_decap_8 FILLER_62_70 ();
 sg13g2_decap_8 FILLER_62_77 ();
 sg13g2_decap_8 FILLER_62_84 ();
 sg13g2_fill_2 FILLER_62_91 ();
 sg13g2_fill_1 FILLER_62_93 ();
 sg13g2_decap_4 FILLER_62_98 ();
 sg13g2_fill_2 FILLER_62_102 ();
 sg13g2_fill_2 FILLER_62_109 ();
 sg13g2_fill_1 FILLER_62_111 ();
 sg13g2_fill_1 FILLER_62_120 ();
 sg13g2_fill_2 FILLER_62_133 ();
 sg13g2_fill_1 FILLER_62_135 ();
 sg13g2_fill_1 FILLER_62_144 ();
 sg13g2_fill_1 FILLER_62_155 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_201 ();
 sg13g2_fill_2 FILLER_62_207 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_4 FILLER_62_224 ();
 sg13g2_fill_2 FILLER_62_228 ();
 sg13g2_fill_1 FILLER_62_246 ();
 sg13g2_fill_1 FILLER_62_252 ();
 sg13g2_fill_2 FILLER_62_262 ();
 sg13g2_fill_2 FILLER_62_272 ();
 sg13g2_fill_1 FILLER_62_307 ();
 sg13g2_fill_1 FILLER_62_336 ();
 sg13g2_decap_4 FILLER_62_349 ();
 sg13g2_fill_1 FILLER_62_353 ();
 sg13g2_decap_8 FILLER_62_362 ();
 sg13g2_fill_2 FILLER_62_369 ();
 sg13g2_decap_4 FILLER_62_380 ();
 sg13g2_decap_4 FILLER_62_400 ();
 sg13g2_decap_4 FILLER_62_408 ();
 sg13g2_fill_2 FILLER_62_412 ();
 sg13g2_fill_2 FILLER_62_427 ();
 sg13g2_fill_1 FILLER_62_429 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_4 FILLER_63_77 ();
 sg13g2_fill_1 FILLER_63_81 ();
 sg13g2_decap_8 FILLER_63_86 ();
 sg13g2_decap_8 FILLER_63_93 ();
 sg13g2_decap_4 FILLER_63_100 ();
 sg13g2_fill_2 FILLER_63_104 ();
 sg13g2_decap_8 FILLER_63_114 ();
 sg13g2_fill_1 FILLER_63_127 ();
 sg13g2_fill_2 FILLER_63_133 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_141 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_fill_1 FILLER_63_159 ();
 sg13g2_fill_2 FILLER_63_164 ();
 sg13g2_decap_4 FILLER_63_170 ();
 sg13g2_fill_2 FILLER_63_179 ();
 sg13g2_fill_1 FILLER_63_181 ();
 sg13g2_fill_2 FILLER_63_222 ();
 sg13g2_fill_1 FILLER_63_232 ();
 sg13g2_fill_1 FILLER_63_244 ();
 sg13g2_decap_4 FILLER_63_250 ();
 sg13g2_fill_2 FILLER_63_254 ();
 sg13g2_decap_4 FILLER_63_260 ();
 sg13g2_fill_2 FILLER_63_268 ();
 sg13g2_fill_1 FILLER_63_270 ();
 sg13g2_decap_8 FILLER_63_275 ();
 sg13g2_decap_8 FILLER_63_282 ();
 sg13g2_decap_4 FILLER_63_289 ();
 sg13g2_fill_2 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_300 ();
 sg13g2_decap_4 FILLER_63_305 ();
 sg13g2_fill_1 FILLER_63_309 ();
 sg13g2_decap_8 FILLER_63_314 ();
 sg13g2_fill_2 FILLER_63_338 ();
 sg13g2_fill_1 FILLER_63_340 ();
 sg13g2_decap_8 FILLER_63_345 ();
 sg13g2_decap_8 FILLER_63_352 ();
 sg13g2_decap_8 FILLER_63_359 ();
 sg13g2_fill_2 FILLER_63_366 ();
 sg13g2_fill_1 FILLER_63_368 ();
 sg13g2_decap_8 FILLER_63_382 ();
 sg13g2_decap_8 FILLER_63_389 ();
 sg13g2_decap_8 FILLER_63_396 ();
 sg13g2_decap_4 FILLER_63_403 ();
 sg13g2_fill_1 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_8 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_21 ();
 sg13g2_decap_8 FILLER_64_28 ();
 sg13g2_decap_8 FILLER_64_35 ();
 sg13g2_decap_8 FILLER_64_42 ();
 sg13g2_decap_8 FILLER_64_49 ();
 sg13g2_decap_8 FILLER_64_56 ();
 sg13g2_decap_8 FILLER_64_63 ();
 sg13g2_decap_4 FILLER_64_70 ();
 sg13g2_fill_1 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_105 ();
 sg13g2_decap_4 FILLER_64_111 ();
 sg13g2_fill_2 FILLER_64_115 ();
 sg13g2_fill_1 FILLER_64_145 ();
 sg13g2_fill_1 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_166 ();
 sg13g2_decap_8 FILLER_64_173 ();
 sg13g2_fill_1 FILLER_64_199 ();
 sg13g2_decap_4 FILLER_64_226 ();
 sg13g2_fill_1 FILLER_64_230 ();
 sg13g2_decap_8 FILLER_64_235 ();
 sg13g2_decap_4 FILLER_64_242 ();
 sg13g2_decap_8 FILLER_64_251 ();
 sg13g2_fill_1 FILLER_64_258 ();
 sg13g2_fill_1 FILLER_64_267 ();
 sg13g2_decap_8 FILLER_64_272 ();
 sg13g2_fill_2 FILLER_64_279 ();
 sg13g2_fill_2 FILLER_64_290 ();
 sg13g2_fill_2 FILLER_64_296 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_314 ();
 sg13g2_fill_2 FILLER_64_321 ();
 sg13g2_fill_1 FILLER_64_323 ();
 sg13g2_decap_4 FILLER_64_333 ();
 sg13g2_decap_8 FILLER_64_342 ();
 sg13g2_decap_8 FILLER_64_349 ();
 sg13g2_decap_8 FILLER_64_356 ();
 sg13g2_decap_4 FILLER_64_363 ();
 sg13g2_fill_1 FILLER_64_367 ();
 sg13g2_decap_4 FILLER_64_373 ();
 sg13g2_decap_8 FILLER_64_381 ();
 sg13g2_decap_8 FILLER_64_388 ();
 sg13g2_fill_2 FILLER_64_395 ();
 sg13g2_fill_1 FILLER_64_397 ();
 sg13g2_decap_4 FILLER_64_424 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_fill_2 FILLER_65_77 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_fill_1 FILLER_65_115 ();
 sg13g2_decap_8 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_131 ();
 sg13g2_fill_1 FILLER_65_138 ();
 sg13g2_fill_2 FILLER_65_152 ();
 sg13g2_decap_8 FILLER_65_164 ();
 sg13g2_decap_8 FILLER_65_171 ();
 sg13g2_decap_8 FILLER_65_178 ();
 sg13g2_fill_2 FILLER_65_185 ();
 sg13g2_fill_1 FILLER_65_187 ();
 sg13g2_fill_2 FILLER_65_220 ();
 sg13g2_decap_4 FILLER_65_252 ();
 sg13g2_fill_1 FILLER_65_256 ();
 sg13g2_fill_1 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_314 ();
 sg13g2_decap_8 FILLER_65_321 ();
 sg13g2_decap_8 FILLER_65_328 ();
 sg13g2_decap_8 FILLER_65_335 ();
 sg13g2_decap_8 FILLER_65_342 ();
 sg13g2_decap_8 FILLER_65_349 ();
 sg13g2_decap_8 FILLER_65_356 ();
 sg13g2_decap_4 FILLER_65_363 ();
 sg13g2_decap_8 FILLER_65_384 ();
 sg13g2_decap_8 FILLER_65_417 ();
 sg13g2_decap_4 FILLER_65_424 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_14 ();
 sg13g2_decap_8 FILLER_66_21 ();
 sg13g2_decap_8 FILLER_66_28 ();
 sg13g2_decap_8 FILLER_66_35 ();
 sg13g2_decap_8 FILLER_66_42 ();
 sg13g2_decap_8 FILLER_66_49 ();
 sg13g2_decap_8 FILLER_66_56 ();
 sg13g2_decap_8 FILLER_66_63 ();
 sg13g2_decap_8 FILLER_66_70 ();
 sg13g2_decap_8 FILLER_66_77 ();
 sg13g2_fill_2 FILLER_66_84 ();
 sg13g2_fill_1 FILLER_66_86 ();
 sg13g2_decap_4 FILLER_66_91 ();
 sg13g2_fill_2 FILLER_66_95 ();
 sg13g2_decap_8 FILLER_66_101 ();
 sg13g2_fill_2 FILLER_66_108 ();
 sg13g2_decap_8 FILLER_66_118 ();
 sg13g2_decap_8 FILLER_66_125 ();
 sg13g2_decap_8 FILLER_66_132 ();
 sg13g2_decap_8 FILLER_66_143 ();
 sg13g2_decap_8 FILLER_66_150 ();
 sg13g2_decap_8 FILLER_66_157 ();
 sg13g2_decap_8 FILLER_66_164 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_fill_2 FILLER_66_190 ();
 sg13g2_decap_8 FILLER_66_196 ();
 sg13g2_decap_8 FILLER_66_203 ();
 sg13g2_decap_8 FILLER_66_210 ();
 sg13g2_decap_8 FILLER_66_227 ();
 sg13g2_decap_8 FILLER_66_234 ();
 sg13g2_decap_8 FILLER_66_241 ();
 sg13g2_decap_8 FILLER_66_248 ();
 sg13g2_decap_8 FILLER_66_255 ();
 sg13g2_decap_8 FILLER_66_262 ();
 sg13g2_decap_8 FILLER_66_269 ();
 sg13g2_decap_8 FILLER_66_276 ();
 sg13g2_decap_8 FILLER_66_296 ();
 sg13g2_decap_4 FILLER_66_303 ();
 sg13g2_fill_1 FILLER_66_307 ();
 sg13g2_decap_8 FILLER_66_325 ();
 sg13g2_decap_8 FILLER_66_332 ();
 sg13g2_fill_2 FILLER_66_339 ();
 sg13g2_fill_1 FILLER_66_341 ();
 sg13g2_decap_8 FILLER_66_350 ();
 sg13g2_decap_8 FILLER_66_357 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_decap_8 FILLER_66_370 ();
 sg13g2_decap_8 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_418 ();
 sg13g2_decap_4 FILLER_66_425 ();
 sg13g2_fill_1 FILLER_66_429 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_8 FILLER_67_28 ();
 sg13g2_decap_8 FILLER_67_35 ();
 sg13g2_decap_8 FILLER_67_42 ();
 sg13g2_decap_8 FILLER_67_49 ();
 sg13g2_decap_8 FILLER_67_56 ();
 sg13g2_decap_8 FILLER_67_63 ();
 sg13g2_fill_1 FILLER_67_70 ();
 sg13g2_fill_2 FILLER_67_97 ();
 sg13g2_fill_2 FILLER_67_107 ();
 sg13g2_fill_1 FILLER_67_109 ();
 sg13g2_fill_2 FILLER_67_114 ();
 sg13g2_fill_2 FILLER_67_131 ();
 sg13g2_fill_1 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_152 ();
 sg13g2_fill_1 FILLER_67_159 ();
 sg13g2_fill_2 FILLER_67_163 ();
 sg13g2_decap_8 FILLER_67_205 ();
 sg13g2_decap_8 FILLER_67_227 ();
 sg13g2_fill_2 FILLER_67_234 ();
 sg13g2_decap_8 FILLER_67_257 ();
 sg13g2_decap_4 FILLER_67_294 ();
 sg13g2_fill_1 FILLER_67_298 ();
 sg13g2_fill_2 FILLER_67_303 ();
 sg13g2_fill_2 FILLER_67_329 ();
 sg13g2_fill_1 FILLER_67_331 ();
 sg13g2_fill_1 FILLER_67_362 ();
 sg13g2_decap_8 FILLER_67_386 ();
 sg13g2_fill_1 FILLER_67_393 ();
 sg13g2_decap_8 FILLER_67_402 ();
 sg13g2_decap_8 FILLER_67_409 ();
 sg13g2_decap_8 FILLER_67_416 ();
 sg13g2_decap_8 FILLER_67_423 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_decap_8 FILLER_68_21 ();
 sg13g2_decap_8 FILLER_68_28 ();
 sg13g2_decap_8 FILLER_68_35 ();
 sg13g2_decap_8 FILLER_68_42 ();
 sg13g2_decap_8 FILLER_68_49 ();
 sg13g2_decap_8 FILLER_68_56 ();
 sg13g2_decap_8 FILLER_68_63 ();
 sg13g2_decap_8 FILLER_68_70 ();
 sg13g2_decap_4 FILLER_68_81 ();
 sg13g2_fill_2 FILLER_68_124 ();
 sg13g2_fill_2 FILLER_68_134 ();
 sg13g2_fill_1 FILLER_68_162 ();
 sg13g2_fill_1 FILLER_68_172 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_2 FILLER_68_210 ();
 sg13g2_fill_2 FILLER_68_354 ();
 sg13g2_fill_1 FILLER_68_356 ();
 sg13g2_decap_4 FILLER_68_360 ();
 sg13g2_fill_2 FILLER_68_364 ();
 sg13g2_fill_1 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_402 ();
 sg13g2_decap_8 FILLER_68_409 ();
 sg13g2_decap_4 FILLER_68_416 ();
 sg13g2_fill_1 FILLER_68_420 ();
 sg13g2_decap_4 FILLER_68_426 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_8 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_63 ();
 sg13g2_decap_8 FILLER_69_70 ();
 sg13g2_decap_8 FILLER_69_77 ();
 sg13g2_decap_8 FILLER_69_84 ();
 sg13g2_fill_1 FILLER_69_91 ();
 sg13g2_decap_8 FILLER_69_101 ();
 sg13g2_decap_8 FILLER_69_108 ();
 sg13g2_fill_2 FILLER_69_115 ();
 sg13g2_fill_1 FILLER_69_131 ();
 sg13g2_decap_4 FILLER_69_161 ();
 sg13g2_fill_1 FILLER_69_170 ();
 sg13g2_decap_4 FILLER_69_175 ();
 sg13g2_fill_2 FILLER_69_188 ();
 sg13g2_decap_8 FILLER_69_194 ();
 sg13g2_decap_8 FILLER_69_201 ();
 sg13g2_decap_8 FILLER_69_208 ();
 sg13g2_fill_2 FILLER_69_215 ();
 sg13g2_decap_4 FILLER_69_232 ();
 sg13g2_fill_1 FILLER_69_236 ();
 sg13g2_fill_1 FILLER_69_249 ();
 sg13g2_decap_8 FILLER_69_254 ();
 sg13g2_fill_1 FILLER_69_265 ();
 sg13g2_fill_1 FILLER_69_270 ();
 sg13g2_fill_1 FILLER_69_274 ();
 sg13g2_decap_8 FILLER_69_279 ();
 sg13g2_fill_2 FILLER_69_290 ();
 sg13g2_decap_8 FILLER_69_296 ();
 sg13g2_decap_8 FILLER_69_303 ();
 sg13g2_fill_2 FILLER_69_310 ();
 sg13g2_fill_2 FILLER_69_354 ();
 sg13g2_fill_1 FILLER_69_356 ();
 sg13g2_decap_4 FILLER_69_362 ();
 sg13g2_fill_1 FILLER_69_366 ();
 sg13g2_fill_1 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_69_382 ();
 sg13g2_decap_8 FILLER_69_389 ();
 sg13g2_fill_1 FILLER_69_396 ();
 sg13g2_decap_4 FILLER_69_402 ();
 sg13g2_fill_1 FILLER_69_406 ();
 sg13g2_decap_8 FILLER_69_411 ();
 sg13g2_decap_8 FILLER_69_418 ();
 sg13g2_decap_4 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_69_429 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_fill_2 FILLER_70_63 ();
 sg13g2_fill_1 FILLER_70_65 ();
 sg13g2_decap_4 FILLER_70_92 ();
 sg13g2_fill_2 FILLER_70_96 ();
 sg13g2_fill_1 FILLER_70_113 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_4 FILLER_70_133 ();
 sg13g2_fill_1 FILLER_70_137 ();
 sg13g2_fill_1 FILLER_70_142 ();
 sg13g2_fill_1 FILLER_70_147 ();
 sg13g2_fill_1 FILLER_70_153 ();
 sg13g2_fill_1 FILLER_70_158 ();
 sg13g2_fill_2 FILLER_70_163 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_191 ();
 sg13g2_fill_2 FILLER_70_207 ();
 sg13g2_decap_8 FILLER_70_213 ();
 sg13g2_decap_8 FILLER_70_225 ();
 sg13g2_decap_8 FILLER_70_232 ();
 sg13g2_decap_8 FILLER_70_239 ();
 sg13g2_decap_8 FILLER_70_246 ();
 sg13g2_fill_2 FILLER_70_253 ();
 sg13g2_decap_8 FILLER_70_258 ();
 sg13g2_decap_8 FILLER_70_265 ();
 sg13g2_decap_4 FILLER_70_272 ();
 sg13g2_fill_2 FILLER_70_276 ();
 sg13g2_decap_4 FILLER_70_283 ();
 sg13g2_decap_4 FILLER_70_292 ();
 sg13g2_decap_4 FILLER_70_300 ();
 sg13g2_fill_1 FILLER_70_304 ();
 sg13g2_decap_8 FILLER_70_321 ();
 sg13g2_fill_2 FILLER_70_328 ();
 sg13g2_fill_1 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_384 ();
 sg13g2_decap_8 FILLER_70_391 ();
 sg13g2_fill_2 FILLER_70_398 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_decap_8 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_42 ();
 sg13g2_decap_8 FILLER_71_49 ();
 sg13g2_decap_8 FILLER_71_56 ();
 sg13g2_decap_8 FILLER_71_63 ();
 sg13g2_fill_2 FILLER_71_70 ();
 sg13g2_fill_1 FILLER_71_72 ();
 sg13g2_decap_4 FILLER_71_77 ();
 sg13g2_fill_2 FILLER_71_81 ();
 sg13g2_decap_4 FILLER_71_113 ();
 sg13g2_decap_8 FILLER_71_125 ();
 sg13g2_fill_2 FILLER_71_132 ();
 sg13g2_decap_4 FILLER_71_138 ();
 sg13g2_fill_2 FILLER_71_142 ();
 sg13g2_decap_8 FILLER_71_162 ();
 sg13g2_decap_8 FILLER_71_169 ();
 sg13g2_decap_8 FILLER_71_176 ();
 sg13g2_decap_8 FILLER_71_183 ();
 sg13g2_decap_4 FILLER_71_190 ();
 sg13g2_fill_2 FILLER_71_224 ();
 sg13g2_decap_8 FILLER_71_235 ();
 sg13g2_decap_4 FILLER_71_242 ();
 sg13g2_fill_2 FILLER_71_246 ();
 sg13g2_decap_8 FILLER_71_252 ();
 sg13g2_decap_8 FILLER_71_259 ();
 sg13g2_decap_4 FILLER_71_266 ();
 sg13g2_fill_1 FILLER_71_270 ();
 sg13g2_decap_8 FILLER_71_275 ();
 sg13g2_decap_4 FILLER_71_282 ();
 sg13g2_fill_2 FILLER_71_299 ();
 sg13g2_fill_2 FILLER_71_314 ();
 sg13g2_decap_8 FILLER_71_320 ();
 sg13g2_decap_8 FILLER_71_327 ();
 sg13g2_fill_2 FILLER_71_334 ();
 sg13g2_fill_1 FILLER_71_340 ();
 sg13g2_fill_2 FILLER_71_349 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_368 ();
 sg13g2_fill_2 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_fill_1 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_4 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_92 ();
 sg13g2_decap_8 FILLER_72_99 ();
 sg13g2_decap_8 FILLER_72_106 ();
 sg13g2_decap_8 FILLER_72_113 ();
 sg13g2_fill_1 FILLER_72_120 ();
 sg13g2_decap_8 FILLER_72_150 ();
 sg13g2_decap_8 FILLER_72_157 ();
 sg13g2_decap_8 FILLER_72_164 ();
 sg13g2_decap_4 FILLER_72_181 ();
 sg13g2_fill_1 FILLER_72_185 ();
 sg13g2_fill_2 FILLER_72_242 ();
 sg13g2_fill_2 FILLER_72_269 ();
 sg13g2_fill_1 FILLER_72_276 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_fill_2 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_367 ();
 sg13g2_decap_8 FILLER_72_374 ();
 sg13g2_decap_4 FILLER_72_381 ();
 sg13g2_fill_2 FILLER_72_389 ();
 sg13g2_fill_1 FILLER_72_391 ();
 sg13g2_fill_1 FILLER_72_398 ();
 sg13g2_fill_1 FILLER_72_403 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_decap_8 FILLER_73_14 ();
 sg13g2_decap_8 FILLER_73_21 ();
 sg13g2_decap_8 FILLER_73_28 ();
 sg13g2_decap_8 FILLER_73_35 ();
 sg13g2_decap_8 FILLER_73_42 ();
 sg13g2_decap_8 FILLER_73_49 ();
 sg13g2_decap_8 FILLER_73_56 ();
 sg13g2_decap_8 FILLER_73_63 ();
 sg13g2_decap_8 FILLER_73_70 ();
 sg13g2_decap_8 FILLER_73_77 ();
 sg13g2_decap_8 FILLER_73_84 ();
 sg13g2_decap_4 FILLER_73_91 ();
 sg13g2_fill_2 FILLER_73_110 ();
 sg13g2_fill_2 FILLER_73_148 ();
 sg13g2_fill_2 FILLER_73_207 ();
 sg13g2_fill_1 FILLER_73_230 ();
 sg13g2_fill_1 FILLER_73_265 ();
 sg13g2_decap_4 FILLER_73_274 ();
 sg13g2_decap_4 FILLER_73_308 ();
 sg13g2_decap_4 FILLER_73_316 ();
 sg13g2_fill_1 FILLER_73_320 ();
 sg13g2_decap_4 FILLER_73_358 ();
 sg13g2_fill_1 FILLER_73_362 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_fill_1 FILLER_73_379 ();
 sg13g2_fill_1 FILLER_73_395 ();
 sg13g2_fill_2 FILLER_73_409 ();
 sg13g2_decap_8 FILLER_73_422 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_8 FILLER_74_49 ();
 sg13g2_decap_8 FILLER_74_56 ();
 sg13g2_decap_8 FILLER_74_63 ();
 sg13g2_decap_8 FILLER_74_70 ();
 sg13g2_decap_8 FILLER_74_77 ();
 sg13g2_decap_4 FILLER_74_84 ();
 sg13g2_fill_1 FILLER_74_88 ();
 sg13g2_decap_4 FILLER_74_156 ();
 sg13g2_fill_2 FILLER_74_160 ();
 sg13g2_fill_2 FILLER_74_171 ();
 sg13g2_decap_8 FILLER_74_185 ();
 sg13g2_decap_4 FILLER_74_192 ();
 sg13g2_decap_8 FILLER_74_199 ();
 sg13g2_decap_8 FILLER_74_206 ();
 sg13g2_decap_8 FILLER_74_213 ();
 sg13g2_fill_2 FILLER_74_220 ();
 sg13g2_decap_4 FILLER_74_242 ();
 sg13g2_fill_2 FILLER_74_250 ();
 sg13g2_decap_4 FILLER_74_256 ();
 sg13g2_decap_4 FILLER_74_264 ();
 sg13g2_fill_2 FILLER_74_280 ();
 sg13g2_fill_1 FILLER_74_282 ();
 sg13g2_fill_1 FILLER_74_291 ();
 sg13g2_decap_4 FILLER_74_296 ();
 sg13g2_decap_8 FILLER_74_319 ();
 sg13g2_decap_4 FILLER_74_326 ();
 sg13g2_fill_1 FILLER_74_330 ();
 sg13g2_fill_2 FILLER_74_343 ();
 sg13g2_fill_1 FILLER_74_345 ();
 sg13g2_fill_1 FILLER_74_359 ();
 sg13g2_decap_4 FILLER_74_373 ();
 sg13g2_fill_2 FILLER_74_377 ();
 sg13g2_fill_1 FILLER_74_407 ();
 sg13g2_fill_1 FILLER_74_413 ();
 sg13g2_decap_8 FILLER_74_422 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_decap_4 FILLER_75_56 ();
 sg13g2_fill_2 FILLER_75_90 ();
 sg13g2_fill_1 FILLER_75_97 ();
 sg13g2_fill_2 FILLER_75_124 ();
 sg13g2_fill_1 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_131 ();
 sg13g2_fill_1 FILLER_75_138 ();
 sg13g2_decap_8 FILLER_75_142 ();
 sg13g2_decap_4 FILLER_75_149 ();
 sg13g2_fill_2 FILLER_75_153 ();
 sg13g2_fill_2 FILLER_75_167 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_4 FILLER_75_189 ();
 sg13g2_fill_1 FILLER_75_193 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_4 FILLER_75_232 ();
 sg13g2_fill_2 FILLER_75_236 ();
 sg13g2_decap_8 FILLER_75_246 ();
 sg13g2_decap_8 FILLER_75_253 ();
 sg13g2_decap_4 FILLER_75_260 ();
 sg13g2_fill_2 FILLER_75_264 ();
 sg13g2_decap_8 FILLER_75_269 ();
 sg13g2_decap_8 FILLER_75_276 ();
 sg13g2_decap_8 FILLER_75_283 ();
 sg13g2_fill_1 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_304 ();
 sg13g2_decap_4 FILLER_75_315 ();
 sg13g2_fill_2 FILLER_75_324 ();
 sg13g2_fill_1 FILLER_75_326 ();
 sg13g2_decap_4 FILLER_75_331 ();
 sg13g2_decap_4 FILLER_75_341 ();
 sg13g2_fill_1 FILLER_75_345 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_fill_1 FILLER_75_378 ();
 sg13g2_fill_1 FILLER_75_385 ();
 sg13g2_fill_2 FILLER_75_390 ();
 sg13g2_decap_8 FILLER_75_418 ();
 sg13g2_decap_4 FILLER_75_425 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_decap_8 FILLER_76_56 ();
 sg13g2_decap_8 FILLER_76_63 ();
 sg13g2_decap_8 FILLER_76_70 ();
 sg13g2_decap_8 FILLER_76_77 ();
 sg13g2_decap_4 FILLER_76_84 ();
 sg13g2_fill_1 FILLER_76_93 ();
 sg13g2_decap_8 FILLER_76_102 ();
 sg13g2_decap_4 FILLER_76_109 ();
 sg13g2_fill_1 FILLER_76_121 ();
 sg13g2_fill_2 FILLER_76_134 ();
 sg13g2_decap_8 FILLER_76_144 ();
 sg13g2_decap_4 FILLER_76_151 ();
 sg13g2_fill_1 FILLER_76_155 ();
 sg13g2_decap_8 FILLER_76_182 ();
 sg13g2_decap_8 FILLER_76_219 ();
 sg13g2_fill_2 FILLER_76_226 ();
 sg13g2_decap_8 FILLER_76_232 ();
 sg13g2_decap_8 FILLER_76_239 ();
 sg13g2_decap_8 FILLER_76_246 ();
 sg13g2_decap_4 FILLER_76_253 ();
 sg13g2_fill_1 FILLER_76_257 ();
 sg13g2_fill_2 FILLER_76_280 ();
 sg13g2_fill_1 FILLER_76_288 ();
 sg13g2_decap_4 FILLER_76_347 ();
 sg13g2_fill_1 FILLER_76_351 ();
 sg13g2_fill_1 FILLER_76_355 ();
 sg13g2_decap_4 FILLER_76_370 ();
 sg13g2_fill_1 FILLER_76_374 ();
 sg13g2_fill_1 FILLER_76_383 ();
 sg13g2_fill_1 FILLER_76_406 ();
 sg13g2_fill_2 FILLER_76_412 ();
 sg13g2_fill_1 FILLER_76_414 ();
 sg13g2_decap_8 FILLER_76_419 ();
 sg13g2_decap_4 FILLER_76_426 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_4 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_137 ();
 sg13g2_decap_8 FILLER_77_144 ();
 sg13g2_decap_8 FILLER_77_151 ();
 sg13g2_decap_4 FILLER_77_158 ();
 sg13g2_fill_2 FILLER_77_166 ();
 sg13g2_fill_1 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_174 ();
 sg13g2_decap_4 FILLER_77_181 ();
 sg13g2_fill_1 FILLER_77_204 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_4 FILLER_77_217 ();
 sg13g2_fill_2 FILLER_77_221 ();
 sg13g2_fill_2 FILLER_77_233 ();
 sg13g2_fill_1 FILLER_77_235 ();
 sg13g2_decap_4 FILLER_77_241 ();
 sg13g2_decap_8 FILLER_77_290 ();
 sg13g2_decap_4 FILLER_77_297 ();
 sg13g2_decap_4 FILLER_77_308 ();
 sg13g2_fill_1 FILLER_77_312 ();
 sg13g2_decap_4 FILLER_77_317 ();
 sg13g2_fill_1 FILLER_77_340 ();
 sg13g2_fill_2 FILLER_77_352 ();
 sg13g2_fill_1 FILLER_77_359 ();
 sg13g2_fill_1 FILLER_77_364 ();
 sg13g2_fill_1 FILLER_77_375 ();
 sg13g2_decap_4 FILLER_77_386 ();
 sg13g2_decap_8 FILLER_77_416 ();
 sg13g2_decap_8 FILLER_77_423 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_decap_8 FILLER_78_56 ();
 sg13g2_decap_8 FILLER_78_63 ();
 sg13g2_decap_8 FILLER_78_70 ();
 sg13g2_decap_8 FILLER_78_77 ();
 sg13g2_fill_1 FILLER_78_84 ();
 sg13g2_decap_4 FILLER_78_109 ();
 sg13g2_fill_2 FILLER_78_121 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_decap_4 FILLER_78_160 ();
 sg13g2_fill_1 FILLER_78_164 ();
 sg13g2_fill_2 FILLER_78_180 ();
 sg13g2_fill_1 FILLER_78_182 ();
 sg13g2_fill_2 FILLER_78_214 ();
 sg13g2_fill_2 FILLER_78_271 ();
 sg13g2_decap_4 FILLER_78_278 ();
 sg13g2_decap_4 FILLER_78_308 ();
 sg13g2_decap_8 FILLER_78_325 ();
 sg13g2_decap_8 FILLER_78_337 ();
 sg13g2_decap_8 FILLER_78_344 ();
 sg13g2_decap_8 FILLER_78_351 ();
 sg13g2_fill_2 FILLER_78_358 ();
 sg13g2_decap_8 FILLER_78_403 ();
 sg13g2_decap_8 FILLER_78_410 ();
 sg13g2_decap_8 FILLER_78_417 ();
 sg13g2_decap_4 FILLER_78_424 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_8 FILLER_79_63 ();
 sg13g2_fill_2 FILLER_79_70 ();
 sg13g2_decap_8 FILLER_79_102 ();
 sg13g2_decap_8 FILLER_79_109 ();
 sg13g2_fill_2 FILLER_79_116 ();
 sg13g2_fill_1 FILLER_79_126 ();
 sg13g2_decap_8 FILLER_79_184 ();
 sg13g2_decap_4 FILLER_79_191 ();
 sg13g2_decap_4 FILLER_79_327 ();
 sg13g2_fill_2 FILLER_79_331 ();
 sg13g2_decap_8 FILLER_79_338 ();
 sg13g2_decap_8 FILLER_79_345 ();
 sg13g2_decap_8 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_359 ();
 sg13g2_decap_8 FILLER_79_366 ();
 sg13g2_decap_4 FILLER_79_373 ();
 sg13g2_fill_2 FILLER_79_381 ();
 sg13g2_fill_1 FILLER_79_383 ();
 sg13g2_decap_8 FILLER_79_388 ();
 sg13g2_decap_8 FILLER_79_395 ();
 sg13g2_decap_8 FILLER_79_402 ();
 sg13g2_decap_8 FILLER_79_409 ();
 sg13g2_decap_8 FILLER_79_416 ();
 sg13g2_decap_8 FILLER_79_423 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_fill_2 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_99 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_1 FILLER_80_118 ();
 sg13g2_fill_1 FILLER_80_127 ();
 sg13g2_fill_1 FILLER_80_136 ();
 sg13g2_fill_1 FILLER_80_141 ();
 sg13g2_fill_1 FILLER_80_146 ();
 sg13g2_fill_1 FILLER_80_151 ();
 sg13g2_fill_1 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_185 ();
 sg13g2_fill_2 FILLER_80_206 ();
 sg13g2_fill_2 FILLER_80_220 ();
 sg13g2_fill_1 FILLER_80_226 ();
 sg13g2_decap_4 FILLER_80_248 ();
 sg13g2_fill_1 FILLER_80_256 ();
 sg13g2_fill_2 FILLER_80_269 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_fill_1 FILLER_80_281 ();
 sg13g2_decap_4 FILLER_80_286 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_fill_1 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_313 ();
 sg13g2_decap_4 FILLER_80_337 ();
 sg13g2_fill_1 FILLER_80_341 ();
 sg13g2_fill_2 FILLER_80_363 ();
 sg13g2_decap_4 FILLER_80_378 ();
 sg13g2_fill_1 FILLER_80_386 ();
 sg13g2_decap_8 FILLER_80_391 ();
 sg13g2_decap_8 FILLER_80_398 ();
 sg13g2_decap_8 FILLER_80_405 ();
 sg13g2_decap_8 FILLER_80_412 ();
 sg13g2_decap_8 FILLER_80_419 ();
 sg13g2_decap_4 FILLER_80_426 ();
endmodule
