module tt_um_a1k0n_nyancat (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire clknet_0_clk;
 wire net154;
 wire audio_pwm;
 wire \audio_pwm_accum[0] ;
 wire \audio_pwm_accum[1] ;
 wire \audio_pwm_accum[2] ;
 wire \audio_pwm_accum[3] ;
 wire \audio_pwm_accum[4] ;
 wire \audio_pwm_accum[5] ;
 wire \audio_pwm_accum[6] ;
 wire \audio_pwm_accum[7] ;
 wire \audio_pwm_accum[8] ;
 wire \audio_pwm_accum[9] ;
 wire \audio_pwm_accum_next[0] ;
 wire \audio_pwm_accum_next[1] ;
 wire \audio_pwm_accum_next[2] ;
 wire \audio_pwm_accum_next[3] ;
 wire \audio_pwm_accum_next[4] ;
 wire \audio_pwm_accum_next[5] ;
 wire \audio_pwm_accum_next[6] ;
 wire \audio_pwm_accum_next[7] ;
 wire \audio_pwm_accum_next[8] ;
 wire \audio_pwm_accum_next[9] ;
 wire \audio_sample_lpf[0] ;
 wire \audio_sample_lpf[1] ;
 wire \audio_sample_lpf[2] ;
 wire \audio_sample_lpf[3] ;
 wire \audio_sample_lpf[4] ;
 wire \audio_sample_lpf[5] ;
 wire \audio_sample_lpf[6] ;
 wire \audio_sample_lpf[7] ;
 wire \audio_sample_lpf[8] ;
 wire \audio_sample_lpf[9] ;
 wire \bass_pha[0] ;
 wire \bass_pha[10] ;
 wire \bass_pha[11] ;
 wire \bass_pha[12] ;
 wire \bass_pha[13] ;
 wire \bass_pha[14] ;
 wire \bass_pha[15] ;
 wire \bass_pha[1] ;
 wire \bass_pha[2] ;
 wire \bass_pha[3] ;
 wire \bass_pha[4] ;
 wire \bass_pha[5] ;
 wire \bass_pha[6] ;
 wire \bass_pha[7] ;
 wire \bass_pha[8] ;
 wire \bass_pha[9] ;
 wire \bass_vol[0] ;
 wire \bass_vol[1] ;
 wire \bass_vol[2] ;
 wire \bass_vol[3] ;
 wire \bass_vol[4] ;
 wire \bass_vol[5] ;
 wire \cos[0] ;
 wire \cos[1] ;
 wire \cos[2] ;
 wire \cos[3] ;
 wire \cos[4] ;
 wire \cos[5] ;
 wire \cos[6] ;
 wire \frame_count[0] ;
 wire \frame_count[1] ;
 wire \frame_count[2] ;
 wire \frame_count[3] ;
 wire \frame_count[4] ;
 wire \frame_count[5] ;
 wire \frame_count[6] ;
 wire \frame_count[7] ;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \kick_ctr[0] ;
 wire \kick_ctr[1] ;
 wire \kick_osci[0] ;
 wire \kick_osci[1] ;
 wire \kick_osci[2] ;
 wire \kick_osci[3] ;
 wire \kick_osci[4] ;
 wire \kick_osci[5] ;
 wire \kick_osci[6] ;
 wire \kick_osci[7] ;
 wire \kick_osci[8] ;
 wire \line_lfsr[0] ;
 wire \line_lfsr[1] ;
 wire \line_lfsr[2] ;
 wire \line_lfsr[3] ;
 wire \line_lfsr[4] ;
 wire \line_lfsr[5] ;
 wire \line_lfsr[6] ;
 wire \nyan_x_offset[0] ;
 wire \nyan_x_offset[1] ;
 wire \nyan_x_offset[2] ;
 wire \nyan_x_offset[3] ;
 wire \nyan_x_offset[4] ;
 wire \nyanframe[0] ;
 wire \nyanframe[1] ;
 wire \nyanframe[2] ;
 wire \sample_beat_ctr[0] ;
 wire \sample_beat_ctr[1] ;
 wire \sample_beat_ctr[2] ;
 wire \sin[0] ;
 wire \sin[6] ;
 wire song_loops;
 wire \songpos[0] ;
 wire \songpos[1] ;
 wire \songpos[2] ;
 wire \songpos[3] ;
 wire \songpos[4] ;
 wire \songpos[5] ;
 wire \songpos[6] ;
 wire \songpos[7] ;
 wire \songpos[8] ;
 wire \sqr_pha[0] ;
 wire \sqr_pha[10] ;
 wire \sqr_pha[11] ;
 wire \sqr_pha[12] ;
 wire \sqr_pha[1] ;
 wire \sqr_pha[2] ;
 wire \sqr_pha[3] ;
 wire \sqr_pha[4] ;
 wire \sqr_pha[5] ;
 wire \sqr_pha[6] ;
 wire \sqr_pha[7] ;
 wire \sqr_pha[8] ;
 wire \sqr_pha[9] ;
 wire \sqr_vol[0] ;
 wire \sqr_vol[1] ;
 wire \sqr_vol[2] ;
 wire \sqr_vol[3] ;
 wire \sqr_vol[4] ;
 wire \sqr_vol[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_dfrbp_1 \B[0]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net138),
    .D(_0000_),
    .Q_N(_3038_),
    .Q(net9));
 sg13g2_dfrbp_1 \B[1]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_0001_),
    .Q_N(_3039_),
    .Q(net5));
 sg13g2_dfrbp_1 \G[0]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net138),
    .D(_0002_),
    .Q_N(_3040_),
    .Q(net8));
 sg13g2_dfrbp_1 \G[1]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_0003_),
    .Q_N(_3041_),
    .Q(net4));
 sg13g2_dfrbp_1 \R[0]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net138),
    .D(_0004_),
    .Q_N(_3042_),
    .Q(net7));
 sg13g2_dfrbp_1 \R[1]$_DFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_0005_),
    .Q_N(_3043_),
    .Q(net3));
 sg13g2_buf_1 _3057_ (.A(\hvsync_gen.vpos[3] ),
    .X(_2302_));
 sg13g2_buf_1 _3058_ (.A(_2302_),
    .X(_2303_));
 sg13g2_buf_2 _3059_ (.A(\songpos[1] ),
    .X(_2304_));
 sg13g2_inv_4 _3060_ (.A(_2304_),
    .Y(_2305_));
 sg13g2_buf_1 _3061_ (.A(\hvsync_gen.vpos[4] ),
    .X(_2306_));
 sg13g2_buf_2 _3062_ (.A(\songpos[2] ),
    .X(_2307_));
 sg13g2_xnor2_1 _3063_ (.Y(_2308_),
    .A(net122),
    .B(_2307_));
 sg13g2_nor3_1 _3064_ (.A(net111),
    .B(net110),
    .C(_2308_),
    .Y(_2309_));
 sg13g2_inv_2 _3065_ (.Y(_2310_),
    .A(net111));
 sg13g2_buf_1 _3066_ (.A(_2304_),
    .X(_2311_));
 sg13g2_inv_1 _3067_ (.Y(_2312_),
    .A(_2308_));
 sg13g2_a21oi_1 _3068_ (.A1(net100),
    .A2(net109),
    .Y(_2313_),
    .B1(_2312_));
 sg13g2_nor2_1 _3069_ (.A(_2309_),
    .B(_2313_),
    .Y(_2314_));
 sg13g2_buf_2 _3070_ (.A(\hvsync_gen.vpos[2] ),
    .X(_2315_));
 sg13g2_buf_1 _3071_ (.A(\songpos[0] ),
    .X(_2316_));
 sg13g2_inv_1 _3072_ (.Y(_2317_),
    .A(net121));
 sg13g2_xor2_1 _3073_ (.B(net109),
    .A(_2302_),
    .X(_2318_));
 sg13g2_nor3_1 _3074_ (.A(_2315_),
    .B(_2317_),
    .C(_2318_),
    .Y(_2319_));
 sg13g2_inv_1 _3075_ (.Y(_2320_),
    .A(_2315_));
 sg13g2_buf_1 _3076_ (.A(net121),
    .X(_2321_));
 sg13g2_inv_1 _3077_ (.Y(_2322_),
    .A(_2318_));
 sg13g2_a21oi_1 _3078_ (.A1(_2320_),
    .A2(net108),
    .Y(_2323_),
    .B1(_2322_));
 sg13g2_inv_1 _3079_ (.Y(_2324_),
    .A(_2323_));
 sg13g2_xor2_1 _3080_ (.B(net121),
    .A(_2315_),
    .X(_2325_));
 sg13g2_nand3b_1 _3081_ (.B(_2324_),
    .C(_2325_),
    .Y(_2326_),
    .A_N(_2319_));
 sg13g2_inv_1 _3082_ (.Y(_2327_),
    .A(_0036_));
 sg13g2_buf_1 _3083_ (.A(\hvsync_gen.vpos[1] ),
    .X(_2328_));
 sg13g2_xnor2_1 _3084_ (.Y(_2329_),
    .A(_2328_),
    .B(_2325_));
 sg13g2_o21ai_1 _3085_ (.B1(_2324_),
    .Y(_2330_),
    .A1(_2327_),
    .A2(_2329_));
 sg13g2_nand2b_1 _3086_ (.Y(_2331_),
    .B(_2330_),
    .A_N(_2319_));
 sg13g2_o21ai_1 _3087_ (.B1(_2331_),
    .Y(_2332_),
    .A1(_0036_),
    .A2(_2326_));
 sg13g2_xnor2_1 _3088_ (.Y(_2333_),
    .A(_2314_),
    .B(_2332_));
 sg13g2_buf_2 _3089_ (.A(song_loops),
    .X(_2334_));
 sg13g2_inv_1 _3090_ (.Y(_2335_),
    .A(_2334_));
 sg13g2_nand2_1 _3091_ (.Y(_2336_),
    .A(_2333_),
    .B(net107));
 sg13g2_buf_2 _3092_ (.A(\songpos[7] ),
    .X(_2337_));
 sg13g2_buf_1 _3093_ (.A(\songpos[6] ),
    .X(_2338_));
 sg13g2_nand2_1 _3094_ (.Y(_2339_),
    .A(_2337_),
    .B(net120));
 sg13g2_inv_2 _3095_ (.Y(_2340_),
    .A(_2339_));
 sg13g2_buf_1 _3096_ (.A(\songpos[5] ),
    .X(_2341_));
 sg13g2_buf_1 _3097_ (.A(\songpos[8] ),
    .X(_2342_));
 sg13g2_a21oi_1 _3098_ (.A1(_2340_),
    .A2(_2341_),
    .Y(_2343_),
    .B1(net118));
 sg13g2_buf_2 _3099_ (.A(_2343_),
    .X(_2344_));
 sg13g2_inv_2 _3100_ (.Y(_2345_),
    .A(net122));
 sg13g2_buf_1 _3101_ (.A(\nyanframe[1] ),
    .X(_2346_));
 sg13g2_inv_1 _3102_ (.Y(_2347_),
    .A(_0035_));
 sg13g2_nor2_1 _3103_ (.A(_2346_),
    .B(_2347_),
    .Y(_2348_));
 sg13g2_nand2_1 _3104_ (.Y(_2349_),
    .A(_2348_),
    .B(net111));
 sg13g2_xnor2_1 _3105_ (.Y(_2350_),
    .A(_2345_),
    .B(_2349_));
 sg13g2_nand2_1 _3106_ (.Y(_2351_),
    .A(_2350_),
    .B(_2334_));
 sg13g2_nor2_2 _3107_ (.A(net107),
    .B(_2344_),
    .Y(_2352_));
 sg13g2_nand2_1 _3108_ (.Y(_2353_),
    .A(_2315_),
    .B(_2316_));
 sg13g2_nor2_1 _3109_ (.A(_2353_),
    .B(_2322_),
    .Y(_2354_));
 sg13g2_nand2_1 _3110_ (.Y(_2355_),
    .A(_2302_),
    .B(net109));
 sg13g2_xnor2_1 _3111_ (.Y(_2356_),
    .A(_2355_),
    .B(_2308_));
 sg13g2_xnor2_1 _3112_ (.Y(_2357_),
    .A(_2354_),
    .B(_2356_));
 sg13g2_a22oi_1 _3113_ (.Y(_2358_),
    .B1(_2352_),
    .B2(_2357_),
    .A2(_2351_),
    .A1(_2344_));
 sg13g2_and2_1 _3114_ (.A(_2336_),
    .B(_2358_),
    .X(_2359_));
 sg13g2_buf_1 _3115_ (.A(_2359_),
    .X(_2360_));
 sg13g2_inv_1 _3116_ (.Y(_2361_),
    .A(_2325_));
 sg13g2_xnor2_1 _3117_ (.Y(_2362_),
    .A(_2327_),
    .B(_2329_));
 sg13g2_inv_1 _3118_ (.Y(_2363_),
    .A(_0037_));
 sg13g2_inv_1 _3119_ (.Y(_2364_),
    .A(_2344_));
 sg13g2_a21oi_1 _3120_ (.A1(_2334_),
    .A2(_2363_),
    .Y(_2365_),
    .B1(_2364_));
 sg13g2_a221oi_1 _3121_ (.B2(net107),
    .C1(_2365_),
    .B1(_2362_),
    .A1(_2361_),
    .Y(_2366_),
    .A2(_2352_));
 sg13g2_buf_1 _3122_ (.A(_2366_),
    .X(_2367_));
 sg13g2_nand2_1 _3123_ (.Y(_2368_),
    .A(_2322_),
    .B(_2353_));
 sg13g2_nand3b_1 _3124_ (.B(_2364_),
    .C(_2368_),
    .Y(_2369_),
    .A_N(_2354_));
 sg13g2_xnor2_1 _3125_ (.Y(_2370_),
    .A(net100),
    .B(_2348_));
 sg13g2_a21oi_1 _3126_ (.A1(_2370_),
    .A2(_2344_),
    .Y(_2371_),
    .B1(net107));
 sg13g2_a21oi_1 _3127_ (.A1(_2318_),
    .A2(_2361_),
    .Y(_2372_),
    .B1(_2344_));
 sg13g2_a21oi_1 _3128_ (.A1(_2326_),
    .A2(_2372_),
    .Y(_2373_),
    .B1(_2334_));
 sg13g2_a21oi_2 _3129_ (.B1(_2373_),
    .Y(_2374_),
    .A2(_2371_),
    .A1(_2369_));
 sg13g2_nor2b_1 _3130_ (.A(_2367_),
    .B_N(_2374_),
    .Y(_2375_));
 sg13g2_buf_8 _3131_ (.A(\hvsync_gen.hpos[4] ),
    .X(_2376_));
 sg13g2_buf_8 _3132_ (.A(\nyan_x_offset[4] ),
    .X(_2377_));
 sg13g2_xor2_1 _3133_ (.B(_2377_),
    .A(net117),
    .X(_2378_));
 sg13g2_buf_8 _3134_ (.A(\hvsync_gen.hpos[3] ),
    .X(_2379_));
 sg13g2_buf_8 _3135_ (.A(\nyan_x_offset[3] ),
    .X(_2380_));
 sg13g2_nand2_1 _3136_ (.Y(_2381_),
    .A(net116),
    .B(net115));
 sg13g2_inv_2 _3137_ (.Y(_2382_),
    .A(_2381_));
 sg13g2_nand2_1 _3138_ (.Y(_2383_),
    .A(_2378_),
    .B(_2382_));
 sg13g2_nand2_1 _3139_ (.Y(_2384_),
    .A(net117),
    .B(_2377_));
 sg13g2_buf_8 _3140_ (.A(\sin[6] ),
    .X(_2385_));
 sg13g2_xnor2_1 _3141_ (.Y(_2386_),
    .A(\hvsync_gen.hpos[5] ),
    .B(net114));
 sg13g2_a21oi_1 _3142_ (.A1(_2383_),
    .A2(_2384_),
    .Y(_2387_),
    .B1(_2386_));
 sg13g2_buf_1 _3143_ (.A(\hvsync_gen.hpos[1] ),
    .X(_2388_));
 sg13g2_nor2_1 _3144_ (.A(_2388_),
    .B(\nyan_x_offset[1] ),
    .Y(_2389_));
 sg13g2_buf_8 _3145_ (.A(\hvsync_gen.hpos[2] ),
    .X(_2390_));
 sg13g2_buf_8 _3146_ (.A(\nyan_x_offset[2] ),
    .X(_2391_));
 sg13g2_xnor2_1 _3147_ (.Y(_2392_),
    .A(_2390_),
    .B(_2391_));
 sg13g2_nor2_1 _3148_ (.A(_2389_),
    .B(_2392_),
    .Y(_2393_));
 sg13g2_xor2_1 _3149_ (.B(net115),
    .A(net116),
    .X(_2394_));
 sg13g2_nand2_1 _3150_ (.Y(_2395_),
    .A(_2390_),
    .B(_2391_));
 sg13g2_nand2b_1 _3151_ (.Y(_2396_),
    .B(_2394_),
    .A_N(_2395_));
 sg13g2_inv_1 _3152_ (.Y(_2397_),
    .A(_2396_));
 sg13g2_a21oi_1 _3153_ (.A1(_2393_),
    .A2(_2394_),
    .Y(_2398_),
    .B1(_2397_));
 sg13g2_inv_1 _3154_ (.Y(_2399_),
    .A(_2384_));
 sg13g2_xnor2_1 _3155_ (.Y(_2400_),
    .A(_2399_),
    .B(_2386_));
 sg13g2_xnor2_1 _3156_ (.Y(_2401_),
    .A(_2376_),
    .B(_2377_));
 sg13g2_xnor2_1 _3157_ (.Y(_2402_),
    .A(_2382_),
    .B(_2401_));
 sg13g2_nand2_1 _3158_ (.Y(_2403_),
    .A(_2400_),
    .B(_2402_));
 sg13g2_nor2_1 _3159_ (.A(_2398_),
    .B(_2403_),
    .Y(_2404_));
 sg13g2_nor2_1 _3160_ (.A(_2387_),
    .B(_2404_),
    .Y(_2405_));
 sg13g2_xor2_1 _3161_ (.B(_2391_),
    .A(_2390_),
    .X(_2406_));
 sg13g2_inv_2 _3162_ (.Y(_2407_),
    .A(_2389_));
 sg13g2_nand2_1 _3163_ (.Y(_2408_),
    .A(_2406_),
    .B(_2407_));
 sg13g2_nand2_1 _3164_ (.Y(_2409_),
    .A(_2392_),
    .B(_2389_));
 sg13g2_nand2_1 _3165_ (.Y(_2410_),
    .A(_2408_),
    .B(_2409_));
 sg13g2_xnor2_1 _3166_ (.Y(_2411_),
    .A(_2379_),
    .B(_2380_));
 sg13g2_nand2_1 _3167_ (.Y(_2412_),
    .A(_2411_),
    .B(_2395_));
 sg13g2_nand2_2 _3168_ (.Y(_2413_),
    .A(_2396_),
    .B(_2412_));
 sg13g2_nor2_1 _3169_ (.A(_2410_),
    .B(_2413_),
    .Y(_2414_));
 sg13g2_buf_1 _3170_ (.A(\hvsync_gen.hpos[5] ),
    .X(_2415_));
 sg13g2_xor2_1 _3171_ (.B(net114),
    .A(net113),
    .X(_2416_));
 sg13g2_nand2_1 _3172_ (.Y(_2417_),
    .A(_2416_),
    .B(_2399_));
 sg13g2_nand2_1 _3173_ (.Y(_2418_),
    .A(_2386_),
    .B(_2384_));
 sg13g2_nand2_1 _3174_ (.Y(_2419_),
    .A(_2417_),
    .B(_2418_));
 sg13g2_nand2_1 _3175_ (.Y(_2420_),
    .A(_2401_),
    .B(_2381_));
 sg13g2_nand2_2 _3176_ (.Y(_2421_),
    .A(_2383_),
    .B(_2420_));
 sg13g2_nor2_1 _3177_ (.A(_2419_),
    .B(_2421_),
    .Y(_2422_));
 sg13g2_buf_2 _3178_ (.A(\hvsync_gen.hpos[0] ),
    .X(_2423_));
 sg13g2_nand2_1 _3179_ (.Y(_2424_),
    .A(_2423_),
    .B(\nyan_x_offset[0] ));
 sg13g2_xnor2_1 _3180_ (.Y(_2425_),
    .A(_2388_),
    .B(\nyan_x_offset[1] ));
 sg13g2_nand2b_1 _3181_ (.Y(_2426_),
    .B(_2425_),
    .A_N(_2424_));
 sg13g2_inv_1 _3182_ (.Y(_2427_),
    .A(_2426_));
 sg13g2_nand3_1 _3183_ (.B(_2422_),
    .C(_2427_),
    .A(_2414_),
    .Y(_2428_));
 sg13g2_nand2_1 _3184_ (.Y(_2429_),
    .A(_2405_),
    .B(_2428_));
 sg13g2_inv_8 _3185_ (.Y(_2430_),
    .A(net114));
 sg13g2_buf_2 _3186_ (.A(\hvsync_gen.hpos[6] ),
    .X(_2431_));
 sg13g2_o21ai_1 _3187_ (.B1(_2431_),
    .Y(_2432_),
    .A1(net113),
    .A2(_2430_));
 sg13g2_inv_1 _3188_ (.Y(_2433_),
    .A(net113));
 sg13g2_inv_2 _3189_ (.Y(_2434_),
    .A(_2431_));
 sg13g2_nand3_1 _3190_ (.B(_2434_),
    .C(_2385_),
    .A(_2433_),
    .Y(_2435_));
 sg13g2_nand2_2 _3191_ (.Y(_2436_),
    .A(_2432_),
    .B(_2435_));
 sg13g2_inv_1 _3192_ (.Y(_2437_),
    .A(_2436_));
 sg13g2_nand2_1 _3193_ (.Y(_2438_),
    .A(_2429_),
    .B(_2437_));
 sg13g2_nand3_1 _3194_ (.B(_2428_),
    .C(_2436_),
    .A(_2405_),
    .Y(_2439_));
 sg13g2_nand2_1 _3195_ (.Y(_2440_),
    .A(_2438_),
    .B(_2439_));
 sg13g2_buf_8 _3196_ (.A(_2440_),
    .X(_2441_));
 sg13g2_buf_8 _3197_ (.A(net52),
    .X(_2442_));
 sg13g2_buf_8 _3198_ (.A(net46),
    .X(_2443_));
 sg13g2_buf_8 _3199_ (.A(net35),
    .X(_2444_));
 sg13g2_nor2_1 _3200_ (.A(_2426_),
    .B(_2410_),
    .Y(_2445_));
 sg13g2_inv_4 _3201_ (.A(_2413_),
    .Y(_2446_));
 sg13g2_nand2_1 _3202_ (.Y(_2447_),
    .A(_2445_),
    .B(_2446_));
 sg13g2_nand2_1 _3203_ (.Y(_2448_),
    .A(_2447_),
    .B(_2398_));
 sg13g2_nand2_2 _3204_ (.Y(_2449_),
    .A(_2448_),
    .B(_2402_));
 sg13g2_nand3_1 _3205_ (.B(_2398_),
    .C(_2421_),
    .A(_2447_),
    .Y(_2450_));
 sg13g2_buf_1 _3206_ (.A(_2450_),
    .X(_2451_));
 sg13g2_a21oi_1 _3207_ (.A1(_2427_),
    .A2(_2409_),
    .Y(_2452_),
    .B1(_2393_));
 sg13g2_xnor2_1 _3208_ (.Y(_2453_),
    .A(_2446_),
    .B(_2452_));
 sg13g2_a21oi_2 _3209_ (.B1(_2453_),
    .Y(_2454_),
    .A2(_2451_),
    .A1(_2449_));
 sg13g2_xnor2_1 _3210_ (.Y(_2455_),
    .A(_2427_),
    .B(_2410_));
 sg13g2_buf_2 _3211_ (.A(_2455_),
    .X(_2456_));
 sg13g2_inv_2 _3212_ (.Y(_2457_),
    .A(_2456_));
 sg13g2_nor2_1 _3213_ (.A(_2407_),
    .B(_2406_),
    .Y(_2458_));
 sg13g2_o21ai_1 _3214_ (.B1(_2408_),
    .Y(_2459_),
    .A1(_2426_),
    .A2(_2458_));
 sg13g2_nor2_1 _3215_ (.A(_2421_),
    .B(_2413_),
    .Y(_2460_));
 sg13g2_nand2_1 _3216_ (.Y(_2461_),
    .A(_2459_),
    .B(_2460_));
 sg13g2_a21oi_1 _3217_ (.A1(_2396_),
    .A2(_2381_),
    .Y(_2462_),
    .B1(_2401_));
 sg13g2_inv_1 _3218_ (.Y(_2463_),
    .A(_2462_));
 sg13g2_nand2_1 _3219_ (.Y(_2464_),
    .A(_2461_),
    .B(_2463_));
 sg13g2_nand2_1 _3220_ (.Y(_2465_),
    .A(_2464_),
    .B(_2400_));
 sg13g2_nand3_1 _3221_ (.B(_2419_),
    .C(_2463_),
    .A(_2461_),
    .Y(_2466_));
 sg13g2_nand2_1 _3222_ (.Y(_2467_),
    .A(_2465_),
    .B(_2466_));
 sg13g2_buf_8 _3223_ (.A(_2467_),
    .X(_2468_));
 sg13g2_buf_8 _3224_ (.A(net51),
    .X(_2469_));
 sg13g2_a21oi_1 _3225_ (.A1(_2454_),
    .A2(_2457_),
    .Y(_2470_),
    .B1(net45));
 sg13g2_xnor2_1 _3226_ (.Y(_2471_),
    .A(net28),
    .B(_2470_));
 sg13g2_xnor2_1 _3227_ (.Y(_2472_),
    .A(_2413_),
    .B(_2452_));
 sg13g2_buf_1 _3228_ (.A(_2472_),
    .X(_2473_));
 sg13g2_nand2_1 _3229_ (.Y(_2474_),
    .A(net65),
    .B(_2457_));
 sg13g2_nand2_1 _3230_ (.Y(_2475_),
    .A(_2449_),
    .B(_2451_));
 sg13g2_buf_8 _3231_ (.A(_2475_),
    .X(_2476_));
 sg13g2_xnor2_1 _3232_ (.Y(_2477_),
    .A(_2474_),
    .B(net50));
 sg13g2_buf_2 _3233_ (.A(\nyanframe[2] ),
    .X(_2478_));
 sg13g2_inv_1 _3234_ (.Y(_2479_),
    .A(_2346_));
 sg13g2_nor2_1 _3235_ (.A(_2478_),
    .B(_2479_),
    .Y(_2480_));
 sg13g2_buf_1 _3236_ (.A(\nyanframe[0] ),
    .X(_2481_));
 sg13g2_inv_2 _3237_ (.Y(_2482_),
    .A(_2481_));
 sg13g2_nor2_1 _3238_ (.A(_2346_),
    .B(_2482_),
    .Y(_2483_));
 sg13g2_inv_1 _3239_ (.Y(_2484_),
    .A(_2483_));
 sg13g2_nor2_1 _3240_ (.A(_2347_),
    .B(_2484_),
    .Y(_2485_));
 sg13g2_nor2_1 _3241_ (.A(_2480_),
    .B(_2485_),
    .Y(_2486_));
 sg13g2_nand2_1 _3242_ (.Y(_2487_),
    .A(_2486_),
    .B(_2334_));
 sg13g2_xnor2_1 _3243_ (.Y(_2488_),
    .A(_2456_),
    .B(net65));
 sg13g2_or2_1 _3244_ (.X(_2489_),
    .B(_2488_),
    .A(_2487_));
 sg13g2_buf_1 _3245_ (.A(_2489_),
    .X(_2490_));
 sg13g2_nor2_1 _3246_ (.A(_2477_),
    .B(_2490_),
    .Y(_2491_));
 sg13g2_inv_2 _3247_ (.Y(_2492_),
    .A(_2491_));
 sg13g2_nand2_1 _3248_ (.Y(_2493_),
    .A(_2464_),
    .B(_2419_));
 sg13g2_nand3_1 _3249_ (.B(_2400_),
    .C(_2463_),
    .A(_2461_),
    .Y(_2494_));
 sg13g2_nand2_1 _3250_ (.Y(_2495_),
    .A(_2493_),
    .B(_2494_));
 sg13g2_buf_8 _3251_ (.A(_2495_),
    .X(_2496_));
 sg13g2_nand2_1 _3252_ (.Y(_2497_),
    .A(net50),
    .B(net65));
 sg13g2_buf_8 _3253_ (.A(_2497_),
    .X(_2498_));
 sg13g2_nor2_2 _3254_ (.A(_2496_),
    .B(_2498_),
    .Y(_2499_));
 sg13g2_a21oi_1 _3255_ (.A1(_2457_),
    .A2(_2499_),
    .Y(_2500_),
    .B1(_2470_));
 sg13g2_inv_1 _3256_ (.Y(_2501_),
    .A(_2500_));
 sg13g2_nor2_1 _3257_ (.A(_2492_),
    .B(_2501_),
    .Y(_2502_));
 sg13g2_xnor2_1 _3258_ (.Y(_2503_),
    .A(_2471_),
    .B(_2502_));
 sg13g2_buf_1 _3259_ (.A(_2503_),
    .X(_2504_));
 sg13g2_nand2_1 _3260_ (.Y(_2505_),
    .A(_2490_),
    .B(_2477_));
 sg13g2_nand2_2 _3261_ (.Y(_2506_),
    .A(_2492_),
    .B(_2505_));
 sg13g2_nor2_1 _3262_ (.A(_2457_),
    .B(_2506_),
    .Y(_2507_));
 sg13g2_inv_1 _3263_ (.Y(_2508_),
    .A(_2507_));
 sg13g2_inv_2 _3264_ (.Y(_2509_),
    .A(_2506_));
 sg13g2_nor2_1 _3265_ (.A(_2457_),
    .B(_2509_),
    .Y(_2510_));
 sg13g2_nand2_1 _3266_ (.Y(_2511_),
    .A(net14),
    .B(_2510_));
 sg13g2_o21ai_1 _3267_ (.B1(_2511_),
    .Y(_2512_),
    .A1(net14),
    .A2(_2508_));
 sg13g2_inv_1 _3268_ (.Y(_2513_),
    .A(_2502_));
 sg13g2_nand2_1 _3269_ (.Y(_2514_),
    .A(_2501_),
    .B(_2492_));
 sg13g2_nand2_1 _3270_ (.Y(_2515_),
    .A(_2513_),
    .B(_2514_));
 sg13g2_buf_1 _3271_ (.A(_2515_),
    .X(_2516_));
 sg13g2_nand3_1 _3272_ (.B(net13),
    .C(_2374_),
    .A(_2512_),
    .Y(_2517_));
 sg13g2_nand2b_1 _3273_ (.Y(_2518_),
    .B(_2517_),
    .A_N(_2375_));
 sg13g2_nand2_1 _3274_ (.Y(_2519_),
    .A(net50),
    .B(_2453_));
 sg13g2_nand3_1 _3275_ (.B(_2451_),
    .C(_2473_),
    .A(_2449_),
    .Y(_2520_));
 sg13g2_buf_2 _3276_ (.A(_2520_),
    .X(_2521_));
 sg13g2_nand2_1 _3277_ (.Y(_2522_),
    .A(_2519_),
    .B(_2521_));
 sg13g2_nand2_1 _3278_ (.Y(_2523_),
    .A(_2488_),
    .B(_2487_));
 sg13g2_nand2_1 _3279_ (.Y(_2524_),
    .A(_2490_),
    .B(_2523_));
 sg13g2_nor2_1 _3280_ (.A(_2456_),
    .B(_2524_),
    .Y(_2525_));
 sg13g2_inv_1 _3281_ (.Y(_2526_),
    .A(_2525_));
 sg13g2_nor2_1 _3282_ (.A(_2522_),
    .B(_2526_),
    .Y(_2527_));
 sg13g2_nor2_1 _3283_ (.A(_2527_),
    .B(net13),
    .Y(_2528_));
 sg13g2_nor2_1 _3284_ (.A(_2477_),
    .B(_2524_),
    .Y(_2529_));
 sg13g2_inv_1 _3285_ (.Y(_2530_),
    .A(_2524_));
 sg13g2_nor2_1 _3286_ (.A(_2530_),
    .B(_2509_),
    .Y(_2531_));
 sg13g2_nor2_1 _3287_ (.A(_2529_),
    .B(_2531_),
    .Y(_2532_));
 sg13g2_inv_1 _3288_ (.Y(_2533_),
    .A(_2532_));
 sg13g2_o21ai_1 _3289_ (.B1(net13),
    .Y(_2534_),
    .A1(_2456_),
    .A2(_2533_));
 sg13g2_nand2b_1 _3290_ (.Y(_2535_),
    .B(_2534_),
    .A_N(_2528_));
 sg13g2_nand3_1 _3291_ (.B(_2457_),
    .C(_2524_),
    .A(_2506_),
    .Y(_2536_));
 sg13g2_inv_4 _3292_ (.A(net13),
    .Y(_2537_));
 sg13g2_nor2_1 _3293_ (.A(_2536_),
    .B(_2537_),
    .Y(_2538_));
 sg13g2_a21oi_1 _3294_ (.A1(_2538_),
    .A2(net14),
    .Y(_2539_),
    .B1(_2367_));
 sg13g2_o21ai_1 _3295_ (.B1(_2539_),
    .Y(_2540_),
    .A1(net14),
    .A2(_2535_));
 sg13g2_nand2_1 _3296_ (.Y(_2541_),
    .A(_2530_),
    .B(_2456_));
 sg13g2_nor2_1 _3297_ (.A(net50),
    .B(_2541_),
    .Y(_2542_));
 sg13g2_nor2_1 _3298_ (.A(_2457_),
    .B(_2537_),
    .Y(_2543_));
 sg13g2_a22oi_1 _3299_ (.Y(_2544_),
    .B1(_2532_),
    .B2(_2543_),
    .A2(_2542_),
    .A1(_2537_));
 sg13g2_inv_1 _3300_ (.Y(_2545_),
    .A(_2503_));
 sg13g2_nand2b_1 _3301_ (.Y(_2546_),
    .B(_2545_),
    .A_N(_2544_));
 sg13g2_nor2_1 _3302_ (.A(_2457_),
    .B(_2530_),
    .Y(_2547_));
 sg13g2_nand2_1 _3303_ (.Y(_2548_),
    .A(_2506_),
    .B(_2547_));
 sg13g2_inv_1 _3304_ (.Y(_2549_),
    .A(_2548_));
 sg13g2_nand3_1 _3305_ (.B(net13),
    .C(_2549_),
    .A(net14),
    .Y(_2550_));
 sg13g2_nand2_1 _3306_ (.Y(_2551_),
    .A(_2546_),
    .B(_2550_));
 sg13g2_nor2b_1 _3307_ (.A(_2374_),
    .B_N(_2367_),
    .Y(_2552_));
 sg13g2_a22oi_1 _3308_ (.Y(_2553_),
    .B1(_2551_),
    .B2(_2552_),
    .A2(_2540_),
    .A1(_2518_));
 sg13g2_nor2_1 _3309_ (.A(_2436_),
    .B(_2419_),
    .Y(_2554_));
 sg13g2_o21ai_1 _3310_ (.B1(_2432_),
    .Y(_2555_),
    .A1(_2417_),
    .A2(_2436_));
 sg13g2_a21oi_1 _3311_ (.A1(_2462_),
    .A2(_2554_),
    .Y(_2556_),
    .B1(_2555_));
 sg13g2_nand3_1 _3312_ (.B(_2460_),
    .C(_2554_),
    .A(_2459_),
    .Y(_2557_));
 sg13g2_nand2_1 _3313_ (.Y(_2558_),
    .A(_2556_),
    .B(_2557_));
 sg13g2_buf_2 _3314_ (.A(\hvsync_gen.hpos[7] ),
    .X(_2559_));
 sg13g2_nand2_1 _3315_ (.Y(_2560_),
    .A(_2558_),
    .B(_2559_));
 sg13g2_inv_1 _3316_ (.Y(_2561_),
    .A(_2559_));
 sg13g2_nand3_1 _3317_ (.B(_2557_),
    .C(_2561_),
    .A(_2556_),
    .Y(_2562_));
 sg13g2_nand2_1 _3318_ (.Y(_2563_),
    .A(_2560_),
    .B(_2562_));
 sg13g2_buf_8 _3319_ (.A(_2563_),
    .X(_2564_));
 sg13g2_buf_8 _3320_ (.A(_2564_),
    .X(_2565_));
 sg13g2_buf_8 _3321_ (.A(net44),
    .X(_2566_));
 sg13g2_buf_8 _3322_ (.A(net34),
    .X(_2567_));
 sg13g2_buf_8 _3323_ (.A(net27),
    .X(_2568_));
 sg13g2_buf_8 _3324_ (.A(net21),
    .X(_2569_));
 sg13g2_nand2_1 _3325_ (.Y(_2570_),
    .A(_2429_),
    .B(_2436_));
 sg13g2_nand3_1 _3326_ (.B(_2428_),
    .C(_2437_),
    .A(_2405_),
    .Y(_2571_));
 sg13g2_nand2_1 _3327_ (.Y(_2572_),
    .A(_2570_),
    .B(_2571_));
 sg13g2_buf_8 _3328_ (.A(_2572_),
    .X(_2573_));
 sg13g2_buf_8 _3329_ (.A(_2573_),
    .X(_2574_));
 sg13g2_buf_8 _3330_ (.A(net43),
    .X(_2575_));
 sg13g2_buf_8 _3331_ (.A(net33),
    .X(_2576_));
 sg13g2_buf_8 _3332_ (.A(net26),
    .X(_2577_));
 sg13g2_nor2_1 _3333_ (.A(net20),
    .B(_2470_),
    .Y(_2578_));
 sg13g2_xnor2_1 _3334_ (.Y(_2579_),
    .A(net17),
    .B(_2578_));
 sg13g2_nand2_1 _3335_ (.Y(_2580_),
    .A(_2502_),
    .B(net28));
 sg13g2_nor2_1 _3336_ (.A(_2579_),
    .B(_2580_),
    .Y(_2581_));
 sg13g2_buf_2 _3337_ (.A(\hvsync_gen.hpos[8] ),
    .X(_2582_));
 sg13g2_inv_2 _3338_ (.Y(_2583_),
    .A(_2582_));
 sg13g2_nor2_1 _3339_ (.A(_0038_),
    .B(_2436_),
    .Y(_2584_));
 sg13g2_nor2b_1 _3340_ (.A(_2403_),
    .B_N(_2584_),
    .Y(_2585_));
 sg13g2_nand2_1 _3341_ (.Y(_2586_),
    .A(_2448_),
    .B(_2585_));
 sg13g2_nor2_1 _3342_ (.A(_0038_),
    .B(_2432_),
    .Y(_2587_));
 sg13g2_a21oi_1 _3343_ (.A1(_2387_),
    .A2(_2584_),
    .Y(_2588_),
    .B1(_2587_));
 sg13g2_nand2_1 _3344_ (.Y(_2589_),
    .A(_2586_),
    .B(_2588_));
 sg13g2_xnor2_1 _3345_ (.Y(_2590_),
    .A(_2583_),
    .B(_2589_));
 sg13g2_buf_8 _3346_ (.A(_2590_),
    .X(_2591_));
 sg13g2_buf_8 _3347_ (.A(net42),
    .X(_2592_));
 sg13g2_buf_1 _3348_ (.A(net32),
    .X(_2593_));
 sg13g2_buf_1 _3349_ (.A(net25),
    .X(_2594_));
 sg13g2_nor3_1 _3350_ (.A(net19),
    .B(net17),
    .C(_2578_),
    .Y(_2595_));
 sg13g2_o21ai_1 _3351_ (.B1(net19),
    .Y(_2596_),
    .A1(net17),
    .A2(_2578_));
 sg13g2_nand2b_1 _3352_ (.Y(_2597_),
    .B(_2596_),
    .A_N(_2595_));
 sg13g2_buf_2 _3353_ (.A(\hvsync_gen.hpos[9] ),
    .X(_2598_));
 sg13g2_nand2_1 _3354_ (.Y(_2599_),
    .A(_2560_),
    .B(_2583_));
 sg13g2_xnor2_1 _3355_ (.Y(_2600_),
    .A(_2598_),
    .B(_2599_));
 sg13g2_inv_1 _3356_ (.Y(_2601_),
    .A(_2600_));
 sg13g2_xnor2_1 _3357_ (.Y(_2602_),
    .A(_2601_),
    .B(_2596_));
 sg13g2_a21oi_1 _3358_ (.A1(_2581_),
    .A2(_2597_),
    .Y(_2603_),
    .B1(_2602_));
 sg13g2_buf_2 _3359_ (.A(\hvsync_gen.vpos[7] ),
    .X(_2604_));
 sg13g2_inv_1 _3360_ (.Y(_2605_),
    .A(net119));
 sg13g2_buf_1 _3361_ (.A(_2605_),
    .X(_2606_));
 sg13g2_nor2_1 _3362_ (.A(_2604_),
    .B(_2606_),
    .Y(_2607_));
 sg13g2_buf_2 _3363_ (.A(\hvsync_gen.vpos[8] ),
    .X(_2608_));
 sg13g2_nor2_1 _3364_ (.A(_2608_),
    .B(net120),
    .Y(_2609_));
 sg13g2_inv_1 _3365_ (.Y(_2610_),
    .A(_2609_));
 sg13g2_nand2_1 _3366_ (.Y(_2611_),
    .A(_2608_),
    .B(net120));
 sg13g2_nand2_1 _3367_ (.Y(_2612_),
    .A(_2610_),
    .B(_2611_));
 sg13g2_xor2_1 _3368_ (.B(_2612_),
    .A(_2607_),
    .X(_2613_));
 sg13g2_buf_1 _3369_ (.A(\songpos[4] ),
    .X(_2614_));
 sg13g2_buf_1 _3370_ (.A(_2614_),
    .X(_2615_));
 sg13g2_inv_1 _3371_ (.Y(_2616_),
    .A(net106));
 sg13g2_buf_1 _3372_ (.A(_2616_),
    .X(_2617_));
 sg13g2_buf_1 _3373_ (.A(net91),
    .X(_2618_));
 sg13g2_buf_2 _3374_ (.A(\hvsync_gen.vpos[6] ),
    .X(_2619_));
 sg13g2_nand2_1 _3375_ (.Y(_2620_),
    .A(_2618_),
    .B(_2619_));
 sg13g2_xnor2_1 _3376_ (.Y(_2621_),
    .A(_2604_),
    .B(net119));
 sg13g2_nor2_1 _3377_ (.A(_2620_),
    .B(_2621_),
    .Y(_2622_));
 sg13g2_buf_1 _3378_ (.A(\hvsync_gen.vpos[5] ),
    .X(_2623_));
 sg13g2_inv_1 _3379_ (.Y(_2624_),
    .A(net112));
 sg13g2_buf_1 _3380_ (.A(\songpos[3] ),
    .X(_2625_));
 sg13g2_buf_1 _3381_ (.A(_2625_),
    .X(_2626_));
 sg13g2_buf_1 _3382_ (.A(net104),
    .X(_2627_));
 sg13g2_xor2_1 _3383_ (.B(_2615_),
    .A(_2619_),
    .X(_2628_));
 sg13g2_nor3_1 _3384_ (.A(net105),
    .B(_2627_),
    .C(_2628_),
    .Y(_2629_));
 sg13g2_nor2_1 _3385_ (.A(_2622_),
    .B(_2629_),
    .Y(_2630_));
 sg13g2_nand2_1 _3386_ (.Y(_2631_),
    .A(_2332_),
    .B(_2314_));
 sg13g2_buf_1 _3387_ (.A(_2307_),
    .X(_2632_));
 sg13g2_xor2_1 _3388_ (.B(net104),
    .A(net112),
    .X(_2633_));
 sg13g2_nor3_1 _3389_ (.A(_2345_),
    .B(net103),
    .C(_2633_),
    .Y(_2634_));
 sg13g2_nor2_1 _3390_ (.A(_2313_),
    .B(_2634_),
    .Y(_2635_));
 sg13g2_inv_1 _3391_ (.Y(_2636_),
    .A(_2307_));
 sg13g2_buf_8 _3392_ (.A(_2636_),
    .X(_2637_));
 sg13g2_inv_1 _3393_ (.Y(_2638_),
    .A(_2633_));
 sg13g2_a21oi_1 _3394_ (.A1(net122),
    .A2(_2637_),
    .Y(_2639_),
    .B1(_2638_));
 sg13g2_a21oi_1 _3395_ (.A1(_2631_),
    .A2(_2635_),
    .Y(_2640_),
    .B1(_2639_));
 sg13g2_inv_2 _3396_ (.Y(_2641_),
    .A(_2625_));
 sg13g2_buf_1 _3397_ (.A(_2641_),
    .X(_2642_));
 sg13g2_inv_1 _3398_ (.Y(_2643_),
    .A(_2628_));
 sg13g2_a21oi_1 _3399_ (.A1(net112),
    .A2(_2642_),
    .Y(_2644_),
    .B1(_2643_));
 sg13g2_nor2_1 _3400_ (.A(_2629_),
    .B(_2644_),
    .Y(_2645_));
 sg13g2_nand2_1 _3401_ (.Y(_2646_),
    .A(_2640_),
    .B(_2645_));
 sg13g2_a22oi_1 _3402_ (.Y(_2647_),
    .B1(_2630_),
    .B2(_2646_),
    .A2(_2621_),
    .A1(_2620_));
 sg13g2_xnor2_1 _3403_ (.Y(_2648_),
    .A(_2613_),
    .B(_2647_));
 sg13g2_inv_1 _3404_ (.Y(_2649_),
    .A(_2608_));
 sg13g2_nand2_1 _3405_ (.Y(_2650_),
    .A(_2649_),
    .B(_2338_));
 sg13g2_buf_1 _3406_ (.A(\hvsync_gen.vpos[9] ),
    .X(_2651_));
 sg13g2_xnor2_1 _3407_ (.Y(_2652_),
    .A(_2651_),
    .B(_2337_));
 sg13g2_xnor2_1 _3408_ (.Y(_2653_),
    .A(_2650_),
    .B(_2652_));
 sg13g2_nor2_1 _3409_ (.A(_2607_),
    .B(_2612_),
    .Y(_2654_));
 sg13g2_nor2_1 _3410_ (.A(_2622_),
    .B(_2654_),
    .Y(_2655_));
 sg13g2_nor2_1 _3411_ (.A(_2313_),
    .B(_2323_),
    .Y(_2656_));
 sg13g2_a21oi_1 _3412_ (.A1(_2326_),
    .A2(_2656_),
    .Y(_2657_),
    .B1(_2309_));
 sg13g2_nor2_1 _3413_ (.A(_2634_),
    .B(_2639_),
    .Y(_2658_));
 sg13g2_nand2_1 _3414_ (.Y(_2659_),
    .A(_2657_),
    .B(_2658_));
 sg13g2_nor2_1 _3415_ (.A(_2634_),
    .B(_2629_),
    .Y(_2660_));
 sg13g2_a21oi_1 _3416_ (.A1(_2659_),
    .A2(_2660_),
    .Y(_2661_),
    .B1(_2644_));
 sg13g2_xor2_1 _3417_ (.B(_2621_),
    .A(_2620_),
    .X(_2662_));
 sg13g2_nand2_1 _3418_ (.Y(_2663_),
    .A(_2661_),
    .B(_2662_));
 sg13g2_a22oi_1 _3419_ (.Y(_2664_),
    .B1(_2655_),
    .B2(_2663_),
    .A2(_2612_),
    .A1(_2607_));
 sg13g2_xnor2_1 _3420_ (.Y(_2665_),
    .A(_2653_),
    .B(_2664_));
 sg13g2_a21oi_1 _3421_ (.A1(_2648_),
    .A2(_2665_),
    .Y(_2666_),
    .B1(_2334_));
 sg13g2_inv_2 _3422_ (.Y(_2667_),
    .A(_2604_));
 sg13g2_nand2_1 _3423_ (.Y(_2668_),
    .A(net112),
    .B(_2619_));
 sg13g2_nand2_1 _3424_ (.Y(_2669_),
    .A(_2349_),
    .B(_0039_));
 sg13g2_nand2b_1 _3425_ (.Y(_2670_),
    .B(_2669_),
    .A_N(_2668_));
 sg13g2_xnor2_1 _3426_ (.Y(_2671_),
    .A(_2667_),
    .B(_2670_));
 sg13g2_nand2_1 _3427_ (.Y(_2672_),
    .A(_2349_),
    .B(_2345_));
 sg13g2_nand2_1 _3428_ (.Y(_2673_),
    .A(_2672_),
    .B(net112));
 sg13g2_xnor2_1 _3429_ (.Y(_2674_),
    .A(_0040_),
    .B(_2673_));
 sg13g2_nand3_1 _3430_ (.B(_2674_),
    .C(_2344_),
    .A(_2671_),
    .Y(_2675_));
 sg13g2_nand2_1 _3431_ (.Y(_2676_),
    .A(net112),
    .B(net98));
 sg13g2_xnor2_1 _3432_ (.Y(_2677_),
    .A(_2676_),
    .B(_2628_));
 sg13g2_nor2_1 _3433_ (.A(_2355_),
    .B(_2312_),
    .Y(_2678_));
 sg13g2_a21oi_1 _3434_ (.A1(_2356_),
    .A2(_2354_),
    .Y(_2679_),
    .B1(_2678_));
 sg13g2_nand2_1 _3435_ (.Y(_2680_),
    .A(_2345_),
    .B(_2637_));
 sg13g2_xor2_1 _3436_ (.B(_2633_),
    .A(_2680_),
    .X(_2681_));
 sg13g2_nand2b_1 _3437_ (.Y(_2682_),
    .B(_2681_),
    .A_N(_2679_));
 sg13g2_nand2_1 _3438_ (.Y(_2683_),
    .A(_2633_),
    .B(_2680_));
 sg13g2_nand2_1 _3439_ (.Y(_2684_),
    .A(_2682_),
    .B(_2683_));
 sg13g2_xor2_1 _3440_ (.B(_2684_),
    .A(_2677_),
    .X(_2685_));
 sg13g2_buf_1 _3441_ (.A(net106),
    .X(_2686_));
 sg13g2_nand2_1 _3442_ (.Y(_2687_),
    .A(_2619_),
    .B(net95));
 sg13g2_xnor2_1 _3443_ (.Y(_2688_),
    .A(_2687_),
    .B(_2621_));
 sg13g2_nand2_1 _3444_ (.Y(_2689_),
    .A(_2684_),
    .B(_2677_));
 sg13g2_o21ai_1 _3445_ (.B1(_2689_),
    .Y(_2690_),
    .A1(_2643_),
    .A2(_2676_));
 sg13g2_xor2_1 _3446_ (.B(_2690_),
    .A(_2688_),
    .X(_2691_));
 sg13g2_nor3_1 _3447_ (.A(_2335_),
    .B(_2685_),
    .C(_2691_),
    .Y(_2692_));
 sg13g2_or2_1 _3448_ (.X(_2693_),
    .B(_2661_),
    .A(_2662_));
 sg13g2_or2_1 _3449_ (.X(_2694_),
    .B(_2640_),
    .A(_2645_));
 sg13g2_a221oi_1 _3450_ (.B2(_2646_),
    .C1(_2334_),
    .B1(_2694_),
    .A1(_2663_),
    .Y(_2695_),
    .A2(_2693_));
 sg13g2_o21ai_1 _3451_ (.B1(_2364_),
    .Y(_2696_),
    .A1(_2692_),
    .A2(_2695_));
 sg13g2_o21ai_1 _3452_ (.B1(_2696_),
    .Y(_2697_),
    .A1(net107),
    .A2(_2675_));
 sg13g2_xnor2_1 _3453_ (.Y(_2698_),
    .A(_2609_),
    .B(_2652_));
 sg13g2_inv_1 _3454_ (.Y(_2699_),
    .A(_2621_));
 sg13g2_nand2_1 _3455_ (.Y(_2700_),
    .A(_2690_),
    .B(_2688_));
 sg13g2_o21ai_1 _3456_ (.B1(_2700_),
    .Y(_2701_),
    .A1(_2699_),
    .A2(_2687_));
 sg13g2_a22oi_1 _3457_ (.Y(_2702_),
    .B1(_2611_),
    .B2(_2610_),
    .A2(_2606_),
    .A1(_2667_));
 sg13g2_nor3_1 _3458_ (.A(_2604_),
    .B(net119),
    .C(_2612_),
    .Y(_2703_));
 sg13g2_nor2_1 _3459_ (.A(_2702_),
    .B(_2703_),
    .Y(_2704_));
 sg13g2_a21oi_1 _3460_ (.A1(_2701_),
    .A2(_2704_),
    .Y(_2705_),
    .B1(_2702_));
 sg13g2_nor2_1 _3461_ (.A(_2698_),
    .B(_2705_),
    .Y(_2706_));
 sg13g2_nor2b_1 _3462_ (.A(_2702_),
    .B_N(_2698_),
    .Y(_2707_));
 sg13g2_nor3_1 _3463_ (.A(_2704_),
    .B(_2707_),
    .C(_2701_),
    .Y(_2708_));
 sg13g2_a21oi_1 _3464_ (.A1(_2701_),
    .A2(_2704_),
    .Y(_2709_),
    .B1(_2708_));
 sg13g2_o21ai_1 _3465_ (.B1(_2352_),
    .Y(_2710_),
    .A1(_2706_),
    .A2(_2709_));
 sg13g2_nor2_1 _3466_ (.A(_2471_),
    .B(net13),
    .Y(_2711_));
 sg13g2_inv_1 _3467_ (.Y(_2712_),
    .A(_2360_));
 sg13g2_nor2_1 _3468_ (.A(_2374_),
    .B(_2367_),
    .Y(_2713_));
 sg13g2_o21ai_1 _3469_ (.B1(_2649_),
    .Y(_2714_),
    .A1(_2667_),
    .A2(_2670_));
 sg13g2_inv_1 _3470_ (.Y(_2715_),
    .A(_2619_));
 sg13g2_inv_2 _3471_ (.Y(_2716_),
    .A(_2651_));
 sg13g2_nor3_1 _3472_ (.A(_2667_),
    .B(_2715_),
    .C(_2716_),
    .Y(_2717_));
 sg13g2_nor2_1 _3473_ (.A(_2717_),
    .B(_2714_),
    .Y(_2718_));
 sg13g2_a21oi_1 _3474_ (.A1(_2651_),
    .A2(_2714_),
    .Y(_2719_),
    .B1(_2718_));
 sg13g2_inv_1 _3475_ (.Y(_2720_),
    .A(_0041_));
 sg13g2_xnor2_1 _3476_ (.Y(_2721_),
    .A(_2720_),
    .B(_2669_));
 sg13g2_nor3_2 _3477_ (.A(_2667_),
    .B(_2649_),
    .C(_2668_),
    .Y(_2722_));
 sg13g2_a221oi_1 _3478_ (.B2(_2649_),
    .C1(net107),
    .B1(_2673_),
    .A1(_2722_),
    .Y(_2723_),
    .A2(_2672_));
 sg13g2_nand3_1 _3479_ (.B(_2721_),
    .C(_2723_),
    .A(_2719_),
    .Y(_2724_));
 sg13g2_xnor2_1 _3480_ (.Y(_2725_),
    .A(_2658_),
    .B(_2657_));
 sg13g2_nand2_1 _3481_ (.Y(_2726_),
    .A(_2725_),
    .B(_2364_));
 sg13g2_inv_1 _3482_ (.Y(_2727_),
    .A(_2681_));
 sg13g2_nand2_1 _3483_ (.Y(_2728_),
    .A(_2682_),
    .B(_2352_));
 sg13g2_a21oi_1 _3484_ (.A1(_2727_),
    .A2(_2679_),
    .Y(_2729_),
    .B1(_2728_));
 sg13g2_a221oi_1 _3485_ (.B2(net107),
    .C1(_2729_),
    .B1(_2726_),
    .A1(_2724_),
    .Y(_2730_),
    .A2(_2344_));
 sg13g2_o21ai_1 _3486_ (.B1(_2730_),
    .Y(_2731_),
    .A1(_2712_),
    .A2(_2713_));
 sg13g2_nor2_1 _3487_ (.A(_2711_),
    .B(_2731_),
    .Y(_2732_));
 sg13g2_nand3_1 _3488_ (.B(_2710_),
    .C(_2732_),
    .A(_2697_),
    .Y(_2733_));
 sg13g2_nor3_1 _3489_ (.A(_2603_),
    .B(_2666_),
    .C(_2733_),
    .Y(_2734_));
 sg13g2_nand3b_1 _3490_ (.B(_2580_),
    .C(_2579_),
    .Y(_2735_),
    .A_N(_2597_));
 sg13g2_nand2_1 _3491_ (.Y(_2736_),
    .A(_2735_),
    .B(_2602_));
 sg13g2_nand2_1 _3492_ (.Y(_2737_),
    .A(_2734_),
    .B(_2736_));
 sg13g2_nor3_2 _3493_ (.A(_2360_),
    .B(_2553_),
    .C(_2737_),
    .Y(_2738_));
 sg13g2_nor2_1 _3494_ (.A(_2547_),
    .B(_2506_),
    .Y(_2739_));
 sg13g2_nor3_1 _3495_ (.A(_2739_),
    .B(_2537_),
    .C(_2545_),
    .Y(_2740_));
 sg13g2_nor2_1 _3496_ (.A(_2525_),
    .B(_2509_),
    .Y(_2741_));
 sg13g2_a221oi_1 _3497_ (.B2(_2548_),
    .C1(net14),
    .B1(_2528_),
    .A1(_2516_),
    .Y(_2742_),
    .A2(_2741_));
 sg13g2_nor3_1 _3498_ (.A(_2712_),
    .B(_2740_),
    .C(_2742_),
    .Y(_2743_));
 sg13g2_nor2_1 _3499_ (.A(_2743_),
    .B(_2737_),
    .Y(_2744_));
 sg13g2_a21oi_1 _3500_ (.A1(_2504_),
    .A2(_2549_),
    .Y(_2745_),
    .B1(_2374_));
 sg13g2_nand2_1 _3501_ (.Y(_2746_),
    .A(_2546_),
    .B(_2745_));
 sg13g2_nand2_1 _3502_ (.Y(_2747_),
    .A(net13),
    .B(_2508_));
 sg13g2_a21oi_1 _3503_ (.A1(_2537_),
    .A2(_2533_),
    .Y(_2748_),
    .B1(net14));
 sg13g2_o21ai_1 _3504_ (.B1(_2748_),
    .Y(_2749_),
    .A1(_2531_),
    .A2(_2747_));
 sg13g2_o21ai_1 _3505_ (.B1(net14),
    .Y(_2750_),
    .A1(_2529_),
    .A2(_2510_));
 sg13g2_nand3_1 _3506_ (.B(_2374_),
    .C(_2750_),
    .A(_2749_),
    .Y(_2751_));
 sg13g2_nand3_1 _3507_ (.B(_2367_),
    .C(_2751_),
    .A(_2746_),
    .Y(_2752_));
 sg13g2_nor2_1 _3508_ (.A(_2530_),
    .B(_2507_),
    .Y(_2753_));
 sg13g2_o21ai_1 _3509_ (.B1(net13),
    .Y(_2754_),
    .A1(_2456_),
    .A2(_2509_));
 sg13g2_o21ai_1 _3510_ (.B1(_2541_),
    .Y(_2755_),
    .A1(_2753_),
    .A2(_2754_));
 sg13g2_a21oi_1 _3511_ (.A1(_2753_),
    .A2(_2754_),
    .Y(_2756_),
    .B1(_2755_));
 sg13g2_nand2b_1 _3512_ (.Y(_2757_),
    .B(_2536_),
    .A_N(_2527_));
 sg13g2_o21ai_1 _3513_ (.B1(_2375_),
    .Y(_2758_),
    .A1(_2757_),
    .A2(_2545_));
 sg13g2_nand2b_1 _3514_ (.Y(_2759_),
    .B(_2758_),
    .A_N(_2711_));
 sg13g2_o21ai_1 _3515_ (.B1(_2759_),
    .Y(_2760_),
    .A1(_2504_),
    .A2(_2756_));
 sg13g2_a21o_1 _3516_ (.A2(_2760_),
    .A1(_2752_),
    .B1(_2360_),
    .X(_2761_));
 sg13g2_nand2_2 _3517_ (.Y(_2762_),
    .A(_2744_),
    .B(_2761_));
 sg13g2_inv_2 _3518_ (.Y(_2763_),
    .A(_2762_));
 sg13g2_nor2_1 _3519_ (.A(_2738_),
    .B(_2763_),
    .Y(_2764_));
 sg13g2_buf_1 _3520_ (.A(\hvsync_gen.vpos[0] ),
    .X(_2765_));
 sg13g2_xnor2_1 _3521_ (.Y(_2766_),
    .A(_2765_),
    .B(_2423_));
 sg13g2_inv_1 _3522_ (.Y(_2767_),
    .A(_2766_));
 sg13g2_nand2_1 _3523_ (.Y(_2768_),
    .A(_2302_),
    .B(net122));
 sg13g2_buf_1 _3524_ (.A(_2768_),
    .X(_2769_));
 sg13g2_xnor2_1 _3525_ (.Y(_2770_),
    .A(net105),
    .B(net94));
 sg13g2_inv_2 _3526_ (.Y(_2771_),
    .A(_2770_));
 sg13g2_inv_1 _3527_ (.Y(_2772_),
    .A(net94));
 sg13g2_a21oi_1 _3528_ (.A1(_2772_),
    .A2(_2624_),
    .Y(_2773_),
    .B1(_2720_));
 sg13g2_nand2b_1 _3529_ (.Y(_2774_),
    .B(_2619_),
    .A_N(_2773_));
 sg13g2_nand2_1 _3530_ (.Y(_2775_),
    .A(_2773_),
    .B(_2715_));
 sg13g2_nand2_1 _3531_ (.Y(_2776_),
    .A(_2774_),
    .B(_2775_));
 sg13g2_buf_2 _3532_ (.A(_2776_),
    .X(_2777_));
 sg13g2_nor2_1 _3533_ (.A(_2771_),
    .B(_2777_),
    .Y(_2778_));
 sg13g2_buf_1 _3534_ (.A(_2778_),
    .X(_2779_));
 sg13g2_inv_2 _3535_ (.Y(_2780_),
    .A(net57));
 sg13g2_nand3_1 _3536_ (.B(_2521_),
    .C(net51),
    .A(_2519_),
    .Y(_2781_));
 sg13g2_buf_2 _3537_ (.A(_2781_),
    .X(_2782_));
 sg13g2_nand2_1 _3538_ (.Y(_2783_),
    .A(_2782_),
    .B(net46));
 sg13g2_nor2_2 _3539_ (.A(net65),
    .B(net50),
    .Y(_2784_));
 sg13g2_nand2_1 _3540_ (.Y(_2785_),
    .A(_2784_),
    .B(net51));
 sg13g2_buf_8 _3541_ (.A(_2785_),
    .X(_2786_));
 sg13g2_buf_8 _3542_ (.A(_2573_),
    .X(_2787_));
 sg13g2_nand2_1 _3543_ (.Y(_2788_),
    .A(_2786_),
    .B(net41));
 sg13g2_nand2_1 _3544_ (.Y(_2789_),
    .A(_2783_),
    .B(_2788_));
 sg13g2_xnor2_1 _3545_ (.Y(_2790_),
    .A(_2561_),
    .B(_2558_));
 sg13g2_buf_1 _3546_ (.A(_2790_),
    .X(_2791_));
 sg13g2_buf_8 _3547_ (.A(net56),
    .X(_2792_));
 sg13g2_nand2_1 _3548_ (.Y(_2793_),
    .A(_2789_),
    .B(net49));
 sg13g2_nand3_1 _3549_ (.B(_2451_),
    .C(_2453_),
    .A(_2449_),
    .Y(_2794_));
 sg13g2_buf_2 _3550_ (.A(_2794_),
    .X(_2795_));
 sg13g2_nor2_1 _3551_ (.A(_2467_),
    .B(_2795_),
    .Y(_2796_));
 sg13g2_nand2_1 _3552_ (.Y(_2797_),
    .A(_2796_),
    .B(_2440_));
 sg13g2_nand2_1 _3553_ (.Y(_2798_),
    .A(_2797_),
    .B(_2564_));
 sg13g2_nand2_2 _3554_ (.Y(_2799_),
    .A(_2798_),
    .B(net42));
 sg13g2_inv_2 _3555_ (.Y(_2800_),
    .A(_2799_));
 sg13g2_nand2_1 _3556_ (.Y(_2801_),
    .A(_2793_),
    .B(_2800_));
 sg13g2_buf_1 _3557_ (.A(_2772_),
    .X(_2802_));
 sg13g2_nand2_1 _3558_ (.Y(_2803_),
    .A(_2801_),
    .B(net83));
 sg13g2_buf_8 _3559_ (.A(_2796_),
    .X(_2804_));
 sg13g2_a21oi_1 _3560_ (.A1(net31),
    .A2(net46),
    .Y(_2805_),
    .B1(net56));
 sg13g2_nor2_1 _3561_ (.A(_2441_),
    .B(_2786_),
    .Y(_2806_));
 sg13g2_inv_2 _3562_ (.Y(_2807_),
    .A(_2806_));
 sg13g2_nand2_1 _3563_ (.Y(_2808_),
    .A(_2805_),
    .B(_2807_));
 sg13g2_nor2_1 _3564_ (.A(net44),
    .B(_2806_),
    .Y(_2809_));
 sg13g2_inv_2 _3565_ (.Y(_2810_),
    .A(_2809_));
 sg13g2_nand3_1 _3566_ (.B(net32),
    .C(_2810_),
    .A(_2808_),
    .Y(_2811_));
 sg13g2_nor2_1 _3567_ (.A(net111),
    .B(_2306_),
    .Y(_2812_));
 sg13g2_buf_1 _3568_ (.A(_2812_),
    .X(_2813_));
 sg13g2_nand2_1 _3569_ (.Y(_2814_),
    .A(_2811_),
    .B(net90));
 sg13g2_nand2_1 _3570_ (.Y(_2815_),
    .A(_2803_),
    .B(_2814_));
 sg13g2_nand2_2 _3571_ (.Y(_2816_),
    .A(_2454_),
    .B(_2496_));
 sg13g2_nand2_1 _3572_ (.Y(_2817_),
    .A(_2816_),
    .B(net43));
 sg13g2_buf_8 _3573_ (.A(_2496_),
    .X(_2818_));
 sg13g2_nand2_1 _3574_ (.Y(_2819_),
    .A(_2784_),
    .B(net40));
 sg13g2_nand2_2 _3575_ (.Y(_2820_),
    .A(_2819_),
    .B(net52));
 sg13g2_nand2_1 _3576_ (.Y(_2821_),
    .A(_2817_),
    .B(_2820_));
 sg13g2_nand2_2 _3577_ (.Y(_2822_),
    .A(_2795_),
    .B(_2468_));
 sg13g2_nand2_1 _3578_ (.Y(_2823_),
    .A(_2821_),
    .B(_2822_));
 sg13g2_nand2_1 _3579_ (.Y(_2824_),
    .A(net42),
    .B(net56));
 sg13g2_buf_1 _3580_ (.A(_2824_),
    .X(_2825_));
 sg13g2_inv_2 _3581_ (.Y(_2826_),
    .A(net24));
 sg13g2_nand2_1 _3582_ (.Y(_2827_),
    .A(_2823_),
    .B(_2826_));
 sg13g2_nor2_1 _3583_ (.A(_2573_),
    .B(net56),
    .Y(_2828_));
 sg13g2_nand2_2 _3584_ (.Y(_2829_),
    .A(_2828_),
    .B(_2499_));
 sg13g2_inv_2 _3585_ (.Y(_2830_),
    .A(_2829_));
 sg13g2_inv_8 _3586_ (.Y(_2831_),
    .A(net42));
 sg13g2_nand2_1 _3587_ (.Y(_2832_),
    .A(_2830_),
    .B(_2831_));
 sg13g2_nand2_1 _3588_ (.Y(_2833_),
    .A(_2832_),
    .B(_2799_));
 sg13g2_nand2_1 _3589_ (.Y(_2834_),
    .A(_2827_),
    .B(_2833_));
 sg13g2_nor2_1 _3590_ (.A(net111),
    .B(_2345_),
    .Y(_2835_));
 sg13g2_buf_1 _3591_ (.A(_2835_),
    .X(_2836_));
 sg13g2_nand2_1 _3592_ (.Y(_2837_),
    .A(_2834_),
    .B(net89));
 sg13g2_nor2_2 _3593_ (.A(net50),
    .B(net51),
    .Y(_2838_));
 sg13g2_nor2_2 _3594_ (.A(net52),
    .B(_2838_),
    .Y(_2839_));
 sg13g2_nand2_1 _3595_ (.Y(_2840_),
    .A(_2839_),
    .B(_2786_));
 sg13g2_nand2_1 _3596_ (.Y(_2841_),
    .A(_2521_),
    .B(_2496_));
 sg13g2_nand2_1 _3597_ (.Y(_2842_),
    .A(_2841_),
    .B(net46));
 sg13g2_nand2_1 _3598_ (.Y(_2843_),
    .A(_2840_),
    .B(_2842_));
 sg13g2_buf_1 _3599_ (.A(net56),
    .X(_2844_));
 sg13g2_nand2_1 _3600_ (.Y(_2845_),
    .A(_2843_),
    .B(net48));
 sg13g2_nand2_1 _3601_ (.Y(_2846_),
    .A(_2845_),
    .B(_2800_));
 sg13g2_nor2_1 _3602_ (.A(net122),
    .B(net100),
    .Y(_2847_));
 sg13g2_buf_1 _3603_ (.A(_2847_),
    .X(_2848_));
 sg13g2_nand2_1 _3604_ (.Y(_2849_),
    .A(_2846_),
    .B(net82));
 sg13g2_nand2_1 _3605_ (.Y(_2850_),
    .A(_2837_),
    .B(_2849_));
 sg13g2_nor2_1 _3606_ (.A(_2815_),
    .B(_2850_),
    .Y(_2851_));
 sg13g2_nor2_1 _3607_ (.A(_2780_),
    .B(_2851_),
    .Y(_2852_));
 sg13g2_nand2_2 _3608_ (.Y(_2853_),
    .A(_2454_),
    .B(net51));
 sg13g2_a21oi_2 _3609_ (.B1(net56),
    .Y(_2854_),
    .A2(net33),
    .A1(_2853_));
 sg13g2_nand2_1 _3610_ (.Y(_2855_),
    .A(_2468_),
    .B(net50));
 sg13g2_nand3_1 _3611_ (.B(_2855_),
    .C(net43),
    .A(net56),
    .Y(_2856_));
 sg13g2_nand2_1 _3612_ (.Y(_2857_),
    .A(_2856_),
    .B(net42));
 sg13g2_nor2_1 _3613_ (.A(_2854_),
    .B(_2857_),
    .Y(_2858_));
 sg13g2_buf_1 _3614_ (.A(net100),
    .X(_2859_));
 sg13g2_nor2_1 _3615_ (.A(_2812_),
    .B(net83),
    .Y(_2860_));
 sg13g2_buf_2 _3616_ (.A(_2860_),
    .X(_2861_));
 sg13g2_a21oi_1 _3617_ (.A1(_2858_),
    .A2(net88),
    .Y(_2862_),
    .B1(_2861_));
 sg13g2_inv_1 _3618_ (.Y(_2863_),
    .A(net89));
 sg13g2_nor2_1 _3619_ (.A(_2809_),
    .B(_2799_),
    .Y(_2864_));
 sg13g2_nor2_1 _3620_ (.A(_2863_),
    .B(_2864_),
    .Y(_2865_));
 sg13g2_inv_1 _3621_ (.Y(_2866_),
    .A(_2847_));
 sg13g2_nor2_1 _3622_ (.A(net52),
    .B(_2853_),
    .Y(_2867_));
 sg13g2_nand2_1 _3623_ (.Y(_2868_),
    .A(_2867_),
    .B(_2591_));
 sg13g2_nor2_2 _3624_ (.A(net40),
    .B(_2521_),
    .Y(_2869_));
 sg13g2_a21oi_2 _3625_ (.B1(_2565_),
    .Y(_2870_),
    .A2(net41),
    .A1(_2869_));
 sg13g2_a21oi_1 _3626_ (.A1(_2868_),
    .A2(net24),
    .Y(_2871_),
    .B1(_2870_));
 sg13g2_nor2_1 _3627_ (.A(_2866_),
    .B(_2871_),
    .Y(_2872_));
 sg13g2_nor2_1 _3628_ (.A(_2865_),
    .B(_2872_),
    .Y(_2873_));
 sg13g2_nand2b_1 _3629_ (.Y(_2874_),
    .B(_2873_),
    .A_N(_2862_));
 sg13g2_nor2_1 _3630_ (.A(_2770_),
    .B(_2777_),
    .Y(_2875_));
 sg13g2_buf_1 _3631_ (.A(_2875_),
    .X(_2876_));
 sg13g2_nand2_1 _3632_ (.Y(_2877_),
    .A(_2874_),
    .B(net55));
 sg13g2_nor2b_1 _3633_ (.A(_2852_),
    .B_N(_2877_),
    .Y(_2878_));
 sg13g2_buf_8 _3634_ (.A(_2831_),
    .X(_2879_));
 sg13g2_buf_8 _3635_ (.A(net23),
    .X(_2880_));
 sg13g2_nor2_1 _3636_ (.A(net49),
    .B(_2804_),
    .Y(_2881_));
 sg13g2_nor2_1 _3637_ (.A(net18),
    .B(_2881_),
    .Y(_2882_));
 sg13g2_nor2_2 _3638_ (.A(_2591_),
    .B(_2829_),
    .Y(_2883_));
 sg13g2_a21oi_1 _3639_ (.A1(_2822_),
    .A2(_2882_),
    .Y(_2884_),
    .B1(_2883_));
 sg13g2_buf_1 _3640_ (.A(net83),
    .X(_2885_));
 sg13g2_buf_1 _3641_ (.A(net90),
    .X(_2886_));
 sg13g2_nor2_1 _3642_ (.A(_2574_),
    .B(_2822_),
    .Y(_2887_));
 sg13g2_inv_1 _3643_ (.Y(_2888_),
    .A(_2887_));
 sg13g2_nor2_1 _3644_ (.A(_2566_),
    .B(_2888_),
    .Y(_2889_));
 sg13g2_nand2_1 _3645_ (.Y(_2890_),
    .A(_2889_),
    .B(net32));
 sg13g2_nand2_1 _3646_ (.Y(_2891_),
    .A(_2833_),
    .B(_2890_));
 sg13g2_a22oi_1 _3647_ (.Y(_2892_),
    .B1(net81),
    .B2(_2891_),
    .A2(net75),
    .A1(_2884_));
 sg13g2_nand2_2 _3648_ (.Y(_2893_),
    .A(net42),
    .B(_2564_));
 sg13g2_inv_2 _3649_ (.Y(_2894_),
    .A(_2893_));
 sg13g2_nand2_1 _3650_ (.Y(_2895_),
    .A(_2821_),
    .B(_2894_));
 sg13g2_nand2_1 _3651_ (.Y(_2896_),
    .A(_2829_),
    .B(_2831_));
 sg13g2_buf_2 _3652_ (.A(_2896_),
    .X(_2897_));
 sg13g2_nand3_1 _3653_ (.B(_2895_),
    .C(_2897_),
    .A(_2890_),
    .Y(_2898_));
 sg13g2_nand2_1 _3654_ (.Y(_2899_),
    .A(_2898_),
    .B(net82));
 sg13g2_xnor2_1 _3655_ (.Y(_2900_),
    .A(_2421_),
    .B(_2448_));
 sg13g2_nor2_1 _3656_ (.A(net65),
    .B(_2900_),
    .Y(_2901_));
 sg13g2_nand2_1 _3657_ (.Y(_2902_),
    .A(_2901_),
    .B(net51));
 sg13g2_nor3_2 _3658_ (.A(net41),
    .B(net44),
    .C(_2902_),
    .Y(_2903_));
 sg13g2_nand2_1 _3659_ (.Y(_2904_),
    .A(_2498_),
    .B(net40));
 sg13g2_nor2_1 _3660_ (.A(net41),
    .B(_2904_),
    .Y(_2905_));
 sg13g2_nor2_2 _3661_ (.A(net49),
    .B(_2905_),
    .Y(_2906_));
 sg13g2_inv_1 _3662_ (.Y(_2907_),
    .A(_2906_));
 sg13g2_nand2_1 _3663_ (.Y(_2908_),
    .A(_2907_),
    .B(net25));
 sg13g2_buf_1 _3664_ (.A(_2863_),
    .X(_2909_));
 sg13g2_nor2_1 _3665_ (.A(_2900_),
    .B(_2496_),
    .Y(_2910_));
 sg13g2_buf_8 _3666_ (.A(_2910_),
    .X(_2911_));
 sg13g2_nand2_1 _3667_ (.Y(_2912_),
    .A(_2911_),
    .B(net52));
 sg13g2_nor3_1 _3668_ (.A(net49),
    .B(net32),
    .C(_2912_),
    .Y(_2913_));
 sg13g2_nor2_1 _3669_ (.A(net74),
    .B(_2913_),
    .Y(_2914_));
 sg13g2_o21ai_1 _3670_ (.B1(_2914_),
    .Y(_2915_),
    .A1(_2903_),
    .A2(_2908_));
 sg13g2_nand3_1 _3671_ (.B(_2899_),
    .C(_2915_),
    .A(_2892_),
    .Y(_2916_));
 sg13g2_inv_1 _3672_ (.Y(_2917_),
    .A(_2777_));
 sg13g2_nor2_1 _3673_ (.A(_2770_),
    .B(_2917_),
    .Y(_2918_));
 sg13g2_buf_2 _3674_ (.A(_2918_),
    .X(_2919_));
 sg13g2_nand2_1 _3675_ (.Y(_2920_),
    .A(_2916_),
    .B(_2919_));
 sg13g2_nor2_2 _3676_ (.A(_2771_),
    .B(_2917_),
    .Y(_2921_));
 sg13g2_inv_1 _3677_ (.Y(_2922_),
    .A(_2921_));
 sg13g2_nor2_1 _3678_ (.A(net44),
    .B(_2912_),
    .Y(_2923_));
 sg13g2_nor2_2 _3679_ (.A(net23),
    .B(_2923_),
    .Y(_2924_));
 sg13g2_inv_4 _3680_ (.A(_2924_),
    .Y(_2925_));
 sg13g2_inv_1 _3681_ (.Y(_2926_),
    .A(_2869_));
 sg13g2_nand2_1 _3682_ (.Y(_2927_),
    .A(_2926_),
    .B(_2576_));
 sg13g2_a21oi_1 _3683_ (.A1(_2888_),
    .A2(_2927_),
    .Y(_2928_),
    .B1(net48));
 sg13g2_nor2_1 _3684_ (.A(net88),
    .B(_2913_),
    .Y(_2929_));
 sg13g2_o21ai_1 _3685_ (.B1(_2929_),
    .Y(_2930_),
    .A1(_2925_),
    .A2(_2928_));
 sg13g2_inv_1 _3686_ (.Y(_2931_),
    .A(_2861_));
 sg13g2_buf_1 _3687_ (.A(_2931_),
    .X(_2932_));
 sg13g2_nand2_1 _3688_ (.Y(_2933_),
    .A(_2930_),
    .B(net61));
 sg13g2_nor2_1 _3689_ (.A(net52),
    .B(_2564_),
    .Y(_2934_));
 sg13g2_inv_2 _3690_ (.Y(_2935_),
    .A(_2934_));
 sg13g2_nor2_1 _3691_ (.A(net43),
    .B(_2911_),
    .Y(_2936_));
 sg13g2_inv_1 _3692_ (.Y(_2937_),
    .A(_2936_));
 sg13g2_nand3_1 _3693_ (.B(_2937_),
    .C(_2592_),
    .A(_2935_),
    .Y(_2938_));
 sg13g2_o21ai_1 _3694_ (.B1(_2879_),
    .Y(_2939_),
    .A1(net48),
    .A2(_2912_));
 sg13g2_nand2_1 _3695_ (.Y(_2940_),
    .A(_2938_),
    .B(_2939_));
 sg13g2_buf_1 _3696_ (.A(_2345_),
    .X(_2941_));
 sg13g2_nand2_1 _3697_ (.Y(_2942_),
    .A(_2940_),
    .B(net93));
 sg13g2_nor2b_1 _3698_ (.A(_2933_),
    .B_N(_2942_),
    .Y(_2943_));
 sg13g2_nor2_1 _3699_ (.A(_2922_),
    .B(_2943_),
    .Y(_2944_));
 sg13g2_nand3_1 _3700_ (.B(net43),
    .C(_2791_),
    .A(net31),
    .Y(_2945_));
 sg13g2_buf_1 _3701_ (.A(_2945_),
    .X(_2946_));
 sg13g2_nor2_1 _3702_ (.A(_2573_),
    .B(_2564_),
    .Y(_2947_));
 sg13g2_buf_1 _3703_ (.A(_2947_),
    .X(_2948_));
 sg13g2_nand2_1 _3704_ (.Y(_2949_),
    .A(net30),
    .B(net50));
 sg13g2_nand2_1 _3705_ (.Y(_2950_),
    .A(_2946_),
    .B(_2949_));
 sg13g2_nor2_1 _3706_ (.A(_2787_),
    .B(_2902_),
    .Y(_2951_));
 sg13g2_a21oi_1 _3707_ (.A1(_2951_),
    .A2(net34),
    .Y(_2952_),
    .B1(_2592_));
 sg13g2_a21oi_1 _3708_ (.A1(net32),
    .A2(_2950_),
    .Y(_2953_),
    .B1(_2952_));
 sg13g2_nor2_1 _3709_ (.A(_2787_),
    .B(_2499_),
    .Y(_2954_));
 sg13g2_nand3_1 _3710_ (.B(_2795_),
    .C(net40),
    .A(_2498_),
    .Y(_2955_));
 sg13g2_buf_1 _3711_ (.A(_2955_),
    .X(_2956_));
 sg13g2_nand2_1 _3712_ (.Y(_2957_),
    .A(_2954_),
    .B(_2956_));
 sg13g2_nand3_1 _3713_ (.B(_2894_),
    .C(_2807_),
    .A(_2957_),
    .Y(_2958_));
 sg13g2_a21oi_1 _3714_ (.A1(_2953_),
    .A2(_2958_),
    .Y(_2959_),
    .B1(net93));
 sg13g2_nor2_1 _3715_ (.A(_2453_),
    .B(_2476_),
    .Y(_2960_));
 sg13g2_nand2_2 _3716_ (.Y(_2961_),
    .A(_2960_),
    .B(_2818_));
 sg13g2_nor2_1 _3717_ (.A(net46),
    .B(_2961_),
    .Y(_2962_));
 sg13g2_nor2_1 _3718_ (.A(net23),
    .B(_2962_),
    .Y(_0188_));
 sg13g2_inv_1 _3719_ (.Y(_0189_),
    .A(_2954_));
 sg13g2_nand3_1 _3720_ (.B(_2567_),
    .C(_0189_),
    .A(_0188_),
    .Y(_0190_));
 sg13g2_nand3_1 _3721_ (.B(_2861_),
    .C(_0190_),
    .A(_2953_),
    .Y(_0191_));
 sg13g2_nand2_1 _3722_ (.Y(_0192_),
    .A(_0191_),
    .B(_2909_));
 sg13g2_nand2b_1 _3723_ (.Y(_0193_),
    .B(_0192_),
    .A_N(_2959_));
 sg13g2_nand2_1 _3724_ (.Y(_0194_),
    .A(_2944_),
    .B(_0193_));
 sg13g2_nand3_1 _3725_ (.B(_2920_),
    .C(_0194_),
    .A(_2878_),
    .Y(_0195_));
 sg13g2_nand3_1 _3726_ (.B(net105),
    .C(_2715_),
    .A(net94),
    .Y(_0196_));
 sg13g2_xnor2_1 _3727_ (.Y(_0197_),
    .A(_2667_),
    .B(_0196_));
 sg13g2_inv_2 _3728_ (.Y(_0198_),
    .A(_0197_));
 sg13g2_nand2_1 _3729_ (.Y(_0199_),
    .A(_0195_),
    .B(_0198_));
 sg13g2_buf_1 _3730_ (.A(_0009_),
    .X(_0200_));
 sg13g2_nand2_1 _3731_ (.Y(_0201_),
    .A(net57),
    .B(_2931_));
 sg13g2_a21oi_1 _3732_ (.A1(_2522_),
    .A2(net45),
    .Y(_0202_),
    .B1(net46));
 sg13g2_inv_1 _3733_ (.Y(_0203_),
    .A(_0202_));
 sg13g2_a21oi_1 _3734_ (.A1(_2838_),
    .A2(net28),
    .Y(_0204_),
    .B1(net27));
 sg13g2_o21ai_1 _3735_ (.B1(_0204_),
    .Y(_0205_),
    .A1(_2838_),
    .A2(_0203_));
 sg13g2_nand2_2 _3736_ (.Y(_0206_),
    .A(_2498_),
    .B(net51));
 sg13g2_nand2_1 _3737_ (.Y(_0207_),
    .A(_0206_),
    .B(net33));
 sg13g2_nand2_1 _3738_ (.Y(_0208_),
    .A(_2838_),
    .B(_2441_));
 sg13g2_nand2_2 _3739_ (.Y(_0209_),
    .A(_0208_),
    .B(net44));
 sg13g2_inv_1 _3740_ (.Y(_0210_),
    .A(_0209_));
 sg13g2_o21ai_1 _3741_ (.B1(_0210_),
    .Y(_0211_),
    .A1(net31),
    .A2(_0207_));
 sg13g2_nand3_1 _3742_ (.B(net19),
    .C(_0211_),
    .A(_0205_),
    .Y(_0212_));
 sg13g2_nor3_1 _3743_ (.A(_0200_),
    .B(_0201_),
    .C(_0212_),
    .Y(_0213_));
 sg13g2_nand3_1 _3744_ (.B(_2494_),
    .C(net65),
    .A(_2493_),
    .Y(_0214_));
 sg13g2_nand2_1 _3745_ (.Y(_0215_),
    .A(_2573_),
    .B(_0214_));
 sg13g2_nor2_1 _3746_ (.A(_2838_),
    .B(_2911_),
    .Y(_0216_));
 sg13g2_nand2_1 _3747_ (.Y(_0217_),
    .A(_2904_),
    .B(net35));
 sg13g2_o21ai_1 _3748_ (.B1(_0217_),
    .Y(_0218_),
    .A1(_0215_),
    .A2(_0216_));
 sg13g2_nor2_1 _3749_ (.A(net31),
    .B(_2869_),
    .Y(_0219_));
 sg13g2_inv_1 _3750_ (.Y(_0220_),
    .A(_0219_));
 sg13g2_nand2_1 _3751_ (.Y(_0221_),
    .A(_2496_),
    .B(_2900_));
 sg13g2_nand2_1 _3752_ (.Y(_0222_),
    .A(_0221_),
    .B(net35));
 sg13g2_inv_1 _3753_ (.Y(_0223_),
    .A(_0222_));
 sg13g2_a21oi_1 _3754_ (.A1(_0220_),
    .A2(net20),
    .Y(_0224_),
    .B1(_0223_));
 sg13g2_nand2_1 _3755_ (.Y(_0225_),
    .A(_0224_),
    .B(_2894_));
 sg13g2_o21ai_1 _3756_ (.B1(_0225_),
    .Y(_0226_),
    .A1(net24),
    .A2(_0218_));
 sg13g2_buf_1 _3757_ (.A(_2836_),
    .X(_0227_));
 sg13g2_buf_1 _3758_ (.A(net80),
    .X(_0228_));
 sg13g2_nand2b_1 _3759_ (.Y(_0229_),
    .B(net73),
    .A_N(_0226_));
 sg13g2_nand3_1 _3760_ (.B(net32),
    .C(_2820_),
    .A(_2854_),
    .Y(_0230_));
 sg13g2_nand2_1 _3761_ (.Y(_0231_),
    .A(_0230_),
    .B(net90));
 sg13g2_nand2_1 _3762_ (.Y(_0232_),
    .A(_0231_),
    .B(net55));
 sg13g2_nor2_1 _3763_ (.A(net40),
    .B(net26),
    .Y(_0233_));
 sg13g2_nor2_1 _3764_ (.A(_0233_),
    .B(net24),
    .Y(_0234_));
 sg13g2_nand2_1 _3765_ (.Y(_0235_),
    .A(_0234_),
    .B(net55));
 sg13g2_nand2_1 _3766_ (.Y(_0236_),
    .A(_0232_),
    .B(_0235_));
 sg13g2_inv_1 _3767_ (.Y(_0237_),
    .A(_2946_));
 sg13g2_buf_8 _3768_ (.A(net49),
    .X(_0238_));
 sg13g2_buf_8 _3769_ (.A(net39),
    .X(_0239_));
 sg13g2_o21ai_1 _3770_ (.B1(net25),
    .Y(_0240_),
    .A1(net29),
    .A2(_0222_));
 sg13g2_buf_1 _3771_ (.A(net82),
    .X(_0241_));
 sg13g2_o21ai_1 _3772_ (.B1(net72),
    .Y(_0242_),
    .A1(_0237_),
    .A2(_0240_));
 sg13g2_a21oi_1 _3773_ (.A1(_2888_),
    .A2(_2844_),
    .Y(_0243_),
    .B1(_2879_));
 sg13g2_nand2_1 _3774_ (.Y(_0244_),
    .A(net45),
    .B(_2900_));
 sg13g2_nand2_1 _3775_ (.Y(_0245_),
    .A(_0244_),
    .B(_2795_));
 sg13g2_nand2_1 _3776_ (.Y(_0246_),
    .A(_2828_),
    .B(_0245_));
 sg13g2_nand2_1 _3777_ (.Y(_0247_),
    .A(_0243_),
    .B(_0246_));
 sg13g2_buf_1 _3778_ (.A(net94),
    .X(_0248_));
 sg13g2_a21o_1 _3779_ (.A2(_2897_),
    .A1(_0247_),
    .B1(net87),
    .X(_0249_));
 sg13g2_nand4_1 _3780_ (.B(_0236_),
    .C(_0242_),
    .A(_0229_),
    .Y(_0250_),
    .D(_0249_));
 sg13g2_buf_1 _3781_ (.A(_0197_),
    .X(_0251_));
 sg13g2_nand3b_1 _3782_ (.B(_0250_),
    .C(net71),
    .Y(_0252_),
    .A_N(_0213_));
 sg13g2_buf_1 _3783_ (.A(_2481_),
    .X(_0253_));
 sg13g2_nand2_1 _3784_ (.Y(_0254_),
    .A(net102),
    .B(_2346_));
 sg13g2_a21oi_1 _3785_ (.A1(_0199_),
    .A2(_0252_),
    .Y(_0255_),
    .B1(_0254_));
 sg13g2_nand2_1 _3786_ (.Y(_0256_),
    .A(_2801_),
    .B(_2836_));
 sg13g2_inv_1 _3787_ (.Y(_0257_),
    .A(_2871_));
 sg13g2_nand2_1 _3788_ (.Y(_0258_),
    .A(_0257_),
    .B(net90));
 sg13g2_o21ai_1 _3789_ (.B1(net105),
    .Y(_0259_),
    .A1(_2854_),
    .A2(_2857_));
 sg13g2_nand3_1 _3790_ (.B(_0258_),
    .C(_0259_),
    .A(_0256_),
    .Y(_0260_));
 sg13g2_nand2_1 _3791_ (.Y(_0261_),
    .A(_0260_),
    .B(net55));
 sg13g2_inv_1 _3792_ (.Y(_0262_),
    .A(_2864_));
 sg13g2_buf_1 _3793_ (.A(_2866_),
    .X(_0263_));
 sg13g2_inv_2 _3794_ (.Y(_0264_),
    .A(_2876_));
 sg13g2_nor2_1 _3795_ (.A(net70),
    .B(_0264_),
    .Y(_0265_));
 sg13g2_a21oi_1 _3796_ (.A1(_0262_),
    .A2(_0265_),
    .Y(_0266_),
    .B1(net71));
 sg13g2_nand2_1 _3797_ (.Y(_0267_),
    .A(_0261_),
    .B(_0266_));
 sg13g2_inv_1 _3798_ (.Y(_0268_),
    .A(_2919_));
 sg13g2_nand3_1 _3799_ (.B(_2926_),
    .C(net27),
    .A(_2937_),
    .Y(_0269_));
 sg13g2_nor2_1 _3800_ (.A(net111),
    .B(_2923_),
    .Y(_0270_));
 sg13g2_buf_1 _3801_ (.A(net18),
    .X(_0271_));
 sg13g2_a21oi_1 _3802_ (.A1(_0269_),
    .A2(_0270_),
    .Y(_0272_),
    .B1(net16));
 sg13g2_buf_8 _3803_ (.A(net34),
    .X(_0273_));
 sg13g2_nand2_1 _3804_ (.Y(_0274_),
    .A(_0189_),
    .B(net22));
 sg13g2_nand2_2 _3805_ (.Y(_0275_),
    .A(_2951_),
    .B(net49));
 sg13g2_buf_1 _3806_ (.A(net111),
    .X(_0276_));
 sg13g2_buf_1 _3807_ (.A(net92),
    .X(_0277_));
 sg13g2_nand3_1 _3808_ (.B(_0275_),
    .C(net86),
    .A(_0274_),
    .Y(_0278_));
 sg13g2_buf_1 _3809_ (.A(_2861_),
    .X(_0279_));
 sg13g2_nand2_1 _3810_ (.Y(_0280_),
    .A(_2939_),
    .B(net63));
 sg13g2_a21oi_1 _3811_ (.A1(_0272_),
    .A2(_0278_),
    .Y(_0281_),
    .B1(_0280_));
 sg13g2_nand2_1 _3812_ (.Y(_0282_),
    .A(_2956_),
    .B(_2853_));
 sg13g2_nand2_1 _3813_ (.Y(_0283_),
    .A(_0282_),
    .B(_2444_));
 sg13g2_inv_1 _3814_ (.Y(_0284_),
    .A(_2817_));
 sg13g2_nor2_1 _3815_ (.A(net39),
    .B(_0284_),
    .Y(_0285_));
 sg13g2_nand2_1 _3816_ (.Y(_0286_),
    .A(_0283_),
    .B(_0285_));
 sg13g2_nand2_1 _3817_ (.Y(_0287_),
    .A(_0286_),
    .B(_0243_));
 sg13g2_nand2_1 _3818_ (.Y(_0288_),
    .A(_0287_),
    .B(net90));
 sg13g2_nand2_1 _3819_ (.Y(_0289_),
    .A(_0247_),
    .B(net83));
 sg13g2_inv_4 _3820_ (.A(_2897_),
    .Y(_0290_));
 sg13g2_a21oi_1 _3821_ (.A1(_0288_),
    .A2(_0289_),
    .Y(_0291_),
    .B1(_0290_));
 sg13g2_nor3_1 _3822_ (.A(_0268_),
    .B(_0281_),
    .C(_0291_),
    .Y(_0292_));
 sg13g2_nor2_1 _3823_ (.A(_0267_),
    .B(_0292_),
    .Y(_0293_));
 sg13g2_nand2_1 _3824_ (.Y(_0294_),
    .A(_2961_),
    .B(net26));
 sg13g2_nand2_1 _3825_ (.Y(_0295_),
    .A(net34),
    .B(net100));
 sg13g2_a21oi_1 _3826_ (.A1(_0294_),
    .A2(_0217_),
    .Y(_0296_),
    .B1(_0295_));
 sg13g2_nor2_1 _3827_ (.A(_2950_),
    .B(_0296_),
    .Y(_0297_));
 sg13g2_nor2_1 _3828_ (.A(_2806_),
    .B(_2798_),
    .Y(_0298_));
 sg13g2_nand2_1 _3829_ (.Y(_0299_),
    .A(_0298_),
    .B(net92));
 sg13g2_a21oi_1 _3830_ (.A1(_0297_),
    .A2(_0299_),
    .Y(_0300_),
    .B1(net16));
 sg13g2_o21ai_1 _3831_ (.B1(net93),
    .Y(_0301_),
    .A1(_2952_),
    .A2(_0300_));
 sg13g2_inv_1 _3832_ (.Y(_0302_),
    .A(_0214_));
 sg13g2_a21oi_1 _3833_ (.A1(_0302_),
    .A2(_2894_),
    .Y(_0303_),
    .B1(_2940_));
 sg13g2_nor2_1 _3834_ (.A(net87),
    .B(_0303_),
    .Y(_0304_));
 sg13g2_a21oi_1 _3835_ (.A1(_2891_),
    .A2(net73),
    .Y(_0305_),
    .B1(_0304_));
 sg13g2_nand2_1 _3836_ (.Y(_0306_),
    .A(_0301_),
    .B(_0305_));
 sg13g2_nand2_1 _3837_ (.Y(_0307_),
    .A(_0306_),
    .B(_2921_));
 sg13g2_a22oi_1 _3838_ (.Y(_0308_),
    .B1(net81),
    .B2(_2846_),
    .A2(net80),
    .A1(_2884_));
 sg13g2_nand2_1 _3839_ (.Y(_0309_),
    .A(_2834_),
    .B(_0241_));
 sg13g2_nand2_1 _3840_ (.Y(_0310_),
    .A(_2811_),
    .B(net75));
 sg13g2_nand3_1 _3841_ (.B(_0309_),
    .C(_0310_),
    .A(_0308_),
    .Y(_0311_));
 sg13g2_nand2_1 _3842_ (.Y(_0312_),
    .A(_0311_),
    .B(net57));
 sg13g2_nand3_1 _3843_ (.B(_0307_),
    .C(_0312_),
    .A(_0293_),
    .Y(_0313_));
 sg13g2_nor2_1 _3844_ (.A(net70),
    .B(_0226_),
    .Y(_0314_));
 sg13g2_inv_1 _3845_ (.Y(_0315_),
    .A(_0230_));
 sg13g2_nor3_1 _3846_ (.A(net87),
    .B(_0234_),
    .C(_0315_),
    .Y(_0316_));
 sg13g2_o21ai_1 _3847_ (.B1(net81),
    .Y(_0317_),
    .A1(_0237_),
    .A2(_0240_));
 sg13g2_nand3_1 _3848_ (.B(net71),
    .C(net55),
    .A(_0317_),
    .Y(_0318_));
 sg13g2_nor2b_1 _3849_ (.A(net74),
    .B_N(_0212_),
    .Y(_0319_));
 sg13g2_nor4_1 _3850_ (.A(_0314_),
    .B(_0316_),
    .C(_0318_),
    .D(_0319_),
    .Y(_0320_));
 sg13g2_nor2_1 _3851_ (.A(_2484_),
    .B(_0320_),
    .Y(_0321_));
 sg13g2_nand2_1 _3852_ (.Y(_0322_),
    .A(_0313_),
    .B(_0321_));
 sg13g2_nand3_1 _3853_ (.B(net46),
    .C(_2816_),
    .A(_2782_),
    .Y(_0323_));
 sg13g2_nor2_1 _3854_ (.A(_2565_),
    .B(_2839_),
    .Y(_0324_));
 sg13g2_nand2_1 _3855_ (.Y(_0325_),
    .A(_0323_),
    .B(_0324_));
 sg13g2_buf_1 _3856_ (.A(net88),
    .X(_0326_));
 sg13g2_inv_1 _3857_ (.Y(_0327_),
    .A(_2962_));
 sg13g2_nand2_1 _3858_ (.Y(_0328_),
    .A(_0210_),
    .B(_0327_));
 sg13g2_nand3_1 _3859_ (.B(net79),
    .C(_0328_),
    .A(_0325_),
    .Y(_0329_));
 sg13g2_nand2_1 _3860_ (.Y(_0330_),
    .A(_2499_),
    .B(_2442_));
 sg13g2_inv_1 _3861_ (.Y(_0331_),
    .A(_0330_));
 sg13g2_nor2_1 _3862_ (.A(_2859_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_o21ai_1 _3863_ (.B1(net27),
    .Y(_0333_),
    .A1(net45),
    .A2(net26));
 sg13g2_a21oi_1 _3864_ (.A1(_0332_),
    .A2(_0333_),
    .Y(_0334_),
    .B1(net18));
 sg13g2_nand2_1 _3865_ (.Y(_0335_),
    .A(_0329_),
    .B(_0334_));
 sg13g2_nand2_1 _3866_ (.Y(_0336_),
    .A(_0335_),
    .B(_2897_));
 sg13g2_nand2_1 _3867_ (.Y(_0337_),
    .A(_0336_),
    .B(net61));
 sg13g2_o21ai_1 _3868_ (.B1(net80),
    .Y(_0338_),
    .A1(_2923_),
    .A2(_2799_));
 sg13g2_buf_1 _3869_ (.A(_2770_),
    .X(_0339_));
 sg13g2_nand2_1 _3870_ (.Y(_0340_),
    .A(_0338_),
    .B(net78));
 sg13g2_nor2_2 _3871_ (.A(_2866_),
    .B(_2883_),
    .Y(_0341_));
 sg13g2_inv_2 _3872_ (.Y(_0342_),
    .A(_0341_));
 sg13g2_inv_1 _3873_ (.Y(_0343_),
    .A(_0325_));
 sg13g2_nor2_1 _3874_ (.A(_2880_),
    .B(_0298_),
    .Y(_0344_));
 sg13g2_nor2b_1 _3875_ (.A(_0343_),
    .B_N(_0344_),
    .Y(_0345_));
 sg13g2_nor2_1 _3876_ (.A(_0342_),
    .B(_0345_),
    .Y(_0346_));
 sg13g2_nor2_1 _3877_ (.A(_0340_),
    .B(_0346_),
    .Y(_0347_));
 sg13g2_nand2_1 _3878_ (.Y(_0348_),
    .A(_0337_),
    .B(_0347_));
 sg13g2_inv_1 _3879_ (.Y(_0349_),
    .A(_2961_));
 sg13g2_nand2_1 _3880_ (.Y(_0350_),
    .A(_0349_),
    .B(net21));
 sg13g2_nand3_1 _3881_ (.B(_0274_),
    .C(_0350_),
    .A(_2924_),
    .Y(_0351_));
 sg13g2_inv_1 _3882_ (.Y(_0352_),
    .A(_2816_));
 sg13g2_nand2_1 _3883_ (.Y(_0353_),
    .A(_2564_),
    .B(net43));
 sg13g2_nor2_1 _3884_ (.A(_0352_),
    .B(_0353_),
    .Y(_0354_));
 sg13g2_nor2_1 _3885_ (.A(_0354_),
    .B(_2925_),
    .Y(_0355_));
 sg13g2_nand2_1 _3886_ (.Y(_0356_),
    .A(_0355_),
    .B(_2829_));
 sg13g2_a22oi_1 _3887_ (.Y(_0357_),
    .B1(net81),
    .B2(_0356_),
    .A2(_2885_),
    .A1(_0351_));
 sg13g2_a21oi_1 _3888_ (.A1(net30),
    .A2(_2499_),
    .Y(_0358_),
    .B1(_2880_));
 sg13g2_nor2b_1 _3889_ (.A(_2928_),
    .B_N(_0358_),
    .Y(_0359_));
 sg13g2_nor2_2 _3890_ (.A(_2863_),
    .B(_2883_),
    .Y(_0360_));
 sg13g2_nand2b_1 _3891_ (.Y(_0361_),
    .B(_0360_),
    .A_N(_0359_));
 sg13g2_o21ai_1 _3892_ (.B1(_2897_),
    .Y(_0362_),
    .A1(_2893_),
    .A2(_2936_));
 sg13g2_a21oi_1 _3893_ (.A1(_0362_),
    .A2(net82),
    .Y(_0363_),
    .B1(net78));
 sg13g2_nand3_1 _3894_ (.B(_0361_),
    .C(_0363_),
    .A(_0357_),
    .Y(_0364_));
 sg13g2_nand3_1 _3895_ (.B(_0364_),
    .C(_2777_),
    .A(_0348_),
    .Y(_0365_));
 sg13g2_inv_1 _3896_ (.Y(_0366_),
    .A(_2822_));
 sg13g2_nand2_1 _3897_ (.Y(_0367_),
    .A(_2937_),
    .B(_0366_));
 sg13g2_a21oi_1 _3898_ (.A1(_0367_),
    .A2(_0208_),
    .Y(_0368_),
    .B1(_2567_));
 sg13g2_nor2_1 _3899_ (.A(_2799_),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_a21oi_1 _3900_ (.A1(_0369_),
    .A2(net86),
    .Y(_0370_),
    .B1(_2932_));
 sg13g2_nand2_1 _3901_ (.Y(_0371_),
    .A(net25),
    .B(net88));
 sg13g2_nand2_1 _3902_ (.Y(_0372_),
    .A(_2957_),
    .B(net27));
 sg13g2_nand2_1 _3903_ (.Y(_0373_),
    .A(net31),
    .B(net26));
 sg13g2_nor2b_1 _3904_ (.A(_0372_),
    .B_N(_0373_),
    .Y(_0374_));
 sg13g2_nor2_1 _3905_ (.A(_0371_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nand2_1 _3906_ (.Y(_0376_),
    .A(_0367_),
    .B(_2797_));
 sg13g2_nand2_1 _3907_ (.Y(_0377_),
    .A(_0376_),
    .B(_0238_));
 sg13g2_nand2_1 _3908_ (.Y(_0378_),
    .A(_0375_),
    .B(_0377_));
 sg13g2_nand2_1 _3909_ (.Y(_0379_),
    .A(_0370_),
    .B(_0378_));
 sg13g2_nand2_1 _3910_ (.Y(_0380_),
    .A(_2498_),
    .B(_2795_));
 sg13g2_nor2_2 _3911_ (.A(net45),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_nand2_1 _3912_ (.Y(_0382_),
    .A(_0381_),
    .B(net33));
 sg13g2_nand3_1 _3913_ (.B(net28),
    .C(_2855_),
    .A(_0380_),
    .Y(_0383_));
 sg13g2_nand3_1 _3914_ (.B(_0382_),
    .C(_0383_),
    .A(_2809_),
    .Y(_0384_));
 sg13g2_nand2_1 _3915_ (.Y(_0385_),
    .A(_0384_),
    .B(_2800_));
 sg13g2_a22oi_1 _3916_ (.Y(_0386_),
    .B1(net81),
    .B2(_0385_),
    .A2(_2623_),
    .A1(_2811_));
 sg13g2_a21oi_1 _3917_ (.A1(_0379_),
    .A2(_0386_),
    .Y(_0387_),
    .B1(_2780_));
 sg13g2_nor2_1 _3918_ (.A(_0267_),
    .B(_0387_),
    .Y(_0388_));
 sg13g2_nand2_1 _3919_ (.Y(_0389_),
    .A(_0365_),
    .B(_0388_));
 sg13g2_nor2_1 _3920_ (.A(_0264_),
    .B(_0271_),
    .Y(_0390_));
 sg13g2_nand2_1 _3921_ (.Y(_0391_),
    .A(_0390_),
    .B(net71));
 sg13g2_inv_2 _3922_ (.Y(_0392_),
    .A(_2812_));
 sg13g2_buf_1 _3923_ (.A(_0392_),
    .X(_0393_));
 sg13g2_nor2_1 _3924_ (.A(net52),
    .B(_0221_),
    .Y(_0394_));
 sg13g2_nor2_1 _3925_ (.A(net44),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_inv_1 _3926_ (.Y(_0396_),
    .A(_0217_));
 sg13g2_nor2_1 _3927_ (.A(net29),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_nor3_1 _3928_ (.A(net77),
    .B(_0395_),
    .C(_0397_),
    .Y(_0398_));
 sg13g2_nor2_1 _3929_ (.A(_2900_),
    .B(net51),
    .Y(_0399_));
 sg13g2_inv_1 _3930_ (.Y(_0400_),
    .A(_0399_));
 sg13g2_nand4_1 _3931_ (.B(net20),
    .C(_0400_),
    .A(_2782_),
    .Y(_0401_),
    .D(net17));
 sg13g2_nor2_1 _3932_ (.A(_2476_),
    .B(_2496_),
    .Y(_0402_));
 sg13g2_nor2_1 _3933_ (.A(net28),
    .B(_0402_),
    .Y(_0403_));
 sg13g2_a21oi_1 _3934_ (.A1(net29),
    .A2(_0403_),
    .Y(_0404_),
    .B1(_0396_));
 sg13g2_a21oi_1 _3935_ (.A1(_0401_),
    .A2(_0404_),
    .Y(_0405_),
    .B1(net74));
 sg13g2_nand2_1 _3936_ (.Y(_0406_),
    .A(_0284_),
    .B(_0206_));
 sg13g2_nor2_1 _3937_ (.A(net21),
    .B(_0233_),
    .Y(_0407_));
 sg13g2_nand2_1 _3938_ (.Y(_0408_),
    .A(_0220_),
    .B(net20));
 sg13g2_a221oi_1 _3939_ (.B2(_0397_),
    .C1(net70),
    .B1(_0408_),
    .A1(_0406_),
    .Y(_0409_),
    .A2(_0407_));
 sg13g2_nor4_1 _3940_ (.A(_0391_),
    .B(_0398_),
    .C(_0405_),
    .D(_0409_),
    .Y(_0410_));
 sg13g2_nand2_1 _3941_ (.Y(_0411_),
    .A(_2499_),
    .B(_2574_));
 sg13g2_nand2_1 _3942_ (.Y(_0412_),
    .A(_0411_),
    .B(_0208_));
 sg13g2_nor2_1 _3943_ (.A(_0237_),
    .B(_2889_),
    .Y(_0413_));
 sg13g2_o21ai_1 _3944_ (.B1(_0413_),
    .Y(_0414_),
    .A1(net29),
    .A2(_0412_));
 sg13g2_nand2_1 _3945_ (.Y(_0415_),
    .A(_0414_),
    .B(net75));
 sg13g2_nor2_1 _3946_ (.A(net102),
    .B(_2346_),
    .Y(_0416_));
 sg13g2_inv_1 _3947_ (.Y(_0417_),
    .A(_0416_));
 sg13g2_a21oi_1 _3948_ (.A1(_0410_),
    .A2(_0415_),
    .Y(_0418_),
    .B1(_0417_));
 sg13g2_nand2_1 _3949_ (.Y(_0419_),
    .A(_0389_),
    .B(_0418_));
 sg13g2_nand2_1 _3950_ (.Y(_0420_),
    .A(_2877_),
    .B(_0198_));
 sg13g2_nor2_1 _3951_ (.A(_2852_),
    .B(_0420_),
    .Y(_0421_));
 sg13g2_nor2_1 _3952_ (.A(net23),
    .B(_2903_),
    .Y(_0422_));
 sg13g2_nand2_1 _3953_ (.Y(_0423_),
    .A(_0422_),
    .B(_0209_));
 sg13g2_nand2_1 _3954_ (.Y(_0424_),
    .A(_0423_),
    .B(_2914_));
 sg13g2_nand3_1 _3955_ (.B(_2899_),
    .C(_0424_),
    .A(_2892_),
    .Y(_0425_));
 sg13g2_nand2_1 _3956_ (.Y(_0426_),
    .A(_0425_),
    .B(_2919_));
 sg13g2_a21oi_1 _3957_ (.A1(_2924_),
    .A2(_0274_),
    .Y(_0427_),
    .B1(_2913_));
 sg13g2_nand2_1 _3958_ (.Y(_0428_),
    .A(_0427_),
    .B(net93));
 sg13g2_nor2b_1 _3959_ (.A(_2933_),
    .B_N(_0428_),
    .Y(_0429_));
 sg13g2_nor2_1 _3960_ (.A(_2922_),
    .B(_0429_),
    .Y(_0430_));
 sg13g2_nor2_2 _3961_ (.A(_2576_),
    .B(_2961_),
    .Y(_0431_));
 sg13g2_nor2b_1 _3962_ (.A(_0431_),
    .B_N(_2912_),
    .Y(_0432_));
 sg13g2_a21o_1 _3963_ (.A2(_2788_),
    .A1(_0432_),
    .B1(_2893_),
    .X(_0433_));
 sg13g2_a21oi_1 _3964_ (.A1(_0433_),
    .A2(_2953_),
    .Y(_0434_),
    .B1(net86));
 sg13g2_nand2b_1 _3965_ (.Y(_0435_),
    .B(_0192_),
    .A_N(_0434_));
 sg13g2_nand2_1 _3966_ (.Y(_0436_),
    .A(_0430_),
    .B(_0435_));
 sg13g2_nand3_1 _3967_ (.B(_0426_),
    .C(_0436_),
    .A(_0421_),
    .Y(_0437_));
 sg13g2_nand2_1 _3968_ (.Y(_0438_),
    .A(_2881_),
    .B(_2443_));
 sg13g2_nand2_1 _3969_ (.Y(_0439_),
    .A(_0438_),
    .B(_2946_));
 sg13g2_nand2_1 _3970_ (.Y(_0440_),
    .A(_0439_),
    .B(net93));
 sg13g2_a21oi_1 _3971_ (.A1(_0440_),
    .A2(_2593_),
    .Y(_0441_),
    .B1(net61));
 sg13g2_a21oi_1 _3972_ (.A1(_2833_),
    .A2(_2890_),
    .Y(_0442_),
    .B1(net87));
 sg13g2_nor2_1 _3973_ (.A(_0441_),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_nand2_1 _3974_ (.Y(_0444_),
    .A(_2805_),
    .B(_2788_));
 sg13g2_o21ai_1 _3975_ (.B1(_0444_),
    .Y(_0445_),
    .A1(_2568_),
    .A2(_0224_));
 sg13g2_nand2_1 _3976_ (.Y(_0446_),
    .A(_0445_),
    .B(net73));
 sg13g2_nand3_1 _3977_ (.B(_0446_),
    .C(_0236_),
    .A(_0443_),
    .Y(_0447_));
 sg13g2_nand2_1 _3978_ (.Y(_0448_),
    .A(_2855_),
    .B(net43));
 sg13g2_nor2b_1 _3979_ (.A(_0448_),
    .B_N(_2904_),
    .Y(_0449_));
 sg13g2_nand2_1 _3980_ (.Y(_0450_),
    .A(_0449_),
    .B(net17));
 sg13g2_nor3_1 _3981_ (.A(_0200_),
    .B(_0201_),
    .C(net16),
    .Y(_0451_));
 sg13g2_nor2_1 _3982_ (.A(net44),
    .B(_0448_),
    .Y(_0452_));
 sg13g2_nand2_2 _3983_ (.Y(_0453_),
    .A(_2795_),
    .B(net40));
 sg13g2_nand2_1 _3984_ (.Y(_0454_),
    .A(_0452_),
    .B(_0453_));
 sg13g2_nand4_1 _3985_ (.B(_0451_),
    .C(_0454_),
    .A(_0450_),
    .Y(_0455_),
    .D(_2820_));
 sg13g2_nand2_1 _3986_ (.Y(_0456_),
    .A(_0447_),
    .B(_0455_));
 sg13g2_nor2_1 _3987_ (.A(net102),
    .B(_2479_),
    .Y(_0457_));
 sg13g2_inv_1 _3988_ (.Y(_0458_),
    .A(_0457_));
 sg13g2_a21oi_1 _3989_ (.A1(_0456_),
    .A2(net71),
    .Y(_0459_),
    .B1(_0458_));
 sg13g2_nand2_1 _3990_ (.Y(_0460_),
    .A(_0437_),
    .B(_0459_));
 sg13g2_nand3_1 _3991_ (.B(_0419_),
    .C(_0460_),
    .A(_0322_),
    .Y(_0461_));
 sg13g2_nor2_1 _3992_ (.A(_0255_),
    .B(_0461_),
    .Y(_0462_));
 sg13g2_nor2_1 _3993_ (.A(_2478_),
    .B(_0462_),
    .Y(_0463_));
 sg13g2_nand2_1 _3994_ (.Y(_0464_),
    .A(_2906_),
    .B(_2859_));
 sg13g2_and2_1 _3995_ (.A(_0464_),
    .B(_0358_),
    .X(_0465_));
 sg13g2_nand2b_1 _3996_ (.Y(_0466_),
    .B(_0276_),
    .A_N(_0269_));
 sg13g2_nand2_1 _3997_ (.Y(_0467_),
    .A(_2832_),
    .B(net61));
 sg13g2_a21oi_1 _3998_ (.A1(_0465_),
    .A2(_0466_),
    .Y(_0468_),
    .B1(_0467_));
 sg13g2_inv_4 _3999_ (.A(_0360_),
    .Y(_0469_));
 sg13g2_nor2_1 _4000_ (.A(_0469_),
    .B(_0345_),
    .Y(_0470_));
 sg13g2_nor2_1 _4001_ (.A(_0468_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_a21oi_1 _4002_ (.A1(_2805_),
    .A2(_0188_),
    .Y(_0472_),
    .B1(_0290_));
 sg13g2_nand3_1 _4003_ (.B(net25),
    .C(_0324_),
    .A(_0323_),
    .Y(_0473_));
 sg13g2_a21oi_1 _4004_ (.A1(_0472_),
    .A2(_0473_),
    .Y(_0474_),
    .B1(_0263_));
 sg13g2_nor2_1 _4005_ (.A(_2771_),
    .B(_0474_),
    .Y(_0475_));
 sg13g2_nand2_1 _4006_ (.Y(_0476_),
    .A(_0471_),
    .B(_0475_));
 sg13g2_nand2_1 _4007_ (.Y(_0477_),
    .A(_0377_),
    .B(_2882_));
 sg13g2_nor2_1 _4008_ (.A(net70),
    .B(_0355_),
    .Y(_0478_));
 sg13g2_a21oi_1 _4009_ (.A1(_0477_),
    .A2(_2885_),
    .Y(_0479_),
    .B1(_0478_));
 sg13g2_nand2_1 _4010_ (.Y(_0480_),
    .A(_0372_),
    .B(_2924_));
 sg13g2_a21oi_1 _4011_ (.A1(_0480_),
    .A2(_2886_),
    .Y(_0481_),
    .B1(net78));
 sg13g2_nor2_1 _4012_ (.A(_0353_),
    .B(_2831_),
    .Y(_0482_));
 sg13g2_o21ai_1 _4013_ (.B1(net73),
    .Y(_0483_),
    .A1(_0482_),
    .A2(_0290_));
 sg13g2_nand3_1 _4014_ (.B(_0481_),
    .C(_0483_),
    .A(_0479_),
    .Y(_0484_));
 sg13g2_nand3_1 _4015_ (.B(_0484_),
    .C(_2777_),
    .A(_0476_),
    .Y(_0485_));
 sg13g2_nand2_1 _4016_ (.Y(_0486_),
    .A(_0385_),
    .B(net72));
 sg13g2_o21ai_1 _4017_ (.B1(_0486_),
    .Y(_0487_),
    .A1(_2909_),
    .A2(_0369_));
 sg13g2_o21ai_1 _4018_ (.B1(net57),
    .Y(_0488_),
    .A1(_2815_),
    .A2(_0487_));
 sg13g2_nand2_1 _4019_ (.Y(_0489_),
    .A(_0485_),
    .B(_0488_));
 sg13g2_a21oi_1 _4020_ (.A1(_0489_),
    .A2(_2482_),
    .Y(_0490_),
    .B1(_0420_));
 sg13g2_nor2_1 _4021_ (.A(_2788_),
    .B(_0381_),
    .Y(_0491_));
 sg13g2_o21ai_1 _4022_ (.B1(net29),
    .Y(_0492_),
    .A1(_2905_),
    .A2(_0491_));
 sg13g2_nand3b_1 _4023_ (.B(_0492_),
    .C(_0344_),
    .Y(_0493_),
    .A_N(_2889_));
 sg13g2_nand2_1 _4024_ (.Y(_0494_),
    .A(_0366_),
    .B(net41));
 sg13g2_nand2_1 _4025_ (.Y(_0495_),
    .A(_0432_),
    .B(_0494_));
 sg13g2_nor2_1 _4026_ (.A(net100),
    .B(net34),
    .Y(_0496_));
 sg13g2_a21oi_1 _4027_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(_2799_));
 sg13g2_o21ai_1 _4028_ (.B1(_0497_),
    .Y(_0498_),
    .A1(_2941_),
    .A2(_0377_));
 sg13g2_a22oi_1 _4029_ (.Y(_0499_),
    .B1(net63),
    .B2(_0498_),
    .A2(_2886_),
    .A1(_0493_));
 sg13g2_nand2_1 _4030_ (.Y(_0500_),
    .A(_0499_),
    .B(_2803_));
 sg13g2_nand2_1 _4031_ (.Y(_0501_),
    .A(_0500_),
    .B(net57));
 sg13g2_nor2_1 _4032_ (.A(_0392_),
    .B(_2883_),
    .Y(_0502_));
 sg13g2_o21ai_1 _4033_ (.B1(_0502_),
    .Y(_0503_),
    .A1(_2908_),
    .A2(_0343_));
 sg13g2_nand2_1 _4034_ (.Y(_0504_),
    .A(_0503_),
    .B(_0248_));
 sg13g2_o21ai_1 _4035_ (.B1(_0393_),
    .Y(_0505_),
    .A1(_2883_),
    .A2(_0359_));
 sg13g2_nand2_1 _4036_ (.Y(_0506_),
    .A(_0504_),
    .B(_0505_));
 sg13g2_o21ai_1 _4037_ (.B1(_0228_),
    .Y(_0507_),
    .A1(_0298_),
    .A2(_2925_));
 sg13g2_nand3_1 _4038_ (.B(_0475_),
    .C(_0507_),
    .A(_0506_),
    .Y(_0508_));
 sg13g2_a21oi_1 _4039_ (.A1(_0402_),
    .A2(net28),
    .Y(_0509_),
    .B1(net31));
 sg13g2_nand3_1 _4040_ (.B(net92),
    .C(net21),
    .A(_0509_),
    .Y(_0510_));
 sg13g2_nand2b_1 _4041_ (.Y(_0511_),
    .B(_2957_),
    .A_N(_0295_));
 sg13g2_nand3_1 _4042_ (.B(_0511_),
    .C(_2924_),
    .A(_0510_),
    .Y(_0512_));
 sg13g2_a21oi_1 _4043_ (.A1(_0512_),
    .A2(_2932_),
    .Y(_0513_),
    .B1(net78));
 sg13g2_nand3b_1 _4044_ (.B(net19),
    .C(_0330_),
    .Y(_0514_),
    .A_N(_0354_));
 sg13g2_a22oi_1 _4045_ (.Y(_0515_),
    .B1(_0228_),
    .B2(_0362_),
    .A2(_0341_),
    .A1(_0514_));
 sg13g2_a21oi_1 _4046_ (.A1(_0513_),
    .A2(_0515_),
    .Y(_0516_),
    .B1(_2917_));
 sg13g2_nand2_1 _4047_ (.Y(_0517_),
    .A(_0508_),
    .B(_0516_));
 sg13g2_nand2_1 _4048_ (.Y(_0518_),
    .A(_0501_),
    .B(_0517_));
 sg13g2_nand2_1 _4049_ (.Y(_0519_),
    .A(_0518_),
    .B(_0253_));
 sg13g2_nand2_1 _4050_ (.Y(_0520_),
    .A(_0490_),
    .B(_0519_));
 sg13g2_a21oi_1 _4051_ (.A1(_0413_),
    .A2(_0209_),
    .Y(_0521_),
    .B1(net87));
 sg13g2_a21oi_1 _4052_ (.A1(_2444_),
    .A2(net40),
    .Y(_0522_),
    .B1(_2839_));
 sg13g2_a22oi_1 _4053_ (.Y(_0523_),
    .B1(net29),
    .B2(_0522_),
    .A2(_0411_),
    .A1(_2906_));
 sg13g2_nor2_1 _4054_ (.A(net77),
    .B(_0523_),
    .Y(_0524_));
 sg13g2_nor2_1 _4055_ (.A(_0521_),
    .B(_0524_),
    .Y(_0525_));
 sg13g2_inv_1 _4056_ (.Y(_0526_),
    .A(net30));
 sg13g2_nand2_1 _4057_ (.Y(_0527_),
    .A(_2786_),
    .B(_0453_));
 sg13g2_a22oi_1 _4058_ (.Y(_0528_),
    .B1(_0206_),
    .B2(_0354_),
    .A2(_0233_),
    .A1(net17));
 sg13g2_o21ai_1 _4059_ (.B1(_0528_),
    .Y(_0529_),
    .A1(_0526_),
    .A2(_0527_));
 sg13g2_nand2_1 _4060_ (.Y(_0530_),
    .A(_0529_),
    .B(net73));
 sg13g2_nand2_1 _4061_ (.Y(_0531_),
    .A(_2934_),
    .B(net40));
 sg13g2_nand2_1 _4062_ (.Y(_0532_),
    .A(_0233_),
    .B(net21));
 sg13g2_nand2_1 _4063_ (.Y(_0533_),
    .A(_0531_),
    .B(_0532_));
 sg13g2_nand3_1 _4064_ (.B(_0279_),
    .C(_0295_),
    .A(_0533_),
    .Y(_0534_));
 sg13g2_nand4_1 _4065_ (.B(_0530_),
    .C(_0390_),
    .A(_0525_),
    .Y(_0535_),
    .D(_0534_));
 sg13g2_inv_1 _4066_ (.Y(_0536_),
    .A(_0453_));
 sg13g2_o21ai_1 _4067_ (.B1(_0207_),
    .Y(_0537_),
    .A1(_2577_),
    .A2(_0536_));
 sg13g2_nor2_1 _4068_ (.A(net43),
    .B(_0399_),
    .Y(_0538_));
 sg13g2_nand2_1 _4069_ (.Y(_0539_),
    .A(_0538_),
    .B(_2786_));
 sg13g2_a21oi_1 _4070_ (.A1(_0539_),
    .A2(_0207_),
    .Y(_0540_),
    .B1(net17));
 sg13g2_a21oi_1 _4071_ (.A1(_2569_),
    .A2(_0537_),
    .Y(_0541_),
    .B1(_0540_));
 sg13g2_a21oi_1 _4072_ (.A1(_0541_),
    .A2(_0451_),
    .Y(_0542_),
    .B1(_2482_));
 sg13g2_a21oi_1 _4073_ (.A1(_0535_),
    .A2(_0542_),
    .Y(_0543_),
    .B1(_0198_));
 sg13g2_nand2_1 _4074_ (.Y(_0544_),
    .A(_2924_),
    .B(_0209_));
 sg13g2_o21ai_1 _4075_ (.B1(_0413_),
    .Y(_0545_),
    .A1(_2907_),
    .A2(_2867_));
 sg13g2_a22oi_1 _4076_ (.Y(_0546_),
    .B1(_2941_),
    .B2(_0545_),
    .A2(_0544_),
    .A1(_0371_));
 sg13g2_nand4_1 _4077_ (.B(_0326_),
    .C(_2594_),
    .A(_0531_),
    .Y(_0547_),
    .D(net55));
 sg13g2_nand2_1 _4078_ (.Y(_0548_),
    .A(_0394_),
    .B(_0239_));
 sg13g2_nand3_1 _4079_ (.B(_0532_),
    .C(_2594_),
    .A(_0548_),
    .Y(_0549_));
 sg13g2_nor2_1 _4080_ (.A(net89),
    .B(_0264_),
    .Y(_0550_));
 sg13g2_inv_1 _4081_ (.Y(_0551_),
    .A(_0550_));
 sg13g2_a21o_1 _4082_ (.A2(_0241_),
    .A1(_0549_),
    .B1(_0551_),
    .X(_0552_));
 sg13g2_o21ai_1 _4083_ (.B1(_0552_),
    .Y(_0553_),
    .A1(_0547_),
    .A2(_0529_));
 sg13g2_o21ai_1 _4084_ (.B1(_0553_),
    .Y(_0554_),
    .A1(net63),
    .A2(_0546_));
 sg13g2_o21ai_1 _4085_ (.B1(_2569_),
    .Y(_0555_),
    .A1(net20),
    .A2(_0453_));
 sg13g2_o21ai_1 _4086_ (.B1(_0451_),
    .Y(_0556_),
    .A1(_0449_),
    .A2(_0555_));
 sg13g2_a21o_1 _4087_ (.A2(_0537_),
    .A1(net29),
    .B1(_0556_),
    .X(_0557_));
 sg13g2_nand3_1 _4088_ (.B(_2482_),
    .C(_0557_),
    .A(_0554_),
    .Y(_0558_));
 sg13g2_inv_1 _4089_ (.Y(_0559_),
    .A(_2478_));
 sg13g2_a21oi_1 _4090_ (.A1(_0543_),
    .A2(_0558_),
    .Y(_0560_),
    .B1(_0559_));
 sg13g2_nor4_1 _4091_ (.A(net20),
    .B(net19),
    .C(net29),
    .D(_2600_),
    .Y(_0561_));
 sg13g2_a22oi_1 _4092_ (.Y(_0562_),
    .B1(_2911_),
    .B2(_0561_),
    .A2(_2601_),
    .A1(net19));
 sg13g2_nor2_1 _4093_ (.A(_0393_),
    .B(_2780_),
    .Y(_0563_));
 sg13g2_nor2_1 _4094_ (.A(_0198_),
    .B(net55),
    .Y(_0564_));
 sg13g2_nand2_1 _4095_ (.Y(_0565_),
    .A(_0196_),
    .B(_2604_));
 sg13g2_nor2_1 _4096_ (.A(_2608_),
    .B(_2716_),
    .Y(_0566_));
 sg13g2_nand2_1 _4097_ (.Y(_0567_),
    .A(_2775_),
    .B(_2604_));
 sg13g2_inv_1 _4098_ (.Y(_0568_),
    .A(_0567_));
 sg13g2_a21oi_1 _4099_ (.A1(_0568_),
    .A2(_0196_),
    .Y(_0569_),
    .B1(_2608_));
 sg13g2_inv_1 _4100_ (.Y(_0570_),
    .A(_0569_));
 sg13g2_a22oi_1 _4101_ (.Y(_0571_),
    .B1(_2716_),
    .B2(_0570_),
    .A2(_0566_),
    .A1(_0565_));
 sg13g2_xnor2_1 _4102_ (.Y(_0572_),
    .A(_2608_),
    .B(_0567_));
 sg13g2_nor2b_1 _4103_ (.A(_0571_),
    .B_N(_0572_),
    .Y(_0573_));
 sg13g2_inv_1 _4104_ (.Y(_0574_),
    .A(_0573_));
 sg13g2_a221oi_1 _4105_ (.B2(_0564_),
    .C1(_0574_),
    .B1(_0201_),
    .A1(net71),
    .Y(_0575_),
    .A2(_0563_));
 sg13g2_nor2b_1 _4106_ (.A(_0562_),
    .B_N(_0575_),
    .Y(_0576_));
 sg13g2_inv_1 _4107_ (.Y(_0577_),
    .A(_0576_));
 sg13g2_a21oi_1 _4108_ (.A1(_0520_),
    .A2(_0560_),
    .Y(_0578_),
    .B1(_0577_));
 sg13g2_nor2b_1 _4109_ (.A(_0463_),
    .B_N(_0578_),
    .Y(_0579_));
 sg13g2_a21oi_1 _4110_ (.A1(_2782_),
    .A2(net26),
    .Y(_0580_),
    .B1(net48));
 sg13g2_nor3_1 _4111_ (.A(net18),
    .B(_0452_),
    .C(_0580_),
    .Y(_0581_));
 sg13g2_nor2_1 _4112_ (.A(net94),
    .B(_0581_),
    .Y(_0582_));
 sg13g2_nand2_1 _4113_ (.Y(_0583_),
    .A(net30),
    .B(_2960_));
 sg13g2_nand2_1 _4114_ (.Y(_0584_),
    .A(_0454_),
    .B(_0583_));
 sg13g2_nand2_1 _4115_ (.Y(_0585_),
    .A(_2853_),
    .B(_2573_));
 sg13g2_nand2_1 _4116_ (.Y(_0586_),
    .A(_0585_),
    .B(_2564_));
 sg13g2_buf_2 _4117_ (.A(_0586_),
    .X(_0587_));
 sg13g2_nand2_1 _4118_ (.Y(_0588_),
    .A(net31),
    .B(net34));
 sg13g2_nand3_1 _4119_ (.B(net32),
    .C(_0588_),
    .A(_0587_),
    .Y(_0589_));
 sg13g2_nor2_1 _4120_ (.A(_0584_),
    .B(_0589_),
    .Y(_0590_));
 sg13g2_nor2_1 _4121_ (.A(net74),
    .B(_0590_),
    .Y(_0591_));
 sg13g2_nor2_1 _4122_ (.A(_0582_),
    .B(_0591_),
    .Y(_0592_));
 sg13g2_nor3_1 _4123_ (.A(net22),
    .B(_2911_),
    .C(_2522_),
    .Y(_0593_));
 sg13g2_nor3_1 _4124_ (.A(_0593_),
    .B(_2854_),
    .C(_2857_),
    .Y(_0594_));
 sg13g2_nand2b_1 _4125_ (.Y(_0595_),
    .B(net81),
    .A_N(_0594_));
 sg13g2_nor2_2 _4126_ (.A(net45),
    .B(_2519_),
    .Y(_0596_));
 sg13g2_nor2_1 _4127_ (.A(_2869_),
    .B(_0596_),
    .Y(_0597_));
 sg13g2_nor2_1 _4128_ (.A(_0526_),
    .B(_0597_),
    .Y(_0598_));
 sg13g2_nand2_2 _4129_ (.Y(_0599_),
    .A(_0587_),
    .B(net42));
 sg13g2_nor2_1 _4130_ (.A(_0598_),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_nor2_1 _4131_ (.A(_2911_),
    .B(_0381_),
    .Y(_0601_));
 sg13g2_nand3_1 _4132_ (.B(net20),
    .C(net39),
    .A(_0601_),
    .Y(_0602_));
 sg13g2_nand2_1 _4133_ (.Y(_0603_),
    .A(_0600_),
    .B(_0602_));
 sg13g2_nand2_1 _4134_ (.Y(_0604_),
    .A(_0603_),
    .B(net72));
 sg13g2_nand3_1 _4135_ (.B(_0595_),
    .C(_0604_),
    .A(_0592_),
    .Y(_0605_));
 sg13g2_a21oi_1 _4136_ (.A1(_2822_),
    .A2(_2575_),
    .Y(_0606_),
    .B1(_2792_));
 sg13g2_nor2_1 _4137_ (.A(net23),
    .B(_0606_),
    .Y(_0607_));
 sg13g2_nand2_1 _4138_ (.Y(_0608_),
    .A(_0607_),
    .B(_2935_));
 sg13g2_nor2_1 _4139_ (.A(net70),
    .B(_0608_),
    .Y(_0609_));
 sg13g2_nand3_1 _4140_ (.B(net39),
    .C(_0411_),
    .A(_2783_),
    .Y(_0610_));
 sg13g2_a21oi_1 _4141_ (.A1(_0448_),
    .A2(net22),
    .Y(_0611_),
    .B1(net18));
 sg13g2_and3_1 _4142_ (.X(_0612_),
    .A(_0610_),
    .B(net80),
    .C(_0611_));
 sg13g2_nor3_1 _4143_ (.A(_0264_),
    .B(_0609_),
    .C(_0612_),
    .Y(_0613_));
 sg13g2_a21oi_1 _4144_ (.A1(_0605_),
    .A2(net57),
    .Y(_0614_),
    .B1(_0613_));
 sg13g2_nand2_1 _4145_ (.Y(_0615_),
    .A(_0215_),
    .B(_2564_));
 sg13g2_nor2_1 _4146_ (.A(_0402_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_nor2_1 _4147_ (.A(net100),
    .B(_0616_),
    .Y(_0617_));
 sg13g2_nand2_1 _4148_ (.Y(_0618_),
    .A(_2911_),
    .B(net33));
 sg13g2_nand2_1 _4149_ (.Y(_0619_),
    .A(_0219_),
    .B(_0618_));
 sg13g2_nand2_1 _4150_ (.Y(_0620_),
    .A(_0619_),
    .B(net48));
 sg13g2_a21oi_1 _4151_ (.A1(_0617_),
    .A2(_0620_),
    .Y(_0621_),
    .B1(_2861_));
 sg13g2_nand2_1 _4152_ (.Y(_0622_),
    .A(net30),
    .B(_2869_));
 sg13g2_nand2_1 _4153_ (.Y(_0623_),
    .A(_2946_),
    .B(_0622_));
 sg13g2_nor2_1 _4154_ (.A(net111),
    .B(_0623_),
    .Y(_0624_));
 sg13g2_nand2_1 _4155_ (.Y(_0625_),
    .A(_2816_),
    .B(_2786_));
 sg13g2_nand2_1 _4156_ (.Y(_0626_),
    .A(_0625_),
    .B(net46));
 sg13g2_a21oi_1 _4157_ (.A1(net41),
    .A2(_2498_),
    .Y(_0627_),
    .B1(net56));
 sg13g2_nand2_1 _4158_ (.Y(_0628_),
    .A(_0626_),
    .B(_0627_));
 sg13g2_nand2_1 _4159_ (.Y(_0629_),
    .A(_0624_),
    .B(_0628_));
 sg13g2_nand2_1 _4160_ (.Y(_0630_),
    .A(net41),
    .B(_2498_));
 sg13g2_nand2_1 _4161_ (.Y(_0631_),
    .A(_0630_),
    .B(net34));
 sg13g2_nand2_1 _4162_ (.Y(_0632_),
    .A(_2949_),
    .B(_0631_));
 sg13g2_nand3_1 _4163_ (.B(_0400_),
    .C(net82),
    .A(_0632_),
    .Y(_0633_));
 sg13g2_nand2_1 _4164_ (.Y(_0634_),
    .A(_0633_),
    .B(net19));
 sg13g2_a21oi_1 _4165_ (.A1(_0621_),
    .A2(_0629_),
    .Y(_0635_),
    .B1(_0634_));
 sg13g2_nor2_1 _4166_ (.A(_0381_),
    .B(_0615_),
    .Y(_0636_));
 sg13g2_nand3_1 _4167_ (.B(_2575_),
    .C(_2792_),
    .A(_0596_),
    .Y(_0637_));
 sg13g2_nand2_1 _4168_ (.Y(_0638_),
    .A(_2948_),
    .B(_0349_));
 sg13g2_nand3_1 _4169_ (.B(_0637_),
    .C(_0638_),
    .A(_0275_),
    .Y(_0639_));
 sg13g2_o21ai_1 _4170_ (.B1(net80),
    .Y(_0640_),
    .A1(_0636_),
    .A2(_0639_));
 sg13g2_a21oi_1 _4171_ (.A1(_0635_),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0268_));
 sg13g2_a21oi_1 _4172_ (.A1(_2902_),
    .A2(_2816_),
    .Y(_0642_),
    .B1(_2935_));
 sg13g2_nand2_1 _4173_ (.Y(_0643_),
    .A(_0275_),
    .B(_0638_));
 sg13g2_nor2_1 _4174_ (.A(_0642_),
    .B(_0643_),
    .Y(_0644_));
 sg13g2_nand2_1 _4175_ (.Y(_0645_),
    .A(_2521_),
    .B(_2469_));
 sg13g2_a21oi_1 _4176_ (.A1(_0645_),
    .A2(net33),
    .Y(_0646_),
    .B1(net49));
 sg13g2_nor2_1 _4177_ (.A(net23),
    .B(_0646_),
    .Y(_0647_));
 sg13g2_a21oi_1 _4178_ (.A1(_0644_),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net70));
 sg13g2_nand2_1 _4179_ (.Y(_0649_),
    .A(_2956_),
    .B(net33));
 sg13g2_nand2_1 _4180_ (.Y(_0650_),
    .A(_0538_),
    .B(_0645_));
 sg13g2_nand2_1 _4181_ (.Y(_0651_),
    .A(_0649_),
    .B(_0650_));
 sg13g2_nand2_1 _4182_ (.Y(_0652_),
    .A(_0651_),
    .B(_2844_));
 sg13g2_nand2_1 _4183_ (.Y(_0653_),
    .A(_0652_),
    .B(_0607_));
 sg13g2_nand2_1 _4184_ (.Y(_0654_),
    .A(_0653_),
    .B(net89));
 sg13g2_nor2_1 _4185_ (.A(_2573_),
    .B(_0402_),
    .Y(_0655_));
 sg13g2_nand2_1 _4186_ (.Y(_0656_),
    .A(_0655_),
    .B(_2522_));
 sg13g2_nand2_1 _4187_ (.Y(_0657_),
    .A(_2839_),
    .B(_0645_));
 sg13g2_nand2_1 _4188_ (.Y(_0658_),
    .A(_0656_),
    .B(_0657_));
 sg13g2_nand2_1 _4189_ (.Y(_0659_),
    .A(_0658_),
    .B(net49));
 sg13g2_inv_2 _4190_ (.Y(_0660_),
    .A(_0599_));
 sg13g2_nand2_1 _4191_ (.Y(_0661_),
    .A(_0659_),
    .B(_0660_));
 sg13g2_nand2_1 _4192_ (.Y(_0662_),
    .A(_0661_),
    .B(net83));
 sg13g2_nand2_1 _4193_ (.Y(_0663_),
    .A(_0206_),
    .B(_2841_));
 sg13g2_nand2_1 _4194_ (.Y(_0664_),
    .A(_0663_),
    .B(net41));
 sg13g2_nand2_1 _4195_ (.Y(_0665_),
    .A(_0664_),
    .B(net34));
 sg13g2_nand2_1 _4196_ (.Y(_0666_),
    .A(_0422_),
    .B(_0665_));
 sg13g2_nand2_1 _4197_ (.Y(_0667_),
    .A(_0666_),
    .B(net90));
 sg13g2_nand3_1 _4198_ (.B(_0662_),
    .C(_0667_),
    .A(_0654_),
    .Y(_0668_));
 sg13g2_nor2_1 _4199_ (.A(_0648_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nor2_1 _4200_ (.A(_2922_),
    .B(_0669_),
    .Y(_0670_));
 sg13g2_nor2_1 _4201_ (.A(_0641_),
    .B(_0670_),
    .Y(_0671_));
 sg13g2_nand2_1 _4202_ (.Y(_0672_),
    .A(_0614_),
    .B(_0671_));
 sg13g2_a21oi_1 _4203_ (.A1(_0672_),
    .A2(_0416_),
    .Y(_0673_),
    .B1(net71));
 sg13g2_nand3_1 _4204_ (.B(net35),
    .C(_2855_),
    .A(_2904_),
    .Y(_0674_));
 sg13g2_nand3_1 _4205_ (.B(_0674_),
    .C(net27),
    .A(_0664_),
    .Y(_0675_));
 sg13g2_inv_1 _4206_ (.Y(_0676_),
    .A(_0622_));
 sg13g2_nor2_1 _4207_ (.A(_2931_),
    .B(_0676_),
    .Y(_0677_));
 sg13g2_a21oi_1 _4208_ (.A1(_0675_),
    .A2(_0677_),
    .Y(_0678_),
    .B1(net18));
 sg13g2_o21ai_1 _4209_ (.B1(_0327_),
    .Y(_0679_),
    .A1(net26),
    .A2(_0219_));
 sg13g2_nand2_1 _4210_ (.Y(_0680_),
    .A(_0679_),
    .B(net48));
 sg13g2_a21oi_1 _4211_ (.A1(_0215_),
    .A2(net27),
    .Y(_0681_),
    .B1(_2861_));
 sg13g2_nand2_1 _4212_ (.Y(_0682_),
    .A(_0680_),
    .B(_0681_));
 sg13g2_nand2_1 _4213_ (.Y(_0683_),
    .A(_0678_),
    .B(_0682_));
 sg13g2_nand2_1 _4214_ (.Y(_0684_),
    .A(_0683_),
    .B(_2897_));
 sg13g2_nand2_1 _4215_ (.Y(_0685_),
    .A(_0684_),
    .B(net86));
 sg13g2_nand3_1 _4216_ (.B(_2807_),
    .C(_0650_),
    .A(_0382_),
    .Y(_0686_));
 sg13g2_nand2_1 _4217_ (.Y(_0687_),
    .A(_0686_),
    .B(net39));
 sg13g2_nand4_1 _4218_ (.B(_2786_),
    .C(_0453_),
    .A(_0630_),
    .Y(_0688_),
    .D(net44));
 sg13g2_nand3_1 _4219_ (.B(net25),
    .C(_0688_),
    .A(_0687_),
    .Y(_0689_));
 sg13g2_nor2_1 _4220_ (.A(_2935_),
    .B(_0597_),
    .Y(_0690_));
 sg13g2_a21oi_1 _4221_ (.A1(net30),
    .A2(_0220_),
    .Y(_0691_),
    .B1(_0690_));
 sg13g2_and2_1 _4222_ (.A(_0691_),
    .B(_0647_),
    .X(_0692_));
 sg13g2_nor2_1 _4223_ (.A(_0469_),
    .B(_0692_),
    .Y(_0693_));
 sg13g2_a21oi_1 _4224_ (.A1(_0689_),
    .A2(_0502_),
    .Y(_0694_),
    .B1(_0693_));
 sg13g2_nand2_1 _4225_ (.Y(_0695_),
    .A(_0685_),
    .B(_0694_));
 sg13g2_nand2_1 _4226_ (.Y(_0696_),
    .A(_0695_),
    .B(_0457_));
 sg13g2_nand3_1 _4227_ (.B(_2469_),
    .C(_2521_),
    .A(net33),
    .Y(_0697_));
 sg13g2_nand2b_1 _4228_ (.Y(_0698_),
    .B(_0697_),
    .A_N(_0655_));
 sg13g2_a21oi_1 _4229_ (.A1(_0698_),
    .A2(net21),
    .Y(_0699_),
    .B1(net92));
 sg13g2_a21oi_1 _4230_ (.A1(_0699_),
    .A2(_0691_),
    .Y(_0700_),
    .B1(net61));
 sg13g2_nor2_1 _4231_ (.A(net52),
    .B(_0663_),
    .Y(_0701_));
 sg13g2_o21ai_1 _4232_ (.B1(net21),
    .Y(_0702_),
    .A1(_0655_),
    .A2(_0701_));
 sg13g2_nand3_1 _4233_ (.B(net86),
    .C(_0622_),
    .A(_0702_),
    .Y(_0703_));
 sg13g2_a21oi_1 _4234_ (.A1(_0700_),
    .A2(_0703_),
    .Y(_0704_),
    .B1(net16));
 sg13g2_nand3_1 _4235_ (.B(net79),
    .C(_0688_),
    .A(_0687_),
    .Y(_0705_));
 sg13g2_nor2_1 _4236_ (.A(net100),
    .B(_0636_),
    .Y(_0706_));
 sg13g2_a21oi_1 _4237_ (.A1(_0680_),
    .A2(_0706_),
    .Y(_0707_),
    .B1(net63));
 sg13g2_nand2_1 _4238_ (.Y(_0708_),
    .A(_0705_),
    .B(_0707_));
 sg13g2_nand2_1 _4239_ (.Y(_0709_),
    .A(_0704_),
    .B(_0708_));
 sg13g2_nor2_1 _4240_ (.A(_0254_),
    .B(_2883_),
    .Y(_0710_));
 sg13g2_nand2_1 _4241_ (.Y(_0711_),
    .A(_0709_),
    .B(_0710_));
 sg13g2_nand2_1 _4242_ (.Y(_0712_),
    .A(_0696_),
    .B(_0711_));
 sg13g2_nor2_1 _4243_ (.A(_2818_),
    .B(_2935_),
    .Y(_0713_));
 sg13g2_inv_1 _4244_ (.Y(_0714_),
    .A(_2786_));
 sg13g2_nand2_1 _4245_ (.Y(_0715_),
    .A(net30),
    .B(_0714_));
 sg13g2_nand2_1 _4246_ (.Y(_0716_),
    .A(_0715_),
    .B(net32));
 sg13g2_nor3_1 _4247_ (.A(_0713_),
    .B(_2854_),
    .C(_0716_),
    .Y(_0717_));
 sg13g2_nor2_1 _4248_ (.A(net77),
    .B(_0717_),
    .Y(_0718_));
 sg13g2_o21ai_1 _4249_ (.B1(net82),
    .Y(_0719_),
    .A1(_0627_),
    .A2(_0716_));
 sg13g2_nand2_1 _4250_ (.Y(_0720_),
    .A(_2948_),
    .B(_0302_));
 sg13g2_nand3_1 _4251_ (.B(_2593_),
    .C(_0720_),
    .A(_0587_),
    .Y(_0721_));
 sg13g2_nand2_1 _4252_ (.Y(_0722_),
    .A(_0721_),
    .B(_0360_));
 sg13g2_nand2_1 _4253_ (.Y(_0723_),
    .A(_0719_),
    .B(_0722_));
 sg13g2_nor2_1 _4254_ (.A(_0718_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_a22oi_1 _4255_ (.Y(_0725_),
    .B1(net39),
    .B2(_0449_),
    .A2(net30),
    .A1(_2784_));
 sg13g2_nand2b_1 _4256_ (.Y(_0726_),
    .B(_0725_),
    .A_N(_0589_));
 sg13g2_nand2_1 _4257_ (.Y(_0727_),
    .A(_0726_),
    .B(net75));
 sg13g2_nand2_1 _4258_ (.Y(_0728_),
    .A(_0724_),
    .B(_0727_));
 sg13g2_o21ai_1 _4259_ (.B1(_2771_),
    .Y(_0729_),
    .A1(net74),
    .A2(_0608_));
 sg13g2_nor2_1 _4260_ (.A(_2777_),
    .B(_0729_),
    .Y(_0730_));
 sg13g2_a21oi_1 _4261_ (.A1(_0728_),
    .A2(_2919_),
    .Y(_0731_),
    .B1(_0730_));
 sg13g2_a21oi_1 _4262_ (.A1(_0610_),
    .A2(_0611_),
    .Y(_0732_),
    .B1(net94));
 sg13g2_nor2_1 _4263_ (.A(_0392_),
    .B(_0581_),
    .Y(_0733_));
 sg13g2_nor2_1 _4264_ (.A(_0732_),
    .B(_0733_),
    .Y(_0734_));
 sg13g2_nor2_1 _4265_ (.A(_2838_),
    .B(_0448_),
    .Y(_0735_));
 sg13g2_o21ai_1 _4266_ (.B1(net39),
    .Y(_0736_),
    .A1(_0431_),
    .A2(_0735_));
 sg13g2_inv_1 _4267_ (.Y(_0737_),
    .A(_0716_));
 sg13g2_nand3_1 _4268_ (.B(_0587_),
    .C(_0737_),
    .A(_0736_),
    .Y(_0738_));
 sg13g2_nand2_1 _4269_ (.Y(_0739_),
    .A(_0738_),
    .B(net80));
 sg13g2_o21ai_1 _4270_ (.B1(_2858_),
    .Y(_0740_),
    .A1(net21),
    .A2(_2841_));
 sg13g2_nand2_1 _4271_ (.Y(_0741_),
    .A(_0740_),
    .B(net72));
 sg13g2_nand3_1 _4272_ (.B(_0739_),
    .C(_0741_),
    .A(_0734_),
    .Y(_0742_));
 sg13g2_nand2_1 _4273_ (.Y(_0743_),
    .A(_0742_),
    .B(net57));
 sg13g2_a21oi_1 _4274_ (.A1(_0731_),
    .A2(_0743_),
    .Y(_0744_),
    .B1(_2479_));
 sg13g2_a21oi_1 _4275_ (.A1(_0712_),
    .A2(_2921_),
    .Y(_0745_),
    .B1(_0744_));
 sg13g2_nand2_1 _4276_ (.Y(_0746_),
    .A(_2956_),
    .B(net35));
 sg13g2_nand3_1 _4277_ (.B(_2303_),
    .C(_2853_),
    .A(_0746_),
    .Y(_0747_));
 sg13g2_nand2b_1 _4278_ (.Y(_0748_),
    .B(_0747_),
    .A_N(_0496_));
 sg13g2_nand2_1 _4279_ (.Y(_0749_),
    .A(_0687_),
    .B(_0748_));
 sg13g2_nor2_1 _4280_ (.A(net92),
    .B(_0676_),
    .Y(_0750_));
 sg13g2_a21oi_1 _4281_ (.A1(_0750_),
    .A2(_0665_),
    .Y(_0751_),
    .B1(net16));
 sg13g2_nand2_1 _4282_ (.Y(_0752_),
    .A(_0749_),
    .B(_0751_));
 sg13g2_nand2_1 _4283_ (.Y(_0753_),
    .A(_0752_),
    .B(_2897_));
 sg13g2_nand2_1 _4284_ (.Y(_0754_),
    .A(_0753_),
    .B(net61));
 sg13g2_nor2_1 _4285_ (.A(_0342_),
    .B(_0692_),
    .Y(_0755_));
 sg13g2_o21ai_1 _4286_ (.B1(_0395_),
    .Y(_0756_),
    .A1(_2577_),
    .A2(_2784_));
 sg13g2_and2_1 _4287_ (.A(_0756_),
    .B(_0607_),
    .X(_0757_));
 sg13g2_o21ai_1 _4288_ (.B1(net78),
    .Y(_0758_),
    .A1(net74),
    .A2(_0757_));
 sg13g2_nor2_1 _4289_ (.A(_0755_),
    .B(_0758_),
    .Y(_0759_));
 sg13g2_nand2_1 _4290_ (.Y(_0760_),
    .A(_0754_),
    .B(_0759_));
 sg13g2_a21oi_1 _4291_ (.A1(_0617_),
    .A2(_0720_),
    .Y(_0761_),
    .B1(net18));
 sg13g2_nor2_1 _4292_ (.A(net65),
    .B(net35),
    .Y(_0762_));
 sg13g2_nor3_1 _4293_ (.A(net48),
    .B(_0762_),
    .C(_0527_),
    .Y(_0763_));
 sg13g2_nor2_1 _4294_ (.A(net92),
    .B(_0763_),
    .Y(_0764_));
 sg13g2_nand2_1 _4295_ (.Y(_0765_),
    .A(_0680_),
    .B(_0764_));
 sg13g2_nand2_1 _4296_ (.Y(_0766_),
    .A(_0761_),
    .B(_0765_));
 sg13g2_nand2_1 _4297_ (.Y(_0767_),
    .A(_0766_),
    .B(_2897_));
 sg13g2_nand2_1 _4298_ (.Y(_0768_),
    .A(_0767_),
    .B(net63));
 sg13g2_nand2_1 _4299_ (.Y(_0769_),
    .A(_0627_),
    .B(_0244_));
 sg13g2_a21oi_1 _4300_ (.A1(_0737_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(net77));
 sg13g2_nor2_1 _4301_ (.A(net87),
    .B(_0717_),
    .Y(_0771_));
 sg13g2_nor3_1 _4302_ (.A(net78),
    .B(_0770_),
    .C(_0771_),
    .Y(_0772_));
 sg13g2_nand2_1 _4303_ (.Y(_0773_),
    .A(_0768_),
    .B(_0772_));
 sg13g2_nand3_1 _4304_ (.B(_0773_),
    .C(_2777_),
    .A(_0760_),
    .Y(_0774_));
 sg13g2_a22oi_1 _4305_ (.Y(_0775_),
    .B1(net73),
    .B2(_0726_),
    .A2(net81),
    .A1(_0740_));
 sg13g2_a21oi_1 _4306_ (.A1(_0738_),
    .A2(net72),
    .Y(_0776_),
    .B1(_0582_));
 sg13g2_nand2_1 _4307_ (.Y(_0777_),
    .A(_0775_),
    .B(_0776_));
 sg13g2_a21oi_1 _4308_ (.A1(_0777_),
    .A2(net57),
    .Y(_0778_),
    .B1(_0613_));
 sg13g2_nand2_1 _4309_ (.Y(_0779_),
    .A(_0774_),
    .B(_0778_));
 sg13g2_nand2_1 _4310_ (.Y(_0780_),
    .A(_0779_),
    .B(_2483_));
 sg13g2_nand3_1 _4311_ (.B(_0745_),
    .C(_0780_),
    .A(_0673_),
    .Y(_0781_));
 sg13g2_nor2_1 _4312_ (.A(net24),
    .B(_0522_),
    .Y(_0782_));
 sg13g2_nor2_1 _4313_ (.A(net87),
    .B(_0782_),
    .Y(_0783_));
 sg13g2_a21oi_1 _4314_ (.A1(_0412_),
    .A2(_2894_),
    .Y(_0784_),
    .B1(net77));
 sg13g2_nor3_1 _4315_ (.A(net45),
    .B(_2900_),
    .C(net28),
    .Y(_0785_));
 sg13g2_nor2_1 _4316_ (.A(_0785_),
    .B(_0209_),
    .Y(_0786_));
 sg13g2_nor3_1 _4317_ (.A(_0200_),
    .B(_0271_),
    .C(_0786_),
    .Y(_0787_));
 sg13g2_nand2b_1 _4318_ (.Y(_0788_),
    .B(_0746_),
    .A_N(_0403_));
 sg13g2_nand2_1 _4319_ (.Y(_0789_),
    .A(_0788_),
    .B(_0239_));
 sg13g2_a21oi_1 _4320_ (.A1(_0787_),
    .A2(_0789_),
    .Y(_0790_),
    .B1(net61));
 sg13g2_nor3_1 _4321_ (.A(_0783_),
    .B(_0784_),
    .C(_0790_),
    .Y(_0791_));
 sg13g2_a21oi_1 _4322_ (.A1(_0791_),
    .A2(net55),
    .Y(_0792_),
    .B1(_0417_));
 sg13g2_nand3_1 _4323_ (.B(_0217_),
    .C(_0373_),
    .A(_2826_),
    .Y(_0793_));
 sg13g2_nand2_1 _4324_ (.Y(_0794_),
    .A(_0793_),
    .B(net81));
 sg13g2_o21ai_1 _4325_ (.B1(_0794_),
    .Y(_0795_),
    .A1(net87),
    .A2(_0757_));
 sg13g2_nor2_1 _4326_ (.A(_0264_),
    .B(_0795_),
    .Y(_0796_));
 sg13g2_o21ai_1 _4327_ (.B1(_2820_),
    .Y(_0797_),
    .A1(_0399_),
    .A2(_0585_));
 sg13g2_nand2_1 _4328_ (.Y(_0798_),
    .A(_0797_),
    .B(net17));
 sg13g2_nand2_1 _4329_ (.Y(_0799_),
    .A(_0625_),
    .B(net20));
 sg13g2_a21oi_1 _4330_ (.A1(_0799_),
    .A2(_0204_),
    .Y(_0800_),
    .B1(net16));
 sg13g2_nand2_1 _4331_ (.Y(_0801_),
    .A(_0798_),
    .B(_0800_));
 sg13g2_a22oi_1 _4332_ (.Y(_0802_),
    .B1(net73),
    .B2(_0801_),
    .A2(_0230_),
    .A1(net72));
 sg13g2_a21oi_1 _4333_ (.A1(_0796_),
    .A2(_0802_),
    .Y(_0803_),
    .B1(_0254_));
 sg13g2_nor2_1 _4334_ (.A(_0411_),
    .B(_2893_),
    .Y(_0804_));
 sg13g2_inv_2 _4335_ (.Y(_0805_),
    .A(_0804_));
 sg13g2_inv_1 _4336_ (.Y(_0806_),
    .A(_0482_));
 sg13g2_nor2_1 _4337_ (.A(_0806_),
    .B(_0601_),
    .Y(_0807_));
 sg13g2_nor2_1 _4338_ (.A(net24),
    .B(_0797_),
    .Y(_0808_));
 sg13g2_nor2_1 _4339_ (.A(_0807_),
    .B(_0808_),
    .Y(_0809_));
 sg13g2_a22oi_1 _4340_ (.Y(_0810_),
    .B1(net73),
    .B2(_0809_),
    .A2(_0805_),
    .A1(net72));
 sg13g2_a21oi_1 _4341_ (.A1(_0796_),
    .A2(_0810_),
    .Y(_0811_),
    .B1(_0458_));
 sg13g2_nor3_1 _4342_ (.A(_0792_),
    .B(_0803_),
    .C(_0811_),
    .Y(_0812_));
 sg13g2_o21ai_1 _4343_ (.B1(_0279_),
    .Y(_0813_),
    .A1(_0200_),
    .A2(_0801_));
 sg13g2_a21oi_1 _4344_ (.A1(net75),
    .A2(_0793_),
    .Y(_0814_),
    .B1(_0232_));
 sg13g2_a21oi_1 _4345_ (.A1(_0813_),
    .A2(_0814_),
    .Y(_0815_),
    .B1(_2484_));
 sg13g2_nor2_1 _4346_ (.A(_0198_),
    .B(_0815_),
    .Y(_0816_));
 sg13g2_a21oi_1 _4347_ (.A1(_0812_),
    .A2(_0816_),
    .Y(_0817_),
    .B1(_2478_));
 sg13g2_nand2_1 _4348_ (.Y(_0818_),
    .A(_0781_),
    .B(_0817_));
 sg13g2_a21oi_1 _4349_ (.A1(_0660_),
    .A2(_0620_),
    .Y(_0819_),
    .B1(net77));
 sg13g2_nor2_1 _4350_ (.A(net112),
    .B(_0590_),
    .Y(_0820_));
 sg13g2_nor2_1 _4351_ (.A(_0819_),
    .B(_0820_),
    .Y(_0821_));
 sg13g2_nor2b_1 _4352_ (.A(_0631_),
    .B_N(_0206_),
    .Y(_0822_));
 sg13g2_o21ai_1 _4353_ (.B1(net92),
    .Y(_0823_),
    .A1(_0822_),
    .A2(_0623_));
 sg13g2_nor2_1 _4354_ (.A(net92),
    .B(_0216_),
    .Y(_0824_));
 sg13g2_a21oi_1 _4355_ (.A1(_0632_),
    .A2(_0824_),
    .Y(_0825_),
    .B1(net16));
 sg13g2_nand2_1 _4356_ (.Y(_0826_),
    .A(_0823_),
    .B(_0825_));
 sg13g2_nand2_1 _4357_ (.Y(_0827_),
    .A(_0826_),
    .B(net63));
 sg13g2_nor2_1 _4358_ (.A(_2481_),
    .B(_0339_),
    .Y(_0828_));
 sg13g2_inv_1 _4359_ (.Y(_0829_),
    .A(_0828_));
 sg13g2_a21oi_1 _4360_ (.A1(_0821_),
    .A2(_0827_),
    .Y(_0830_),
    .B1(_0829_));
 sg13g2_o21ai_1 _4361_ (.B1(net25),
    .Y(_0831_),
    .A1(_0431_),
    .A2(_0615_));
 sg13g2_nor2_1 _4362_ (.A(_0831_),
    .B(_0639_),
    .Y(_0832_));
 sg13g2_nor2_1 _4363_ (.A(net94),
    .B(_0832_),
    .Y(_0833_));
 sg13g2_a21oi_1 _4364_ (.A1(_0644_),
    .A2(_0647_),
    .Y(_0834_),
    .B1(net74));
 sg13g2_nand2_1 _4365_ (.Y(_0835_),
    .A(_0661_),
    .B(net90));
 sg13g2_nand2_1 _4366_ (.Y(_0836_),
    .A(_0666_),
    .B(net82));
 sg13g2_nand2_1 _4367_ (.Y(_0837_),
    .A(_0835_),
    .B(_0836_));
 sg13g2_nor3_1 _4368_ (.A(_0833_),
    .B(_0834_),
    .C(_0837_),
    .Y(_0838_));
 sg13g2_nor2_1 _4369_ (.A(net102),
    .B(_2771_),
    .Y(_0839_));
 sg13g2_nor2b_1 _4370_ (.A(_0838_),
    .B_N(_0839_),
    .Y(_0840_));
 sg13g2_nor3_1 _4371_ (.A(_2917_),
    .B(_0830_),
    .C(_0840_),
    .Y(_0841_));
 sg13g2_nand2_1 _4372_ (.Y(_0842_),
    .A(_0659_),
    .B(_0706_));
 sg13g2_nand3_1 _4373_ (.B(_0587_),
    .C(_2310_),
    .A(_0275_),
    .Y(_0843_));
 sg13g2_nand2_1 _4374_ (.Y(_0844_),
    .A(_0842_),
    .B(_0843_));
 sg13g2_nand2_1 _4375_ (.Y(_0845_),
    .A(_0844_),
    .B(_2931_));
 sg13g2_nand2b_1 _4376_ (.Y(_0846_),
    .B(net89),
    .A_N(_0646_));
 sg13g2_a21oi_1 _4377_ (.A1(_0238_),
    .A2(_0651_),
    .Y(_0847_),
    .B1(_0846_));
 sg13g2_nand2_1 _4378_ (.Y(_0848_),
    .A(_0665_),
    .B(_2847_));
 sg13g2_nor2b_1 _4379_ (.A(_2903_),
    .B_N(_0638_),
    .Y(_0849_));
 sg13g2_inv_1 _4380_ (.Y(_0850_),
    .A(_0642_));
 sg13g2_nand2_1 _4381_ (.Y(_0851_),
    .A(_0849_),
    .B(_0850_));
 sg13g2_nor2_1 _4382_ (.A(_0848_),
    .B(_0851_),
    .Y(_0852_));
 sg13g2_nor2_1 _4383_ (.A(_0847_),
    .B(_0852_),
    .Y(_0853_));
 sg13g2_nand2_1 _4384_ (.Y(_0854_),
    .A(_0845_),
    .B(_0853_));
 sg13g2_nand2_1 _4385_ (.Y(_0855_),
    .A(_0854_),
    .B(net78));
 sg13g2_nand2_1 _4386_ (.Y(_0856_),
    .A(_0270_),
    .B(_0638_));
 sg13g2_nand2_1 _4387_ (.Y(_0857_),
    .A(_0688_),
    .B(_0637_));
 sg13g2_nor2_1 _4388_ (.A(_0856_),
    .B(_0857_),
    .Y(_0858_));
 sg13g2_nand3_1 _4389_ (.B(_0275_),
    .C(_2303_),
    .A(_0769_),
    .Y(_0859_));
 sg13g2_nand2_1 _4390_ (.Y(_0860_),
    .A(_0859_),
    .B(_2861_));
 sg13g2_nor2_1 _4391_ (.A(_0858_),
    .B(_0860_),
    .Y(_0861_));
 sg13g2_nor2_1 _4392_ (.A(net78),
    .B(_0861_),
    .Y(_0862_));
 sg13g2_a21oi_1 _4393_ (.A1(_2804_),
    .A2(net22),
    .Y(_0863_),
    .B1(net88));
 sg13g2_nand3_1 _4394_ (.B(_0587_),
    .C(_0863_),
    .A(_0620_),
    .Y(_0864_));
 sg13g2_nand2b_1 _4395_ (.Y(_0865_),
    .B(_0624_),
    .A_N(_0616_));
 sg13g2_nand3_1 _4396_ (.B(_0865_),
    .C(_2931_),
    .A(_0864_),
    .Y(_0866_));
 sg13g2_nand2_1 _4397_ (.Y(_0867_),
    .A(_0862_),
    .B(_0866_));
 sg13g2_nand2_1 _4398_ (.Y(_0868_),
    .A(_0855_),
    .B(_0867_));
 sg13g2_nand2_1 _4399_ (.Y(_0869_),
    .A(_0868_),
    .B(net19));
 sg13g2_nand2_1 _4400_ (.Y(_0870_),
    .A(_0869_),
    .B(net102));
 sg13g2_nand2_1 _4401_ (.Y(_0871_),
    .A(_0841_),
    .B(_0870_));
 sg13g2_nor2_1 _4402_ (.A(net70),
    .B(_0594_),
    .Y(_0872_));
 sg13g2_a21oi_1 _4403_ (.A1(_0603_),
    .A2(net80),
    .Y(_0873_),
    .B1(_0872_));
 sg13g2_nand2_1 _4404_ (.Y(_0874_),
    .A(_0873_),
    .B(_0734_));
 sg13g2_nand2_1 _4405_ (.Y(_0875_),
    .A(_0729_),
    .B(_2917_));
 sg13g2_a21oi_1 _4406_ (.A1(_0874_),
    .A2(_0839_),
    .Y(_0876_),
    .B1(_0875_));
 sg13g2_nor2_1 _4407_ (.A(net65),
    .B(net45),
    .Y(_0877_));
 sg13g2_o21ai_1 _4408_ (.B1(net35),
    .Y(_0878_),
    .A1(_0877_),
    .A2(_2869_));
 sg13g2_o21ai_1 _4409_ (.B1(_0878_),
    .Y(_0879_),
    .A1(_2911_),
    .A2(_0649_));
 sg13g2_nand2_1 _4410_ (.Y(_0880_),
    .A(_0879_),
    .B(_0496_));
 sg13g2_nand2_1 _4411_ (.Y(_0881_),
    .A(_0584_),
    .B(net122));
 sg13g2_nand3_1 _4412_ (.B(_0660_),
    .C(_0881_),
    .A(_0880_),
    .Y(_0882_));
 sg13g2_nand2_1 _4413_ (.Y(_0883_),
    .A(_0882_),
    .B(net63));
 sg13g2_nor2_1 _4414_ (.A(_0392_),
    .B(net27),
    .Y(_0884_));
 sg13g2_and2_1 _4415_ (.A(_0625_),
    .B(_0884_),
    .X(_0885_));
 sg13g2_nor3_1 _4416_ (.A(_0885_),
    .B(_0732_),
    .C(_0733_),
    .Y(_0886_));
 sg13g2_nand2_1 _4417_ (.Y(_0887_),
    .A(_0883_),
    .B(_0886_));
 sg13g2_nor2_1 _4418_ (.A(_2482_),
    .B(_2771_),
    .Y(_0888_));
 sg13g2_nand2_1 _4419_ (.Y(_0889_),
    .A(_0887_),
    .B(_0888_));
 sg13g2_a21oi_1 _4420_ (.A1(_0876_),
    .A2(_0889_),
    .Y(_0890_),
    .B1(net71));
 sg13g2_nand2_1 _4421_ (.Y(_0891_),
    .A(_0871_),
    .B(_0890_));
 sg13g2_nor2_1 _4422_ (.A(net77),
    .B(_0782_),
    .Y(_0892_));
 sg13g2_nand2_1 _4423_ (.Y(_0893_),
    .A(_0653_),
    .B(net75));
 sg13g2_a21oi_1 _4424_ (.A1(_2894_),
    .A2(_2905_),
    .Y(_0894_),
    .B1(net70));
 sg13g2_nor3_1 _4425_ (.A(net102),
    .B(_0264_),
    .C(_0894_),
    .Y(_0895_));
 sg13g2_nand2_1 _4426_ (.Y(_0896_),
    .A(_0893_),
    .B(_0895_));
 sg13g2_nand3b_1 _4427_ (.B(_0548_),
    .C(_0715_),
    .Y(_0897_),
    .A_N(_0606_));
 sg13g2_nand2_1 _4428_ (.Y(_0898_),
    .A(_0897_),
    .B(net75));
 sg13g2_nor2_1 _4429_ (.A(net77),
    .B(_0431_),
    .Y(_0899_));
 sg13g2_nor3_1 _4430_ (.A(_2482_),
    .B(_0884_),
    .C(_0899_),
    .Y(_0900_));
 sg13g2_o21ai_1 _4431_ (.B1(net72),
    .Y(_0901_),
    .A1(_2870_),
    .A2(_2906_));
 sg13g2_nand4_1 _4432_ (.B(_0900_),
    .C(_0390_),
    .A(_0898_),
    .Y(_0902_),
    .D(_0901_));
 sg13g2_o21ai_1 _4433_ (.B1(_0902_),
    .Y(_0903_),
    .A1(_0892_),
    .A2(_0896_));
 sg13g2_nor3_1 _4434_ (.A(net24),
    .B(_0538_),
    .C(_0202_),
    .Y(_0904_));
 sg13g2_nor2_1 _4435_ (.A(net74),
    .B(_0904_),
    .Y(_0905_));
 sg13g2_o21ai_1 _4436_ (.B1(_0905_),
    .Y(_0906_),
    .A1(_2893_),
    .A2(_0788_));
 sg13g2_a21o_1 _4437_ (.A2(_0906_),
    .A1(_0903_),
    .B1(_0198_),
    .X(_0907_));
 sg13g2_nand2_1 _4438_ (.Y(_0908_),
    .A(_0891_),
    .B(_0907_));
 sg13g2_a21oi_1 _4439_ (.A1(_0908_),
    .A2(_2478_),
    .Y(_0909_),
    .B1(_0577_));
 sg13g2_nand2_2 _4440_ (.Y(_0910_),
    .A(_0818_),
    .B(_0909_));
 sg13g2_a21oi_1 _4441_ (.A1(_2826_),
    .A2(_0331_),
    .Y(_0911_),
    .B1(_0804_));
 sg13g2_nor2_1 _4442_ (.A(_2498_),
    .B(_0806_),
    .Y(_0912_));
 sg13g2_nor2_1 _4443_ (.A(net88),
    .B(_0912_),
    .Y(_0913_));
 sg13g2_a21oi_1 _4444_ (.A1(_0911_),
    .A2(net79),
    .Y(_0914_),
    .B1(_0913_));
 sg13g2_o21ai_1 _4445_ (.B1(net22),
    .Y(_0915_),
    .A1(_0536_),
    .A2(_0207_));
 sg13g2_nor2_1 _4446_ (.A(net23),
    .B(_2870_),
    .Y(_0916_));
 sg13g2_nand2_1 _4447_ (.Y(_0917_),
    .A(_0915_),
    .B(_0916_));
 sg13g2_nor2_1 _4448_ (.A(_0392_),
    .B(_0804_),
    .Y(_0918_));
 sg13g2_a21oi_1 _4449_ (.A1(_0917_),
    .A2(net83),
    .Y(_0919_),
    .B1(_0918_));
 sg13g2_o21ai_1 _4450_ (.B1(_0919_),
    .Y(_0920_),
    .A1(net61),
    .A2(_0914_));
 sg13g2_nand2_1 _4451_ (.Y(_0921_),
    .A(_0701_),
    .B(net42));
 sg13g2_nand2_1 _4452_ (.Y(_0922_),
    .A(_0921_),
    .B(net24));
 sg13g2_nand2_1 _4453_ (.Y(_0923_),
    .A(_0626_),
    .B(_0395_));
 sg13g2_nand2_1 _4454_ (.Y(_0924_),
    .A(_0922_),
    .B(_0923_));
 sg13g2_nor2_1 _4455_ (.A(net88),
    .B(_0924_),
    .Y(_0925_));
 sg13g2_nor2_1 _4456_ (.A(_2931_),
    .B(_0925_),
    .Y(_0926_));
 sg13g2_a21oi_1 _4457_ (.A1(_0697_),
    .A2(_2566_),
    .Y(_0927_),
    .B1(net23));
 sg13g2_nand3_1 _4458_ (.B(_0923_),
    .C(_0326_),
    .A(_0927_),
    .Y(_0928_));
 sg13g2_nand2_1 _4459_ (.Y(_0929_),
    .A(_0926_),
    .B(_0928_));
 sg13g2_inv_1 _4460_ (.Y(_0930_),
    .A(_0596_));
 sg13g2_a21oi_1 _4461_ (.A1(net28),
    .A2(_0930_),
    .Y(_0931_),
    .B1(_0284_));
 sg13g2_nor2_1 _4462_ (.A(_0214_),
    .B(_2442_),
    .Y(_0932_));
 sg13g2_inv_1 _4463_ (.Y(_0933_),
    .A(_0932_));
 sg13g2_a21oi_1 _4464_ (.A1(_0933_),
    .A2(net22),
    .Y(_0934_),
    .B1(net18));
 sg13g2_o21ai_1 _4465_ (.B1(_0934_),
    .Y(_0935_),
    .A1(_2568_),
    .A2(_0931_));
 sg13g2_a21oi_1 _4466_ (.A1(_0935_),
    .A2(net75),
    .Y(_0936_),
    .B1(_0918_));
 sg13g2_nand2_1 _4467_ (.Y(_0937_),
    .A(_0929_),
    .B(_0936_));
 sg13g2_a22oi_1 _4468_ (.Y(_0938_),
    .B1(_0839_),
    .B2(_0937_),
    .A2(_0828_),
    .A1(_0920_));
 sg13g2_nor3_1 _4469_ (.A(net16),
    .B(_0295_),
    .C(_0697_),
    .Y(_0939_));
 sg13g2_nand2b_1 _4470_ (.Y(_0940_),
    .B(_0926_),
    .A_N(_0939_));
 sg13g2_a21oi_1 _4471_ (.A1(_2894_),
    .A2(_0932_),
    .Y(_0941_),
    .B1(net94));
 sg13g2_nand2_1 _4472_ (.Y(_0942_),
    .A(_2868_),
    .B(_2825_));
 sg13g2_a21oi_1 _4473_ (.A1(_0923_),
    .A2(_0942_),
    .Y(_0943_),
    .B1(_0392_));
 sg13g2_nor3_1 _4474_ (.A(_2771_),
    .B(_0941_),
    .C(_0943_),
    .Y(_0944_));
 sg13g2_nand2_1 _4475_ (.Y(_0945_),
    .A(_0940_),
    .B(_0944_));
 sg13g2_a21oi_1 _4476_ (.A1(_2954_),
    .A2(_0930_),
    .Y(_0946_),
    .B1(_0284_));
 sg13g2_nand2_1 _4477_ (.Y(_0947_),
    .A(_0805_),
    .B(net88));
 sg13g2_a21oi_1 _4478_ (.A1(_0946_),
    .A2(_2826_),
    .Y(_0948_),
    .B1(_0947_));
 sg13g2_o21ai_1 _4479_ (.B1(net63),
    .Y(_0949_),
    .A1(_0913_),
    .A2(_0948_));
 sg13g2_nand2_1 _4480_ (.Y(_0950_),
    .A(_2853_),
    .B(_2819_));
 sg13g2_a21oi_1 _4481_ (.A1(_0482_),
    .A2(_0950_),
    .Y(_0951_),
    .B1(_2769_));
 sg13g2_nor3_1 _4482_ (.A(_0339_),
    .B(_0918_),
    .C(_0951_),
    .Y(_0952_));
 sg13g2_nand2_1 _4483_ (.Y(_0953_),
    .A(_0949_),
    .B(_0952_));
 sg13g2_nand3_1 _4484_ (.B(_0253_),
    .C(_0953_),
    .A(_0945_),
    .Y(_0954_));
 sg13g2_nand2_1 _4485_ (.Y(_0955_),
    .A(_0938_),
    .B(_0954_));
 sg13g2_nand2_1 _4486_ (.Y(_0956_),
    .A(_0955_),
    .B(_2777_));
 sg13g2_o21ai_1 _4487_ (.B1(_0273_),
    .Y(_0957_),
    .A1(_2443_),
    .A2(_2782_));
 sg13g2_nand2_1 _4488_ (.Y(_0958_),
    .A(_0957_),
    .B(_0916_));
 sg13g2_nand2_1 _4489_ (.Y(_0959_),
    .A(_0203_),
    .B(_2783_));
 sg13g2_nand2_1 _4490_ (.Y(_0960_),
    .A(_0959_),
    .B(net48));
 sg13g2_nand2_1 _4491_ (.Y(_0961_),
    .A(_0618_),
    .B(net22));
 sg13g2_nand3_1 _4492_ (.B(net25),
    .C(_0961_),
    .A(_0960_),
    .Y(_0962_));
 sg13g2_a22oi_1 _4493_ (.Y(_0963_),
    .B1(_2802_),
    .B2(_0962_),
    .A2(_0958_),
    .A1(_2813_));
 sg13g2_nand2_1 _4494_ (.Y(_0964_),
    .A(_2870_),
    .B(_2797_));
 sg13g2_nand2_1 _4495_ (.Y(_0965_),
    .A(_0942_),
    .B(_0964_));
 sg13g2_nor2_1 _4496_ (.A(_0276_),
    .B(_2871_),
    .Y(_0966_));
 sg13g2_o21ai_1 _4497_ (.B1(_2861_),
    .Y(_0967_),
    .A1(_0965_),
    .A2(_0966_));
 sg13g2_nand2_1 _4498_ (.Y(_0968_),
    .A(_0963_),
    .B(_0967_));
 sg13g2_nor2_1 _4499_ (.A(_2831_),
    .B(_0494_),
    .Y(_0969_));
 sg13g2_a221oi_1 _4500_ (.B2(net82),
    .C1(_0264_),
    .B1(_2858_),
    .A1(net89),
    .Y(_0970_),
    .A2(_0969_));
 sg13g2_nand2b_1 _4501_ (.Y(_0971_),
    .B(_0198_),
    .A_N(_0970_));
 sg13g2_a21oi_1 _4502_ (.A1(_0968_),
    .A2(_2779_),
    .Y(_0972_),
    .B1(_0971_));
 sg13g2_nand2_1 _4503_ (.Y(_0973_),
    .A(_0956_),
    .B(_0972_));
 sg13g2_nand2_1 _4504_ (.Y(_0974_),
    .A(_0243_),
    .B(_0587_));
 sg13g2_nor2_1 _4505_ (.A(_0407_),
    .B(_0599_),
    .Y(_0975_));
 sg13g2_a21oi_1 _4506_ (.A1(_0975_),
    .A2(net102),
    .Y(_0976_),
    .B1(_0277_));
 sg13g2_o21ai_1 _4507_ (.B1(_0976_),
    .Y(_0977_),
    .A1(net102),
    .A2(_0974_));
 sg13g2_nand2_1 _4508_ (.Y(_0978_),
    .A(_0969_),
    .B(net22));
 sg13g2_nand3_1 _4509_ (.B(_0197_),
    .C(_2866_),
    .A(_0550_),
    .Y(_0979_));
 sg13g2_a21oi_1 _4510_ (.A1(_0978_),
    .A2(_0277_),
    .Y(_0980_),
    .B1(_0979_));
 sg13g2_a21oi_1 _4511_ (.A1(_0977_),
    .A2(_0980_),
    .Y(_0981_),
    .B1(_0559_));
 sg13g2_a21oi_1 _4512_ (.A1(_0973_),
    .A2(_0981_),
    .Y(_0982_),
    .B1(_0577_));
 sg13g2_a21oi_1 _4513_ (.A1(_0596_),
    .A2(net26),
    .Y(_0983_),
    .B1(_0273_));
 sg13g2_nand2b_1 _4514_ (.Y(_0984_),
    .B(_0983_),
    .A_N(_0431_));
 sg13g2_nand2_1 _4515_ (.Y(_0985_),
    .A(_0984_),
    .B(_0934_));
 sg13g2_nor2_1 _4516_ (.A(net35),
    .B(net31),
    .Y(_0986_));
 sg13g2_o21ai_1 _4517_ (.B1(net39),
    .Y(_0987_),
    .A1(_0538_),
    .A2(_0986_));
 sg13g2_nand2_1 _4518_ (.Y(_0988_),
    .A(_0987_),
    .B(_0927_));
 sg13g2_a22oi_1 _4519_ (.Y(_0989_),
    .B1(_0360_),
    .B2(_0988_),
    .A2(_2802_),
    .A1(_0985_));
 sg13g2_nand2_1 _4520_ (.Y(_0990_),
    .A(_0922_),
    .B(_0987_));
 sg13g2_nand2_1 _4521_ (.Y(_0991_),
    .A(_0990_),
    .B(_0341_));
 sg13g2_nand3b_1 _4522_ (.B(_0989_),
    .C(_0991_),
    .Y(_0992_),
    .A_N(_0918_));
 sg13g2_a22oi_1 _4523_ (.Y(_0993_),
    .B1(_2921_),
    .B2(_0992_),
    .A2(_2919_),
    .A1(_0920_));
 sg13g2_nand2_1 _4524_ (.Y(_0994_),
    .A(_0972_),
    .B(_0993_));
 sg13g2_o21ai_1 _4525_ (.B1(net79),
    .Y(_0995_),
    .A1(_0407_),
    .A2(_0599_));
 sg13g2_a21oi_1 _4526_ (.A1(_0995_),
    .A2(_0980_),
    .Y(_0996_),
    .B1(_2479_));
 sg13g2_nand2_1 _4527_ (.Y(_0997_),
    .A(_0994_),
    .B(_0996_));
 sg13g2_a22oi_1 _4528_ (.Y(_0998_),
    .B1(net89),
    .B2(_0917_),
    .A2(_2813_),
    .A1(_0965_));
 sg13g2_a21oi_1 _4529_ (.A1(net83),
    .A2(_0958_),
    .Y(_0999_),
    .B1(_2872_));
 sg13g2_a21oi_1 _4530_ (.A1(_0998_),
    .A2(_0999_),
    .Y(_1000_),
    .B1(_2780_));
 sg13g2_inv_1 _4531_ (.Y(_1001_),
    .A(_0969_));
 sg13g2_a21oi_1 _4532_ (.A1(_2848_),
    .A2(_1001_),
    .Y(_1002_),
    .B1(_2862_));
 sg13g2_nand2_1 _4533_ (.Y(_1003_),
    .A(_0962_),
    .B(net80));
 sg13g2_a21oi_1 _4534_ (.A1(_1002_),
    .A2(_1003_),
    .Y(_1004_),
    .B1(_0264_));
 sg13g2_nor3_1 _4535_ (.A(_0251_),
    .B(_1000_),
    .C(_1004_),
    .Y(_1005_));
 sg13g2_nand2_1 _4536_ (.Y(_1006_),
    .A(_0805_),
    .B(net83));
 sg13g2_o21ai_1 _4537_ (.B1(_1006_),
    .Y(_1007_),
    .A1(_0392_),
    .A2(_0912_));
 sg13g2_a21oi_1 _4538_ (.A1(_2848_),
    .A2(_0911_),
    .Y(_1008_),
    .B1(_1007_));
 sg13g2_nand2_1 _4539_ (.Y(_1009_),
    .A(_0985_),
    .B(_0227_));
 sg13g2_nand2_1 _4540_ (.Y(_1010_),
    .A(_1008_),
    .B(_1009_));
 sg13g2_nand2_1 _4541_ (.Y(_1011_),
    .A(_0978_),
    .B(net89));
 sg13g2_nand2_1 _4542_ (.Y(_1012_),
    .A(_1011_),
    .B(_1006_));
 sg13g2_a22oi_1 _4543_ (.Y(_1013_),
    .B1(_0502_),
    .B2(_0990_),
    .A2(_0341_),
    .A1(_0988_));
 sg13g2_nand2b_1 _4544_ (.Y(_1014_),
    .B(_1013_),
    .A_N(_1012_));
 sg13g2_a22oi_1 _4545_ (.Y(_1015_),
    .B1(_2921_),
    .B2(_1014_),
    .A2(_2919_),
    .A1(_1010_));
 sg13g2_nand2_1 _4546_ (.Y(_1016_),
    .A(_1005_),
    .B(_1015_));
 sg13g2_nor2_1 _4547_ (.A(_0200_),
    .B(_0979_),
    .Y(_1017_));
 sg13g2_a21oi_1 _4548_ (.A1(_0975_),
    .A2(_1017_),
    .Y(_1018_),
    .B1(_2484_));
 sg13g2_nand2_1 _4549_ (.Y(_1019_),
    .A(_1016_),
    .B(_1018_));
 sg13g2_a21oi_1 _4550_ (.A1(_0924_),
    .A2(net90),
    .Y(_1020_),
    .B1(_1012_));
 sg13g2_a21o_1 _4551_ (.A2(_0923_),
    .A1(_0927_),
    .B1(_0263_),
    .X(_1021_));
 sg13g2_nand2_1 _4552_ (.Y(_1022_),
    .A(_1020_),
    .B(_1021_));
 sg13g2_nand2_1 _4553_ (.Y(_1023_),
    .A(_0935_),
    .B(_0227_));
 sg13g2_nand2_1 _4554_ (.Y(_1024_),
    .A(_1008_),
    .B(_1023_));
 sg13g2_a22oi_1 _4555_ (.Y(_1025_),
    .B1(_2919_),
    .B2(_1024_),
    .A2(_2921_),
    .A1(_1022_));
 sg13g2_nand2_1 _4556_ (.Y(_1026_),
    .A(_1005_),
    .B(_1025_));
 sg13g2_nor2b_1 _4557_ (.A(_0974_),
    .B_N(_1017_),
    .Y(_1027_));
 sg13g2_nor2_1 _4558_ (.A(_0417_),
    .B(_1027_),
    .Y(_1028_));
 sg13g2_nand2_1 _4559_ (.Y(_1029_),
    .A(_1026_),
    .B(_1028_));
 sg13g2_nand3_1 _4560_ (.B(_1019_),
    .C(_1029_),
    .A(_0997_),
    .Y(_1030_));
 sg13g2_nand2_1 _4561_ (.Y(_1031_),
    .A(_1030_),
    .B(_0559_));
 sg13g2_nand2_1 _4562_ (.Y(_1032_),
    .A(_0982_),
    .B(_1031_));
 sg13g2_buf_2 _4563_ (.A(_1032_),
    .X(_1033_));
 sg13g2_nand2_1 _4564_ (.Y(_1034_),
    .A(_0910_),
    .B(_1033_));
 sg13g2_nor2_1 _4565_ (.A(_0579_),
    .B(_1034_),
    .Y(_1035_));
 sg13g2_nor2_1 _4566_ (.A(_2582_),
    .B(_2598_),
    .Y(_1036_));
 sg13g2_inv_1 _4567_ (.Y(_1037_),
    .A(_1036_));
 sg13g2_nor3_1 _4568_ (.A(_2559_),
    .B(_2431_),
    .C(_2583_),
    .Y(_1038_));
 sg13g2_nand3_1 _4569_ (.B(_2390_),
    .C(net113),
    .A(net116),
    .Y(_1039_));
 sg13g2_inv_1 _4570_ (.Y(_1040_),
    .A(_2598_));
 sg13g2_nand2_1 _4571_ (.Y(_1041_),
    .A(net117),
    .B(net113));
 sg13g2_nand4_1 _4572_ (.B(_1039_),
    .C(_1040_),
    .A(_1038_),
    .Y(_1042_),
    .D(_1041_));
 sg13g2_a21oi_1 _4573_ (.A1(_1037_),
    .A2(_1042_),
    .Y(_1043_),
    .B1(_0574_));
 sg13g2_o21ai_1 _4574_ (.B1(_0251_),
    .Y(_1044_),
    .A1(_0265_),
    .A2(_0551_));
 sg13g2_and2_1 _4575_ (.A(_1043_),
    .B(_1044_),
    .X(_1045_));
 sg13g2_nand2_1 _4576_ (.Y(_1046_),
    .A(_1035_),
    .B(_1045_));
 sg13g2_buf_8 _4577_ (.A(_1046_),
    .X(_1047_));
 sg13g2_buf_1 _4578_ (.A(\frame_count[0] ),
    .X(_1048_));
 sg13g2_xnor2_1 _4579_ (.Y(_1049_),
    .A(_2423_),
    .B(_1048_));
 sg13g2_inv_1 _4580_ (.Y(_1050_),
    .A(_2764_));
 sg13g2_nor2_1 _4581_ (.A(_1049_),
    .B(_1050_),
    .Y(_1051_));
 sg13g2_a22oi_1 _4582_ (.Y(_1052_),
    .B1(_1047_),
    .B2(_1051_),
    .A2(_2767_),
    .A1(_2764_));
 sg13g2_inv_2 _4583_ (.Y(_1053_),
    .A(_0910_));
 sg13g2_nand2_1 _4584_ (.Y(_1054_),
    .A(_0579_),
    .B(_1053_));
 sg13g2_inv_1 _4585_ (.Y(_1055_),
    .A(_1054_));
 sg13g2_nand2_1 _4586_ (.Y(_1056_),
    .A(_1055_),
    .B(_1033_));
 sg13g2_xor2_1 _4587_ (.B(\frame_count[4] ),
    .A(_2431_),
    .X(_1057_));
 sg13g2_inv_1 _4588_ (.Y(_1058_),
    .A(\frame_count[3] ));
 sg13g2_inv_1 _4589_ (.Y(_1059_),
    .A(net117));
 sg13g2_inv_1 _4590_ (.Y(_1060_),
    .A(\frame_count[2] ));
 sg13g2_nand2_1 _4591_ (.Y(_1061_),
    .A(_2390_),
    .B(_1048_));
 sg13g2_buf_1 _4592_ (.A(\frame_count[1] ),
    .X(_1062_));
 sg13g2_xnor2_1 _4593_ (.Y(_1063_),
    .A(net116),
    .B(_1062_));
 sg13g2_nand2_1 _4594_ (.Y(_1064_),
    .A(net116),
    .B(_1062_));
 sg13g2_o21ai_1 _4595_ (.B1(_1064_),
    .Y(_1065_),
    .A1(_1061_),
    .A2(_1063_));
 sg13g2_xor2_1 _4596_ (.B(\frame_count[2] ),
    .A(net117),
    .X(_1066_));
 sg13g2_nand2_1 _4597_ (.Y(_1067_),
    .A(_1065_),
    .B(_1066_));
 sg13g2_o21ai_1 _4598_ (.B1(_1067_),
    .Y(_1068_),
    .A1(_1059_),
    .A2(_1060_));
 sg13g2_xor2_1 _4599_ (.B(\frame_count[3] ),
    .A(net113),
    .X(_1069_));
 sg13g2_nand2_1 _4600_ (.Y(_1070_),
    .A(_1068_),
    .B(_1069_));
 sg13g2_o21ai_1 _4601_ (.B1(_1070_),
    .Y(_1071_),
    .A1(_2433_),
    .A2(_1058_));
 sg13g2_xnor2_1 _4602_ (.Y(_1072_),
    .A(_1057_),
    .B(_1071_));
 sg13g2_nand2_1 _4603_ (.Y(_1073_),
    .A(_1072_),
    .B(net79));
 sg13g2_nor2_1 _4604_ (.A(net122),
    .B(_1073_),
    .Y(_1074_));
 sg13g2_nor2_1 _4605_ (.A(net105),
    .B(_1074_),
    .Y(_1075_));
 sg13g2_inv_1 _4606_ (.Y(_1076_),
    .A(_1075_));
 sg13g2_nand2_1 _4607_ (.Y(_1077_),
    .A(_1074_),
    .B(net105));
 sg13g2_nand2_1 _4608_ (.Y(_1078_),
    .A(_1076_),
    .B(_1077_));
 sg13g2_inv_1 _4609_ (.Y(_1079_),
    .A(_1078_));
 sg13g2_inv_1 _4610_ (.Y(_1080_),
    .A(_0040_));
 sg13g2_xnor2_1 _4611_ (.Y(_1081_),
    .A(_1080_),
    .B(_1075_));
 sg13g2_xor2_1 _4612_ (.B(_1073_),
    .A(_0039_),
    .X(_1082_));
 sg13g2_inv_1 _4613_ (.Y(_1083_),
    .A(_1082_));
 sg13g2_nand2_1 _4614_ (.Y(_1084_),
    .A(_1081_),
    .B(_1083_));
 sg13g2_nor2_1 _4615_ (.A(_1079_),
    .B(_1084_),
    .Y(_1085_));
 sg13g2_nor2_1 _4616_ (.A(_1085_),
    .B(_1047_),
    .Y(_1086_));
 sg13g2_a21oi_1 _4617_ (.A1(_1047_),
    .A2(_1056_),
    .Y(_1087_),
    .B1(_1086_));
 sg13g2_nor2b_1 _4618_ (.A(_1052_),
    .B_N(_1087_),
    .Y(_1088_));
 sg13g2_inv_1 _4619_ (.Y(_1089_),
    .A(_1033_));
 sg13g2_inv_1 _4620_ (.Y(_1090_),
    .A(\line_lfsr[4] ));
 sg13g2_buf_1 _4621_ (.A(\frame_count[5] ),
    .X(_1091_));
 sg13g2_xor2_1 _4622_ (.B(_1091_),
    .A(_2559_),
    .X(_1092_));
 sg13g2_inv_1 _4623_ (.Y(_1093_),
    .A(\frame_count[4] ));
 sg13g2_nand2_1 _4624_ (.Y(_1094_),
    .A(_1071_),
    .B(_1057_));
 sg13g2_o21ai_1 _4625_ (.B1(_1094_),
    .Y(_1095_),
    .A1(_2434_),
    .A2(_1093_));
 sg13g2_xor2_1 _4626_ (.B(_1095_),
    .A(_1092_),
    .X(_1096_));
 sg13g2_nor2_1 _4627_ (.A(_1090_),
    .B(_1096_),
    .Y(_1097_));
 sg13g2_nor2b_1 _4628_ (.A(\line_lfsr[4] ),
    .B_N(_1096_),
    .Y(_1098_));
 sg13g2_inv_1 _4629_ (.Y(_1099_),
    .A(\line_lfsr[5] ));
 sg13g2_nor2_1 _4630_ (.A(_2582_),
    .B(\frame_count[6] ),
    .Y(_1100_));
 sg13g2_nand2_1 _4631_ (.Y(_1101_),
    .A(_2582_),
    .B(\frame_count[6] ));
 sg13g2_nor2b_1 _4632_ (.A(_1100_),
    .B_N(_1101_),
    .Y(_1102_));
 sg13g2_and2_1 _4633_ (.A(_1095_),
    .B(_1092_),
    .X(_1103_));
 sg13g2_a21oi_1 _4634_ (.A1(_2559_),
    .A2(_1091_),
    .Y(_1104_),
    .B1(_1103_));
 sg13g2_xnor2_1 _4635_ (.Y(_1105_),
    .A(_1102_),
    .B(_1104_));
 sg13g2_nor2_1 _4636_ (.A(_1099_),
    .B(_1105_),
    .Y(_1106_));
 sg13g2_nor2b_1 _4637_ (.A(\line_lfsr[5] ),
    .B_N(_1105_),
    .Y(_1107_));
 sg13g2_nor4_1 _4638_ (.A(_1097_),
    .B(_1098_),
    .C(_1106_),
    .D(_1107_),
    .Y(_1108_));
 sg13g2_inv_1 _4639_ (.Y(_1109_),
    .A(\line_lfsr[6] ));
 sg13g2_xor2_1 _4640_ (.B(\frame_count[7] ),
    .A(_2598_),
    .X(_1110_));
 sg13g2_o21ai_1 _4641_ (.B1(_1101_),
    .Y(_1111_),
    .A1(_1100_),
    .A2(_1104_));
 sg13g2_xnor2_1 _4642_ (.Y(_1112_),
    .A(_1110_),
    .B(_1111_));
 sg13g2_xnor2_1 _4643_ (.Y(_1113_),
    .A(_1109_),
    .B(_1112_));
 sg13g2_inv_1 _4644_ (.Y(_1114_),
    .A(\line_lfsr[1] ));
 sg13g2_xnor2_1 _4645_ (.Y(_1115_),
    .A(_1066_),
    .B(_1065_));
 sg13g2_xnor2_1 _4646_ (.Y(_1116_),
    .A(_1114_),
    .B(_1115_));
 sg13g2_inv_1 _4647_ (.Y(_1117_),
    .A(\line_lfsr[0] ));
 sg13g2_xnor2_1 _4648_ (.Y(_1118_),
    .A(_1061_),
    .B(_1063_));
 sg13g2_xnor2_1 _4649_ (.Y(_1119_),
    .A(_1117_),
    .B(_1118_));
 sg13g2_nand2_1 _4650_ (.Y(_1120_),
    .A(_1116_),
    .B(_1119_));
 sg13g2_xnor2_1 _4651_ (.Y(_1121_),
    .A(_1069_),
    .B(_1068_));
 sg13g2_xnor2_1 _4652_ (.Y(_1122_),
    .A(\line_lfsr[2] ),
    .B(_1121_));
 sg13g2_nor2_1 _4653_ (.A(\line_lfsr[3] ),
    .B(_1072_),
    .Y(_1123_));
 sg13g2_inv_1 _4654_ (.Y(_1124_),
    .A(\line_lfsr[3] ));
 sg13g2_nor2b_1 _4655_ (.A(_1124_),
    .B_N(_1072_),
    .Y(_1125_));
 sg13g2_nor4_1 _4656_ (.A(_1120_),
    .B(_1122_),
    .C(_1123_),
    .D(_1125_),
    .Y(_1126_));
 sg13g2_nand3_1 _4657_ (.B(_1113_),
    .C(_1126_),
    .A(_1108_),
    .Y(_1127_));
 sg13g2_inv_1 _4658_ (.Y(_1128_),
    .A(_1127_));
 sg13g2_o21ai_1 _4659_ (.B1(_1035_),
    .Y(_1129_),
    .A1(_1045_),
    .A2(_1128_));
 sg13g2_buf_8 _4660_ (.A(_1129_),
    .X(_1130_));
 sg13g2_nand2_1 _4661_ (.Y(_1131_),
    .A(_1130_),
    .B(_0910_));
 sg13g2_nand2_1 _4662_ (.Y(_1132_),
    .A(_1079_),
    .B(_1083_));
 sg13g2_nor2_1 _4663_ (.A(_1082_),
    .B(_1079_),
    .Y(_1133_));
 sg13g2_nor2_1 _4664_ (.A(_1081_),
    .B(_1133_),
    .Y(_1134_));
 sg13g2_inv_4 _4665_ (.A(_1047_),
    .Y(_1135_));
 sg13g2_nand2b_1 _4666_ (.Y(_1136_),
    .B(_1135_),
    .A_N(_1134_));
 sg13g2_nand2_1 _4667_ (.Y(_1137_),
    .A(_1136_),
    .B(_2762_));
 sg13g2_o21ai_1 _4668_ (.B1(_1137_),
    .Y(_1138_),
    .A1(_2763_),
    .A2(_1132_));
 sg13g2_o21ai_1 _4669_ (.B1(_1138_),
    .Y(_1139_),
    .A1(_1089_),
    .A2(_1131_));
 sg13g2_inv_1 _4670_ (.Y(_1140_),
    .A(_2738_));
 sg13g2_nand2_1 _4671_ (.Y(_1141_),
    .A(_1139_),
    .B(_1140_));
 sg13g2_a21oi_1 _4672_ (.A1(_2583_),
    .A2(_0038_),
    .Y(_1142_),
    .B1(_1040_));
 sg13g2_nor3_2 _4673_ (.A(_2651_),
    .B(_1142_),
    .C(_2722_),
    .Y(_1143_));
 sg13g2_o21ai_1 _4674_ (.B1(_1143_),
    .Y(_1144_),
    .A1(_1088_),
    .A2(_1141_));
 sg13g2_nand2_1 _4675_ (.Y(_1145_),
    .A(_1141_),
    .B(_1088_));
 sg13g2_nor2b_1 _4676_ (.A(_1144_),
    .B_N(_1145_),
    .Y(_0004_));
 sg13g2_o21ai_1 _4677_ (.B1(_0559_),
    .Y(_1146_),
    .A1(_0255_),
    .A2(_0461_));
 sg13g2_nand2_1 _4678_ (.Y(_1147_),
    .A(_1146_),
    .B(_0578_));
 sg13g2_a21oi_1 _4679_ (.A1(_1131_),
    .A2(_1147_),
    .Y(_1148_),
    .B1(_1089_));
 sg13g2_nor2_1 _4680_ (.A(_1137_),
    .B(_1148_),
    .Y(_1149_));
 sg13g2_nor2_1 _4681_ (.A(_2738_),
    .B(_1149_),
    .Y(_1150_));
 sg13g2_inv_1 _4682_ (.Y(_1151_),
    .A(_1143_));
 sg13g2_a21oi_1 _4683_ (.A1(_1145_),
    .A2(_1150_),
    .Y(_0005_),
    .B1(_1151_));
 sg13g2_nand2_1 _4684_ (.Y(_1152_),
    .A(_1147_),
    .B(_0910_));
 sg13g2_nand2_1 _4685_ (.Y(_1153_),
    .A(_1152_),
    .B(_1054_));
 sg13g2_nand2_1 _4686_ (.Y(_1154_),
    .A(_1153_),
    .B(_1089_));
 sg13g2_nand3_1 _4687_ (.B(_1033_),
    .C(_0910_),
    .A(_0579_),
    .Y(_1155_));
 sg13g2_nand3_1 _4688_ (.B(_1130_),
    .C(_1155_),
    .A(_1154_),
    .Y(_1156_));
 sg13g2_a21oi_1 _4689_ (.A1(_1072_),
    .A2(net79),
    .Y(_1157_),
    .B1(net93));
 sg13g2_inv_1 _4690_ (.Y(_1158_),
    .A(_1081_));
 sg13g2_o21ai_1 _4691_ (.B1(_1158_),
    .Y(_1159_),
    .A1(_1074_),
    .A2(_1157_));
 sg13g2_nand2_1 _4692_ (.Y(_1160_),
    .A(_1086_),
    .B(_1159_));
 sg13g2_nand2_1 _4693_ (.Y(_1161_),
    .A(_1156_),
    .B(_1160_));
 sg13g2_nand2_1 _4694_ (.Y(_1162_),
    .A(_1161_),
    .B(_2764_));
 sg13g2_nand2_1 _4695_ (.Y(_1163_),
    .A(_1159_),
    .B(_1084_));
 sg13g2_inv_1 _4696_ (.Y(_1164_),
    .A(_1051_));
 sg13g2_a21oi_1 _4697_ (.A1(_1135_),
    .A2(_1163_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_a21oi_1 _4698_ (.A1(_1053_),
    .A2(_1033_),
    .Y(_1166_),
    .B1(_1147_));
 sg13g2_nor3_1 _4699_ (.A(_1127_),
    .B(_0579_),
    .C(_1034_),
    .Y(_1167_));
 sg13g2_o21ai_1 _4700_ (.B1(_1047_),
    .Y(_1168_),
    .A1(_1166_),
    .A2(_1167_));
 sg13g2_nand3_1 _4701_ (.B(_1168_),
    .C(_2767_),
    .A(_1165_),
    .Y(_1169_));
 sg13g2_nand2_1 _4702_ (.Y(_1170_),
    .A(_1162_),
    .B(_1169_));
 sg13g2_nand2_1 _4703_ (.Y(_1171_),
    .A(_1165_),
    .B(_1168_));
 sg13g2_nand2_1 _4704_ (.Y(_1172_),
    .A(_1171_),
    .B(_2766_));
 sg13g2_inv_1 _4705_ (.Y(_1173_),
    .A(_1131_));
 sg13g2_xnor2_1 _4706_ (.Y(_1174_),
    .A(_1080_),
    .B(_1077_));
 sg13g2_o21ai_1 _4707_ (.B1(_2762_),
    .Y(_1175_),
    .A1(_1174_),
    .A2(_1047_));
 sg13g2_o21ai_1 _4708_ (.B1(_1140_),
    .Y(_1176_),
    .A1(_1173_),
    .A2(_1175_));
 sg13g2_a21oi_1 _4709_ (.A1(_1170_),
    .A2(_1172_),
    .Y(_1177_),
    .B1(_1176_));
 sg13g2_nand3_1 _4710_ (.B(_1176_),
    .C(_1172_),
    .A(_1170_),
    .Y(_1178_));
 sg13g2_nand2_1 _4711_ (.Y(_1179_),
    .A(_1178_),
    .B(_1143_));
 sg13g2_nor2_1 _4712_ (.A(_1177_),
    .B(_1179_),
    .Y(_0002_));
 sg13g2_a21oi_1 _4713_ (.A1(_1154_),
    .A2(_1130_),
    .Y(_1180_),
    .B1(_2763_));
 sg13g2_nor2_1 _4714_ (.A(_1083_),
    .B(_1078_),
    .Y(_1181_));
 sg13g2_inv_1 _4715_ (.Y(_1182_),
    .A(_1181_));
 sg13g2_o21ai_1 _4716_ (.B1(_1086_),
    .Y(_1183_),
    .A1(_1081_),
    .A2(_1182_));
 sg13g2_nand2_1 _4717_ (.Y(_1184_),
    .A(_1180_),
    .B(_1183_));
 sg13g2_nand2_1 _4718_ (.Y(_1185_),
    .A(_1184_),
    .B(_1140_));
 sg13g2_inv_1 _4719_ (.Y(_1186_),
    .A(_1185_));
 sg13g2_nand2_1 _4720_ (.Y(_1187_),
    .A(_1178_),
    .B(_1186_));
 sg13g2_nand2_1 _4721_ (.Y(_1188_),
    .A(_1187_),
    .B(_1143_));
 sg13g2_nand4_1 _4722_ (.B(_1185_),
    .C(_1176_),
    .A(_1170_),
    .Y(_1189_),
    .D(_1172_));
 sg13g2_nor2b_1 _4723_ (.A(_1188_),
    .B_N(_1189_),
    .Y(_0003_));
 sg13g2_o21ai_1 _4724_ (.B1(_1135_),
    .Y(_1190_),
    .A1(_1134_),
    .A2(_1085_));
 sg13g2_nand3_1 _4725_ (.B(_2762_),
    .C(_1155_),
    .A(_1190_),
    .Y(_1191_));
 sg13g2_nor2_1 _4726_ (.A(_1181_),
    .B(_1158_),
    .Y(_1192_));
 sg13g2_xnor2_1 _4727_ (.Y(_1193_),
    .A(_1033_),
    .B(_1054_));
 sg13g2_nand2_1 _4728_ (.Y(_1194_),
    .A(_1193_),
    .B(_1152_));
 sg13g2_nand2_1 _4729_ (.Y(_1195_),
    .A(_1194_),
    .B(_1130_));
 sg13g2_o21ai_1 _4730_ (.B1(_1195_),
    .Y(_1196_),
    .A1(_1136_),
    .A2(_1192_));
 sg13g2_o21ai_1 _4731_ (.B1(_2766_),
    .Y(_1197_),
    .A1(_1164_),
    .A2(_1193_));
 sg13g2_nand3_1 _4732_ (.B(_2764_),
    .C(_1197_),
    .A(_1196_),
    .Y(_1198_));
 sg13g2_nand2_1 _4733_ (.Y(_1199_),
    .A(_1198_),
    .B(_1143_));
 sg13g2_a21oi_1 _4734_ (.A1(_1140_),
    .A2(_1191_),
    .Y(_0000_),
    .B1(_1199_));
 sg13g2_nor2_1 _4735_ (.A(_1033_),
    .B(_1055_),
    .Y(_1200_));
 sg13g2_inv_1 _4736_ (.Y(_1201_),
    .A(_1133_));
 sg13g2_a21oi_1 _4737_ (.A1(_1201_),
    .A2(_1192_),
    .Y(_1202_),
    .B1(_1047_));
 sg13g2_nor4_1 _4738_ (.A(_2763_),
    .B(_1200_),
    .C(_1202_),
    .D(_1148_),
    .Y(_1203_));
 sg13g2_nor2_1 _4739_ (.A(_2738_),
    .B(_1203_),
    .Y(_1204_));
 sg13g2_a21oi_1 _4740_ (.A1(_1204_),
    .A2(_1198_),
    .Y(_0001_),
    .B1(_1151_));
 sg13g2_inv_1 _4741_ (.Y(_1205_),
    .A(_2328_));
 sg13g2_nor3_1 _4742_ (.A(_2315_),
    .B(_1205_),
    .C(net79),
    .Y(_1206_));
 sg13g2_nand4_1 _4743_ (.B(_1206_),
    .C(net93),
    .A(_2722_),
    .Y(_0007_),
    .D(_2716_));
 sg13g2_nor3_1 _4744_ (.A(_2582_),
    .B(_2561_),
    .C(_1040_),
    .Y(_1207_));
 sg13g2_nor2_1 _4745_ (.A(net117),
    .B(net113),
    .Y(_1208_));
 sg13g2_nand2_1 _4746_ (.Y(_1209_),
    .A(_1208_),
    .B(_2434_));
 sg13g2_nand3_1 _4747_ (.B(net113),
    .C(_2431_),
    .A(net117),
    .Y(_1210_));
 sg13g2_nand3_1 _4748_ (.B(_1209_),
    .C(_1210_),
    .A(_1207_),
    .Y(_0006_));
 sg13g2_buf_1 _4749_ (.A(\audio_sample_lpf[0] ),
    .X(_1211_));
 sg13g2_inv_1 _4750_ (.Y(_1212_),
    .A(_1211_));
 sg13g2_inv_1 _4751_ (.Y(_1213_),
    .A(net130));
 sg13g2_nor2_1 _4752_ (.A(_2388_),
    .B(_2423_),
    .Y(_1214_));
 sg13g2_nand4_1 _4753_ (.B(_1214_),
    .C(_2561_),
    .A(_1208_),
    .Y(_1215_),
    .D(_2434_));
 sg13g2_nor4_1 _4754_ (.A(net116),
    .B(_2390_),
    .C(_1037_),
    .D(_1215_),
    .Y(_1216_));
 sg13g2_buf_2 _4755_ (.A(_1216_),
    .X(_1217_));
 sg13g2_inv_1 _4756_ (.Y(_1218_),
    .A(_1217_));
 sg13g2_nor2_1 _4757_ (.A(_1213_),
    .B(_1218_),
    .Y(_1219_));
 sg13g2_buf_1 _4758_ (.A(_1219_),
    .X(_1220_));
 sg13g2_buf_1 _4759_ (.A(net62),
    .X(_1221_));
 sg13g2_buf_1 _4760_ (.A(\audio_sample_lpf[3] ),
    .X(_1222_));
 sg13g2_nor2_1 _4761_ (.A(net119),
    .B(net120),
    .Y(_1223_));
 sg13g2_inv_1 _4762_ (.Y(_1224_),
    .A(_2337_));
 sg13g2_nand2_1 _4763_ (.Y(_1225_),
    .A(_1223_),
    .B(_1224_));
 sg13g2_nor2_1 _4764_ (.A(net118),
    .B(_1225_),
    .Y(_1226_));
 sg13g2_inv_1 _4765_ (.Y(_1227_),
    .A(_1226_));
 sg13g2_xor2_1 _4766_ (.B(_2304_),
    .A(net121),
    .X(_1228_));
 sg13g2_nand2_1 _4767_ (.Y(_1229_),
    .A(_1228_),
    .B(net97));
 sg13g2_nand2_2 _4768_ (.Y(_1230_),
    .A(_2625_),
    .B(_2614_));
 sg13g2_inv_1 _4769_ (.Y(_1231_),
    .A(_1230_));
 sg13g2_nand2_2 _4770_ (.Y(_1232_),
    .A(net121),
    .B(_2307_));
 sg13g2_nand2_2 _4771_ (.Y(_1233_),
    .A(_1232_),
    .B(net104));
 sg13g2_nand2_1 _4772_ (.Y(_1234_),
    .A(net110),
    .B(net97));
 sg13g2_nand2_1 _4773_ (.Y(_1235_),
    .A(net109),
    .B(_2307_));
 sg13g2_nand2_1 _4774_ (.Y(_1236_),
    .A(_1234_),
    .B(_1235_));
 sg13g2_nor2_1 _4775_ (.A(_1233_),
    .B(_1236_),
    .Y(_1237_));
 sg13g2_a22oi_1 _4776_ (.Y(_1238_),
    .B1(_2617_),
    .B2(_1237_),
    .A2(_1231_),
    .A1(_1229_));
 sg13g2_nor2_1 _4777_ (.A(_1227_),
    .B(_1238_),
    .Y(_1239_));
 sg13g2_inv_1 _4778_ (.Y(_1240_),
    .A(_1239_));
 sg13g2_nand2_1 _4779_ (.Y(_1241_),
    .A(\sqr_pha[9] ),
    .B(\sqr_pha[10] ));
 sg13g2_nand2_1 _4780_ (.Y(_1242_),
    .A(net110),
    .B(_2307_));
 sg13g2_nand2_1 _4781_ (.Y(_1243_),
    .A(_1242_),
    .B(net104));
 sg13g2_inv_1 _4782_ (.Y(_1244_),
    .A(_1243_));
 sg13g2_nor2_1 _4783_ (.A(net109),
    .B(_2317_),
    .Y(_1245_));
 sg13g2_inv_1 _4784_ (.Y(_1246_),
    .A(_1245_));
 sg13g2_a21oi_2 _4785_ (.B1(_2616_),
    .Y(_1247_),
    .A2(_1246_),
    .A1(_1244_));
 sg13g2_nand2_2 _4786_ (.Y(_1248_),
    .A(_2636_),
    .B(_2304_));
 sg13g2_nor2_1 _4787_ (.A(net121),
    .B(_1248_),
    .Y(_1249_));
 sg13g2_inv_1 _4788_ (.Y(_1250_),
    .A(_1249_));
 sg13g2_nand2_1 _4789_ (.Y(_1251_),
    .A(_1250_),
    .B(_2641_));
 sg13g2_nand2_1 _4790_ (.Y(_1252_),
    .A(_1247_),
    .B(_1251_));
 sg13g2_nand2_1 _4791_ (.Y(_1253_),
    .A(_1242_),
    .B(_1232_));
 sg13g2_nor2_1 _4792_ (.A(_2307_),
    .B(_1245_),
    .Y(_1254_));
 sg13g2_nor3_1 _4793_ (.A(_2641_),
    .B(_1253_),
    .C(_1254_),
    .Y(_1255_));
 sg13g2_nand2_1 _4794_ (.Y(_1256_),
    .A(_1255_),
    .B(net91));
 sg13g2_nor2_1 _4795_ (.A(_2337_),
    .B(net120),
    .Y(_1257_));
 sg13g2_nor2_1 _4796_ (.A(_1257_),
    .B(_2340_),
    .Y(_1258_));
 sg13g2_nand3_1 _4797_ (.B(_1256_),
    .C(_1258_),
    .A(_1252_),
    .Y(_1259_));
 sg13g2_nor2_1 _4798_ (.A(net103),
    .B(_1230_),
    .Y(_1260_));
 sg13g2_nor2_1 _4799_ (.A(_2614_),
    .B(_2641_),
    .Y(_1261_));
 sg13g2_inv_1 _4800_ (.Y(_1262_),
    .A(_1261_));
 sg13g2_nor2_1 _4801_ (.A(_1248_),
    .B(_1262_),
    .Y(_1263_));
 sg13g2_o21ai_1 _4802_ (.B1(_2340_),
    .Y(_1264_),
    .A1(_1260_),
    .A2(_1263_));
 sg13g2_nand2_1 _4803_ (.Y(_1265_),
    .A(_1238_),
    .B(_1257_));
 sg13g2_nand3_1 _4804_ (.B(_1264_),
    .C(_1265_),
    .A(_1259_),
    .Y(_1266_));
 sg13g2_nand2_1 _4805_ (.Y(_1267_),
    .A(_1266_),
    .B(net99));
 sg13g2_nand2_1 _4806_ (.Y(_1268_),
    .A(net121),
    .B(_2311_));
 sg13g2_buf_2 _4807_ (.A(_1268_),
    .X(_1269_));
 sg13g2_nor2_1 _4808_ (.A(net97),
    .B(_1269_),
    .Y(_1270_));
 sg13g2_nor2_1 _4809_ (.A(net98),
    .B(_1270_),
    .Y(_1271_));
 sg13g2_nor2b_1 _4810_ (.A(_1243_),
    .B_N(_1248_),
    .Y(_1272_));
 sg13g2_inv_1 _4811_ (.Y(_1273_),
    .A(_1272_));
 sg13g2_nand3b_1 _4812_ (.B(_1273_),
    .C(net84),
    .Y(_1274_),
    .A_N(_1271_));
 sg13g2_nor2_2 _4813_ (.A(net121),
    .B(net97),
    .Y(_1275_));
 sg13g2_a21oi_1 _4814_ (.A1(_1275_),
    .A2(net110),
    .Y(_1276_),
    .B1(net104));
 sg13g2_inv_1 _4815_ (.Y(_1277_),
    .A(_1276_));
 sg13g2_nand3_1 _4816_ (.B(net95),
    .C(_1233_),
    .A(_1277_),
    .Y(_1278_));
 sg13g2_nor2_1 _4817_ (.A(_2337_),
    .B(net99),
    .Y(_1279_));
 sg13g2_nand3_1 _4818_ (.B(_1278_),
    .C(_1279_),
    .A(_1274_),
    .Y(_1280_));
 sg13g2_inv_2 _4819_ (.Y(_1281_),
    .A(_1228_));
 sg13g2_nor2_1 _4820_ (.A(net103),
    .B(net106),
    .Y(_1282_));
 sg13g2_nand2_1 _4821_ (.Y(_1283_),
    .A(net119),
    .B(_2337_));
 sg13g2_a21oi_1 _4822_ (.A1(_1281_),
    .A2(_1282_),
    .Y(_1284_),
    .B1(_1283_));
 sg13g2_nand2_1 _4823_ (.Y(_1285_),
    .A(net97),
    .B(net98));
 sg13g2_inv_1 _4824_ (.Y(_1286_),
    .A(_1269_));
 sg13g2_o21ai_1 _4825_ (.B1(_1262_),
    .Y(_1287_),
    .A1(_1285_),
    .A2(_1286_));
 sg13g2_a21oi_1 _4826_ (.A1(_1284_),
    .A2(_1287_),
    .Y(_1288_),
    .B1(net118));
 sg13g2_nand3_1 _4827_ (.B(_1280_),
    .C(_1288_),
    .A(_1267_),
    .Y(_1289_));
 sg13g2_inv_2 _4828_ (.Y(_1290_),
    .A(net118));
 sg13g2_nor2_1 _4829_ (.A(_1290_),
    .B(_1263_),
    .Y(_1291_));
 sg13g2_nor2_1 _4830_ (.A(net91),
    .B(_1243_),
    .Y(_1292_));
 sg13g2_inv_1 _4831_ (.Y(_1293_),
    .A(_1292_));
 sg13g2_nand2_1 _4832_ (.Y(_1294_),
    .A(_1291_),
    .B(_1293_));
 sg13g2_nand2_1 _4833_ (.Y(_1295_),
    .A(_1289_),
    .B(_1294_));
 sg13g2_o21ai_1 _4834_ (.B1(_1295_),
    .Y(_1296_),
    .A1(_0027_),
    .A2(_1239_));
 sg13g2_inv_1 _4835_ (.Y(_1297_),
    .A(_0026_));
 sg13g2_nand3_1 _4836_ (.B(_0025_),
    .C(_1294_),
    .A(_1289_),
    .Y(_1298_));
 sg13g2_nand3_1 _4837_ (.B(_1297_),
    .C(_1298_),
    .A(_1296_),
    .Y(_1299_));
 sg13g2_o21ai_1 _4838_ (.B1(_1299_),
    .Y(_1300_),
    .A1(_1240_),
    .A2(_1241_));
 sg13g2_buf_1 _4839_ (.A(_1300_),
    .X(_1301_));
 sg13g2_nand2_1 _4840_ (.Y(_1302_),
    .A(net15),
    .B(\sqr_vol[0] ));
 sg13g2_xnor2_1 _4841_ (.Y(_1303_),
    .A(_1211_),
    .B(_1302_));
 sg13g2_inv_1 _4842_ (.Y(_1304_),
    .A(_1225_));
 sg13g2_nor2_1 _4843_ (.A(net110),
    .B(_1231_),
    .Y(_1305_));
 sg13g2_nand2_1 _4844_ (.Y(_1306_),
    .A(_1231_),
    .B(net110));
 sg13g2_nand2b_1 _4845_ (.Y(_1307_),
    .B(_1306_),
    .A_N(_1305_));
 sg13g2_inv_1 _4846_ (.Y(_1308_),
    .A(_1283_));
 sg13g2_nor3_1 _4847_ (.A(net118),
    .B(_2340_),
    .C(_1308_),
    .Y(_1309_));
 sg13g2_buf_2 _4848_ (.A(_1309_),
    .X(_1310_));
 sg13g2_nor3_1 _4849_ (.A(net109),
    .B(net103),
    .C(_1230_),
    .Y(_1311_));
 sg13g2_nor2_1 _4850_ (.A(net95),
    .B(_1235_),
    .Y(_1312_));
 sg13g2_nor3_1 _4851_ (.A(_1311_),
    .B(_1312_),
    .C(_1310_),
    .Y(_1313_));
 sg13g2_a221oi_1 _4852_ (.B2(_1310_),
    .C1(_1313_),
    .B1(_1307_),
    .A1(_1290_),
    .Y(_1314_),
    .A2(_1304_));
 sg13g2_inv_1 _4853_ (.Y(_1315_),
    .A(_0021_));
 sg13g2_nor2_1 _4854_ (.A(net118),
    .B(_2340_),
    .Y(_1316_));
 sg13g2_a21oi_1 _4855_ (.A1(_1305_),
    .A2(_1316_),
    .Y(_1317_),
    .B1(_1226_));
 sg13g2_o21ai_1 _4856_ (.B1(_1317_),
    .Y(_1318_),
    .A1(_1310_),
    .A2(_1311_));
 sg13g2_buf_1 _4857_ (.A(_1318_),
    .X(_1319_));
 sg13g2_nor2_1 _4858_ (.A(_0023_),
    .B(_1319_),
    .Y(_1320_));
 sg13g2_a21oi_1 _4859_ (.A1(_1315_),
    .A2(_1319_),
    .Y(_1321_),
    .B1(_1320_));
 sg13g2_inv_1 _4860_ (.Y(_1322_),
    .A(_0020_));
 sg13g2_nand2_1 _4861_ (.Y(_1323_),
    .A(_1319_),
    .B(_1322_));
 sg13g2_o21ai_1 _4862_ (.B1(_1323_),
    .Y(_1324_),
    .A1(_0022_),
    .A2(_1319_));
 sg13g2_nand2_1 _4863_ (.Y(_1325_),
    .A(_1324_),
    .B(_1314_));
 sg13g2_o21ai_1 _4864_ (.B1(_1325_),
    .Y(_1326_),
    .A1(_1314_),
    .A2(_1321_));
 sg13g2_buf_2 _4865_ (.A(_1326_),
    .X(_1327_));
 sg13g2_nand2_1 _4866_ (.Y(_1328_),
    .A(_1327_),
    .B(\bass_vol[0] ));
 sg13g2_nor2_1 _4867_ (.A(\kick_ctr[1] ),
    .B(\kick_ctr[0] ),
    .Y(_1329_));
 sg13g2_buf_1 _4868_ (.A(_1329_),
    .X(_1330_));
 sg13g2_inv_1 _4869_ (.Y(_1331_),
    .A(_0023_));
 sg13g2_nor2_1 _4870_ (.A(_1331_),
    .B(net101),
    .Y(_1332_));
 sg13g2_a21oi_1 _4871_ (.A1(_1328_),
    .A2(net101),
    .Y(_1333_),
    .B1(_1332_));
 sg13g2_nor2b_1 _4872_ (.A(_1303_),
    .B_N(_1333_),
    .Y(_1334_));
 sg13g2_nand2b_1 _4873_ (.Y(_1335_),
    .B(_1303_),
    .A_N(_1333_));
 sg13g2_nand2b_1 _4874_ (.Y(_1336_),
    .B(_1335_),
    .A_N(_1334_));
 sg13g2_inv_1 _4875_ (.Y(_1337_),
    .A(net62));
 sg13g2_a21oi_1 _4876_ (.A1(_1336_),
    .A2(_1222_),
    .Y(_1338_),
    .B1(_1337_));
 sg13g2_o21ai_1 _4877_ (.B1(_1338_),
    .Y(_1339_),
    .A1(_1222_),
    .A2(_1336_));
 sg13g2_o21ai_1 _4878_ (.B1(_1339_),
    .Y(_0061_),
    .A1(_1212_),
    .A2(net60));
 sg13g2_a21oi_1 _4879_ (.A1(_1335_),
    .A2(_0031_),
    .Y(_1340_),
    .B1(_1334_));
 sg13g2_inv_1 _4880_ (.Y(_1341_),
    .A(_0030_));
 sg13g2_nand2_1 _4881_ (.Y(_1342_),
    .A(_1302_),
    .B(_1212_));
 sg13g2_buf_1 _4882_ (.A(\audio_sample_lpf[1] ),
    .X(_1343_));
 sg13g2_inv_1 _4883_ (.Y(_1344_),
    .A(_1330_));
 sg13g2_a21oi_1 _4884_ (.A1(_1327_),
    .A2(\bass_vol[1] ),
    .Y(_1345_),
    .B1(_1344_));
 sg13g2_inv_1 _4885_ (.Y(_1346_),
    .A(_1332_));
 sg13g2_nand2b_1 _4886_ (.Y(_1347_),
    .B(_1346_),
    .A_N(_1345_));
 sg13g2_xnor2_1 _4887_ (.Y(_1348_),
    .A(_1343_),
    .B(_1347_));
 sg13g2_a21oi_1 _4888_ (.A1(net15),
    .A2(\sqr_vol[1] ),
    .Y(_1349_),
    .B1(_1348_));
 sg13g2_nand3_1 _4889_ (.B(\sqr_vol[1] ),
    .C(_1348_),
    .A(_1300_),
    .Y(_1350_));
 sg13g2_nand2b_1 _4890_ (.Y(_1351_),
    .B(_1350_),
    .A_N(_1349_));
 sg13g2_xor2_1 _4891_ (.B(_1351_),
    .A(_1342_),
    .X(_1352_));
 sg13g2_xnor2_1 _4892_ (.Y(_1353_),
    .A(_1341_),
    .B(_1352_));
 sg13g2_xnor2_1 _4893_ (.Y(_1354_),
    .A(_1340_),
    .B(_1353_));
 sg13g2_nor2_1 _4894_ (.A(_1343_),
    .B(net60),
    .Y(_1355_));
 sg13g2_a21oi_1 _4895_ (.A1(_1354_),
    .A2(net60),
    .Y(_0062_),
    .B1(_1355_));
 sg13g2_nor2_1 _4896_ (.A(_1340_),
    .B(_1353_),
    .Y(_1356_));
 sg13g2_inv_1 _4897_ (.Y(_1357_),
    .A(_0028_));
 sg13g2_nor2b_1 _4898_ (.A(_1347_),
    .B_N(_1343_),
    .Y(_1358_));
 sg13g2_nor2b_1 _4899_ (.A(_1358_),
    .B_N(_1350_),
    .Y(_1359_));
 sg13g2_buf_1 _4900_ (.A(\bass_vol[2] ),
    .X(_1360_));
 sg13g2_buf_1 _4901_ (.A(_1344_),
    .X(_1361_));
 sg13g2_a21oi_1 _4902_ (.A1(_1327_),
    .A2(_1360_),
    .Y(_1362_),
    .B1(net85));
 sg13g2_nand2b_1 _4903_ (.Y(_1363_),
    .B(_1346_),
    .A_N(_1362_));
 sg13g2_xor2_1 _4904_ (.B(_1363_),
    .A(_0029_),
    .X(_1364_));
 sg13g2_a21oi_1 _4905_ (.A1(net15),
    .A2(\sqr_vol[2] ),
    .Y(_1365_),
    .B1(_1364_));
 sg13g2_nand3_1 _4906_ (.B(_1364_),
    .C(\sqr_vol[2] ),
    .A(net15),
    .Y(_1366_));
 sg13g2_nand2b_1 _4907_ (.Y(_1367_),
    .B(_1366_),
    .A_N(_1365_));
 sg13g2_xnor2_1 _4908_ (.Y(_1368_),
    .A(_1359_),
    .B(_1367_));
 sg13g2_xnor2_1 _4909_ (.Y(_1369_),
    .A(_1357_),
    .B(_1368_));
 sg13g2_nor2b_1 _4910_ (.A(_1351_),
    .B_N(_1342_),
    .Y(_1370_));
 sg13g2_nor2_1 _4911_ (.A(_1341_),
    .B(_1352_),
    .Y(_1371_));
 sg13g2_nor2_1 _4912_ (.A(_1370_),
    .B(_1371_),
    .Y(_1372_));
 sg13g2_xor2_1 _4913_ (.B(_1372_),
    .A(_1369_),
    .X(_1373_));
 sg13g2_xnor2_1 _4914_ (.Y(_1374_),
    .A(_1356_),
    .B(_1373_));
 sg13g2_nor2_1 _4915_ (.A(\audio_sample_lpf[2] ),
    .B(net62),
    .Y(_1375_));
 sg13g2_a21oi_1 _4916_ (.A1(_1374_),
    .A2(net60),
    .Y(_0063_),
    .B1(_1375_));
 sg13g2_inv_1 _4917_ (.Y(_1376_),
    .A(_1222_));
 sg13g2_nand2_1 _4918_ (.Y(_1377_),
    .A(_1373_),
    .B(_1356_));
 sg13g2_o21ai_1 _4919_ (.B1(_1377_),
    .Y(_1378_),
    .A1(_1372_),
    .A2(_1369_));
 sg13g2_buf_1 _4920_ (.A(_1378_),
    .X(_1379_));
 sg13g2_nor2_1 _4921_ (.A(_1359_),
    .B(_1367_),
    .Y(_1380_));
 sg13g2_nor2_1 _4922_ (.A(_1357_),
    .B(_1368_),
    .Y(_1381_));
 sg13g2_nor2_1 _4923_ (.A(_1380_),
    .B(_1381_),
    .Y(_1382_));
 sg13g2_nor2_1 _4924_ (.A(_0029_),
    .B(_1363_),
    .Y(_1383_));
 sg13g2_nor2b_1 _4925_ (.A(_1383_),
    .B_N(_1366_),
    .Y(_1384_));
 sg13g2_buf_1 _4926_ (.A(\sqr_vol[3] ),
    .X(_1385_));
 sg13g2_buf_1 _4927_ (.A(\bass_vol[3] ),
    .X(_1386_));
 sg13g2_a21oi_1 _4928_ (.A1(_1327_),
    .A2(_1386_),
    .Y(_1387_),
    .B1(net85));
 sg13g2_nand2b_1 _4929_ (.Y(_1388_),
    .B(_1346_),
    .A_N(_1387_));
 sg13g2_xor2_1 _4930_ (.B(_1388_),
    .A(_0031_),
    .X(_1389_));
 sg13g2_a21oi_1 _4931_ (.A1(net15),
    .A2(_1385_),
    .Y(_1390_),
    .B1(_1389_));
 sg13g2_nand3_1 _4932_ (.B(_1389_),
    .C(_1385_),
    .A(net15),
    .Y(_1391_));
 sg13g2_nand2b_1 _4933_ (.Y(_1392_),
    .B(_1391_),
    .A_N(_1390_));
 sg13g2_nor2_1 _4934_ (.A(_1384_),
    .B(_1392_),
    .Y(_1393_));
 sg13g2_nand2_1 _4935_ (.Y(_1394_),
    .A(_1392_),
    .B(_1384_));
 sg13g2_nor2b_1 _4936_ (.A(_1393_),
    .B_N(_1394_),
    .Y(_1395_));
 sg13g2_xnor2_1 _4937_ (.Y(_1396_),
    .A(_0032_),
    .B(_1395_));
 sg13g2_xor2_1 _4938_ (.B(_1396_),
    .A(_1382_),
    .X(_1397_));
 sg13g2_inv_1 _4939_ (.Y(_1398_),
    .A(_1397_));
 sg13g2_nand2b_1 _4940_ (.Y(_1399_),
    .B(_1398_),
    .A_N(_1379_));
 sg13g2_nand2_1 _4941_ (.Y(_1400_),
    .A(_1379_),
    .B(_1397_));
 sg13g2_nand3_1 _4942_ (.B(net62),
    .C(_1400_),
    .A(_1399_),
    .Y(_1401_));
 sg13g2_o21ai_1 _4943_ (.B1(_1401_),
    .Y(_0064_),
    .A1(_1376_),
    .A2(net60));
 sg13g2_a21oi_1 _4944_ (.A1(_1394_),
    .A2(_0032_),
    .Y(_1402_),
    .B1(_1393_));
 sg13g2_nor2_1 _4945_ (.A(_0031_),
    .B(_1388_),
    .Y(_1403_));
 sg13g2_nor2b_1 _4946_ (.A(_1403_),
    .B_N(_1391_),
    .Y(_1404_));
 sg13g2_buf_2 _4947_ (.A(\sqr_vol[4] ),
    .X(_1405_));
 sg13g2_inv_1 _4948_ (.Y(_1406_),
    .A(_0010_));
 sg13g2_a21oi_1 _4949_ (.A1(_1327_),
    .A2(_1406_),
    .Y(_1407_),
    .B1(_1361_));
 sg13g2_nand2b_1 _4950_ (.Y(_1408_),
    .B(_1346_),
    .A_N(_1407_));
 sg13g2_xnor2_1 _4951_ (.Y(_1409_),
    .A(_1341_),
    .B(_1408_));
 sg13g2_a21oi_1 _4952_ (.A1(net15),
    .A2(_1405_),
    .Y(_1410_),
    .B1(_1409_));
 sg13g2_nand3_1 _4953_ (.B(_1405_),
    .C(_1409_),
    .A(net15),
    .Y(_1411_));
 sg13g2_nand2b_1 _4954_ (.Y(_1412_),
    .B(_1411_),
    .A_N(_1410_));
 sg13g2_xnor2_1 _4955_ (.Y(_1413_),
    .A(_1404_),
    .B(_1412_));
 sg13g2_xor2_1 _4956_ (.B(_1413_),
    .A(_0033_),
    .X(_1414_));
 sg13g2_xor2_1 _4957_ (.B(_1414_),
    .A(_1402_),
    .X(_1415_));
 sg13g2_nor2_1 _4958_ (.A(_1382_),
    .B(_1396_),
    .Y(_1416_));
 sg13g2_nand2b_1 _4959_ (.Y(_1417_),
    .B(_1400_),
    .A_N(_1416_));
 sg13g2_xnor2_1 _4960_ (.Y(_1418_),
    .A(_1415_),
    .B(_1417_));
 sg13g2_nor2_1 _4961_ (.A(\audio_sample_lpf[4] ),
    .B(net62),
    .Y(_1419_));
 sg13g2_a21oi_1 _4962_ (.A1(_1418_),
    .A2(net60),
    .Y(_0065_),
    .B1(_1419_));
 sg13g2_nand2_1 _4963_ (.Y(_1420_),
    .A(_1412_),
    .B(_1404_));
 sg13g2_nor2_1 _4964_ (.A(_1404_),
    .B(_1412_),
    .Y(_1421_));
 sg13g2_a21oi_1 _4965_ (.A1(_1420_),
    .A2(_0033_),
    .Y(_1422_),
    .B1(_1421_));
 sg13g2_nor2_1 _4966_ (.A(_0030_),
    .B(_1408_),
    .Y(_1423_));
 sg13g2_nor2b_1 _4967_ (.A(_1423_),
    .B_N(_1411_),
    .Y(_1424_));
 sg13g2_buf_1 _4968_ (.A(\bass_vol[5] ),
    .X(_1425_));
 sg13g2_a21oi_1 _4969_ (.A1(_1327_),
    .A2(_1425_),
    .Y(_1426_),
    .B1(net85));
 sg13g2_nand2b_1 _4970_ (.Y(_1427_),
    .B(_1346_),
    .A_N(_1426_));
 sg13g2_xnor2_1 _4971_ (.Y(_1428_),
    .A(_1357_),
    .B(_1427_));
 sg13g2_a21oi_1 _4972_ (.A1(_1301_),
    .A2(\sqr_vol[5] ),
    .Y(_1429_),
    .B1(_1428_));
 sg13g2_nand3_1 _4973_ (.B(\sqr_vol[5] ),
    .C(_1428_),
    .A(_1301_),
    .Y(_1430_));
 sg13g2_nand2b_1 _4974_ (.Y(_1431_),
    .B(_1430_),
    .A_N(_1429_));
 sg13g2_xnor2_1 _4975_ (.Y(_1432_),
    .A(_1424_),
    .B(_1431_));
 sg13g2_xor2_1 _4976_ (.B(_1432_),
    .A(_0034_),
    .X(_1433_));
 sg13g2_nor2_1 _4977_ (.A(_1422_),
    .B(_1433_),
    .Y(_1434_));
 sg13g2_inv_1 _4978_ (.Y(_1435_),
    .A(_1434_));
 sg13g2_nand2_1 _4979_ (.Y(_1436_),
    .A(_1433_),
    .B(_1422_));
 sg13g2_nand2_1 _4980_ (.Y(_1437_),
    .A(_1435_),
    .B(_1436_));
 sg13g2_inv_1 _4981_ (.Y(_1438_),
    .A(_1437_));
 sg13g2_nor2b_1 _4982_ (.A(_1398_),
    .B_N(_1415_),
    .Y(_1439_));
 sg13g2_nor2_1 _4983_ (.A(_1402_),
    .B(_1414_),
    .Y(_1440_));
 sg13g2_a21oi_1 _4984_ (.A1(_1415_),
    .A2(_1416_),
    .Y(_1441_),
    .B1(_1440_));
 sg13g2_inv_1 _4985_ (.Y(_1442_),
    .A(_1441_));
 sg13g2_a21o_1 _4986_ (.A2(_1439_),
    .A1(_1379_),
    .B1(_1442_),
    .X(_1443_));
 sg13g2_xnor2_1 _4987_ (.Y(_1444_),
    .A(_1438_),
    .B(_1443_));
 sg13g2_nor2_1 _4988_ (.A(\audio_sample_lpf[5] ),
    .B(net62),
    .Y(_1445_));
 sg13g2_a21oi_1 _4989_ (.A1(_1444_),
    .A2(net60),
    .Y(_0066_),
    .B1(_1445_));
 sg13g2_buf_1 _4990_ (.A(\audio_sample_lpf[6] ),
    .X(_1446_));
 sg13g2_buf_2 _4991_ (.A(\audio_sample_lpf[9] ),
    .X(_1447_));
 sg13g2_xnor2_1 _4992_ (.Y(_1448_),
    .A(_1446_),
    .B(_1447_));
 sg13g2_o21ai_1 _4993_ (.B1(_1430_),
    .Y(_1449_),
    .A1(_0028_),
    .A2(_1427_));
 sg13g2_xor2_1 _4994_ (.B(_1449_),
    .A(_1448_),
    .X(_1450_));
 sg13g2_nand2_1 _4995_ (.Y(_1451_),
    .A(_1431_),
    .B(_1424_));
 sg13g2_nor2_1 _4996_ (.A(_1424_),
    .B(_1431_),
    .Y(_1452_));
 sg13g2_a21oi_1 _4997_ (.A1(_1451_),
    .A2(_0034_),
    .Y(_1453_),
    .B1(_1452_));
 sg13g2_xnor2_1 _4998_ (.Y(_1454_),
    .A(_1450_),
    .B(_1453_));
 sg13g2_inv_1 _4999_ (.Y(_1455_),
    .A(_1454_));
 sg13g2_a21oi_1 _5000_ (.A1(_1443_),
    .A2(_1436_),
    .Y(_1456_),
    .B1(_1434_));
 sg13g2_xnor2_1 _5001_ (.Y(_1457_),
    .A(_1455_),
    .B(_1456_));
 sg13g2_nor2_1 _5002_ (.A(_1446_),
    .B(net62),
    .Y(_1458_));
 sg13g2_a21oi_1 _5003_ (.A1(_1457_),
    .A2(net60),
    .Y(_0067_),
    .B1(_1458_));
 sg13g2_buf_1 _5004_ (.A(\audio_sample_lpf[7] ),
    .X(_1459_));
 sg13g2_inv_1 _5005_ (.Y(_1460_),
    .A(_1459_));
 sg13g2_nor2_1 _5006_ (.A(_1455_),
    .B(_1437_),
    .Y(_1461_));
 sg13g2_nand3_1 _5007_ (.B(_1439_),
    .C(_1461_),
    .A(_1379_),
    .Y(_1462_));
 sg13g2_nand2b_1 _5008_ (.Y(_1463_),
    .B(_1450_),
    .A_N(_1453_));
 sg13g2_o21ai_1 _5009_ (.B1(_1463_),
    .Y(_1464_),
    .A1(_1455_),
    .A2(_1435_));
 sg13g2_a21oi_1 _5010_ (.A1(_1442_),
    .A2(_1461_),
    .Y(_1465_),
    .B1(_1464_));
 sg13g2_inv_1 _5011_ (.Y(_1466_),
    .A(_1446_));
 sg13g2_nor2_1 _5012_ (.A(_1447_),
    .B(_1466_),
    .Y(_1467_));
 sg13g2_nand2_1 _5013_ (.Y(_1468_),
    .A(_1449_),
    .B(_1448_));
 sg13g2_nand2b_1 _5014_ (.Y(_1469_),
    .B(_1468_),
    .A_N(_1467_));
 sg13g2_xnor2_1 _5015_ (.Y(_1470_),
    .A(_1460_),
    .B(_1469_));
 sg13g2_a21oi_1 _5016_ (.A1(_1462_),
    .A2(_1465_),
    .Y(_1471_),
    .B1(_1470_));
 sg13g2_nand3_1 _5017_ (.B(_1465_),
    .C(_1470_),
    .A(_1462_),
    .Y(_1472_));
 sg13g2_nand3b_1 _5018_ (.B(net62),
    .C(_1472_),
    .Y(_1473_),
    .A_N(_1471_));
 sg13g2_o21ai_1 _5019_ (.B1(_1473_),
    .Y(_0068_),
    .A1(_1460_),
    .A2(_1221_));
 sg13g2_buf_2 _5020_ (.A(\audio_sample_lpf[8] ),
    .X(_1474_));
 sg13g2_inv_1 _5021_ (.Y(_1475_),
    .A(_1474_));
 sg13g2_nor2_1 _5022_ (.A(_1470_),
    .B(_1455_),
    .Y(_1476_));
 sg13g2_nand4_1 _5023_ (.B(_1415_),
    .C(_1438_),
    .A(_1417_),
    .Y(_1477_),
    .D(_1476_));
 sg13g2_a21oi_1 _5024_ (.A1(_1440_),
    .A2(_1436_),
    .Y(_1478_),
    .B1(_1434_));
 sg13g2_inv_1 _5025_ (.Y(_1479_),
    .A(_1478_));
 sg13g2_nor2_1 _5026_ (.A(_1459_),
    .B(_1468_),
    .Y(_1480_));
 sg13g2_inv_1 _5027_ (.Y(_1481_),
    .A(_1480_));
 sg13g2_o21ai_1 _5028_ (.B1(_1481_),
    .Y(_1482_),
    .A1(_1470_),
    .A2(_1463_));
 sg13g2_a21oi_1 _5029_ (.A1(_1479_),
    .A2(_1476_),
    .Y(_1483_),
    .B1(_1482_));
 sg13g2_nor2_1 _5030_ (.A(_1459_),
    .B(_1467_),
    .Y(_1484_));
 sg13g2_xnor2_1 _5031_ (.Y(_1485_),
    .A(_1474_),
    .B(_1484_));
 sg13g2_a21oi_1 _5032_ (.A1(_1477_),
    .A2(_1483_),
    .Y(_1486_),
    .B1(_1485_));
 sg13g2_nand3_1 _5033_ (.B(_1483_),
    .C(_1485_),
    .A(_1477_),
    .Y(_1487_));
 sg13g2_nand3b_1 _5034_ (.B(_1220_),
    .C(_1487_),
    .Y(_1488_),
    .A_N(_1486_));
 sg13g2_o21ai_1 _5035_ (.B1(_1488_),
    .Y(_0069_),
    .A1(_1475_),
    .A2(_1221_));
 sg13g2_nor2_1 _5036_ (.A(_1474_),
    .B(_1460_),
    .Y(_1489_));
 sg13g2_xnor2_1 _5037_ (.Y(_1490_),
    .A(_1474_),
    .B(_1447_));
 sg13g2_xor2_1 _5038_ (.B(_1490_),
    .A(_1489_),
    .X(_1491_));
 sg13g2_nor2_1 _5039_ (.A(_1485_),
    .B(_1470_),
    .Y(_1492_));
 sg13g2_nand3_1 _5040_ (.B(_1461_),
    .C(_1492_),
    .A(_1443_),
    .Y(_1493_));
 sg13g2_nand3_1 _5041_ (.B(_1460_),
    .C(_1475_),
    .A(_1467_),
    .Y(_1494_));
 sg13g2_o21ai_1 _5042_ (.B1(_1494_),
    .Y(_1495_),
    .A1(_1485_),
    .A2(_1481_));
 sg13g2_a21oi_1 _5043_ (.A1(_1464_),
    .A2(_1492_),
    .Y(_1496_),
    .B1(_1495_));
 sg13g2_nand2_1 _5044_ (.Y(_1497_),
    .A(_1493_),
    .B(_1496_));
 sg13g2_xnor2_1 _5045_ (.Y(_1498_),
    .A(_1491_),
    .B(_1497_));
 sg13g2_nand2_1 _5046_ (.Y(_1499_),
    .A(_1337_),
    .B(_1447_));
 sg13g2_o21ai_1 _5047_ (.B1(_1499_),
    .Y(_0070_),
    .A1(_1337_),
    .A2(_1498_));
 sg13g2_inv_1 _5048_ (.Y(_1500_),
    .A(\sample_beat_ctr[1] ));
 sg13g2_buf_1 _5049_ (.A(\sample_beat_ctr[0] ),
    .X(_1501_));
 sg13g2_nand3_1 _5050_ (.B(_1501_),
    .C(\sample_beat_ctr[2] ),
    .A(_1500_),
    .Y(_1502_));
 sg13g2_buf_2 _5051_ (.A(_1502_),
    .X(_1503_));
 sg13g2_inv_1 _5052_ (.Y(_1504_),
    .A(_1503_));
 sg13g2_buf_1 _5053_ (.A(_1504_),
    .X(_1505_));
 sg13g2_nand2_1 _5054_ (.Y(_1506_),
    .A(_2649_),
    .B(_2716_));
 sg13g2_nor2_1 _5055_ (.A(_2328_),
    .B(_2765_),
    .Y(_1507_));
 sg13g2_nand2_1 _5056_ (.Y(_1508_),
    .A(_1507_),
    .B(_2320_));
 sg13g2_nand4_1 _5057_ (.B(net93),
    .C(_2667_),
    .A(net105),
    .Y(_1509_),
    .D(_2715_));
 sg13g2_nor4_2 _5058_ (.A(net86),
    .B(_1506_),
    .C(_1508_),
    .Y(_1510_),
    .D(_1509_));
 sg13g2_inv_1 _5059_ (.Y(_1511_),
    .A(_1510_));
 sg13g2_nor2_1 _5060_ (.A(_1511_),
    .B(_1218_),
    .Y(_1512_));
 sg13g2_buf_2 _5061_ (.A(_1512_),
    .X(_1513_));
 sg13g2_inv_1 _5062_ (.Y(_1514_),
    .A(_1513_));
 sg13g2_buf_1 _5063_ (.A(_1514_),
    .X(_1515_));
 sg13g2_nor2_2 _5064_ (.A(net76),
    .B(_1515_),
    .Y(_1516_));
 sg13g2_xnor2_1 _5065_ (.Y(_1517_),
    .A(_1360_),
    .B(\bass_vol[0] ));
 sg13g2_inv_1 _5066_ (.Y(_1518_),
    .A(\bass_vol[0] ));
 sg13g2_inv_1 _5067_ (.Y(_1519_),
    .A(_1270_));
 sg13g2_nor2_1 _5068_ (.A(net96),
    .B(_1519_),
    .Y(_1520_));
 sg13g2_inv_1 _5069_ (.Y(_1521_),
    .A(_1520_));
 sg13g2_nor2_1 _5070_ (.A(net84),
    .B(_1521_),
    .Y(_1522_));
 sg13g2_inv_1 _5071_ (.Y(_1523_),
    .A(_1522_));
 sg13g2_nor3_1 _5072_ (.A(_1290_),
    .B(_1225_),
    .C(_1523_),
    .Y(_1524_));
 sg13g2_nor2_1 _5073_ (.A(net99),
    .B(_1523_),
    .Y(_1525_));
 sg13g2_nand2_1 _5074_ (.Y(_1526_),
    .A(_1525_),
    .B(_2340_));
 sg13g2_xnor2_1 _5075_ (.Y(_1527_),
    .A(net118),
    .B(_1526_));
 sg13g2_nor2b_1 _5076_ (.A(_1524_),
    .B_N(_1527_),
    .Y(_1528_));
 sg13g2_buf_1 _5077_ (.A(_1528_),
    .X(_1529_));
 sg13g2_inv_1 _5078_ (.Y(_1530_),
    .A(_1529_));
 sg13g2_xnor2_1 _5079_ (.Y(_1531_),
    .A(net99),
    .B(_1522_));
 sg13g2_buf_1 _5080_ (.A(_1531_),
    .X(_1532_));
 sg13g2_nor2_1 _5081_ (.A(net120),
    .B(_1525_),
    .Y(_1533_));
 sg13g2_inv_1 _5082_ (.Y(_1534_),
    .A(net120));
 sg13g2_inv_1 _5083_ (.Y(_1535_),
    .A(_1525_));
 sg13g2_nor2_1 _5084_ (.A(_1534_),
    .B(_1535_),
    .Y(_1536_));
 sg13g2_nor2_2 _5085_ (.A(_1533_),
    .B(_1536_),
    .Y(_1537_));
 sg13g2_nor2_1 _5086_ (.A(net47),
    .B(_1537_),
    .Y(_1538_));
 sg13g2_xnor2_1 _5087_ (.Y(_1539_),
    .A(_1224_),
    .B(_1536_));
 sg13g2_inv_1 _5088_ (.Y(_1540_),
    .A(_1539_));
 sg13g2_nand4_1 _5089_ (.B(_1228_),
    .C(_1538_),
    .A(_1530_),
    .Y(_1541_),
    .D(_1540_));
 sg13g2_nand3_1 _5090_ (.B(net108),
    .C(_1513_),
    .A(_1541_),
    .Y(_1542_));
 sg13g2_nor2b_1 _5091_ (.A(_1516_),
    .B_N(_1542_),
    .Y(_1543_));
 sg13g2_buf_1 _5092_ (.A(_1543_),
    .X(_1544_));
 sg13g2_a22oi_1 _5093_ (.Y(_0087_),
    .B1(_1518_),
    .B2(_1544_),
    .A2(_1517_),
    .A1(_1516_));
 sg13g2_inv_1 _5094_ (.Y(_1545_),
    .A(\bass_vol[1] ));
 sg13g2_inv_1 _5095_ (.Y(_1546_),
    .A(_1544_));
 sg13g2_inv_1 _5096_ (.Y(_1547_),
    .A(_1360_));
 sg13g2_nor2_1 _5097_ (.A(\bass_vol[0] ),
    .B(_1547_),
    .Y(_1548_));
 sg13g2_xnor2_1 _5098_ (.Y(_1549_),
    .A(_1386_),
    .B(\bass_vol[1] ));
 sg13g2_xnor2_1 _5099_ (.Y(_1550_),
    .A(_1548_),
    .B(_1549_));
 sg13g2_o21ai_1 _5100_ (.B1(_1546_),
    .Y(_1551_),
    .A1(net76),
    .A2(_1550_));
 sg13g2_o21ai_1 _5101_ (.B1(_1551_),
    .Y(_0088_),
    .A1(_1545_),
    .A2(_1546_));
 sg13g2_xnor2_1 _5102_ (.Y(_1552_),
    .A(_1360_),
    .B(\bass_vol[4] ));
 sg13g2_inv_1 _5103_ (.Y(_1553_),
    .A(_1548_));
 sg13g2_inv_1 _5104_ (.Y(_1554_),
    .A(_1386_));
 sg13g2_nand2_1 _5105_ (.Y(_1555_),
    .A(_1554_),
    .B(\bass_vol[1] ));
 sg13g2_inv_1 _5106_ (.Y(_1556_),
    .A(_1555_));
 sg13g2_a21oi_1 _5107_ (.A1(_1549_),
    .A2(_1553_),
    .Y(_1557_),
    .B1(_1556_));
 sg13g2_xnor2_1 _5108_ (.Y(_1558_),
    .A(_1552_),
    .B(_1557_));
 sg13g2_o21ai_1 _5109_ (.B1(_1546_),
    .Y(_1559_),
    .A1(_1505_),
    .A2(_1558_));
 sg13g2_o21ai_1 _5110_ (.B1(_1559_),
    .Y(_0089_),
    .A1(_1547_),
    .A2(_1546_));
 sg13g2_xnor2_1 _5111_ (.Y(_1560_),
    .A(_1386_),
    .B(_1425_));
 sg13g2_inv_1 _5112_ (.Y(_1561_),
    .A(_1560_));
 sg13g2_inv_1 _5113_ (.Y(_1562_),
    .A(\bass_vol[4] ));
 sg13g2_nor2b_1 _5114_ (.A(_1557_),
    .B_N(_1552_),
    .Y(_1563_));
 sg13g2_a21oi_1 _5115_ (.A1(_1360_),
    .A2(_1562_),
    .Y(_1564_),
    .B1(_1563_));
 sg13g2_nor2_1 _5116_ (.A(_1561_),
    .B(_1564_),
    .Y(_1565_));
 sg13g2_inv_1 _5117_ (.Y(_1566_),
    .A(_1565_));
 sg13g2_nand2_1 _5118_ (.Y(_1567_),
    .A(_1564_),
    .B(_1561_));
 sg13g2_a21oi_1 _5119_ (.A1(_1566_),
    .A2(_1567_),
    .Y(_1568_),
    .B1(_1505_));
 sg13g2_nand2_1 _5120_ (.Y(_1569_),
    .A(_1544_),
    .B(_1386_));
 sg13g2_o21ai_1 _5121_ (.B1(_1569_),
    .Y(_0090_),
    .A1(_1544_),
    .A2(_1568_));
 sg13g2_nor2_1 _5122_ (.A(_1425_),
    .B(_1554_),
    .Y(_1570_));
 sg13g2_nor3_1 _5123_ (.A(_1570_),
    .B(_1565_),
    .C(_1544_),
    .Y(_1571_));
 sg13g2_nand2b_1 _5124_ (.Y(_1572_),
    .B(\bass_vol[4] ),
    .A_N(_1571_));
 sg13g2_nor2_1 _5125_ (.A(_1503_),
    .B(_1515_),
    .Y(_1573_));
 sg13g2_buf_1 _5126_ (.A(_1573_),
    .X(_1574_));
 sg13g2_nand3_1 _5127_ (.B(_2321_),
    .C(net38),
    .A(_1541_),
    .Y(_1575_));
 sg13g2_nand2_1 _5128_ (.Y(_1576_),
    .A(_1571_),
    .B(_1562_));
 sg13g2_nand3_1 _5129_ (.B(_1575_),
    .C(_1576_),
    .A(_1572_),
    .Y(_0091_));
 sg13g2_o21ai_1 _5130_ (.B1(_0010_),
    .Y(_1577_),
    .A1(\bass_vol[4] ),
    .A2(_1566_));
 sg13g2_nor3_1 _5131_ (.A(_1570_),
    .B(_1577_),
    .C(_1544_),
    .Y(_1578_));
 sg13g2_nand2b_1 _5132_ (.Y(_1579_),
    .B(_1425_),
    .A_N(_1578_));
 sg13g2_nand2b_1 _5133_ (.Y(_1580_),
    .B(_1578_),
    .A_N(_1425_));
 sg13g2_nand3_1 _5134_ (.B(_1575_),
    .C(_1580_),
    .A(_1579_),
    .Y(_0092_));
 sg13g2_inv_1 _5135_ (.Y(_1581_),
    .A(_0046_));
 sg13g2_buf_1 _5136_ (.A(_1513_),
    .X(_1582_));
 sg13g2_buf_1 _5137_ (.A(_1513_),
    .X(_1583_));
 sg13g2_nand2b_2 _5138_ (.Y(_1584_),
    .B(net115),
    .A_N(\cos[0] ));
 sg13g2_inv_1 _5139_ (.Y(_1585_),
    .A(net115));
 sg13g2_nand2_1 _5140_ (.Y(_1586_),
    .A(_1585_),
    .B(\cos[0] ));
 sg13g2_nand3_1 _5141_ (.B(_1584_),
    .C(_1586_),
    .A(net58),
    .Y(_1587_));
 sg13g2_o21ai_1 _5142_ (.B1(_1587_),
    .Y(_0093_),
    .A1(_1581_),
    .A2(net59));
 sg13g2_xnor2_1 _5143_ (.Y(_1588_),
    .A(_2377_),
    .B(\cos[1] ));
 sg13g2_xor2_1 _5144_ (.B(_1588_),
    .A(_1584_),
    .X(_1589_));
 sg13g2_nor2_1 _5145_ (.A(_0047_),
    .B(net58),
    .Y(_1590_));
 sg13g2_a21oi_1 _5146_ (.A1(net59),
    .A2(_1589_),
    .Y(_0094_),
    .B1(_1590_));
 sg13g2_nor2_1 _5147_ (.A(\cos[2] ),
    .B(_2430_),
    .Y(_1591_));
 sg13g2_inv_1 _5148_ (.Y(_1592_),
    .A(\cos[2] ));
 sg13g2_nor2_1 _5149_ (.A(net114),
    .B(_1592_),
    .Y(_1593_));
 sg13g2_nor2_1 _5150_ (.A(_1591_),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_nor2b_1 _5151_ (.A(_2377_),
    .B_N(\cos[1] ),
    .Y(_1595_));
 sg13g2_a21oi_2 _5152_ (.B1(_1595_),
    .Y(_1596_),
    .A2(_1584_),
    .A1(_1588_));
 sg13g2_xnor2_1 _5153_ (.Y(_1597_),
    .A(_1594_),
    .B(_1596_));
 sg13g2_nor2_1 _5154_ (.A(_0048_),
    .B(net58),
    .Y(_1598_));
 sg13g2_a21oi_1 _5155_ (.A1(net59),
    .A2(_1597_),
    .Y(_0095_),
    .B1(_1598_));
 sg13g2_nor2_1 _5156_ (.A(\cos[3] ),
    .B(_2430_),
    .Y(_1599_));
 sg13g2_nor2b_1 _5157_ (.A(net114),
    .B_N(\cos[3] ),
    .Y(_1600_));
 sg13g2_nor2_1 _5158_ (.A(_1599_),
    .B(_1600_),
    .Y(_1601_));
 sg13g2_inv_1 _5159_ (.Y(_1602_),
    .A(_1593_));
 sg13g2_o21ai_1 _5160_ (.B1(_1602_),
    .Y(_1603_),
    .A1(_1591_),
    .A2(_1596_));
 sg13g2_xor2_1 _5161_ (.B(_1603_),
    .A(_1601_),
    .X(_1604_));
 sg13g2_nor2_1 _5162_ (.A(_0049_),
    .B(net58),
    .Y(_1605_));
 sg13g2_a21oi_1 _5163_ (.A1(_1604_),
    .A2(net59),
    .Y(_0096_),
    .B1(_1605_));
 sg13g2_inv_1 _5164_ (.Y(_1606_),
    .A(_0050_));
 sg13g2_xnor2_1 _5165_ (.Y(_1607_),
    .A(net114),
    .B(\cos[4] ));
 sg13g2_nand2_1 _5166_ (.Y(_1608_),
    .A(_1601_),
    .B(_1594_));
 sg13g2_nor2_1 _5167_ (.A(_1593_),
    .B(_1600_),
    .Y(_1609_));
 sg13g2_o21ai_1 _5168_ (.B1(_1609_),
    .Y(_1610_),
    .A1(_1608_),
    .A2(_1596_));
 sg13g2_xor2_1 _5169_ (.B(_1610_),
    .A(_1607_),
    .X(_1611_));
 sg13g2_nor2b_1 _5170_ (.A(net54),
    .B_N(_1611_),
    .Y(_1612_));
 sg13g2_a21oi_1 _5171_ (.A1(_1606_),
    .A2(net54),
    .Y(_0097_),
    .B1(_1612_));
 sg13g2_xnor2_1 _5172_ (.Y(_1613_),
    .A(net114),
    .B(\cos[5] ));
 sg13g2_nand3_1 _5173_ (.B(_1601_),
    .C(_1607_),
    .A(_1603_),
    .Y(_1614_));
 sg13g2_nand2_1 _5174_ (.Y(_1615_),
    .A(_2430_),
    .B(\cos[4] ));
 sg13g2_nand3b_1 _5175_ (.B(_1614_),
    .C(_1615_),
    .Y(_1616_),
    .A_N(_1600_));
 sg13g2_xnor2_1 _5176_ (.Y(_1617_),
    .A(_1613_),
    .B(_1616_));
 sg13g2_mux2_1 _5177_ (.A0(_0051_),
    .A1(_1617_),
    .S(net59),
    .X(_0098_));
 sg13g2_nand3_1 _5178_ (.B(_1607_),
    .C(_1613_),
    .A(_1610_),
    .Y(_1618_));
 sg13g2_nand2_1 _5179_ (.Y(_1619_),
    .A(_2430_),
    .B(\cos[5] ));
 sg13g2_nand3_1 _5180_ (.B(_1615_),
    .C(_1619_),
    .A(_1618_),
    .Y(_1620_));
 sg13g2_xor2_1 _5181_ (.B(\cos[6] ),
    .A(net114),
    .X(_1621_));
 sg13g2_nand2b_1 _5182_ (.Y(_1622_),
    .B(_1621_),
    .A_N(_1620_));
 sg13g2_nand2b_1 _5183_ (.Y(_1623_),
    .B(_1620_),
    .A_N(_1621_));
 sg13g2_nand2_2 _5184_ (.Y(_1624_),
    .A(_1622_),
    .B(_1623_));
 sg13g2_nor2_1 _5185_ (.A(\cos[6] ),
    .B(net58),
    .Y(_1625_));
 sg13g2_a21oi_1 _5186_ (.A1(_1624_),
    .A2(net59),
    .Y(_0099_),
    .B1(_1625_));
 sg13g2_mux2_1 _5187_ (.A0(_1048_),
    .A1(_0045_),
    .S(_1583_),
    .X(_0100_));
 sg13g2_nor2_1 _5188_ (.A(_1062_),
    .B(net58),
    .Y(_1626_));
 sg13g2_nor3_1 _5189_ (.A(_1062_),
    .B(_1048_),
    .C(net54),
    .Y(_1627_));
 sg13g2_buf_2 _5190_ (.A(_1627_),
    .X(_1628_));
 sg13g2_and3_1 _5191_ (.X(_1629_),
    .A(_1513_),
    .B(_1062_),
    .C(_1048_));
 sg13g2_buf_1 _5192_ (.A(_1629_),
    .X(_1630_));
 sg13g2_nor3_1 _5193_ (.A(_1626_),
    .B(_1628_),
    .C(_1630_),
    .Y(_0101_));
 sg13g2_xnor2_1 _5194_ (.Y(_0102_),
    .A(_1060_),
    .B(_1630_));
 sg13g2_nand2_1 _5195_ (.Y(_1631_),
    .A(_1630_),
    .B(\frame_count[2] ));
 sg13g2_xnor2_1 _5196_ (.Y(_0103_),
    .A(\frame_count[3] ),
    .B(_1631_));
 sg13g2_nor2_1 _5197_ (.A(_1058_),
    .B(_1631_),
    .Y(_1632_));
 sg13g2_xnor2_1 _5198_ (.Y(_0104_),
    .A(_1093_),
    .B(_1632_));
 sg13g2_nand2_1 _5199_ (.Y(_1633_),
    .A(_1632_),
    .B(\frame_count[4] ));
 sg13g2_xnor2_1 _5200_ (.Y(_0105_),
    .A(_1091_),
    .B(_1633_));
 sg13g2_nand3_1 _5201_ (.B(\frame_count[4] ),
    .C(_1091_),
    .A(_1632_),
    .Y(_1634_));
 sg13g2_xnor2_1 _5202_ (.Y(_0106_),
    .A(\frame_count[6] ),
    .B(_1634_));
 sg13g2_nor2b_1 _5203_ (.A(_1634_),
    .B_N(\frame_count[6] ),
    .Y(_1635_));
 sg13g2_xor2_1 _5204_ (.B(_1635_),
    .A(\frame_count[7] ),
    .X(_0107_));
 sg13g2_inv_1 _5205_ (.Y(_1636_),
    .A(_2765_));
 sg13g2_nand2_1 _5206_ (.Y(_1637_),
    .A(_2388_),
    .B(_2423_));
 sg13g2_inv_1 _5207_ (.Y(_1638_),
    .A(_1637_));
 sg13g2_nand2_1 _5208_ (.Y(_1639_),
    .A(_1638_),
    .B(_2390_));
 sg13g2_inv_1 _5209_ (.Y(_1640_),
    .A(_1639_));
 sg13g2_nand2_1 _5210_ (.Y(_1641_),
    .A(_1640_),
    .B(net116));
 sg13g2_nor2_1 _5211_ (.A(_1059_),
    .B(_1641_),
    .Y(_1642_));
 sg13g2_nand4_1 _5212_ (.B(_2433_),
    .C(_2598_),
    .A(_1642_),
    .Y(_1643_),
    .D(_1038_));
 sg13g2_nand2_1 _5213_ (.Y(_1644_),
    .A(_1643_),
    .B(net130));
 sg13g2_buf_1 _5214_ (.A(_1644_),
    .X(_1645_));
 sg13g2_inv_1 _5215_ (.Y(_1646_),
    .A(_1507_));
 sg13g2_nand2_1 _5216_ (.Y(_1647_),
    .A(net86),
    .B(_2315_));
 sg13g2_nor3_1 _5217_ (.A(_1646_),
    .B(_1647_),
    .C(_1509_),
    .Y(_1648_));
 sg13g2_a21oi_1 _5218_ (.A1(_1648_),
    .A2(_0566_),
    .Y(_1649_),
    .B1(_1213_));
 sg13g2_nand3_1 _5219_ (.B(_0043_),
    .C(_1649_),
    .A(_1645_),
    .Y(_1650_));
 sg13g2_o21ai_1 _5220_ (.B1(_1650_),
    .Y(_0118_),
    .A1(_1636_),
    .A2(net53));
 sg13g2_nand2_1 _5221_ (.Y(_1651_),
    .A(_2328_),
    .B(_2765_));
 sg13g2_nand4_1 _5222_ (.B(_1649_),
    .C(_1646_),
    .A(_1644_),
    .Y(_1652_),
    .D(_1651_));
 sg13g2_o21ai_1 _5223_ (.B1(_1652_),
    .Y(_0119_),
    .A1(_1205_),
    .A2(_1645_));
 sg13g2_inv_1 _5224_ (.Y(_1653_),
    .A(_1644_));
 sg13g2_o21ai_1 _5225_ (.B1(_2320_),
    .Y(_1654_),
    .A1(_1651_),
    .A2(_1653_));
 sg13g2_nor3_1 _5226_ (.A(_2320_),
    .B(_1651_),
    .C(_1653_),
    .Y(_1655_));
 sg13g2_inv_1 _5227_ (.Y(_1656_),
    .A(_1655_));
 sg13g2_nor2_1 _5228_ (.A(_1649_),
    .B(_1653_),
    .Y(_1657_));
 sg13g2_buf_2 _5229_ (.A(_1657_),
    .X(_1658_));
 sg13g2_inv_1 _5230_ (.Y(_1659_),
    .A(_1658_));
 sg13g2_and3_1 _5231_ (.X(_0120_),
    .A(_1654_),
    .B(_1656_),
    .C(_1659_));
 sg13g2_nor2_1 _5232_ (.A(net86),
    .B(_1655_),
    .Y(_1660_));
 sg13g2_nor2_1 _5233_ (.A(net79),
    .B(_1656_),
    .Y(_1661_));
 sg13g2_nor3_1 _5234_ (.A(_1658_),
    .B(_1660_),
    .C(_1661_),
    .Y(_0121_));
 sg13g2_nor2_1 _5235_ (.A(_0248_),
    .B(_1656_),
    .Y(_1662_));
 sg13g2_nor2_1 _5236_ (.A(net122),
    .B(_1661_),
    .Y(_1663_));
 sg13g2_nor3_1 _5237_ (.A(_1658_),
    .B(_1662_),
    .C(_1663_),
    .Y(_0122_));
 sg13g2_nor2_1 _5238_ (.A(net112),
    .B(_1662_),
    .Y(_1664_));
 sg13g2_inv_1 _5239_ (.Y(_1665_),
    .A(_1662_));
 sg13g2_nor2_1 _5240_ (.A(net105),
    .B(_1665_),
    .Y(_1666_));
 sg13g2_nor3_1 _5241_ (.A(_1658_),
    .B(_1664_),
    .C(_1666_),
    .Y(_0123_));
 sg13g2_nor2_1 _5242_ (.A(_2668_),
    .B(_1665_),
    .Y(_1667_));
 sg13g2_nor2_1 _5243_ (.A(_2619_),
    .B(_1666_),
    .Y(_1668_));
 sg13g2_nor3_1 _5244_ (.A(_1658_),
    .B(_1667_),
    .C(_1668_),
    .Y(_0124_));
 sg13g2_nor3_1 _5245_ (.A(_2667_),
    .B(_2668_),
    .C(_1665_),
    .Y(_1669_));
 sg13g2_nor2_1 _5246_ (.A(_2604_),
    .B(_1667_),
    .Y(_1670_));
 sg13g2_nor3_1 _5247_ (.A(_1658_),
    .B(_1669_),
    .C(_1670_),
    .Y(_0125_));
 sg13g2_nor2_1 _5248_ (.A(_2608_),
    .B(_1669_),
    .Y(_1671_));
 sg13g2_nand2_1 _5249_ (.Y(_1672_),
    .A(_1669_),
    .B(_2608_));
 sg13g2_inv_1 _5250_ (.Y(_1673_),
    .A(_1672_));
 sg13g2_nor3_1 _5251_ (.A(_1658_),
    .B(_1671_),
    .C(_1673_),
    .Y(_0126_));
 sg13g2_o21ai_1 _5252_ (.B1(_1659_),
    .Y(_1674_),
    .A1(_2716_),
    .A2(_1672_));
 sg13g2_a21oi_1 _5253_ (.A1(_2716_),
    .A2(_1672_),
    .Y(_0127_),
    .B1(_1674_));
 sg13g2_inv_1 _5254_ (.Y(_1675_),
    .A(\kick_ctr[0] ));
 sg13g2_nor2_1 _5255_ (.A(_1271_),
    .B(_1520_),
    .Y(_1676_));
 sg13g2_inv_1 _5256_ (.Y(_1677_),
    .A(_1676_));
 sg13g2_nor2_2 _5257_ (.A(net84),
    .B(_1677_),
    .Y(_1678_));
 sg13g2_inv_1 _5258_ (.Y(_1679_),
    .A(_1235_));
 sg13g2_nor2_1 _5259_ (.A(_1679_),
    .B(_1286_),
    .Y(_1680_));
 sg13g2_inv_1 _5260_ (.Y(_1681_),
    .A(_1680_));
 sg13g2_o21ai_1 _5261_ (.B1(_1681_),
    .Y(_1682_),
    .A1(_1270_),
    .A2(_1678_));
 sg13g2_nor2_1 _5262_ (.A(_2317_),
    .B(_1236_),
    .Y(_1683_));
 sg13g2_inv_1 _5263_ (.Y(_1684_),
    .A(_1683_));
 sg13g2_a21oi_1 _5264_ (.A1(_1677_),
    .A2(_1228_),
    .Y(_1685_),
    .B1(_1684_));
 sg13g2_inv_1 _5265_ (.Y(_1686_),
    .A(_1537_));
 sg13g2_o21ai_1 _5266_ (.B1(_1686_),
    .Y(_1687_),
    .A1(net47),
    .A2(_1685_));
 sg13g2_a21oi_1 _5267_ (.A1(net47),
    .A2(_1682_),
    .Y(_1688_),
    .B1(_1687_));
 sg13g2_nand2_1 _5268_ (.Y(_1689_),
    .A(_1521_),
    .B(net84));
 sg13g2_nand2_1 _5269_ (.Y(_1690_),
    .A(_1523_),
    .B(_1689_));
 sg13g2_buf_2 _5270_ (.A(_1690_),
    .X(_1691_));
 sg13g2_inv_1 _5271_ (.Y(_1692_),
    .A(_1691_));
 sg13g2_nor2_1 _5272_ (.A(net97),
    .B(_1281_),
    .Y(_1693_));
 sg13g2_nand2_1 _5273_ (.Y(_1694_),
    .A(_1677_),
    .B(net108));
 sg13g2_nand3_1 _5274_ (.B(_1693_),
    .C(_1694_),
    .A(_1692_),
    .Y(_1695_));
 sg13g2_nor2_1 _5275_ (.A(net108),
    .B(net110),
    .Y(_1696_));
 sg13g2_inv_1 _5276_ (.Y(_1697_),
    .A(_1275_));
 sg13g2_nand2_1 _5277_ (.Y(_1698_),
    .A(_1684_),
    .B(_1697_));
 sg13g2_nand3_1 _5278_ (.B(_1696_),
    .C(_1698_),
    .A(_1691_),
    .Y(_1699_));
 sg13g2_inv_1 _5279_ (.Y(_1700_),
    .A(_1531_));
 sg13g2_nand4_1 _5280_ (.B(_1699_),
    .C(_1519_),
    .A(_1695_),
    .Y(_1701_),
    .D(_1700_));
 sg13g2_nand2_1 _5281_ (.Y(_1702_),
    .A(_1685_),
    .B(_1692_));
 sg13g2_nor2_1 _5282_ (.A(_2632_),
    .B(_1269_),
    .Y(_1703_));
 sg13g2_nand2_1 _5283_ (.Y(_1704_),
    .A(_1691_),
    .B(_1703_));
 sg13g2_nand3_1 _5284_ (.B(net47),
    .C(_1704_),
    .A(_1702_),
    .Y(_1705_));
 sg13g2_nand3_1 _5285_ (.B(_1537_),
    .C(_1705_),
    .A(_1701_),
    .Y(_1706_));
 sg13g2_nand3b_1 _5286_ (.B(_1539_),
    .C(_1706_),
    .Y(_1707_),
    .A_N(_1688_));
 sg13g2_nand2_1 _5287_ (.Y(_1708_),
    .A(_1678_),
    .B(_1683_));
 sg13g2_a21oi_1 _5288_ (.A1(_1708_),
    .A2(_1269_),
    .Y(_1709_),
    .B1(net47));
 sg13g2_o21ai_1 _5289_ (.B1(net47),
    .Y(_1710_),
    .A1(_1681_),
    .A2(_1678_));
 sg13g2_a21oi_1 _5290_ (.A1(_1269_),
    .A2(_1678_),
    .Y(_1711_),
    .B1(_1710_));
 sg13g2_o21ai_1 _5291_ (.B1(_1537_),
    .Y(_1712_),
    .A1(_1709_),
    .A2(_1711_));
 sg13g2_nor3_1 _5292_ (.A(net97),
    .B(_1230_),
    .C(_1281_),
    .Y(_1713_));
 sg13g2_nor2b_1 _5293_ (.A(net47),
    .B_N(_1713_),
    .Y(_1714_));
 sg13g2_nor2_1 _5294_ (.A(_1269_),
    .B(_1700_),
    .Y(_1715_));
 sg13g2_o21ai_1 _5295_ (.B1(_1686_),
    .Y(_1716_),
    .A1(_1714_),
    .A2(_1715_));
 sg13g2_nand3_1 _5296_ (.B(_1540_),
    .C(_1716_),
    .A(_1712_),
    .Y(_1717_));
 sg13g2_nand3_1 _5297_ (.B(_1530_),
    .C(_1717_),
    .A(_1707_),
    .Y(_1718_));
 sg13g2_nor2_2 _5298_ (.A(net108),
    .B(_2632_),
    .Y(_1719_));
 sg13g2_inv_1 _5299_ (.Y(_1720_),
    .A(_1719_));
 sg13g2_nand3_1 _5300_ (.B(_1720_),
    .C(_1678_),
    .A(_1529_),
    .Y(_1721_));
 sg13g2_nand3_1 _5301_ (.B(net76),
    .C(_1721_),
    .A(_1718_),
    .Y(_1722_));
 sg13g2_o21ai_1 _5302_ (.B1(net135),
    .Y(_1723_),
    .A1(_1361_),
    .A2(_1504_));
 sg13g2_nor2_1 _5303_ (.A(_1723_),
    .B(_1514_),
    .Y(_1724_));
 sg13g2_nand2_2 _5304_ (.Y(_1725_),
    .A(_1722_),
    .B(_1724_));
 sg13g2_inv_1 _5305_ (.Y(_1726_),
    .A(_1725_));
 sg13g2_buf_1 _5306_ (.A(_1726_),
    .X(_1727_));
 sg13g2_o21ai_1 _5307_ (.B1(net11),
    .Y(_1728_),
    .A1(_0044_),
    .A2(net76));
 sg13g2_o21ai_1 _5308_ (.B1(_1728_),
    .Y(_0128_),
    .A1(_1675_),
    .A2(net11));
 sg13g2_a21oi_1 _5309_ (.A1(_1726_),
    .A2(\kick_ctr[0] ),
    .Y(_1729_),
    .B1(\kick_ctr[1] ));
 sg13g2_nor2_1 _5310_ (.A(_1503_),
    .B(_1725_),
    .Y(_1730_));
 sg13g2_and3_1 _5311_ (.X(_1731_),
    .A(_1726_),
    .B(\kick_ctr[1] ),
    .C(\kick_ctr[0] ));
 sg13g2_nor3_1 _5312_ (.A(_1729_),
    .B(_1730_),
    .C(_1731_),
    .Y(_0129_));
 sg13g2_a21oi_1 _5313_ (.A1(_1726_),
    .A2(\kick_osci[3] ),
    .Y(_1732_),
    .B1(\kick_osci[0] ));
 sg13g2_and3_1 _5314_ (.X(_1733_),
    .A(_1726_),
    .B(\kick_osci[3] ),
    .C(\kick_osci[0] ));
 sg13g2_nor3_1 _5315_ (.A(_1730_),
    .B(_1732_),
    .C(_1733_),
    .Y(_0130_));
 sg13g2_inv_1 _5316_ (.Y(_1734_),
    .A(\kick_osci[3] ));
 sg13g2_nor2_1 _5317_ (.A(\kick_osci[0] ),
    .B(_1734_),
    .Y(_1735_));
 sg13g2_xnor2_1 _5318_ (.Y(_1736_),
    .A(\kick_osci[4] ),
    .B(\kick_osci[1] ));
 sg13g2_inv_1 _5319_ (.Y(_1737_),
    .A(_1736_));
 sg13g2_nor2_1 _5320_ (.A(_1735_),
    .B(_1737_),
    .Y(_1738_));
 sg13g2_a21oi_1 _5321_ (.A1(_1737_),
    .A2(_1735_),
    .Y(_1739_),
    .B1(net76));
 sg13g2_nand2b_1 _5322_ (.Y(_1740_),
    .B(_1739_),
    .A_N(_1738_));
 sg13g2_nand2_1 _5323_ (.Y(_1741_),
    .A(_1725_),
    .B(\kick_osci[1] ));
 sg13g2_o21ai_1 _5324_ (.B1(_1741_),
    .Y(_0131_),
    .A1(_1725_),
    .A2(_1740_));
 sg13g2_inv_1 _5325_ (.Y(_1742_),
    .A(\kick_osci[2] ));
 sg13g2_buf_1 _5326_ (.A(\kick_osci[5] ),
    .X(_1743_));
 sg13g2_xnor2_1 _5327_ (.Y(_1744_),
    .A(_1743_),
    .B(\kick_osci[2] ));
 sg13g2_inv_1 _5328_ (.Y(_1745_),
    .A(_1744_));
 sg13g2_inv_1 _5329_ (.Y(_1746_),
    .A(\kick_osci[4] ));
 sg13g2_a21oi_1 _5330_ (.A1(_1746_),
    .A2(\kick_osci[1] ),
    .Y(_1747_),
    .B1(_1738_));
 sg13g2_nor2_1 _5331_ (.A(_1745_),
    .B(_1747_),
    .Y(_1748_));
 sg13g2_a21oi_1 _5332_ (.A1(_1747_),
    .A2(_1745_),
    .Y(_1749_),
    .B1(net76));
 sg13g2_nand3b_1 _5333_ (.B(net11),
    .C(_1749_),
    .Y(_1750_),
    .A_N(_1748_));
 sg13g2_o21ai_1 _5334_ (.B1(_1750_),
    .Y(_0132_),
    .A1(_1742_),
    .A2(net11));
 sg13g2_inv_1 _5335_ (.Y(_1751_),
    .A(_1743_));
 sg13g2_a21oi_1 _5336_ (.A1(_1751_),
    .A2(\kick_osci[2] ),
    .Y(_1752_),
    .B1(_1748_));
 sg13g2_xnor2_1 _5337_ (.Y(_1753_),
    .A(\kick_osci[3] ),
    .B(\kick_osci[6] ));
 sg13g2_nand2b_1 _5338_ (.Y(_1754_),
    .B(_1753_),
    .A_N(_1752_));
 sg13g2_nand2b_1 _5339_ (.Y(_1755_),
    .B(_1752_),
    .A_N(_1753_));
 sg13g2_nand4_1 _5340_ (.B(_1503_),
    .C(_1754_),
    .A(_1727_),
    .Y(_1756_),
    .D(_1755_));
 sg13g2_o21ai_1 _5341_ (.B1(_1756_),
    .Y(_0133_),
    .A1(_1734_),
    .A2(_1727_));
 sg13g2_xnor2_1 _5342_ (.Y(_1757_),
    .A(\kick_osci[4] ),
    .B(\kick_osci[7] ));
 sg13g2_o21ai_1 _5343_ (.B1(_1754_),
    .Y(_1758_),
    .A1(_1734_),
    .A2(\kick_osci[6] ));
 sg13g2_o21ai_1 _5344_ (.B1(_1503_),
    .Y(_1759_),
    .A1(_1757_),
    .A2(_1758_));
 sg13g2_nand2_1 _5345_ (.Y(_1760_),
    .A(_1758_),
    .B(_1757_));
 sg13g2_nand3b_1 _5346_ (.B(net11),
    .C(_1760_),
    .Y(_1761_),
    .A_N(_1759_));
 sg13g2_o21ai_1 _5347_ (.B1(_1761_),
    .Y(_0134_),
    .A1(_1746_),
    .A2(net11));
 sg13g2_buf_1 _5348_ (.A(\kick_osci[8] ),
    .X(_1762_));
 sg13g2_xnor2_1 _5349_ (.Y(_1763_),
    .A(_1762_),
    .B(_1743_));
 sg13g2_o21ai_1 _5350_ (.B1(_1760_),
    .Y(_1764_),
    .A1(_1746_),
    .A2(\kick_osci[7] ));
 sg13g2_or2_1 _5351_ (.X(_1765_),
    .B(_1764_),
    .A(_1763_));
 sg13g2_nand2_1 _5352_ (.Y(_1766_),
    .A(_1764_),
    .B(_1763_));
 sg13g2_nand4_1 _5353_ (.B(_1503_),
    .C(_1765_),
    .A(net11),
    .Y(_1767_),
    .D(_1766_));
 sg13g2_o21ai_1 _5354_ (.B1(_1767_),
    .Y(_0135_),
    .A1(_1751_),
    .A2(net11));
 sg13g2_inv_1 _5355_ (.Y(_1768_),
    .A(\kick_osci[6] ));
 sg13g2_inv_1 _5356_ (.Y(_1769_),
    .A(_1762_));
 sg13g2_inv_1 _5357_ (.Y(_1770_),
    .A(_1766_));
 sg13g2_a21oi_1 _5358_ (.A1(_1769_),
    .A2(_1743_),
    .Y(_1771_),
    .B1(_1770_));
 sg13g2_nand2_1 _5359_ (.Y(_1772_),
    .A(_1726_),
    .B(_1771_));
 sg13g2_inv_1 _5360_ (.Y(_1773_),
    .A(_1730_));
 sg13g2_o21ai_1 _5361_ (.B1(_1773_),
    .Y(_1774_),
    .A1(_1768_),
    .A2(_1772_));
 sg13g2_a21oi_1 _5362_ (.A1(_1768_),
    .A2(_1772_),
    .Y(_0136_),
    .B1(_1774_));
 sg13g2_inv_1 _5363_ (.Y(_1775_),
    .A(\kick_osci[7] ));
 sg13g2_a22oi_1 _5364_ (.Y(_1776_),
    .B1(_1768_),
    .B2(_1770_),
    .A2(_1743_),
    .A1(_1769_));
 sg13g2_nand4_1 _5365_ (.B(_0017_),
    .C(_1775_),
    .A(_1726_),
    .Y(_1777_),
    .D(_1776_));
 sg13g2_nand2_1 _5366_ (.Y(_1778_),
    .A(_1776_),
    .B(_0017_));
 sg13g2_o21ai_1 _5367_ (.B1(\kick_osci[7] ),
    .Y(_1779_),
    .A1(_1778_),
    .A2(_1725_));
 sg13g2_nand3_1 _5368_ (.B(_1773_),
    .C(_1779_),
    .A(_1777_),
    .Y(_0137_));
 sg13g2_nand2_1 _5369_ (.Y(_1780_),
    .A(_1768_),
    .B(_1775_));
 sg13g2_o21ai_1 _5370_ (.B1(_1762_),
    .Y(_1781_),
    .A1(_1780_),
    .A2(_1772_));
 sg13g2_nand2_1 _5371_ (.Y(_0138_),
    .A(_1781_),
    .B(_1773_));
 sg13g2_nor2_1 _5372_ (.A(_1508_),
    .B(_1337_),
    .Y(_1782_));
 sg13g2_buf_1 _5373_ (.A(_1782_),
    .X(_1783_));
 sg13g2_buf_1 _5374_ (.A(_1783_),
    .X(_1784_));
 sg13g2_nand3_1 _5375_ (.B(\line_lfsr[1] ),
    .C(_1511_),
    .A(_1783_),
    .Y(_1785_));
 sg13g2_o21ai_1 _5376_ (.B1(_1785_),
    .Y(_0139_),
    .A1(_1117_),
    .A2(net37));
 sg13g2_o21ai_1 _5377_ (.B1(net37),
    .Y(_1786_),
    .A1(\line_lfsr[2] ),
    .A2(_1510_));
 sg13g2_o21ai_1 _5378_ (.B1(_1786_),
    .Y(_0140_),
    .A1(_1114_),
    .A2(_1784_));
 sg13g2_inv_1 _5379_ (.Y(_1787_),
    .A(\line_lfsr[2] ));
 sg13g2_nand3_1 _5380_ (.B(\line_lfsr[3] ),
    .C(_1511_),
    .A(_1783_),
    .Y(_1788_));
 sg13g2_o21ai_1 _5381_ (.B1(_1788_),
    .Y(_0141_),
    .A1(_1787_),
    .A2(_1784_));
 sg13g2_o21ai_1 _5382_ (.B1(net37),
    .Y(_1789_),
    .A1(\line_lfsr[4] ),
    .A2(_1510_));
 sg13g2_o21ai_1 _5383_ (.B1(_1789_),
    .Y(_0142_),
    .A1(_1124_),
    .A2(net37));
 sg13g2_o21ai_1 _5384_ (.B1(net37),
    .Y(_1790_),
    .A1(\line_lfsr[5] ),
    .A2(_1510_));
 sg13g2_o21ai_1 _5385_ (.B1(_1790_),
    .Y(_0143_),
    .A1(_1090_),
    .A2(net37));
 sg13g2_nand2_1 _5386_ (.Y(_1791_),
    .A(_1117_),
    .B(_1109_));
 sg13g2_nand2_1 _5387_ (.Y(_1792_),
    .A(\line_lfsr[0] ),
    .B(\line_lfsr[6] ));
 sg13g2_nand4_1 _5388_ (.B(_1511_),
    .C(_1791_),
    .A(_1783_),
    .Y(_1793_),
    .D(_1792_));
 sg13g2_o21ai_1 _5389_ (.B1(_1793_),
    .Y(_0144_),
    .A1(_1099_),
    .A2(net37));
 sg13g2_o21ai_1 _5390_ (.B1(_1783_),
    .Y(_1794_),
    .A1(\line_lfsr[0] ),
    .A2(_1510_));
 sg13g2_o21ai_1 _5391_ (.B1(_1794_),
    .Y(_0145_),
    .A1(_1109_),
    .A2(net37));
 sg13g2_nand2_1 _5392_ (.Y(_1795_),
    .A(_2483_),
    .B(_2347_));
 sg13g2_nand3_1 _5393_ (.B(_0008_),
    .C(_1795_),
    .A(_1628_),
    .Y(_1796_));
 sg13g2_o21ai_1 _5394_ (.B1(_1796_),
    .Y(_0146_),
    .A1(_2482_),
    .A2(_1628_));
 sg13g2_o21ai_1 _5395_ (.B1(_1628_),
    .Y(_1797_),
    .A1(_2485_),
    .A2(_0457_));
 sg13g2_o21ai_1 _5396_ (.B1(_1797_),
    .Y(_0147_),
    .A1(_2479_),
    .A2(_1628_));
 sg13g2_nor3_1 _5397_ (.A(_2482_),
    .B(_2348_),
    .C(_2480_),
    .Y(_1798_));
 sg13g2_nand2b_1 _5398_ (.Y(_1799_),
    .B(_1628_),
    .A_N(_0254_));
 sg13g2_a22oi_1 _5399_ (.Y(_0148_),
    .B1(_0559_),
    .B2(_1799_),
    .A2(_1798_),
    .A1(_1628_));
 sg13g2_xor2_1 _5400_ (.B(net59),
    .A(_1501_),
    .X(_0149_));
 sg13g2_buf_1 _5401_ (.A(_1573_),
    .X(_1800_));
 sg13g2_a21oi_1 _5402_ (.A1(net58),
    .A2(_1501_),
    .Y(_1801_),
    .B1(\sample_beat_ctr[1] ));
 sg13g2_nand2_1 _5403_ (.Y(_1802_),
    .A(_1513_),
    .B(_1501_));
 sg13g2_nor2_1 _5404_ (.A(_1500_),
    .B(_1802_),
    .Y(_1803_));
 sg13g2_nor3_1 _5405_ (.A(_1800_),
    .B(_1801_),
    .C(_1803_),
    .Y(_0150_));
 sg13g2_mux2_1 _5406_ (.A0(_1803_),
    .A1(_1802_),
    .S(\sample_beat_ctr[2] ),
    .X(_0151_));
 sg13g2_xor2_1 _5407_ (.B(_1612_),
    .A(\sin[0] ),
    .X(_0152_));
 sg13g2_nand2_1 _5408_ (.Y(_1804_),
    .A(_1611_),
    .B(\sin[0] ));
 sg13g2_inv_1 _5409_ (.Y(_1805_),
    .A(\nyan_x_offset[0] ));
 sg13g2_xnor2_1 _5410_ (.Y(_1806_),
    .A(_1805_),
    .B(_1617_));
 sg13g2_xnor2_1 _5411_ (.Y(_1807_),
    .A(_1804_),
    .B(_1806_));
 sg13g2_nor2_1 _5412_ (.A(\nyan_x_offset[0] ),
    .B(_1583_),
    .Y(_1808_));
 sg13g2_a21oi_1 _5413_ (.A1(_1807_),
    .A2(_1582_),
    .Y(_0153_),
    .B1(_1808_));
 sg13g2_inv_1 _5414_ (.Y(_1809_),
    .A(\nyan_x_offset[1] ));
 sg13g2_inv_1 _5415_ (.Y(_1810_),
    .A(_1617_));
 sg13g2_nor2_1 _5416_ (.A(_1804_),
    .B(_1806_),
    .Y(_1811_));
 sg13g2_a21oi_1 _5417_ (.A1(\nyan_x_offset[0] ),
    .A2(_1810_),
    .Y(_1812_),
    .B1(_1811_));
 sg13g2_inv_1 _5418_ (.Y(_1813_),
    .A(_1624_));
 sg13g2_nor2_1 _5419_ (.A(\nyan_x_offset[1] ),
    .B(_1813_),
    .Y(_1814_));
 sg13g2_nor2_1 _5420_ (.A(_1809_),
    .B(_1624_),
    .Y(_1815_));
 sg13g2_inv_1 _5421_ (.Y(_1816_),
    .A(_1815_));
 sg13g2_nand2b_1 _5422_ (.Y(_1817_),
    .B(_1816_),
    .A_N(_1814_));
 sg13g2_a21oi_1 _5423_ (.A1(_1812_),
    .A2(_1817_),
    .Y(_1818_),
    .B1(net54));
 sg13g2_o21ai_1 _5424_ (.B1(_1818_),
    .Y(_1819_),
    .A1(_1812_),
    .A2(_1817_));
 sg13g2_o21ai_1 _5425_ (.B1(_1819_),
    .Y(_0154_),
    .A1(_1809_),
    .A2(_1582_));
 sg13g2_inv_1 _5426_ (.Y(_1820_),
    .A(_2391_));
 sg13g2_nor2_1 _5427_ (.A(_1820_),
    .B(_1624_),
    .Y(_1821_));
 sg13g2_nor2_1 _5428_ (.A(_2391_),
    .B(_1813_),
    .Y(_1822_));
 sg13g2_nor2_1 _5429_ (.A(_1821_),
    .B(_1822_),
    .Y(_1823_));
 sg13g2_o21ai_1 _5430_ (.B1(_1816_),
    .Y(_1824_),
    .A1(_1814_),
    .A2(_1812_));
 sg13g2_xnor2_1 _5431_ (.Y(_1825_),
    .A(_1823_),
    .B(_1824_));
 sg13g2_nand2_1 _5432_ (.Y(_1826_),
    .A(net54),
    .B(_2391_));
 sg13g2_o21ai_1 _5433_ (.B1(_1826_),
    .Y(_0155_),
    .A1(net54),
    .A2(_1825_));
 sg13g2_xnor2_1 _5434_ (.Y(_1827_),
    .A(net115),
    .B(_1624_));
 sg13g2_inv_1 _5435_ (.Y(_1828_),
    .A(_1824_));
 sg13g2_nor2_1 _5436_ (.A(_1822_),
    .B(_1828_),
    .Y(_1829_));
 sg13g2_or2_1 _5437_ (.X(_1830_),
    .B(_1829_),
    .A(_1821_));
 sg13g2_xnor2_1 _5438_ (.Y(_1831_),
    .A(_1827_),
    .B(_1830_));
 sg13g2_nor2_1 _5439_ (.A(net115),
    .B(net58),
    .Y(_1832_));
 sg13g2_a21oi_1 _5440_ (.A1(_1831_),
    .A2(net59),
    .Y(_0156_),
    .B1(_1832_));
 sg13g2_nor2_1 _5441_ (.A(_1585_),
    .B(_1624_),
    .Y(_1833_));
 sg13g2_nor2_1 _5442_ (.A(net115),
    .B(_1828_),
    .Y(_1834_));
 sg13g2_nor4_1 _5443_ (.A(net54),
    .B(_1822_),
    .C(_1833_),
    .D(_1834_),
    .Y(_1835_));
 sg13g2_o21ai_1 _5444_ (.B1(_1835_),
    .Y(_1836_),
    .A1(_1820_),
    .A2(_1824_));
 sg13g2_xnor2_1 _5445_ (.Y(_0157_),
    .A(_2377_),
    .B(_1836_));
 sg13g2_inv_1 _5446_ (.Y(_1837_),
    .A(_2377_));
 sg13g2_a22oi_1 _5447_ (.Y(_1838_),
    .B1(net115),
    .B2(_1829_),
    .A2(_1813_),
    .A1(_1837_));
 sg13g2_and3_1 _5448_ (.X(_1839_),
    .A(_1830_),
    .B(_1837_),
    .C(_1827_));
 sg13g2_nor4_1 _5449_ (.A(net54),
    .B(_1833_),
    .C(_1838_),
    .D(_1839_),
    .Y(_1840_));
 sg13g2_xnor2_1 _5450_ (.Y(_0158_),
    .A(_2430_),
    .B(_1840_));
 sg13g2_nand2_1 _5451_ (.Y(_1841_),
    .A(net38),
    .B(_1524_));
 sg13g2_nor2_1 _5452_ (.A(_2963_),
    .B(_1841_),
    .Y(_1842_));
 sg13g2_a21oi_1 _5453_ (.A1(net107),
    .A2(_1841_),
    .Y(_0159_),
    .B1(_1842_));
 sg13g2_mux2_1 _5454_ (.A0(_0052_),
    .A1(_2321_),
    .S(net36),
    .X(_0160_));
 sg13g2_nor2_1 _5455_ (.A(_0053_),
    .B(net38),
    .Y(_1843_));
 sg13g2_a21oi_1 _5456_ (.A1(_1228_),
    .A2(net36),
    .Y(_0161_),
    .B1(_1843_));
 sg13g2_nor2_1 _5457_ (.A(_0054_),
    .B(_1574_),
    .Y(_1844_));
 sg13g2_a21oi_1 _5458_ (.A1(_1698_),
    .A2(net36),
    .Y(_0162_),
    .B1(_1844_));
 sg13g2_nor2_1 _5459_ (.A(_0055_),
    .B(net38),
    .Y(_1845_));
 sg13g2_a21oi_1 _5460_ (.A1(net36),
    .A2(_1676_),
    .Y(_0163_),
    .B1(_1845_));
 sg13g2_nor2_1 _5461_ (.A(_0056_),
    .B(_1574_),
    .Y(_1846_));
 sg13g2_a21oi_1 _5462_ (.A1(net36),
    .A2(_1692_),
    .Y(_0164_),
    .B1(_1846_));
 sg13g2_nor2_1 _5463_ (.A(_0057_),
    .B(net38),
    .Y(_1847_));
 sg13g2_a21oi_1 _5464_ (.A1(net47),
    .A2(net36),
    .Y(_0165_),
    .B1(_1847_));
 sg13g2_nor2_1 _5465_ (.A(_0058_),
    .B(net38),
    .Y(_1848_));
 sg13g2_a21oi_1 _5466_ (.A1(_1537_),
    .A2(_1800_),
    .Y(_0166_),
    .B1(_1848_));
 sg13g2_nor2_1 _5467_ (.A(_0059_),
    .B(net38),
    .Y(_1849_));
 sg13g2_a21oi_1 _5468_ (.A1(_1539_),
    .A2(net36),
    .Y(_0167_),
    .B1(_1849_));
 sg13g2_nor2_1 _5469_ (.A(_0060_),
    .B(net38),
    .Y(_1850_));
 sg13g2_a21oi_1 _5470_ (.A1(_1529_),
    .A2(net36),
    .Y(_0168_),
    .B1(_1850_));
 sg13g2_nand2b_1 _5471_ (.Y(_1851_),
    .B(_1385_),
    .A_N(\sqr_vol[0] ));
 sg13g2_nand2_1 _5472_ (.Y(_1852_),
    .A(_1719_),
    .B(_2642_));
 sg13g2_inv_1 _5473_ (.Y(_1853_),
    .A(_1234_));
 sg13g2_nor3_1 _5474_ (.A(net108),
    .B(net96),
    .C(_1853_),
    .Y(_1854_));
 sg13g2_inv_1 _5475_ (.Y(_1855_),
    .A(_1854_));
 sg13g2_nor2_2 _5476_ (.A(_2311_),
    .B(net104),
    .Y(_1856_));
 sg13g2_a21oi_1 _5477_ (.A1(_1719_),
    .A2(_1856_),
    .Y(_1857_),
    .B1(_1691_));
 sg13g2_a22oi_1 _5478_ (.Y(_1858_),
    .B1(_1855_),
    .B2(_1857_),
    .A2(_1852_),
    .A1(_1691_));
 sg13g2_nand3b_1 _5479_ (.B(_1537_),
    .C(_1700_),
    .Y(_1859_),
    .A_N(_1858_));
 sg13g2_a21oi_1 _5480_ (.A1(_1691_),
    .A2(_1236_),
    .Y(_1860_),
    .B1(net108));
 sg13g2_o21ai_1 _5481_ (.B1(_1677_),
    .Y(_1861_),
    .A1(_1248_),
    .A2(_1691_));
 sg13g2_nand2_1 _5482_ (.Y(_1862_),
    .A(_1861_),
    .B(_1699_));
 sg13g2_o21ai_1 _5483_ (.B1(_1862_),
    .Y(_1863_),
    .A1(_1676_),
    .A2(_1860_));
 sg13g2_nand2_1 _5484_ (.Y(_1864_),
    .A(_1863_),
    .B(_1538_));
 sg13g2_nor2_1 _5485_ (.A(net109),
    .B(_1232_),
    .Y(_1865_));
 sg13g2_o21ai_1 _5486_ (.B1(_1677_),
    .Y(_1866_),
    .A1(_1865_),
    .A2(_1719_));
 sg13g2_and3_1 _5487_ (.X(_1867_),
    .A(_1866_),
    .B(_1691_),
    .C(_1855_));
 sg13g2_o21ai_1 _5488_ (.B1(_1532_),
    .Y(_1868_),
    .A1(_1857_),
    .A2(_1867_));
 sg13g2_nand3_1 _5489_ (.B(_1864_),
    .C(_1868_),
    .A(_1859_),
    .Y(_1869_));
 sg13g2_a21oi_1 _5490_ (.A1(_2317_),
    .A2(_1856_),
    .Y(_1870_),
    .B1(_1692_));
 sg13g2_inv_1 _5491_ (.Y(_1871_),
    .A(_1870_));
 sg13g2_nand2_1 _5492_ (.Y(_1872_),
    .A(_1692_),
    .B(_1852_));
 sg13g2_a21oi_1 _5493_ (.A1(_1871_),
    .A2(_1872_),
    .Y(_1873_),
    .B1(_1700_));
 sg13g2_nor2b_1 _5494_ (.A(_1858_),
    .B_N(_1538_),
    .Y(_1874_));
 sg13g2_nand2_1 _5495_ (.Y(_1875_),
    .A(_1275_),
    .B(net98));
 sg13g2_a21oi_1 _5496_ (.A1(_1857_),
    .A2(_1875_),
    .Y(_1876_),
    .B1(_1870_));
 sg13g2_nor3_1 _5497_ (.A(_1686_),
    .B(_1532_),
    .C(_1876_),
    .Y(_1877_));
 sg13g2_nor3_1 _5498_ (.A(_1873_),
    .B(_1874_),
    .C(_1877_),
    .Y(_1878_));
 sg13g2_a21oi_1 _5499_ (.A1(_1878_),
    .A2(_1539_),
    .Y(_1879_),
    .B1(_1529_));
 sg13g2_o21ai_1 _5500_ (.B1(_1879_),
    .Y(_1880_),
    .A1(_1539_),
    .A2(_1869_));
 sg13g2_nand2b_1 _5501_ (.Y(_1881_),
    .B(_1529_),
    .A_N(_1876_));
 sg13g2_nand3_1 _5502_ (.B(net76),
    .C(_1881_),
    .A(_1880_),
    .Y(_1882_));
 sg13g2_nand2_1 _5503_ (.Y(_1883_),
    .A(_1882_),
    .B(_1513_));
 sg13g2_buf_1 _5504_ (.A(_1883_),
    .X(_1884_));
 sg13g2_a21oi_1 _5505_ (.A1(_1503_),
    .A2(_1851_),
    .Y(_1885_),
    .B1(net12));
 sg13g2_inv_1 _5506_ (.Y(_1886_),
    .A(_1385_));
 sg13g2_o21ai_1 _5507_ (.B1(\sqr_vol[0] ),
    .Y(_1887_),
    .A1(_1886_),
    .A2(net12));
 sg13g2_nand2b_1 _5508_ (.Y(_0182_),
    .B(_1887_),
    .A_N(_1885_));
 sg13g2_xnor2_1 _5509_ (.Y(_1888_),
    .A(_1405_),
    .B(\sqr_vol[1] ));
 sg13g2_xnor2_1 _5510_ (.Y(_1889_),
    .A(_1851_),
    .B(_1888_));
 sg13g2_inv_1 _5511_ (.Y(_1890_),
    .A(\sqr_vol[1] ));
 sg13g2_a22oi_1 _5512_ (.Y(_0183_),
    .B1(_1890_),
    .B2(net12),
    .A2(_1889_),
    .A1(_1516_));
 sg13g2_inv_1 _5513_ (.Y(_1891_),
    .A(\sqr_vol[2] ));
 sg13g2_nor2_1 _5514_ (.A(\sqr_vol[5] ),
    .B(_1891_),
    .Y(_1892_));
 sg13g2_inv_1 _5515_ (.Y(_1893_),
    .A(\sqr_vol[5] ));
 sg13g2_nor2_1 _5516_ (.A(\sqr_vol[2] ),
    .B(_1893_),
    .Y(_1894_));
 sg13g2_nor2_1 _5517_ (.A(_1892_),
    .B(_1894_),
    .Y(_1895_));
 sg13g2_nor2_1 _5518_ (.A(_1405_),
    .B(_1890_),
    .Y(_1896_));
 sg13g2_nand2_1 _5519_ (.Y(_1897_),
    .A(_1888_),
    .B(_1851_));
 sg13g2_nand2b_1 _5520_ (.Y(_1898_),
    .B(_1897_),
    .A_N(_1896_));
 sg13g2_xnor2_1 _5521_ (.Y(_1899_),
    .A(_1895_),
    .B(_1898_));
 sg13g2_a22oi_1 _5522_ (.Y(_0184_),
    .B1(_1891_),
    .B2(net12),
    .A2(_1899_),
    .A1(_1516_));
 sg13g2_nor2_1 _5523_ (.A(_1896_),
    .B(_1892_),
    .Y(_1900_));
 sg13g2_a21oi_1 _5524_ (.A1(_1897_),
    .A2(_1900_),
    .Y(_1901_),
    .B1(_1894_));
 sg13g2_nor3_1 _5525_ (.A(_1385_),
    .B(_1901_),
    .C(net12),
    .Y(_1902_));
 sg13g2_o21ai_1 _5526_ (.B1(_1385_),
    .Y(_1903_),
    .A1(_1901_),
    .A2(net12));
 sg13g2_nand3_1 _5527_ (.B(_1513_),
    .C(net76),
    .A(_1882_),
    .Y(_1904_));
 sg13g2_nand3b_1 _5528_ (.B(_1903_),
    .C(_1904_),
    .Y(_0185_),
    .A_N(_1902_));
 sg13g2_nand2b_1 _5529_ (.Y(_1905_),
    .B(_1886_),
    .A_N(_1901_));
 sg13g2_nor3_1 _5530_ (.A(_1405_),
    .B(_1905_),
    .C(net12),
    .Y(_1906_));
 sg13g2_o21ai_1 _5531_ (.B1(_1405_),
    .Y(_1907_),
    .A1(_1905_),
    .A2(net12));
 sg13g2_nand3b_1 _5532_ (.B(_1907_),
    .C(_1904_),
    .Y(_0186_),
    .A_N(_1906_));
 sg13g2_nor3_1 _5533_ (.A(_1405_),
    .B(_1905_),
    .C(_1884_),
    .Y(_1908_));
 sg13g2_o21ai_1 _5534_ (.B1(_1904_),
    .Y(_0187_),
    .A1(_1893_),
    .A2(_1908_));
 sg13g2_buf_1 _5535_ (.A(_1218_),
    .X(_1909_));
 sg13g2_inv_1 _5536_ (.Y(_1910_),
    .A(_0011_));
 sg13g2_o21ai_1 _5537_ (.B1(_1230_),
    .Y(_1911_),
    .A1(net103),
    .A2(net95));
 sg13g2_nor2_1 _5538_ (.A(net106),
    .B(_1248_),
    .Y(_1912_));
 sg13g2_inv_1 _5539_ (.Y(_1913_),
    .A(_1912_));
 sg13g2_nor2_1 _5540_ (.A(net109),
    .B(_2616_),
    .Y(_1914_));
 sg13g2_a21oi_1 _5541_ (.A1(_1285_),
    .A2(_1914_),
    .Y(_1915_),
    .B1(_1310_));
 sg13g2_a22oi_1 _5542_ (.Y(_1916_),
    .B1(_1913_),
    .B2(_1915_),
    .A2(_1911_),
    .A1(_1310_));
 sg13g2_nand2_1 _5543_ (.Y(_1917_),
    .A(_1916_),
    .B(_1227_));
 sg13g2_o21ai_1 _5544_ (.B1(net103),
    .Y(_1918_),
    .A1(net106),
    .A2(net110));
 sg13g2_nand3_1 _5545_ (.B(_1918_),
    .C(_1306_),
    .A(_1913_),
    .Y(_1919_));
 sg13g2_inv_1 _5546_ (.Y(_1920_),
    .A(_1310_));
 sg13g2_a21oi_1 _5547_ (.A1(net97),
    .A2(_1230_),
    .Y(_1921_),
    .B1(_1920_));
 sg13g2_a21oi_1 _5548_ (.A1(_1919_),
    .A2(_1920_),
    .Y(_1922_),
    .B1(_1921_));
 sg13g2_nor2b_1 _5549_ (.A(_1226_),
    .B_N(_1922_),
    .Y(_1923_));
 sg13g2_xnor2_1 _5550_ (.Y(_1924_),
    .A(net98),
    .B(_1282_));
 sg13g2_nor2_1 _5551_ (.A(_2626_),
    .B(_1853_),
    .Y(_1925_));
 sg13g2_nor2_1 _5552_ (.A(net91),
    .B(_1925_),
    .Y(_1926_));
 sg13g2_a22oi_1 _5553_ (.Y(_1927_),
    .B1(_1273_),
    .B2(_1926_),
    .A2(_1244_),
    .A1(net91));
 sg13g2_nor2_1 _5554_ (.A(_1310_),
    .B(_1927_),
    .Y(_1928_));
 sg13g2_a21oi_1 _5555_ (.A1(_1310_),
    .A2(_1924_),
    .Y(_1929_),
    .B1(_1928_));
 sg13g2_a21oi_1 _5556_ (.A1(_1923_),
    .A2(_1929_),
    .Y(_1930_),
    .B1(_1344_));
 sg13g2_a22oi_1 _5557_ (.Y(_1931_),
    .B1(_1917_),
    .B2(_1930_),
    .A2(_1344_),
    .A1(_1910_));
 sg13g2_nor2_1 _5558_ (.A(net64),
    .B(_1931_),
    .Y(_1932_));
 sg13g2_xor2_1 _5559_ (.B(_1932_),
    .A(\bass_pha[0] ),
    .X(_0071_));
 sg13g2_buf_1 _5560_ (.A(\bass_pha[10] ),
    .X(_1933_));
 sg13g2_inv_1 _5561_ (.Y(_1934_),
    .A(\bass_pha[8] ));
 sg13g2_nor3_1 _5562_ (.A(_1769_),
    .B(_1934_),
    .C(net101),
    .Y(_1935_));
 sg13g2_a21oi_1 _5563_ (.A1(net85),
    .A2(_1762_),
    .Y(_1936_),
    .B1(\bass_pha[8] ));
 sg13g2_nor2_1 _5564_ (.A(_1935_),
    .B(_1936_),
    .Y(_1937_));
 sg13g2_inv_1 _5565_ (.Y(_1938_),
    .A(_1937_));
 sg13g2_inv_1 _5566_ (.Y(_1939_),
    .A(\bass_pha[4] ));
 sg13g2_a21oi_1 _5567_ (.A1(_1923_),
    .A2(_1917_),
    .Y(_1940_),
    .B1(net85));
 sg13g2_a21o_1 _5568_ (.A2(net85),
    .A1(_0015_),
    .B1(_1940_),
    .X(_1941_));
 sg13g2_nor2_1 _5569_ (.A(_1939_),
    .B(_1941_),
    .Y(_1942_));
 sg13g2_inv_1 _5570_ (.Y(_1943_),
    .A(_1923_));
 sg13g2_inv_1 _5571_ (.Y(_1944_),
    .A(_1917_));
 sg13g2_a21oi_1 _5572_ (.A1(_1943_),
    .A2(_1944_),
    .Y(_1945_),
    .B1(net85));
 sg13g2_a21oi_1 _5573_ (.A1(_0016_),
    .A2(net85),
    .Y(_1946_),
    .B1(_1945_));
 sg13g2_nor2_1 _5574_ (.A(\bass_pha[5] ),
    .B(_1946_),
    .Y(_1947_));
 sg13g2_nand2_1 _5575_ (.Y(_1948_),
    .A(_1946_),
    .B(\bass_pha[5] ));
 sg13g2_nor2b_1 _5576_ (.A(_1947_),
    .B_N(_1948_),
    .Y(_1949_));
 sg13g2_nand2_1 _5577_ (.Y(_1950_),
    .A(_1944_),
    .B(_1929_));
 sg13g2_nand2_1 _5578_ (.Y(_1951_),
    .A(_1950_),
    .B(_1943_));
 sg13g2_nand2_1 _5579_ (.Y(_1952_),
    .A(_1951_),
    .B(_1940_));
 sg13g2_o21ai_1 _5580_ (.B1(_1952_),
    .Y(_1953_),
    .A1(_0014_),
    .A2(net101));
 sg13g2_nor2_1 _5581_ (.A(\bass_pha[3] ),
    .B(_1953_),
    .Y(_1954_));
 sg13g2_inv_1 _5582_ (.Y(_1955_),
    .A(\bass_pha[1] ));
 sg13g2_a21o_1 _5583_ (.A2(_1344_),
    .A1(_0012_),
    .B1(_1930_),
    .X(_1956_));
 sg13g2_nor2_1 _5584_ (.A(_1955_),
    .B(_1956_),
    .Y(_1957_));
 sg13g2_nand2b_1 _5585_ (.Y(_1958_),
    .B(\bass_pha[0] ),
    .A_N(_1931_));
 sg13g2_xnor2_1 _5586_ (.Y(_1959_),
    .A(\bass_pha[1] ),
    .B(_1956_));
 sg13g2_inv_1 _5587_ (.Y(_1960_),
    .A(_1959_));
 sg13g2_nor2_1 _5588_ (.A(_1958_),
    .B(_1960_),
    .Y(_1961_));
 sg13g2_nor2_1 _5589_ (.A(_1957_),
    .B(_1961_),
    .Y(_1962_));
 sg13g2_inv_1 _5590_ (.Y(_1963_),
    .A(_1962_));
 sg13g2_inv_1 _5591_ (.Y(_1964_),
    .A(_0013_));
 sg13g2_nand2_1 _5592_ (.Y(_1965_),
    .A(_1930_),
    .B(_1950_));
 sg13g2_o21ai_1 _5593_ (.B1(_1965_),
    .Y(_1966_),
    .A1(_1964_),
    .A2(net101));
 sg13g2_xnor2_1 _5594_ (.Y(_1967_),
    .A(\bass_pha[2] ),
    .B(_1966_));
 sg13g2_inv_1 _5595_ (.Y(_1968_),
    .A(\bass_pha[2] ));
 sg13g2_nor2_1 _5596_ (.A(_1968_),
    .B(_1966_),
    .Y(_1969_));
 sg13g2_a21oi_1 _5597_ (.A1(_1963_),
    .A2(_1967_),
    .Y(_1970_),
    .B1(_1969_));
 sg13g2_nand2_1 _5598_ (.Y(_1971_),
    .A(_1953_),
    .B(\bass_pha[3] ));
 sg13g2_o21ai_1 _5599_ (.B1(_1971_),
    .Y(_1972_),
    .A1(_1954_),
    .A2(_1970_));
 sg13g2_buf_1 _5600_ (.A(_1972_),
    .X(_1973_));
 sg13g2_inv_1 _5601_ (.Y(_1974_),
    .A(_1949_));
 sg13g2_nand2_1 _5602_ (.Y(_1975_),
    .A(_1941_),
    .B(_1939_));
 sg13g2_inv_1 _5603_ (.Y(_1976_),
    .A(_1975_));
 sg13g2_nor2_1 _5604_ (.A(_1942_),
    .B(_1976_),
    .Y(_1977_));
 sg13g2_nor2b_1 _5605_ (.A(_1974_),
    .B_N(_1977_),
    .Y(_1978_));
 sg13g2_inv_1 _5606_ (.Y(_1979_),
    .A(_1948_));
 sg13g2_a221oi_1 _5607_ (.B2(_1978_),
    .C1(_1979_),
    .B1(_1973_),
    .A1(_1942_),
    .Y(_1980_),
    .A2(_1949_));
 sg13g2_inv_1 _5608_ (.Y(_1981_),
    .A(_1980_));
 sg13g2_inv_1 _5609_ (.Y(_1982_),
    .A(\bass_pha[6] ));
 sg13g2_inv_1 _5610_ (.Y(_1983_),
    .A(_0017_));
 sg13g2_nor2_1 _5611_ (.A(_1226_),
    .B(_1929_),
    .Y(_1984_));
 sg13g2_nor2_1 _5612_ (.A(_1944_),
    .B(_1984_),
    .Y(_1985_));
 sg13g2_nand3_1 _5613_ (.B(net101),
    .C(_1943_),
    .A(_1985_),
    .Y(_1986_));
 sg13g2_o21ai_1 _5614_ (.B1(_1986_),
    .Y(_1987_),
    .A1(_1983_),
    .A2(net101));
 sg13g2_nor2_1 _5615_ (.A(_1982_),
    .B(_1987_),
    .Y(_1988_));
 sg13g2_inv_1 _5616_ (.Y(_1989_),
    .A(_1988_));
 sg13g2_nand2_1 _5617_ (.Y(_1990_),
    .A(_1987_),
    .B(_1982_));
 sg13g2_nand2_1 _5618_ (.Y(_1991_),
    .A(_1989_),
    .B(_1990_));
 sg13g2_o21ai_1 _5619_ (.B1(_1986_),
    .Y(_1992_),
    .A1(_0018_),
    .A2(net101));
 sg13g2_nor2_1 _5620_ (.A(\bass_pha[7] ),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nand2_1 _5621_ (.Y(_1994_),
    .A(_1992_),
    .B(\bass_pha[7] ));
 sg13g2_nand2b_1 _5622_ (.Y(_1995_),
    .B(_1994_),
    .A_N(_1993_));
 sg13g2_nor2_1 _5623_ (.A(_1991_),
    .B(_1995_),
    .Y(_1996_));
 sg13g2_a21oi_1 _5624_ (.A1(_1989_),
    .A2(_1994_),
    .Y(_1997_),
    .B1(_1993_));
 sg13g2_a21oi_1 _5625_ (.A1(_1981_),
    .A2(_1996_),
    .Y(_1998_),
    .B1(_1997_));
 sg13g2_nor2_1 _5626_ (.A(_1938_),
    .B(_1998_),
    .Y(_1999_));
 sg13g2_nor2_1 _5627_ (.A(_1935_),
    .B(_1999_),
    .Y(_2000_));
 sg13g2_nor2_1 _5628_ (.A(_0019_),
    .B(_2000_),
    .Y(_2001_));
 sg13g2_buf_1 _5629_ (.A(_1217_),
    .X(_2002_));
 sg13g2_nand2_1 _5630_ (.Y(_2003_),
    .A(_2001_),
    .B(net69));
 sg13g2_xnor2_1 _5631_ (.Y(_0072_),
    .A(_1933_),
    .B(_2003_));
 sg13g2_nand2_1 _5632_ (.Y(_2004_),
    .A(_1933_),
    .B(\bass_pha[9] ));
 sg13g2_nor2_1 _5633_ (.A(_2004_),
    .B(_2000_),
    .Y(_2005_));
 sg13g2_nand2_1 _5634_ (.Y(_2006_),
    .A(_2005_),
    .B(net69));
 sg13g2_xnor2_1 _5635_ (.Y(_0073_),
    .A(\bass_pha[11] ),
    .B(_2006_));
 sg13g2_inv_1 _5636_ (.Y(_2007_),
    .A(\bass_pha[12] ));
 sg13g2_buf_1 _5637_ (.A(_1217_),
    .X(_2008_));
 sg13g2_nand3_1 _5638_ (.B(_1933_),
    .C(\bass_pha[11] ),
    .A(_2001_),
    .Y(_2009_));
 sg13g2_nand2b_1 _5639_ (.Y(_2010_),
    .B(_1322_),
    .A_N(_2009_));
 sg13g2_nand2_1 _5640_ (.Y(_2011_),
    .A(_2009_),
    .B(_0020_));
 sg13g2_nand3_1 _5641_ (.B(_2011_),
    .C(net69),
    .A(_2010_),
    .Y(_2012_));
 sg13g2_o21ai_1 _5642_ (.B1(_2012_),
    .Y(_0074_),
    .A1(_2007_),
    .A2(net68));
 sg13g2_inv_1 _5643_ (.Y(_2013_),
    .A(\bass_pha[13] ));
 sg13g2_nand2_1 _5644_ (.Y(_2014_),
    .A(\bass_pha[11] ),
    .B(\bass_pha[12] ));
 sg13g2_inv_1 _5645_ (.Y(_2015_),
    .A(_2005_));
 sg13g2_o21ai_1 _5646_ (.B1(_0021_),
    .Y(_2016_),
    .A1(_2014_),
    .A2(_2015_));
 sg13g2_buf_1 _5647_ (.A(_1217_),
    .X(_2017_));
 sg13g2_inv_1 _5648_ (.Y(_2018_),
    .A(_2014_));
 sg13g2_nand3_1 _5649_ (.B(_1315_),
    .C(_2018_),
    .A(_2005_),
    .Y(_2019_));
 sg13g2_nand3_1 _5650_ (.B(net67),
    .C(_2019_),
    .A(_2016_),
    .Y(_2020_));
 sg13g2_o21ai_1 _5651_ (.B1(_2020_),
    .Y(_0075_),
    .A1(_2013_),
    .A2(net68));
 sg13g2_nand3_1 _5652_ (.B(_1933_),
    .C(\bass_pha[13] ),
    .A(_2018_),
    .Y(_2021_));
 sg13g2_inv_1 _5653_ (.Y(_2022_),
    .A(_2001_));
 sg13g2_nor2_1 _5654_ (.A(_2021_),
    .B(_2022_),
    .Y(_2023_));
 sg13g2_xor2_1 _5655_ (.B(_2023_),
    .A(_0022_),
    .X(_2024_));
 sg13g2_nor2_1 _5656_ (.A(\bass_pha[14] ),
    .B(net67),
    .Y(_2025_));
 sg13g2_a21oi_1 _5657_ (.A1(_2024_),
    .A2(net68),
    .Y(_0076_),
    .B1(_2025_));
 sg13g2_nand3_1 _5658_ (.B(\bass_pha[13] ),
    .C(\bass_pha[14] ),
    .A(_2018_),
    .Y(_2026_));
 sg13g2_nor2_1 _5659_ (.A(_2026_),
    .B(_2015_),
    .Y(_2027_));
 sg13g2_xnor2_1 _5660_ (.Y(_2028_),
    .A(_1331_),
    .B(_2027_));
 sg13g2_nor2_1 _5661_ (.A(\bass_pha[15] ),
    .B(net67),
    .Y(_2029_));
 sg13g2_a21oi_1 _5662_ (.A1(_2028_),
    .A2(net68),
    .Y(_0077_),
    .B1(_2029_));
 sg13g2_buf_1 _5663_ (.A(_1217_),
    .X(_2030_));
 sg13g2_nand2_1 _5664_ (.Y(_2031_),
    .A(_1960_),
    .B(_1958_));
 sg13g2_nand3b_1 _5665_ (.B(net69),
    .C(_2031_),
    .Y(_2032_),
    .A_N(_1961_));
 sg13g2_o21ai_1 _5666_ (.B1(_2032_),
    .Y(_0078_),
    .A1(_1955_),
    .A2(net66));
 sg13g2_a21oi_1 _5667_ (.A1(_1963_),
    .A2(_1967_),
    .Y(_2033_),
    .B1(net64));
 sg13g2_o21ai_1 _5668_ (.B1(_2033_),
    .Y(_2034_),
    .A1(_1963_),
    .A2(_1967_));
 sg13g2_o21ai_1 _5669_ (.B1(_2034_),
    .Y(_0079_),
    .A1(_1968_),
    .A2(_2030_));
 sg13g2_nand2b_1 _5670_ (.Y(_2035_),
    .B(_1971_),
    .A_N(_1954_));
 sg13g2_xnor2_1 _5671_ (.Y(_2036_),
    .A(_2035_),
    .B(_1970_));
 sg13g2_nor2_1 _5672_ (.A(\bass_pha[3] ),
    .B(net67),
    .Y(_2037_));
 sg13g2_a21oi_1 _5673_ (.A1(_2036_),
    .A2(net68),
    .Y(_0080_),
    .B1(_2037_));
 sg13g2_a21oi_1 _5674_ (.A1(_1973_),
    .A2(_1977_),
    .Y(_2038_),
    .B1(net64));
 sg13g2_o21ai_1 _5675_ (.B1(_2038_),
    .Y(_2039_),
    .A1(_1977_),
    .A2(_1973_));
 sg13g2_o21ai_1 _5676_ (.B1(_2039_),
    .Y(_0081_),
    .A1(_1939_),
    .A2(net66));
 sg13g2_a21oi_1 _5677_ (.A1(_1973_),
    .A2(_1975_),
    .Y(_2040_),
    .B1(_1942_));
 sg13g2_xnor2_1 _5678_ (.Y(_2041_),
    .A(_1974_),
    .B(_2040_));
 sg13g2_nor2_1 _5679_ (.A(\bass_pha[5] ),
    .B(net67),
    .Y(_2042_));
 sg13g2_a21oi_1 _5680_ (.A1(_2041_),
    .A2(net68),
    .Y(_0082_),
    .B1(_2042_));
 sg13g2_o21ai_1 _5681_ (.B1(_1217_),
    .Y(_2043_),
    .A1(_1991_),
    .A2(_1980_));
 sg13g2_a21oi_1 _5682_ (.A1(_1991_),
    .A2(_1980_),
    .Y(_2044_),
    .B1(_2043_));
 sg13g2_a21o_1 _5683_ (.A2(_1909_),
    .A1(\bass_pha[6] ),
    .B1(_2044_),
    .X(_0083_));
 sg13g2_nor2_1 _5684_ (.A(_1979_),
    .B(_1988_),
    .Y(_2045_));
 sg13g2_o21ai_1 _5685_ (.B1(_2045_),
    .Y(_2046_),
    .A1(_1974_),
    .A2(_2040_));
 sg13g2_nand2_1 _5686_ (.Y(_2047_),
    .A(_2046_),
    .B(_1990_));
 sg13g2_o21ai_1 _5687_ (.B1(_1217_),
    .Y(_2048_),
    .A1(_1995_),
    .A2(_2047_));
 sg13g2_a21oi_1 _5688_ (.A1(_1995_),
    .A2(_2047_),
    .Y(_2049_),
    .B1(_2048_));
 sg13g2_a21o_1 _5689_ (.A2(net64),
    .A1(\bass_pha[7] ),
    .B1(_2049_),
    .X(_0084_));
 sg13g2_nand2_1 _5690_ (.Y(_2050_),
    .A(_1998_),
    .B(_1938_));
 sg13g2_nand3b_1 _5691_ (.B(_2002_),
    .C(_2050_),
    .Y(_2051_),
    .A_N(_1999_));
 sg13g2_o21ai_1 _5692_ (.B1(_2051_),
    .Y(_0085_),
    .A1(_1934_),
    .A2(_2030_));
 sg13g2_inv_1 _5693_ (.Y(_2052_),
    .A(\bass_pha[9] ));
 sg13g2_nand2_1 _5694_ (.Y(_2053_),
    .A(_2000_),
    .B(_0019_));
 sg13g2_nand3_1 _5695_ (.B(_2053_),
    .C(net69),
    .A(_2022_),
    .Y(_2054_));
 sg13g2_o21ai_1 _5696_ (.B1(_2054_),
    .Y(_0086_),
    .A1(_2052_),
    .A2(net66));
 sg13g2_inv_1 _5697_ (.Y(_2055_),
    .A(\sqr_pha[0] ));
 sg13g2_nor2_1 _5698_ (.A(net103),
    .B(_1286_),
    .Y(_2056_));
 sg13g2_inv_1 _5699_ (.Y(_2057_),
    .A(_2056_));
 sg13g2_a22oi_1 _5700_ (.Y(_2058_),
    .B1(net95),
    .B2(_1233_),
    .A2(_1719_),
    .A1(_1914_));
 sg13g2_a21oi_1 _5701_ (.A1(_1276_),
    .A2(_2057_),
    .Y(_2059_),
    .B1(_2058_));
 sg13g2_inv_1 _5702_ (.Y(_2060_),
    .A(_1254_));
 sg13g2_nand2_1 _5703_ (.Y(_2061_),
    .A(_2060_),
    .B(_1244_));
 sg13g2_nor2_1 _5704_ (.A(net106),
    .B(_1856_),
    .Y(_2062_));
 sg13g2_nand2_1 _5705_ (.Y(_2063_),
    .A(_1275_),
    .B(net96));
 sg13g2_nand3_1 _5706_ (.B(_2062_),
    .C(_2063_),
    .A(_2061_),
    .Y(_2064_));
 sg13g2_nor2b_1 _5707_ (.A(_2059_),
    .B_N(_2064_),
    .Y(_2065_));
 sg13g2_and2_1 _5708_ (.A(_1229_),
    .B(_1232_),
    .X(_2066_));
 sg13g2_a21oi_1 _5709_ (.A1(_2066_),
    .A2(_1292_),
    .Y(_2067_),
    .B1(_1283_));
 sg13g2_nor2_1 _5710_ (.A(net104),
    .B(_2305_),
    .Y(_2068_));
 sg13g2_a21oi_1 _5711_ (.A1(_2068_),
    .A2(_2317_),
    .Y(_2069_),
    .B1(net95));
 sg13g2_nor3_1 _5712_ (.A(net84),
    .B(_1270_),
    .C(_1277_),
    .Y(_2070_));
 sg13g2_nand2b_1 _5713_ (.Y(_2071_),
    .B(_1261_),
    .A_N(_2066_));
 sg13g2_o21ai_1 _5714_ (.B1(_2071_),
    .Y(_2072_),
    .A1(_2069_),
    .A2(_2070_));
 sg13g2_a22oi_1 _5715_ (.Y(_2073_),
    .B1(_2067_),
    .B2(_2072_),
    .A2(_2065_),
    .A1(_1279_));
 sg13g2_o21ai_1 _5716_ (.B1(_1247_),
    .Y(_2074_),
    .A1(net98),
    .A2(_2056_));
 sg13g2_nor3_1 _5717_ (.A(net119),
    .B(_1257_),
    .C(_2340_),
    .Y(_2075_));
 sg13g2_nand2_1 _5718_ (.Y(_2076_),
    .A(_1229_),
    .B(_1697_));
 sg13g2_nand3_1 _5719_ (.B(net84),
    .C(_1277_),
    .A(_2076_),
    .Y(_2077_));
 sg13g2_nand3_1 _5720_ (.B(_2075_),
    .C(_2077_),
    .A(_2074_),
    .Y(_2078_));
 sg13g2_nand2b_1 _5721_ (.Y(_2079_),
    .B(_2060_),
    .A_N(_1696_));
 sg13g2_o21ai_1 _5722_ (.B1(_2061_),
    .Y(_2080_),
    .A1(_2627_),
    .A2(_2079_));
 sg13g2_nand2_1 _5723_ (.Y(_2081_),
    .A(_2080_),
    .B(net84));
 sg13g2_a21o_1 _5724_ (.A2(_2626_),
    .A1(_2317_),
    .B1(_2068_),
    .X(_2082_));
 sg13g2_nand4_1 _5725_ (.B(_2686_),
    .C(_1234_),
    .A(_2082_),
    .Y(_2083_),
    .D(_1852_));
 sg13g2_nand3_1 _5726_ (.B(_1304_),
    .C(_2083_),
    .A(_2081_),
    .Y(_2084_));
 sg13g2_nand3_1 _5727_ (.B(_2078_),
    .C(_2084_),
    .A(_2073_),
    .Y(_2085_));
 sg13g2_nand2_1 _5728_ (.Y(_2086_),
    .A(_2340_),
    .B(_2605_));
 sg13g2_nand3_1 _5729_ (.B(net98),
    .C(_1234_),
    .A(_1697_),
    .Y(_2087_));
 sg13g2_a221oi_1 _5730_ (.B2(net96),
    .C1(net84),
    .B1(_1683_),
    .A1(_1244_),
    .Y(_2088_),
    .A2(_1720_));
 sg13g2_a221oi_1 _5731_ (.B2(_2069_),
    .C1(_2088_),
    .B1(_2087_),
    .A1(_1290_),
    .Y(_2089_),
    .A2(_2086_));
 sg13g2_a21oi_2 _5732_ (.B1(_2089_),
    .Y(_2090_),
    .A2(_1290_),
    .A1(_2085_));
 sg13g2_o21ai_1 _5733_ (.B1(_1247_),
    .Y(_2091_),
    .A1(_1865_),
    .A2(_1251_));
 sg13g2_nand3_1 _5734_ (.B(net91),
    .C(_1232_),
    .A(_1925_),
    .Y(_2092_));
 sg13g2_nand3_1 _5735_ (.B(_1256_),
    .C(_2092_),
    .A(_2091_),
    .Y(_2093_));
 sg13g2_nand3_1 _5736_ (.B(net99),
    .C(_1534_),
    .A(_2093_),
    .Y(_2094_));
 sg13g2_a221oi_1 _5737_ (.B2(net99),
    .C1(_1223_),
    .B1(_1263_),
    .A1(_2056_),
    .Y(_2095_),
    .A2(_1231_));
 sg13g2_a21oi_1 _5738_ (.A1(_1281_),
    .A2(_1697_),
    .Y(_2096_),
    .B1(_1262_));
 sg13g2_o21ai_1 _5739_ (.B1(net119),
    .Y(_2097_),
    .A1(_1713_),
    .A2(_2096_));
 sg13g2_a21oi_1 _5740_ (.A1(_2095_),
    .A2(_2097_),
    .Y(_2098_),
    .B1(_1224_));
 sg13g2_a21oi_1 _5741_ (.A1(_2094_),
    .A2(_2098_),
    .Y(_2099_),
    .B1(net118));
 sg13g2_nand3_1 _5742_ (.B(net99),
    .C(net120),
    .A(_2093_),
    .Y(_2100_));
 sg13g2_nand2_1 _5743_ (.Y(_2101_),
    .A(_1253_),
    .B(_1246_));
 sg13g2_nand2_1 _5744_ (.Y(_2102_),
    .A(_2101_),
    .B(_2641_));
 sg13g2_o21ai_1 _5745_ (.B1(_2102_),
    .Y(_2103_),
    .A1(_1233_),
    .A2(_1719_));
 sg13g2_nand3_1 _5746_ (.B(_2641_),
    .C(net103),
    .A(_1269_),
    .Y(_2104_));
 sg13g2_a21oi_1 _5747_ (.A1(_1273_),
    .A2(_2104_),
    .Y(_2105_),
    .B1(net106));
 sg13g2_a21oi_1 _5748_ (.A1(_2103_),
    .A2(net95),
    .Y(_2106_),
    .B1(_2105_));
 sg13g2_a21oi_1 _5749_ (.A1(_2106_),
    .A2(net119),
    .Y(_2107_),
    .B1(_2337_));
 sg13g2_nor2_1 _5750_ (.A(net104),
    .B(_1914_),
    .Y(_2108_));
 sg13g2_nand3_1 _5751_ (.B(_1918_),
    .C(_2108_),
    .A(_1913_),
    .Y(_2109_));
 sg13g2_nand3_1 _5752_ (.B(_1223_),
    .C(_2109_),
    .A(_1238_),
    .Y(_2110_));
 sg13g2_nand3_1 _5753_ (.B(_2107_),
    .C(_2110_),
    .A(_2100_),
    .Y(_2111_));
 sg13g2_nand2_1 _5754_ (.Y(_2112_),
    .A(_2099_),
    .B(_2111_));
 sg13g2_o21ai_1 _5755_ (.B1(_1291_),
    .Y(_2113_),
    .A1(_1703_),
    .A2(_1293_));
 sg13g2_nand2_2 _5756_ (.Y(_2114_),
    .A(_2112_),
    .B(_2113_));
 sg13g2_inv_1 _5757_ (.Y(_2115_),
    .A(_2114_));
 sg13g2_nand2_1 _5758_ (.Y(_2116_),
    .A(_2090_),
    .B(_2115_));
 sg13g2_nand3_1 _5759_ (.B(net96),
    .C(_2615_),
    .A(_1693_),
    .Y(_2117_));
 sg13g2_o21ai_1 _5760_ (.B1(_2062_),
    .Y(_2118_),
    .A1(_1696_),
    .A2(_1233_));
 sg13g2_nand2_1 _5761_ (.Y(_2119_),
    .A(_1681_),
    .B(_1231_));
 sg13g2_nand3_1 _5762_ (.B(_2118_),
    .C(_2119_),
    .A(_2117_),
    .Y(_2120_));
 sg13g2_inv_1 _5763_ (.Y(_2121_),
    .A(_1856_));
 sg13g2_nor2_1 _5764_ (.A(_1275_),
    .B(_2121_),
    .Y(_2122_));
 sg13g2_and3_1 _5765_ (.X(_2123_),
    .A(_1261_),
    .B(_1242_),
    .C(_1232_));
 sg13g2_a22oi_1 _5766_ (.Y(_2124_),
    .B1(_1250_),
    .B2(_2123_),
    .A2(_2122_),
    .A1(_2618_));
 sg13g2_nand2b_1 _5767_ (.Y(_2125_),
    .B(_1247_),
    .A_N(_2101_));
 sg13g2_nand3_1 _5768_ (.B(_1252_),
    .C(_2125_),
    .A(_2124_),
    .Y(_2126_));
 sg13g2_nand2_1 _5769_ (.Y(_2127_),
    .A(_2126_),
    .B(_2075_));
 sg13g2_nor2_1 _5770_ (.A(_1243_),
    .B(_1228_),
    .Y(_2128_));
 sg13g2_o21ai_1 _5771_ (.B1(_2686_),
    .Y(_2129_),
    .A1(_1856_),
    .A2(_2128_));
 sg13g2_nand3_1 _5772_ (.B(net91),
    .C(_1235_),
    .A(_2082_),
    .Y(_2130_));
 sg13g2_nand3_1 _5773_ (.B(_2130_),
    .C(_1304_),
    .A(_2129_),
    .Y(_2131_));
 sg13g2_a21oi_1 _5774_ (.A1(_1703_),
    .A2(_1231_),
    .Y(_2132_),
    .B1(_2086_));
 sg13g2_nand3_1 _5775_ (.B(_2118_),
    .C(_2132_),
    .A(_2117_),
    .Y(_2133_));
 sg13g2_nand3_1 _5776_ (.B(_1290_),
    .C(_2133_),
    .A(_2131_),
    .Y(_2134_));
 sg13g2_nor2_1 _5777_ (.A(net106),
    .B(_1273_),
    .Y(_2135_));
 sg13g2_a21oi_1 _5778_ (.A1(_1275_),
    .A2(_2641_),
    .Y(_2136_),
    .B1(_2617_));
 sg13g2_o21ai_1 _5779_ (.B1(_2136_),
    .Y(_2137_),
    .A1(net96),
    .A2(_2079_));
 sg13g2_a21oi_1 _5780_ (.A1(_1282_),
    .A2(net96),
    .Y(_2138_),
    .B1(_2337_));
 sg13g2_nand2_1 _5781_ (.Y(_2139_),
    .A(_2137_),
    .B(_2138_));
 sg13g2_nor3_1 _5782_ (.A(net99),
    .B(_2135_),
    .C(_2139_),
    .Y(_2140_));
 sg13g2_nor2_1 _5783_ (.A(net96),
    .B(_1249_),
    .Y(_2141_));
 sg13g2_o21ai_1 _5784_ (.B1(net95),
    .Y(_2142_),
    .A1(net98),
    .A2(_1253_));
 sg13g2_a21oi_1 _5785_ (.A1(_2101_),
    .A2(_2141_),
    .Y(_2143_),
    .B1(_2142_));
 sg13g2_a221oi_1 _5786_ (.B2(net108),
    .C1(_1283_),
    .B1(_2135_),
    .A1(net91),
    .Y(_2144_),
    .A2(_2068_));
 sg13g2_nor2b_1 _5787_ (.A(_2143_),
    .B_N(_2144_),
    .Y(_2145_));
 sg13g2_nor3_1 _5788_ (.A(_2134_),
    .B(_2140_),
    .C(_2145_),
    .Y(_2146_));
 sg13g2_a22oi_1 _5789_ (.Y(_2147_),
    .B1(_2127_),
    .B2(_2146_),
    .A2(_2120_),
    .A1(_2342_));
 sg13g2_buf_2 _5790_ (.A(_2147_),
    .X(_2148_));
 sg13g2_nand2_1 _5791_ (.Y(_2149_),
    .A(_2116_),
    .B(_2148_));
 sg13g2_nor2_1 _5792_ (.A(_1909_),
    .B(_2149_),
    .Y(_2150_));
 sg13g2_xnor2_1 _5793_ (.Y(_0169_),
    .A(_2055_),
    .B(_2150_));
 sg13g2_nand2_2 _5794_ (.Y(_2151_),
    .A(_2148_),
    .B(_2090_));
 sg13g2_nor2_2 _5795_ (.A(_2115_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_xnor2_1 _5796_ (.Y(_2153_),
    .A(\sqr_pha[7] ),
    .B(_2152_));
 sg13g2_inv_1 _5797_ (.Y(_2154_),
    .A(\sqr_pha[6] ));
 sg13g2_xnor2_1 _5798_ (.Y(_2155_),
    .A(_2154_),
    .B(_2152_));
 sg13g2_nand2b_1 _5799_ (.Y(_2156_),
    .B(_2148_),
    .A_N(_2090_));
 sg13g2_nand2_1 _5800_ (.Y(_2157_),
    .A(_2148_),
    .B(_2115_));
 sg13g2_nand2_1 _5801_ (.Y(_2158_),
    .A(_2156_),
    .B(_2157_));
 sg13g2_nor2_1 _5802_ (.A(\sqr_pha[4] ),
    .B(_2158_),
    .Y(_2159_));
 sg13g2_inv_1 _5803_ (.Y(_2160_),
    .A(\sqr_pha[1] ));
 sg13g2_nor2_1 _5804_ (.A(_2114_),
    .B(_2151_),
    .Y(_2161_));
 sg13g2_xnor2_1 _5805_ (.Y(_2162_),
    .A(_2160_),
    .B(_2161_));
 sg13g2_nor2_1 _5806_ (.A(_2055_),
    .B(_2149_),
    .Y(_2163_));
 sg13g2_nand2_1 _5807_ (.Y(_2164_),
    .A(_2162_),
    .B(_2163_));
 sg13g2_inv_1 _5808_ (.Y(_2165_),
    .A(_2164_));
 sg13g2_nand2b_1 _5809_ (.Y(_2166_),
    .B(_2090_),
    .A_N(_2148_));
 sg13g2_nand2_1 _5810_ (.Y(_2167_),
    .A(_2166_),
    .B(_2116_));
 sg13g2_nor2_1 _5811_ (.A(\sqr_pha[2] ),
    .B(_2167_),
    .Y(_2168_));
 sg13g2_nand2_1 _5812_ (.Y(_2169_),
    .A(_2167_),
    .B(\sqr_pha[2] ));
 sg13g2_inv_1 _5813_ (.Y(_2170_),
    .A(_2169_));
 sg13g2_nor2_1 _5814_ (.A(_2168_),
    .B(_2170_),
    .Y(_2171_));
 sg13g2_nor3_1 _5815_ (.A(_2160_),
    .B(_2114_),
    .C(_2151_),
    .Y(_2172_));
 sg13g2_nor2_1 _5816_ (.A(_2172_),
    .B(_2170_),
    .Y(_2173_));
 sg13g2_inv_1 _5817_ (.Y(_2174_),
    .A(_2173_));
 sg13g2_a21oi_1 _5818_ (.A1(_2165_),
    .A2(_2171_),
    .Y(_2175_),
    .B1(_2174_));
 sg13g2_inv_1 _5819_ (.Y(_2176_),
    .A(_2175_));
 sg13g2_nand3_1 _5820_ (.B(_2114_),
    .C(_2156_),
    .A(_2166_),
    .Y(_2177_));
 sg13g2_nand2_1 _5821_ (.Y(_2178_),
    .A(_2177_),
    .B(_2157_));
 sg13g2_inv_1 _5822_ (.Y(_2179_),
    .A(\sqr_pha[3] ));
 sg13g2_nand2_1 _5823_ (.Y(_2180_),
    .A(_2178_),
    .B(_2179_));
 sg13g2_nor2_1 _5824_ (.A(_2179_),
    .B(_2178_),
    .Y(_2181_));
 sg13g2_a21oi_1 _5825_ (.A1(_2176_),
    .A2(_2180_),
    .Y(_2182_),
    .B1(_2181_));
 sg13g2_nand2_1 _5826_ (.Y(_2183_),
    .A(_2158_),
    .B(\sqr_pha[4] ));
 sg13g2_o21ai_1 _5827_ (.B1(_2183_),
    .Y(_2184_),
    .A1(_2159_),
    .A2(_2182_));
 sg13g2_inv_1 _5828_ (.Y(_2185_),
    .A(\sqr_pha[5] ));
 sg13g2_nand2_1 _5829_ (.Y(_2186_),
    .A(_2151_),
    .B(_2114_));
 sg13g2_xnor2_1 _5830_ (.Y(_2187_),
    .A(_2185_),
    .B(_2186_));
 sg13g2_inv_1 _5831_ (.Y(_2188_),
    .A(_2187_));
 sg13g2_nand2_1 _5832_ (.Y(_2189_),
    .A(_2184_),
    .B(_2188_));
 sg13g2_nor2_1 _5833_ (.A(_2185_),
    .B(_2186_),
    .Y(_2190_));
 sg13g2_nor2_1 _5834_ (.A(_2154_),
    .B(_2152_),
    .Y(_2191_));
 sg13g2_a21oi_1 _5835_ (.A1(_2190_),
    .A2(_2154_),
    .Y(_2192_),
    .B1(_2191_));
 sg13g2_o21ai_1 _5836_ (.B1(_2192_),
    .Y(_2193_),
    .A1(_2155_),
    .A2(_2189_));
 sg13g2_nand2b_1 _5837_ (.Y(_2194_),
    .B(_2193_),
    .A_N(_2153_));
 sg13g2_inv_1 _5838_ (.Y(_2195_),
    .A(\sqr_pha[7] ));
 sg13g2_inv_1 _5839_ (.Y(_2196_),
    .A(_2152_));
 sg13g2_nor2_1 _5840_ (.A(_2195_),
    .B(_2196_),
    .Y(_2197_));
 sg13g2_inv_1 _5841_ (.Y(_2198_),
    .A(_2197_));
 sg13g2_nand2_1 _5842_ (.Y(_2199_),
    .A(_2194_),
    .B(_2198_));
 sg13g2_nand3_1 _5843_ (.B(\sqr_pha[9] ),
    .C(\sqr_pha[8] ),
    .A(_2199_),
    .Y(_2200_));
 sg13g2_xnor2_1 _5844_ (.Y(_2201_),
    .A(_0025_),
    .B(_2200_));
 sg13g2_nor2_1 _5845_ (.A(\sqr_pha[10] ),
    .B(net67),
    .Y(_2202_));
 sg13g2_a21oi_1 _5846_ (.A1(_2201_),
    .A2(net68),
    .Y(_0170_),
    .B1(_2202_));
 sg13g2_inv_1 _5847_ (.Y(_2203_),
    .A(_2199_));
 sg13g2_nor2_1 _5848_ (.A(_0024_),
    .B(_2203_),
    .Y(_2204_));
 sg13g2_inv_1 _5849_ (.Y(_2205_),
    .A(_2204_));
 sg13g2_nor2_1 _5850_ (.A(_1241_),
    .B(_2205_),
    .Y(_2206_));
 sg13g2_xnor2_1 _5851_ (.Y(_2207_),
    .A(_1297_),
    .B(_2206_));
 sg13g2_nor2_1 _5852_ (.A(\sqr_pha[11] ),
    .B(_2017_),
    .Y(_2208_));
 sg13g2_a21oi_1 _5853_ (.A1(_2207_),
    .A2(_2008_),
    .Y(_0171_),
    .B1(_2208_));
 sg13g2_nand3b_1 _5854_ (.B(\sqr_pha[10] ),
    .C(\sqr_pha[11] ),
    .Y(_2209_),
    .A_N(_2200_));
 sg13g2_xnor2_1 _5855_ (.Y(_2210_),
    .A(_0027_),
    .B(_2209_));
 sg13g2_nor2_1 _5856_ (.A(\sqr_pha[12] ),
    .B(_2017_),
    .Y(_2211_));
 sg13g2_a21oi_1 _5857_ (.A1(_2210_),
    .A2(_2008_),
    .Y(_0172_),
    .B1(_2211_));
 sg13g2_nor2_1 _5858_ (.A(_2163_),
    .B(_2162_),
    .Y(_2212_));
 sg13g2_nand3b_1 _5859_ (.B(_2002_),
    .C(_2164_),
    .Y(_2213_),
    .A_N(_2212_));
 sg13g2_o21ai_1 _5860_ (.B1(_2213_),
    .Y(_0173_),
    .A1(_2160_),
    .A2(net66));
 sg13g2_nor2_1 _5861_ (.A(_2172_),
    .B(_2165_),
    .Y(_2214_));
 sg13g2_xor2_1 _5862_ (.B(_2214_),
    .A(_2171_),
    .X(_2215_));
 sg13g2_nor2_1 _5863_ (.A(\sqr_pha[2] ),
    .B(net67),
    .Y(_2216_));
 sg13g2_a21oi_1 _5864_ (.A1(_2215_),
    .A2(net68),
    .Y(_0174_),
    .B1(_2216_));
 sg13g2_nor2b_1 _5865_ (.A(_2181_),
    .B_N(_2180_),
    .Y(_2217_));
 sg13g2_xor2_1 _5866_ (.B(_2175_),
    .A(_2217_),
    .X(_2218_));
 sg13g2_nand2_1 _5867_ (.Y(_2219_),
    .A(net64),
    .B(\sqr_pha[3] ));
 sg13g2_o21ai_1 _5868_ (.B1(_2219_),
    .Y(_0175_),
    .A1(net64),
    .A2(_2218_));
 sg13g2_inv_1 _5869_ (.Y(_2220_),
    .A(\sqr_pha[4] ));
 sg13g2_inv_1 _5870_ (.Y(_2221_),
    .A(_2183_));
 sg13g2_nor2_1 _5871_ (.A(_2159_),
    .B(_2221_),
    .Y(_2222_));
 sg13g2_inv_1 _5872_ (.Y(_2223_),
    .A(_2182_));
 sg13g2_a21oi_1 _5873_ (.A1(_2223_),
    .A2(_2222_),
    .Y(_2224_),
    .B1(net64));
 sg13g2_o21ai_1 _5874_ (.B1(_2224_),
    .Y(_2225_),
    .A1(_2222_),
    .A2(_2223_));
 sg13g2_o21ai_1 _5875_ (.B1(_2225_),
    .Y(_0176_),
    .A1(_2220_),
    .A2(net66));
 sg13g2_nand2b_1 _5876_ (.Y(_2226_),
    .B(_2187_),
    .A_N(_2184_));
 sg13g2_nand3_1 _5877_ (.B(net67),
    .C(_2189_),
    .A(_2226_),
    .Y(_2227_));
 sg13g2_o21ai_1 _5878_ (.B1(_2227_),
    .Y(_0177_),
    .A1(_2185_),
    .A2(net66));
 sg13g2_nor3_1 _5879_ (.A(_2221_),
    .B(_2159_),
    .C(_2187_),
    .Y(_2228_));
 sg13g2_a221oi_1 _5880_ (.B2(_2228_),
    .C1(_2190_),
    .B1(_2223_),
    .A1(_2221_),
    .Y(_2229_),
    .A2(_2188_));
 sg13g2_o21ai_1 _5881_ (.B1(_1217_),
    .Y(_2230_),
    .A1(_2155_),
    .A2(_2229_));
 sg13g2_a21oi_1 _5882_ (.A1(_2155_),
    .A2(_2229_),
    .Y(_2231_),
    .B1(_2230_));
 sg13g2_a21o_1 _5883_ (.A2(net64),
    .A1(\sqr_pha[6] ),
    .B1(_2231_),
    .X(_0178_));
 sg13g2_nand2b_1 _5884_ (.Y(_2232_),
    .B(_2153_),
    .A_N(_2193_));
 sg13g2_nand3_1 _5885_ (.B(net69),
    .C(_2194_),
    .A(_2232_),
    .Y(_2233_));
 sg13g2_o21ai_1 _5886_ (.B1(_2233_),
    .Y(_0179_),
    .A1(_2195_),
    .A2(net66));
 sg13g2_inv_1 _5887_ (.Y(_2234_),
    .A(\sqr_pha[8] ));
 sg13g2_nand2_1 _5888_ (.Y(_2235_),
    .A(_2203_),
    .B(_0024_));
 sg13g2_nand3_1 _5889_ (.B(net69),
    .C(_2235_),
    .A(_2205_),
    .Y(_2236_));
 sg13g2_o21ai_1 _5890_ (.B1(_2236_),
    .Y(_0180_),
    .A1(_2234_),
    .A2(net66));
 sg13g2_nand2_1 _5891_ (.Y(_2237_),
    .A(_2204_),
    .B(net69));
 sg13g2_xnor2_1 _5892_ (.Y(_0181_),
    .A(\sqr_pha[9] ),
    .B(_2237_));
 sg13g2_nor2b_1 _5893_ (.A(net53),
    .B_N(_0042_),
    .Y(_0108_));
 sg13g2_nand3b_1 _5894_ (.B(_1653_),
    .C(_1637_),
    .Y(_2238_),
    .A_N(_1214_));
 sg13g2_inv_1 _5895_ (.Y(_0109_),
    .A(_2238_));
 sg13g2_nor2_1 _5896_ (.A(_2390_),
    .B(_1638_),
    .Y(_2239_));
 sg13g2_nor3_1 _5897_ (.A(_1640_),
    .B(_2239_),
    .C(net53),
    .Y(_0110_));
 sg13g2_nor2_1 _5898_ (.A(net116),
    .B(_1640_),
    .Y(_2240_));
 sg13g2_inv_1 _5899_ (.Y(_2241_),
    .A(_1641_));
 sg13g2_nor3_1 _5900_ (.A(_1213_),
    .B(_2240_),
    .C(_2241_),
    .Y(_0111_));
 sg13g2_nor2_1 _5901_ (.A(net117),
    .B(_2241_),
    .Y(_2242_));
 sg13g2_nor3_1 _5902_ (.A(_1213_),
    .B(_1642_),
    .C(_2242_),
    .Y(_0112_));
 sg13g2_nand2_1 _5903_ (.Y(_2243_),
    .A(_1642_),
    .B(_2415_));
 sg13g2_inv_1 _5904_ (.Y(_2244_),
    .A(_2243_));
 sg13g2_nor2_1 _5905_ (.A(_2415_),
    .B(_1642_),
    .Y(_2245_));
 sg13g2_nor3_1 _5906_ (.A(_2244_),
    .B(_2245_),
    .C(net53),
    .Y(_0113_));
 sg13g2_nor2_1 _5907_ (.A(_2434_),
    .B(_2243_),
    .Y(_2246_));
 sg13g2_nor2_1 _5908_ (.A(_2431_),
    .B(_2244_),
    .Y(_2247_));
 sg13g2_nor3_1 _5909_ (.A(_2246_),
    .B(_2247_),
    .C(net53),
    .Y(_0114_));
 sg13g2_nor2_1 _5910_ (.A(_2559_),
    .B(_2246_),
    .Y(_2248_));
 sg13g2_nand2_1 _5911_ (.Y(_2249_),
    .A(_2246_),
    .B(_2559_));
 sg13g2_inv_1 _5912_ (.Y(_2250_),
    .A(_2249_));
 sg13g2_nor3_1 _5913_ (.A(_2248_),
    .B(_2250_),
    .C(net53),
    .Y(_0115_));
 sg13g2_nor2_1 _5914_ (.A(_2583_),
    .B(_2249_),
    .Y(_2251_));
 sg13g2_nor2_1 _5915_ (.A(_2582_),
    .B(_2250_),
    .Y(_2252_));
 sg13g2_nor3_1 _5916_ (.A(net53),
    .B(_2251_),
    .C(_2252_),
    .Y(_0116_));
 sg13g2_nor3_1 _5917_ (.A(_2583_),
    .B(_1040_),
    .C(_2249_),
    .Y(_2253_));
 sg13g2_nor2_1 _5918_ (.A(_2598_),
    .B(_2251_),
    .Y(_2254_));
 sg13g2_nor3_1 _5919_ (.A(net53),
    .B(_2253_),
    .C(_2254_),
    .Y(_0117_));
 sg13g2_nor2_1 _5920_ (.A(\audio_pwm_accum[9] ),
    .B(_1447_),
    .Y(_2255_));
 sg13g2_nor2_1 _5921_ (.A(\audio_pwm_accum[7] ),
    .B(_1459_),
    .Y(_2256_));
 sg13g2_nor2_1 _5922_ (.A(\audio_pwm_accum[5] ),
    .B(\audio_sample_lpf[5] ),
    .Y(_2257_));
 sg13g2_nand2_1 _5923_ (.Y(_2258_),
    .A(\audio_pwm_accum[4] ),
    .B(\audio_sample_lpf[4] ));
 sg13g2_nand2_1 _5924_ (.Y(_2259_),
    .A(\audio_pwm_accum[5] ),
    .B(\audio_sample_lpf[5] ));
 sg13g2_nand2_1 _5925_ (.Y(_2260_),
    .A(_2258_),
    .B(_2259_));
 sg13g2_nor2_1 _5926_ (.A(\audio_pwm_accum[4] ),
    .B(\audio_sample_lpf[4] ),
    .Y(_2261_));
 sg13g2_nor2b_1 _5927_ (.A(_2261_),
    .B_N(_2258_),
    .Y(_2262_));
 sg13g2_inv_1 _5928_ (.Y(_2263_),
    .A(_2262_));
 sg13g2_nor2_1 _5929_ (.A(\audio_pwm_accum[3] ),
    .B(_1222_),
    .Y(_2264_));
 sg13g2_nand2_1 _5930_ (.Y(_2265_),
    .A(\audio_pwm_accum[0] ),
    .B(_1211_));
 sg13g2_xor2_1 _5931_ (.B(\audio_pwm_accum[1] ),
    .A(_1343_),
    .X(_2266_));
 sg13g2_inv_1 _5932_ (.Y(_2267_),
    .A(_2266_));
 sg13g2_nand2_1 _5933_ (.Y(_2268_),
    .A(_1343_),
    .B(\audio_pwm_accum[1] ));
 sg13g2_o21ai_1 _5934_ (.B1(_2268_),
    .Y(_2269_),
    .A1(_2265_),
    .A2(_2267_));
 sg13g2_xor2_1 _5935_ (.B(\audio_pwm_accum[2] ),
    .A(\audio_sample_lpf[2] ),
    .X(_2270_));
 sg13g2_and2_1 _5936_ (.A(_2269_),
    .B(_2270_),
    .X(_2271_));
 sg13g2_a21oi_1 _5937_ (.A1(\audio_sample_lpf[2] ),
    .A2(\audio_pwm_accum[2] ),
    .Y(_2272_),
    .B1(_2271_));
 sg13g2_nand2_1 _5938_ (.Y(_2273_),
    .A(\audio_pwm_accum[3] ),
    .B(_1222_));
 sg13g2_o21ai_1 _5939_ (.B1(_2273_),
    .Y(_2274_),
    .A1(_2264_),
    .A2(_2272_));
 sg13g2_inv_1 _5940_ (.Y(_2275_),
    .A(_2274_));
 sg13g2_nor2_1 _5941_ (.A(_2263_),
    .B(_2275_),
    .Y(_2276_));
 sg13g2_nor2_1 _5942_ (.A(_2260_),
    .B(_2276_),
    .Y(_2277_));
 sg13g2_nor2_1 _5943_ (.A(_2257_),
    .B(_2277_),
    .Y(_2278_));
 sg13g2_nor2_1 _5944_ (.A(\audio_pwm_accum[6] ),
    .B(_1446_),
    .Y(_2279_));
 sg13g2_nand2_1 _5945_ (.Y(_2280_),
    .A(\audio_pwm_accum[6] ),
    .B(_1446_));
 sg13g2_nor2b_1 _5946_ (.A(_2279_),
    .B_N(_2280_),
    .Y(_2281_));
 sg13g2_nand2_1 _5947_ (.Y(_2282_),
    .A(_2278_),
    .B(_2281_));
 sg13g2_nand2_1 _5948_ (.Y(_2283_),
    .A(\audio_pwm_accum[7] ),
    .B(_1459_));
 sg13g2_and3_1 _5949_ (.X(_2284_),
    .A(_2282_),
    .B(_2280_),
    .C(_2283_));
 sg13g2_nor2_1 _5950_ (.A(_2256_),
    .B(_2284_),
    .Y(_2285_));
 sg13g2_nor2_1 _5951_ (.A(\audio_pwm_accum[8] ),
    .B(_1474_),
    .Y(_2286_));
 sg13g2_nand2_1 _5952_ (.Y(_2287_),
    .A(\audio_pwm_accum[8] ),
    .B(_1474_));
 sg13g2_inv_1 _5953_ (.Y(_2288_),
    .A(_2287_));
 sg13g2_nor2_1 _5954_ (.A(_2286_),
    .B(_2288_),
    .Y(_2289_));
 sg13g2_a221oi_1 _5955_ (.B2(_2289_),
    .C1(_2288_),
    .B1(_2285_),
    .A1(\audio_pwm_accum[9] ),
    .Y(_2290_),
    .A2(_1447_));
 sg13g2_nor2_1 _5956_ (.A(_2255_),
    .B(_2290_),
    .Y(audio_pwm));
 sg13g2_xor2_1 _5957_ (.B(_1211_),
    .A(\audio_pwm_accum[0] ),
    .X(\audio_pwm_accum_next[0] ));
 sg13g2_xnor2_1 _5958_ (.Y(\audio_pwm_accum_next[1] ),
    .A(_2265_),
    .B(_2266_));
 sg13g2_xor2_1 _5959_ (.B(_2269_),
    .A(_2270_),
    .X(\audio_pwm_accum_next[2] ));
 sg13g2_nor2b_1 _5960_ (.A(_2264_),
    .B_N(_2273_),
    .Y(_2291_));
 sg13g2_xnor2_1 _5961_ (.Y(\audio_pwm_accum_next[3] ),
    .A(_2291_),
    .B(_2272_));
 sg13g2_xnor2_1 _5962_ (.Y(\audio_pwm_accum_next[4] ),
    .A(_2263_),
    .B(_2274_));
 sg13g2_nor2b_1 _5963_ (.A(_2257_),
    .B_N(_2259_),
    .Y(_2292_));
 sg13g2_o21ai_1 _5964_ (.B1(_2258_),
    .Y(_2293_),
    .A1(_2261_),
    .A2(_2275_));
 sg13g2_xor2_1 _5965_ (.B(_2293_),
    .A(_2292_),
    .X(\audio_pwm_accum_next[5] ));
 sg13g2_xor2_1 _5966_ (.B(_2278_),
    .A(_2281_),
    .X(\audio_pwm_accum_next[6] ));
 sg13g2_nor2b_1 _5967_ (.A(_2256_),
    .B_N(_2283_),
    .Y(_2294_));
 sg13g2_nand2_1 _5968_ (.Y(_2295_),
    .A(_2280_),
    .B(_2259_));
 sg13g2_a21oi_1 _5969_ (.A1(_2293_),
    .A2(_2292_),
    .Y(_2296_),
    .B1(_2295_));
 sg13g2_nor2_1 _5970_ (.A(_2279_),
    .B(_2296_),
    .Y(_2297_));
 sg13g2_xor2_1 _5971_ (.B(_2297_),
    .A(_2294_),
    .X(\audio_pwm_accum_next[7] ));
 sg13g2_xor2_1 _5972_ (.B(_2285_),
    .A(_2289_),
    .X(\audio_pwm_accum_next[8] ));
 sg13g2_xor2_1 _5973_ (.B(_1447_),
    .A(\audio_pwm_accum[9] ),
    .X(_2298_));
 sg13g2_nand2_1 _5974_ (.Y(_2299_),
    .A(_2287_),
    .B(_2283_));
 sg13g2_a21oi_1 _5975_ (.A1(_2297_),
    .A2(_2294_),
    .Y(_2300_),
    .B1(_2299_));
 sg13g2_nor2_1 _5976_ (.A(_2286_),
    .B(_2300_),
    .Y(_2301_));
 sg13g2_xor2_1 _5977_ (.B(_2301_),
    .A(_2298_),
    .X(\audio_pwm_accum_next[9] ));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _5987__154 (.L_HI(net154));
 sg13g2_buf_1 _5980_ (.A(net140),
    .X(uio_oe[0]));
 sg13g2_buf_1 _5981_ (.A(net141),
    .X(uio_oe[1]));
 sg13g2_buf_1 _5982_ (.A(net142),
    .X(uio_oe[2]));
 sg13g2_buf_1 _5983_ (.A(net143),
    .X(uio_oe[3]));
 sg13g2_buf_1 _5984_ (.A(net144),
    .X(uio_oe[4]));
 sg13g2_buf_1 _5985_ (.A(net145),
    .X(uio_oe[5]));
 sg13g2_buf_1 _5986_ (.A(net146),
    .X(uio_oe[6]));
 sg13g2_buf_1 _5987_ (.A(net154),
    .X(uio_oe[7]));
 sg13g2_buf_1 _5988_ (.A(net147),
    .X(uio_out[0]));
 sg13g2_buf_1 _5989_ (.A(net148),
    .X(uio_out[1]));
 sg13g2_buf_1 _5990_ (.A(net149),
    .X(uio_out[2]));
 sg13g2_buf_1 _5991_ (.A(net150),
    .X(uio_out[3]));
 sg13g2_buf_1 _5992_ (.A(net151),
    .X(uio_out[4]));
 sg13g2_buf_1 _5993_ (.A(net152),
    .X(uio_out[5]));
 sg13g2_buf_1 _5994_ (.A(net153),
    .X(uio_out[6]));
 sg13g2_buf_1 _5995_ (.A(audio_pwm),
    .X(net2));
 sg13g2_buf_1 _5996_ (.A(\hvsync_gen.vsync ),
    .X(net6));
 sg13g2_buf_1 _5997_ (.A(hsync),
    .X(net10));
 sg13g2_dfrbp_1 \audio_pwm_accum[0]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[0] ),
    .Q_N(_3044_),
    .Q(\audio_pwm_accum[0] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[1]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[1] ),
    .Q_N(_3045_),
    .Q(\audio_pwm_accum[1] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[2]$_DFF_PN0_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[2] ),
    .Q_N(_3046_),
    .Q(\audio_pwm_accum[2] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[3]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[3] ),
    .Q_N(_3047_),
    .Q(\audio_pwm_accum[3] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[4]$_DFF_PN0_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[4] ),
    .Q_N(_3048_),
    .Q(\audio_pwm_accum[4] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[5]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[5] ),
    .Q_N(_3049_),
    .Q(\audio_pwm_accum[5] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[6]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[6] ),
    .Q_N(_3050_),
    .Q(\audio_pwm_accum[6] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[7]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net136),
    .D(\audio_pwm_accum_next[7] ),
    .Q_N(_3051_),
    .Q(\audio_pwm_accum[7] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[8]$_DFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net137),
    .D(\audio_pwm_accum_next[8] ),
    .Q_N(_3052_),
    .Q(\audio_pwm_accum[8] ));
 sg13g2_dfrbp_1 \audio_pwm_accum[9]$_DFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net139),
    .D(\audio_pwm_accum_next[9] ),
    .Q_N(_3037_),
    .Q(\audio_pwm_accum[9] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[0]$_DFFE_PP_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net155),
    .D(_0061_),
    .Q_N(_3036_),
    .Q(\audio_sample_lpf[0] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[1]$_DFFE_PP_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net156),
    .D(_0062_),
    .Q_N(_3035_),
    .Q(\audio_sample_lpf[1] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[2]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net157),
    .D(_0063_),
    .Q_N(_0029_),
    .Q(\audio_sample_lpf[2] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[3]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net158),
    .D(_0064_),
    .Q_N(_0031_),
    .Q(\audio_sample_lpf[3] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[4]$_DFFE_PP_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net159),
    .D(_0065_),
    .Q_N(_0030_),
    .Q(\audio_sample_lpf[4] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[5]$_DFFE_PP_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net160),
    .D(_0066_),
    .Q_N(_0028_),
    .Q(\audio_sample_lpf[5] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[6]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net161),
    .D(_0067_),
    .Q_N(_0032_),
    .Q(\audio_sample_lpf[6] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[7]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net162),
    .D(_0068_),
    .Q_N(_0033_),
    .Q(\audio_sample_lpf[7] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[8]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net163),
    .D(_0069_),
    .Q_N(_0034_),
    .Q(\audio_sample_lpf[8] ));
 sg13g2_dfrbp_1 \audio_sample_lpf[9]$_DFFE_PP_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net164),
    .D(_0070_),
    .Q_N(_3034_),
    .Q(\audio_sample_lpf[9] ));
 sg13g2_dfrbp_1 \bass_pha[0]$_DFFE_PN0N_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net130),
    .D(_0071_),
    .Q_N(_3033_),
    .Q(\bass_pha[0] ));
 sg13g2_dfrbp_1 \bass_pha[10]$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net123),
    .D(_0072_),
    .Q_N(_3032_),
    .Q(\bass_pha[10] ));
 sg13g2_dfrbp_1 \bass_pha[11]$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net123),
    .D(_0073_),
    .Q_N(_3031_),
    .Q(\bass_pha[11] ));
 sg13g2_dfrbp_1 \bass_pha[12]$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net123),
    .D(_0074_),
    .Q_N(_0020_),
    .Q(\bass_pha[12] ));
 sg13g2_dfrbp_1 \bass_pha[13]$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net123),
    .D(_0075_),
    .Q_N(_0021_),
    .Q(\bass_pha[13] ));
 sg13g2_dfrbp_1 \bass_pha[14]$_DFFE_PN0N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net124),
    .D(_0076_),
    .Q_N(_0022_),
    .Q(\bass_pha[14] ));
 sg13g2_dfrbp_1 \bass_pha[15]$_DFFE_PN0N_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net124),
    .D(_0077_),
    .Q_N(_0023_),
    .Q(\bass_pha[15] ));
 sg13g2_dfrbp_1 \bass_pha[1]$_DFFE_PN0N_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net130),
    .D(_0078_),
    .Q_N(_3030_),
    .Q(\bass_pha[1] ));
 sg13g2_dfrbp_1 \bass_pha[2]$_DFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0079_),
    .Q_N(_3029_),
    .Q(\bass_pha[2] ));
 sg13g2_dfrbp_1 \bass_pha[3]$_DFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net124),
    .D(_0080_),
    .Q_N(_3028_),
    .Q(\bass_pha[3] ));
 sg13g2_dfrbp_1 \bass_pha[4]$_DFFE_PN0N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net123),
    .D(_0081_),
    .Q_N(_3027_),
    .Q(\bass_pha[4] ));
 sg13g2_dfrbp_1 \bass_pha[5]$_DFFE_PN0N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net124),
    .D(_0082_),
    .Q_N(_3026_),
    .Q(\bass_pha[5] ));
 sg13g2_dfrbp_1 \bass_pha[6]$_DFFE_PN0N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net124),
    .D(_0083_),
    .Q_N(_3025_),
    .Q(\bass_pha[6] ));
 sg13g2_dfrbp_1 \bass_pha[7]$_DFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net124),
    .D(_0084_),
    .Q_N(_3024_),
    .Q(\bass_pha[7] ));
 sg13g2_dfrbp_1 \bass_pha[8]$_DFFE_PN0N_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net130),
    .D(_0085_),
    .Q_N(_3023_),
    .Q(\bass_pha[8] ));
 sg13g2_dfrbp_1 \bass_pha[9]$_DFFE_PN0N_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net123),
    .D(_0086_),
    .Q_N(_0019_),
    .Q(\bass_pha[9] ));
 sg13g2_dfrbp_1 \bass_vol[0]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net135),
    .D(_0087_),
    .Q_N(_3022_),
    .Q(\bass_vol[0] ));
 sg13g2_dfrbp_1 \bass_vol[1]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net133),
    .D(_0088_),
    .Q_N(_3021_),
    .Q(\bass_vol[1] ));
 sg13g2_dfrbp_1 \bass_vol[2]$_DFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net135),
    .D(_0089_),
    .Q_N(_3020_),
    .Q(\bass_vol[2] ));
 sg13g2_dfrbp_1 \bass_vol[3]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net133),
    .D(_0090_),
    .Q_N(_3019_),
    .Q(\bass_vol[3] ));
 sg13g2_dfrbp_1 \bass_vol[4]$_DFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net133),
    .D(_0091_),
    .Q_N(_0010_),
    .Q(\bass_vol[4] ));
 sg13g2_dfrbp_1 \bass_vol[5]$_DFFE_PN0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net133),
    .D(_0092_),
    .Q_N(_3018_),
    .Q(\bass_vol[5] ));
 sg13g2_dfrbp_1 \cos[0]$_DFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net127),
    .D(_0093_),
    .Q_N(\cos[0] ),
    .Q(_0046_));
 sg13g2_dfrbp_1 \cos[1]$_DFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net127),
    .D(_0094_),
    .Q_N(\cos[1] ),
    .Q(_0047_));
 sg13g2_dfrbp_1 \cos[2]$_DFFE_PN1P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net127),
    .D(_0095_),
    .Q_N(\cos[2] ),
    .Q(_0048_));
 sg13g2_dfrbp_1 \cos[3]$_DFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net127),
    .D(_0096_),
    .Q_N(\cos[3] ),
    .Q(_0049_));
 sg13g2_dfrbp_1 \cos[4]$_DFFE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net128),
    .D(_0097_),
    .Q_N(\cos[4] ),
    .Q(_0050_));
 sg13g2_dfrbp_1 \cos[5]$_DFFE_PN1P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net127),
    .D(_0098_),
    .Q_N(\cos[5] ),
    .Q(_0051_));
 sg13g2_dfrbp_1 \cos[6]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net128),
    .D(_0099_),
    .Q_N(_3017_),
    .Q(\cos[6] ));
 sg13g2_dfrbp_1 \frame_count[0]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net131),
    .D(_0100_),
    .Q_N(_0045_),
    .Q(\frame_count[0] ));
 sg13g2_dfrbp_1 \frame_count[1]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net131),
    .D(_0101_),
    .Q_N(_3016_),
    .Q(\frame_count[1] ));
 sg13g2_dfrbp_1 \frame_count[2]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net131),
    .D(_0102_),
    .Q_N(_3015_),
    .Q(\frame_count[2] ));
 sg13g2_dfrbp_1 \frame_count[3]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net128),
    .D(_0103_),
    .Q_N(_3014_),
    .Q(\frame_count[3] ));
 sg13g2_dfrbp_1 \frame_count[4]$_DFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net128),
    .D(_0104_),
    .Q_N(_3013_),
    .Q(\frame_count[4] ));
 sg13g2_dfrbp_1 \frame_count[5]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net127),
    .D(_0105_),
    .Q_N(_3012_),
    .Q(\frame_count[5] ));
 sg13g2_dfrbp_1 \frame_count[6]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net127),
    .D(_0106_),
    .Q_N(_3011_),
    .Q(\frame_count[6] ));
 sg13g2_dfrbp_1 \frame_count[7]$_DFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net127),
    .D(_0107_),
    .Q_N(_3010_),
    .Q(\frame_count[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net165),
    .D(_0108_),
    .Q_N(_0042_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net166),
    .D(_0109_),
    .Q_N(_3009_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net167),
    .D(_0110_),
    .Q_N(_3008_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net168),
    .D(_0111_),
    .Q_N(_3007_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net169),
    .D(_0112_),
    .Q_N(_3006_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net170),
    .D(_0113_),
    .Q_N(_3005_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net171),
    .D(_0114_),
    .Q_N(_3004_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net172),
    .D(_0115_),
    .Q_N(_0038_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net173),
    .D(_0116_),
    .Q_N(_3003_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net174),
    .D(_0117_),
    .Q_N(_3053_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net175),
    .D(_0006_),
    .Q_N(_3002_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net176),
    .D(_0118_),
    .Q_N(_0043_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net177),
    .D(_0119_),
    .Q_N(_0036_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net178),
    .D(_0120_),
    .Q_N(_0037_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net179),
    .D(_0121_),
    .Q_N(_0009_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net180),
    .D(_0122_),
    .Q_N(_0039_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net181),
    .D(_0123_),
    .Q_N(_0041_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net182),
    .D(_0124_),
    .Q_N(_0040_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net183),
    .D(_0125_),
    .Q_N(_3001_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net184),
    .D(_0126_),
    .Q_N(_3000_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net185),
    .D(_0127_),
    .Q_N(_3054_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net186),
    .D(_0007_),
    .Q_N(_2999_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \kick_ctr[0]$_SDFFCE_PP1P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net187),
    .D(_0128_),
    .Q_N(_0044_),
    .Q(\kick_ctr[0] ));
 sg13g2_dfrbp_1 \kick_ctr[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net188),
    .D(_0129_),
    .Q_N(_2998_),
    .Q(\kick_ctr[1] ));
 sg13g2_dfrbp_1 \kick_osci[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net189),
    .D(_0130_),
    .Q_N(_0011_),
    .Q(\kick_osci[0] ));
 sg13g2_dfrbp_1 \kick_osci[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net190),
    .D(_0131_),
    .Q_N(_0012_),
    .Q(\kick_osci[1] ));
 sg13g2_dfrbp_1 \kick_osci[2]$_SDFFCE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net191),
    .D(_0132_),
    .Q_N(_0013_),
    .Q(\kick_osci[2] ));
 sg13g2_dfrbp_1 \kick_osci[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net192),
    .D(_0133_),
    .Q_N(_0014_),
    .Q(\kick_osci[3] ));
 sg13g2_dfrbp_1 \kick_osci[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net193),
    .D(_0134_),
    .Q_N(_0015_),
    .Q(\kick_osci[4] ));
 sg13g2_dfrbp_1 \kick_osci[5]$_SDFFCE_PP0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net194),
    .D(_0135_),
    .Q_N(_0016_),
    .Q(\kick_osci[5] ));
 sg13g2_dfrbp_1 \kick_osci[6]$_SDFFCE_PP0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net195),
    .D(_0136_),
    .Q_N(_0017_),
    .Q(\kick_osci[6] ));
 sg13g2_dfrbp_1 \kick_osci[7]$_SDFFCE_PP1P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net196),
    .D(_0137_),
    .Q_N(_0018_),
    .Q(\kick_osci[7] ));
 sg13g2_dfrbp_1 \kick_osci[8]$_SDFFCE_PP1P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net197),
    .D(_0138_),
    .Q_N(_2997_),
    .Q(\kick_osci[8] ));
 sg13g2_dfrbp_1 \line_lfsr[0]$_SDFFCE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net198),
    .D(_0139_),
    .Q_N(_2996_),
    .Q(\line_lfsr[0] ));
 sg13g2_dfrbp_1 \line_lfsr[1]$_SDFFCE_PN1P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net199),
    .D(_0140_),
    .Q_N(_2995_),
    .Q(\line_lfsr[1] ));
 sg13g2_dfrbp_1 \line_lfsr[2]$_SDFFCE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net200),
    .D(_0141_),
    .Q_N(_2994_),
    .Q(\line_lfsr[2] ));
 sg13g2_dfrbp_1 \line_lfsr[3]$_SDFFCE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net201),
    .D(_0142_),
    .Q_N(_2993_),
    .Q(\line_lfsr[3] ));
 sg13g2_dfrbp_1 \line_lfsr[4]$_SDFFCE_PN1P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net202),
    .D(_0143_),
    .Q_N(_2992_),
    .Q(\line_lfsr[4] ));
 sg13g2_dfrbp_1 \line_lfsr[5]$_SDFFCE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net203),
    .D(_0144_),
    .Q_N(_2991_),
    .Q(\line_lfsr[5] ));
 sg13g2_dfrbp_1 \line_lfsr[6]$_SDFFCE_PN1P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net204),
    .D(_0145_),
    .Q_N(_2990_),
    .Q(\line_lfsr[6] ));
 sg13g2_dfrbp_1 \nyanframe[0]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net138),
    .D(_0146_),
    .Q_N(_0008_),
    .Q(\nyanframe[0] ));
 sg13g2_dfrbp_1 \nyanframe[1]$_DFFE_PN0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net139),
    .D(_0147_),
    .Q_N(_2989_),
    .Q(\nyanframe[1] ));
 sg13g2_dfrbp_1 \nyanframe[2]$_DFFE_PN0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net138),
    .D(_0148_),
    .Q_N(_0035_),
    .Q(\nyanframe[2] ));
 sg13g2_dfrbp_1 \sample_beat_ctr[0]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net125),
    .D(_0149_),
    .Q_N(_2988_),
    .Q(\sample_beat_ctr[0] ));
 sg13g2_dfrbp_1 \sample_beat_ctr[1]$_DFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net130),
    .D(_0150_),
    .Q_N(_2987_),
    .Q(\sample_beat_ctr[1] ));
 sg13g2_dfrbp_1 \sample_beat_ctr[2]$_DFFE_PN0P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net131),
    .D(_0151_),
    .Q_N(_2986_),
    .Q(\sample_beat_ctr[2] ));
 sg13g2_dfrbp_1 \sin[0]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net128),
    .D(_0152_),
    .Q_N(_2985_),
    .Q(\sin[0] ));
 sg13g2_dfrbp_1 \sin[1]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net129),
    .D(_0153_),
    .Q_N(_2984_),
    .Q(\nyan_x_offset[0] ));
 sg13g2_dfrbp_1 \sin[2]$_DFFE_PN0P_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net129),
    .D(_0154_),
    .Q_N(_2983_),
    .Q(\nyan_x_offset[1] ));
 sg13g2_dfrbp_1 \sin[3]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net129),
    .D(_0155_),
    .Q_N(_2982_),
    .Q(\nyan_x_offset[2] ));
 sg13g2_dfrbp_1 \sin[4]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net128),
    .D(_0156_),
    .Q_N(_2981_),
    .Q(\nyan_x_offset[3] ));
 sg13g2_dfrbp_1 \sin[5]$_DFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net129),
    .D(_0157_),
    .Q_N(_2980_),
    .Q(\nyan_x_offset[4] ));
 sg13g2_dfrbp_1 \sin[6]$_DFFE_PN0P_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net128),
    .D(_0158_),
    .Q_N(_2979_),
    .Q(\sin[6] ));
 sg13g2_dfrbp_1 \song_loops$_DFFE_PN0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net134),
    .D(_0159_),
    .Q_N(_2963_),
    .Q(song_loops));
 sg13g2_dfrbp_1 \songpos[0]$_DFFE_PN1P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net137),
    .D(_0160_),
    .Q_N(\songpos[0] ),
    .Q(_0052_));
 sg13g2_dfrbp_1 \songpos[1]$_DFFE_PN1P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net134),
    .D(_0161_),
    .Q_N(\songpos[1] ),
    .Q(_0053_));
 sg13g2_dfrbp_1 \songpos[2]$_DFFE_PN1P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net134),
    .D(_0162_),
    .Q_N(\songpos[2] ),
    .Q(_0054_));
 sg13g2_dfrbp_1 \songpos[3]$_DFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net135),
    .D(_0163_),
    .Q_N(\songpos[3] ),
    .Q(_0055_));
 sg13g2_dfrbp_1 \songpos[4]$_DFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net134),
    .D(_0164_),
    .Q_N(\songpos[4] ),
    .Q(_0056_));
 sg13g2_dfrbp_1 \songpos[5]$_DFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net133),
    .D(_0165_),
    .Q_N(\songpos[5] ),
    .Q(_0057_));
 sg13g2_dfrbp_1 \songpos[6]$_DFFE_PN1P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net133),
    .D(_0166_),
    .Q_N(\songpos[6] ),
    .Q(_0058_));
 sg13g2_dfrbp_1 \songpos[7]$_DFFE_PN1P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net134),
    .D(_0167_),
    .Q_N(\songpos[7] ),
    .Q(_0059_));
 sg13g2_dfrbp_1 \songpos[8]$_DFFE_PN1P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net135),
    .D(_0168_),
    .Q_N(\songpos[8] ),
    .Q(_0060_));
 sg13g2_dfrbp_1 \sqr_pha[0]$_DFFE_PN0N_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net125),
    .D(_0169_),
    .Q_N(_2978_),
    .Q(\sqr_pha[0] ));
 sg13g2_dfrbp_1 \sqr_pha[10]$_DFFE_PN0N_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net125),
    .D(_0170_),
    .Q_N(_0025_),
    .Q(\sqr_pha[10] ));
 sg13g2_dfrbp_1 \sqr_pha[11]$_DFFE_PN0N_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net124),
    .D(_0171_),
    .Q_N(_0026_),
    .Q(\sqr_pha[11] ));
 sg13g2_dfrbp_1 \sqr_pha[12]$_DFFE_PN0N_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net130),
    .D(_0172_),
    .Q_N(_0027_),
    .Q(\sqr_pha[12] ));
 sg13g2_dfrbp_1 \sqr_pha[1]$_DFFE_PN0N_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net125),
    .D(_0173_),
    .Q_N(_2977_),
    .Q(\sqr_pha[1] ));
 sg13g2_dfrbp_1 \sqr_pha[2]$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net125),
    .D(_0174_),
    .Q_N(_2976_),
    .Q(\sqr_pha[2] ));
 sg13g2_dfrbp_1 \sqr_pha[3]$_DFFE_PN0N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net123),
    .D(_0175_),
    .Q_N(_2975_),
    .Q(\sqr_pha[3] ));
 sg13g2_dfrbp_1 \sqr_pha[4]$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net123),
    .D(_0176_),
    .Q_N(_2974_),
    .Q(\sqr_pha[4] ));
 sg13g2_dfrbp_1 \sqr_pha[5]$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net126),
    .D(_0177_),
    .Q_N(_2973_),
    .Q(\sqr_pha[5] ));
 sg13g2_dfrbp_1 \sqr_pha[6]$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net126),
    .D(_0178_),
    .Q_N(_2972_),
    .Q(\sqr_pha[6] ));
 sg13g2_dfrbp_1 \sqr_pha[7]$_DFFE_PN0N_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net126),
    .D(_0179_),
    .Q_N(_2971_),
    .Q(\sqr_pha[7] ));
 sg13g2_dfrbp_1 \sqr_pha[8]$_DFFE_PN0N_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net124),
    .D(_0180_),
    .Q_N(_0024_),
    .Q(\sqr_pha[8] ));
 sg13g2_dfrbp_1 \sqr_pha[9]$_DFFE_PN0N_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net125),
    .D(_0181_),
    .Q_N(_2970_),
    .Q(\sqr_pha[9] ));
 sg13g2_dfrbp_1 \sqr_vol[0]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net137),
    .D(_0182_),
    .Q_N(_2969_),
    .Q(\sqr_vol[0] ));
 sg13g2_dfrbp_1 \sqr_vol[1]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net137),
    .D(_0183_),
    .Q_N(_2968_),
    .Q(\sqr_vol[1] ));
 sg13g2_dfrbp_1 \sqr_vol[2]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net137),
    .D(_0184_),
    .Q_N(_2967_),
    .Q(\sqr_vol[2] ));
 sg13g2_dfrbp_1 \sqr_vol[3]$_DFFE_PN0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net133),
    .D(_0185_),
    .Q_N(_2966_),
    .Q(\sqr_vol[3] ));
 sg13g2_dfrbp_1 \sqr_vol[4]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net133),
    .D(_0186_),
    .Q_N(_2965_),
    .Q(\sqr_vol[4] ));
 sg13g2_dfrbp_1 \sqr_vol[5]$_DFFE_PN0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net134),
    .D(_0187_),
    .Q_N(_2964_),
    .Q(\sqr_vol[5] ));
 sg13g2_buf_1 input1 (.A(rst_n),
    .X(net1));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[7]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uo_out[0]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uo_out[1]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uo_out[2]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[3]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[5]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[6]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout11 (.A(_1727_),
    .X(net11));
 sg13g2_buf_2 fanout12 (.A(_1884_),
    .X(net12));
 sg13g2_buf_2 fanout13 (.A(_2516_),
    .X(net13));
 sg13g2_buf_2 fanout14 (.A(_2504_),
    .X(net14));
 sg13g2_buf_2 fanout15 (.A(_1301_),
    .X(net15));
 sg13g2_buf_2 fanout16 (.A(_0271_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_2569_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_2880_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2594_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2577_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_2568_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0273_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_2879_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_2825_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_2593_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_2576_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_2567_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_2444_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0239_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_2948_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_2804_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_2592_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_2575_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_2566_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2443_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_1800_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_1784_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_1574_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0238_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_2818_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_2787_),
    .X(net41));
 sg13g2_buf_4 fanout42 (.X(net42),
    .A(_2591_));
 sg13g2_buf_2 fanout43 (.A(_2574_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2565_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_2469_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_2442_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_1532_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_2844_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_2792_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_2476_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_2468_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_2441_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_1645_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_1515_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2876_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_2791_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_2779_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1583_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1582_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1221_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_2932_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1220_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_0279_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_1909_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_2473_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2030_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_2017_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_2008_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_2002_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_0263_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_0251_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_0241_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_0228_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_2909_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_2885_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_1505_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_0393_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_0339_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_0326_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_0227_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_2886_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_2848_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_2802_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_2618_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_1361_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_0277_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_0248_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_2859_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_2836_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_2813_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_2617_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_0276_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_2941_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_2769_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_2686_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_2642_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_2637_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_2627_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_2606_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_2310_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_1330_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_0253_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_2632_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_2626_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_2624_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_2615_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_2335_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_2321_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_2311_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_2305_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_2303_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_2623_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_2415_),
    .X(net113));
 sg13g2_buf_4 fanout114 (.X(net114),
    .A(_2385_));
 sg13g2_buf_2 fanout115 (.A(_2380_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_2379_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_2376_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_2342_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_2341_),
    .X(net119));
 sg13g2_buf_2 fanout120 (.A(_2338_),
    .X(net120));
 sg13g2_buf_2 fanout121 (.A(_2316_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_2306_),
    .X(net122));
 sg13g2_buf_4 fanout123 (.X(net123),
    .A(net126));
 sg13g2_buf_4 fanout124 (.X(net124),
    .A(net126));
 sg13g2_buf_2 fanout125 (.A(net126),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(net132),
    .X(net126));
 sg13g2_buf_4 fanout127 (.X(net127),
    .A(net128));
 sg13g2_buf_4 fanout128 (.X(net128),
    .A(net132));
 sg13g2_buf_2 fanout129 (.A(net132),
    .X(net129));
 sg13g2_buf_4 fanout130 (.X(net130),
    .A(net132));
 sg13g2_buf_2 fanout131 (.A(net132),
    .X(net131));
 sg13g2_buf_1 fanout132 (.A(net1),
    .X(net132));
 sg13g2_buf_4 fanout133 (.X(net133),
    .A(net134));
 sg13g2_buf_4 fanout134 (.X(net134),
    .A(net135));
 sg13g2_buf_2 fanout135 (.A(net139),
    .X(net135));
 sg13g2_buf_4 fanout136 (.X(net136),
    .A(net137));
 sg13g2_buf_2 fanout137 (.A(net139),
    .X(net137));
 sg13g2_buf_4 fanout138 (.X(net138),
    .A(net139));
 sg13g2_buf_2 fanout139 (.A(net1),
    .X(net139));
 sg13g2_tielo _5980__140 (.L_LO(net140));
 sg13g2_tielo _5981__141 (.L_LO(net141));
 sg13g2_tielo _5982__142 (.L_LO(net142));
 sg13g2_tielo _5983__143 (.L_LO(net143));
 sg13g2_tielo _5984__144 (.L_LO(net144));
 sg13g2_tielo _5985__145 (.L_LO(net145));
 sg13g2_tielo _5986__146 (.L_LO(net146));
 sg13g2_tielo _5988__147 (.L_LO(net147));
 sg13g2_tielo _5989__148 (.L_LO(net148));
 sg13g2_tielo _5990__149 (.L_LO(net149));
 sg13g2_tielo _5991__150 (.L_LO(net150));
 sg13g2_tielo _5992__151 (.L_LO(net151));
 sg13g2_tielo _5993__152 (.L_LO(net152));
 sg13g2_tielo _5994__153 (.L_LO(net153));
 sg13g2_tiehi \audio_sample_lpf[0]$_DFFE_PP__155  (.L_HI(net155));
 sg13g2_tiehi \audio_sample_lpf[1]$_DFFE_PP__156  (.L_HI(net156));
 sg13g2_tiehi \audio_sample_lpf[2]$_DFFE_PP__157  (.L_HI(net157));
 sg13g2_tiehi \audio_sample_lpf[3]$_DFFE_PP__158  (.L_HI(net158));
 sg13g2_tiehi \audio_sample_lpf[4]$_DFFE_PP__159  (.L_HI(net159));
 sg13g2_tiehi \audio_sample_lpf[5]$_DFFE_PP__160  (.L_HI(net160));
 sg13g2_tiehi \audio_sample_lpf[6]$_DFFE_PP__161  (.L_HI(net161));
 sg13g2_tiehi \audio_sample_lpf[7]$_DFFE_PP__162  (.L_HI(net162));
 sg13g2_tiehi \audio_sample_lpf[8]$_DFFE_PP__163  (.L_HI(net163));
 sg13g2_tiehi \audio_sample_lpf[9]$_DFFE_PP__164  (.L_HI(net164));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__169  (.L_HI(net169));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__170  (.L_HI(net170));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__171  (.L_HI(net171));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__172  (.L_HI(net172));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__173  (.L_HI(net173));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__174  (.L_HI(net174));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__175  (.L_HI(net175));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__179  (.L_HI(net179));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__180  (.L_HI(net180));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__181  (.L_HI(net181));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__182  (.L_HI(net182));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__183  (.L_HI(net183));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__184  (.L_HI(net184));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__185  (.L_HI(net185));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__186  (.L_HI(net186));
 sg13g2_tiehi \kick_ctr[0]$_SDFFCE_PP1P__187  (.L_HI(net187));
 sg13g2_tiehi \kick_ctr[1]$_SDFFCE_PP0P__188  (.L_HI(net188));
 sg13g2_tiehi \kick_osci[0]$_SDFFCE_PP0P__189  (.L_HI(net189));
 sg13g2_tiehi \kick_osci[1]$_SDFFCE_PP0P__190  (.L_HI(net190));
 sg13g2_tiehi \kick_osci[2]$_SDFFCE_PP0P__191  (.L_HI(net191));
 sg13g2_tiehi \kick_osci[3]$_SDFFCE_PP0P__192  (.L_HI(net192));
 sg13g2_tiehi \kick_osci[4]$_SDFFCE_PP0P__193  (.L_HI(net193));
 sg13g2_tiehi \kick_osci[5]$_SDFFCE_PP0P__194  (.L_HI(net194));
 sg13g2_tiehi \kick_osci[6]$_SDFFCE_PP0P__195  (.L_HI(net195));
 sg13g2_tiehi \kick_osci[7]$_SDFFCE_PP1P__196  (.L_HI(net196));
 sg13g2_tiehi \kick_osci[8]$_SDFFCE_PP1P__197  (.L_HI(net197));
 sg13g2_tiehi \line_lfsr[0]$_SDFFCE_PN0P__198  (.L_HI(net198));
 sg13g2_tiehi \line_lfsr[1]$_SDFFCE_PN1P__199  (.L_HI(net199));
 sg13g2_tiehi \line_lfsr[2]$_SDFFCE_PN0P__200  (.L_HI(net200));
 sg13g2_tiehi \line_lfsr[3]$_SDFFCE_PN1P__201  (.L_HI(net201));
 sg13g2_tiehi \line_lfsr[4]$_SDFFCE_PN1P__202  (.L_HI(net202));
 sg13g2_tiehi \line_lfsr[5]$_SDFFCE_PN0P__203  (.L_HI(net203));
 sg13g2_tiehi \line_lfsr[6]$_SDFFCE_PN1P__204  (.L_HI(net204));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_7__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_11__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_15__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_19__leaf_clk));
 sg13g2_inv_1 clkload9 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload10 (.A(clknet_5_23__leaf_clk));
 sg13g2_inv_1 clkload11 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload12 (.A(clknet_5_27__leaf_clk));
 sg13g2_inv_1 clkload13 (.A(clknet_5_29__leaf_clk));
 sg13g2_inv_1 clkload14 (.A(clknet_5_31__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(_0006_));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_antennanp ANTENNA_4 (.A(_0006_));
 sg13g2_antennanp ANTENNA_5 (.A(clk));
 sg13g2_antennanp ANTENNA_6 (.A(_0006_));
 sg13g2_antennanp ANTENNA_7 (.A(clk));
 sg13g2_antennanp ANTENNA_8 (.A(_0006_));
 sg13g2_antennanp ANTENNA_9 (.A(clk));
 sg13g2_antennanp ANTENNA_10 (.A(_0006_));
 sg13g2_antennanp ANTENNA_11 (.A(clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_fill_2 FILLER_0_427 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_263 ();
 sg13g2_decap_8 FILLER_1_270 ();
 sg13g2_decap_8 FILLER_1_277 ();
 sg13g2_decap_8 FILLER_1_284 ();
 sg13g2_decap_8 FILLER_1_291 ();
 sg13g2_decap_8 FILLER_1_298 ();
 sg13g2_decap_8 FILLER_1_305 ();
 sg13g2_decap_8 FILLER_1_312 ();
 sg13g2_decap_8 FILLER_1_319 ();
 sg13g2_decap_8 FILLER_1_326 ();
 sg13g2_decap_8 FILLER_1_333 ();
 sg13g2_decap_8 FILLER_1_340 ();
 sg13g2_decap_8 FILLER_1_347 ();
 sg13g2_decap_8 FILLER_1_354 ();
 sg13g2_decap_8 FILLER_1_361 ();
 sg13g2_decap_8 FILLER_1_368 ();
 sg13g2_decap_8 FILLER_1_375 ();
 sg13g2_decap_8 FILLER_1_382 ();
 sg13g2_decap_8 FILLER_1_389 ();
 sg13g2_decap_8 FILLER_1_396 ();
 sg13g2_decap_8 FILLER_1_403 ();
 sg13g2_decap_8 FILLER_1_410 ();
 sg13g2_decap_8 FILLER_1_417 ();
 sg13g2_decap_4 FILLER_1_424 ();
 sg13g2_fill_2 FILLER_1_428 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_4 FILLER_2_238 ();
 sg13g2_fill_1 FILLER_2_242 ();
 sg13g2_fill_2 FILLER_2_282 ();
 sg13g2_decap_8 FILLER_2_293 ();
 sg13g2_decap_8 FILLER_2_300 ();
 sg13g2_decap_8 FILLER_2_307 ();
 sg13g2_decap_8 FILLER_2_314 ();
 sg13g2_decap_8 FILLER_2_321 ();
 sg13g2_decap_8 FILLER_2_328 ();
 sg13g2_decap_8 FILLER_2_335 ();
 sg13g2_decap_8 FILLER_2_342 ();
 sg13g2_decap_8 FILLER_2_349 ();
 sg13g2_decap_8 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_363 ();
 sg13g2_decap_8 FILLER_2_370 ();
 sg13g2_decap_8 FILLER_2_377 ();
 sg13g2_decap_8 FILLER_2_384 ();
 sg13g2_decap_8 FILLER_2_391 ();
 sg13g2_decap_8 FILLER_2_398 ();
 sg13g2_decap_8 FILLER_2_405 ();
 sg13g2_decap_8 FILLER_2_412 ();
 sg13g2_decap_8 FILLER_2_419 ();
 sg13g2_decap_4 FILLER_2_426 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_fill_2 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_82 ();
 sg13g2_decap_8 FILLER_3_89 ();
 sg13g2_decap_8 FILLER_3_96 ();
 sg13g2_decap_8 FILLER_3_103 ();
 sg13g2_decap_8 FILLER_3_110 ();
 sg13g2_decap_8 FILLER_3_117 ();
 sg13g2_decap_8 FILLER_3_124 ();
 sg13g2_decap_8 FILLER_3_131 ();
 sg13g2_decap_8 FILLER_3_138 ();
 sg13g2_decap_8 FILLER_3_145 ();
 sg13g2_decap_8 FILLER_3_152 ();
 sg13g2_decap_8 FILLER_3_159 ();
 sg13g2_decap_8 FILLER_3_166 ();
 sg13g2_decap_8 FILLER_3_173 ();
 sg13g2_decap_8 FILLER_3_180 ();
 sg13g2_decap_8 FILLER_3_187 ();
 sg13g2_decap_8 FILLER_3_194 ();
 sg13g2_decap_8 FILLER_3_201 ();
 sg13g2_decap_8 FILLER_3_208 ();
 sg13g2_decap_4 FILLER_3_215 ();
 sg13g2_decap_4 FILLER_3_250 ();
 sg13g2_fill_1 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_263 ();
 sg13g2_decap_8 FILLER_3_298 ();
 sg13g2_decap_8 FILLER_3_305 ();
 sg13g2_decap_8 FILLER_3_312 ();
 sg13g2_decap_8 FILLER_3_319 ();
 sg13g2_decap_8 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_333 ();
 sg13g2_decap_8 FILLER_3_340 ();
 sg13g2_decap_8 FILLER_3_347 ();
 sg13g2_decap_8 FILLER_3_354 ();
 sg13g2_decap_8 FILLER_3_361 ();
 sg13g2_decap_8 FILLER_3_368 ();
 sg13g2_decap_8 FILLER_3_375 ();
 sg13g2_decap_8 FILLER_3_382 ();
 sg13g2_decap_8 FILLER_3_389 ();
 sg13g2_decap_8 FILLER_3_396 ();
 sg13g2_decap_8 FILLER_3_403 ();
 sg13g2_decap_8 FILLER_3_410 ();
 sg13g2_decap_8 FILLER_3_417 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_4 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_128 ();
 sg13g2_decap_8 FILLER_4_135 ();
 sg13g2_decap_8 FILLER_4_142 ();
 sg13g2_decap_8 FILLER_4_149 ();
 sg13g2_decap_8 FILLER_4_156 ();
 sg13g2_decap_8 FILLER_4_163 ();
 sg13g2_decap_8 FILLER_4_170 ();
 sg13g2_decap_8 FILLER_4_177 ();
 sg13g2_decap_8 FILLER_4_184 ();
 sg13g2_decap_8 FILLER_4_191 ();
 sg13g2_decap_8 FILLER_4_198 ();
 sg13g2_decap_8 FILLER_4_205 ();
 sg13g2_decap_8 FILLER_4_212 ();
 sg13g2_decap_8 FILLER_4_219 ();
 sg13g2_decap_8 FILLER_4_226 ();
 sg13g2_decap_4 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_237 ();
 sg13g2_fill_2 FILLER_4_266 ();
 sg13g2_fill_1 FILLER_4_271 ();
 sg13g2_decap_4 FILLER_4_276 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_fill_2 FILLER_5_35 ();
 sg13g2_fill_1 FILLER_5_37 ();
 sg13g2_fill_1 FILLER_5_50 ();
 sg13g2_fill_1 FILLER_5_59 ();
 sg13g2_decap_8 FILLER_5_64 ();
 sg13g2_decap_8 FILLER_5_71 ();
 sg13g2_decap_4 FILLER_5_78 ();
 sg13g2_fill_1 FILLER_5_82 ();
 sg13g2_decap_4 FILLER_5_112 ();
 sg13g2_fill_1 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_120 ();
 sg13g2_decap_8 FILLER_5_127 ();
 sg13g2_decap_8 FILLER_5_134 ();
 sg13g2_decap_8 FILLER_5_141 ();
 sg13g2_decap_8 FILLER_5_148 ();
 sg13g2_decap_8 FILLER_5_155 ();
 sg13g2_decap_8 FILLER_5_162 ();
 sg13g2_decap_8 FILLER_5_169 ();
 sg13g2_decap_8 FILLER_5_176 ();
 sg13g2_decap_8 FILLER_5_183 ();
 sg13g2_decap_8 FILLER_5_190 ();
 sg13g2_decap_8 FILLER_5_197 ();
 sg13g2_decap_8 FILLER_5_204 ();
 sg13g2_decap_8 FILLER_5_211 ();
 sg13g2_decap_4 FILLER_5_218 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_227 ();
 sg13g2_decap_8 FILLER_5_234 ();
 sg13g2_fill_2 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_261 ();
 sg13g2_fill_1 FILLER_5_267 ();
 sg13g2_decap_8 FILLER_5_289 ();
 sg13g2_decap_8 FILLER_5_296 ();
 sg13g2_decap_8 FILLER_5_303 ();
 sg13g2_decap_8 FILLER_5_310 ();
 sg13g2_decap_8 FILLER_5_317 ();
 sg13g2_decap_8 FILLER_5_324 ();
 sg13g2_decap_8 FILLER_5_331 ();
 sg13g2_decap_8 FILLER_5_338 ();
 sg13g2_decap_8 FILLER_5_345 ();
 sg13g2_decap_8 FILLER_5_352 ();
 sg13g2_decap_8 FILLER_5_359 ();
 sg13g2_decap_8 FILLER_5_366 ();
 sg13g2_decap_8 FILLER_5_373 ();
 sg13g2_decap_8 FILLER_5_380 ();
 sg13g2_decap_8 FILLER_5_387 ();
 sg13g2_decap_8 FILLER_5_394 ();
 sg13g2_decap_8 FILLER_5_401 ();
 sg13g2_decap_8 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_5_415 ();
 sg13g2_decap_8 FILLER_5_422 ();
 sg13g2_fill_1 FILLER_5_429 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_fill_2 FILLER_6_51 ();
 sg13g2_fill_1 FILLER_6_53 ();
 sg13g2_fill_1 FILLER_6_58 ();
 sg13g2_fill_2 FILLER_6_64 ();
 sg13g2_fill_1 FILLER_6_66 ();
 sg13g2_fill_1 FILLER_6_71 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_4 FILLER_6_91 ();
 sg13g2_fill_2 FILLER_6_109 ();
 sg13g2_fill_1 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_121 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_4 FILLER_6_196 ();
 sg13g2_fill_2 FILLER_6_200 ();
 sg13g2_fill_2 FILLER_6_228 ();
 sg13g2_fill_1 FILLER_6_230 ();
 sg13g2_fill_1 FILLER_6_241 ();
 sg13g2_fill_2 FILLER_6_257 ();
 sg13g2_fill_1 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_286 ();
 sg13g2_decap_4 FILLER_6_292 ();
 sg13g2_fill_2 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_fill_2 FILLER_6_427 ();
 sg13g2_fill_1 FILLER_6_429 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_4 FILLER_7_14 ();
 sg13g2_fill_1 FILLER_7_18 ();
 sg13g2_decap_4 FILLER_7_84 ();
 sg13g2_fill_1 FILLER_7_93 ();
 sg13g2_fill_2 FILLER_7_116 ();
 sg13g2_fill_2 FILLER_7_141 ();
 sg13g2_decap_8 FILLER_7_146 ();
 sg13g2_decap_8 FILLER_7_153 ();
 sg13g2_decap_8 FILLER_7_160 ();
 sg13g2_decap_8 FILLER_7_167 ();
 sg13g2_decap_8 FILLER_7_174 ();
 sg13g2_decap_4 FILLER_7_181 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_decap_4 FILLER_7_213 ();
 sg13g2_fill_2 FILLER_7_217 ();
 sg13g2_decap_8 FILLER_7_258 ();
 sg13g2_decap_4 FILLER_7_265 ();
 sg13g2_fill_1 FILLER_7_269 ();
 sg13g2_decap_8 FILLER_7_274 ();
 sg13g2_fill_1 FILLER_7_281 ();
 sg13g2_decap_8 FILLER_7_308 ();
 sg13g2_decap_8 FILLER_7_315 ();
 sg13g2_decap_8 FILLER_7_322 ();
 sg13g2_decap_8 FILLER_7_329 ();
 sg13g2_decap_8 FILLER_7_336 ();
 sg13g2_decap_8 FILLER_7_343 ();
 sg13g2_decap_8 FILLER_7_350 ();
 sg13g2_decap_8 FILLER_7_357 ();
 sg13g2_decap_8 FILLER_7_364 ();
 sg13g2_decap_8 FILLER_7_371 ();
 sg13g2_decap_8 FILLER_7_378 ();
 sg13g2_decap_8 FILLER_7_385 ();
 sg13g2_decap_8 FILLER_7_392 ();
 sg13g2_decap_8 FILLER_7_399 ();
 sg13g2_decap_8 FILLER_7_406 ();
 sg13g2_decap_8 FILLER_7_413 ();
 sg13g2_decap_8 FILLER_7_420 ();
 sg13g2_fill_2 FILLER_7_427 ();
 sg13g2_fill_1 FILLER_7_429 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_fill_1 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_48 ();
 sg13g2_fill_1 FILLER_8_67 ();
 sg13g2_fill_1 FILLER_8_102 ();
 sg13g2_fill_1 FILLER_8_111 ();
 sg13g2_fill_2 FILLER_8_136 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_decap_8 FILLER_8_153 ();
 sg13g2_decap_8 FILLER_8_160 ();
 sg13g2_decap_8 FILLER_8_167 ();
 sg13g2_decap_8 FILLER_8_174 ();
 sg13g2_decap_8 FILLER_8_181 ();
 sg13g2_decap_8 FILLER_8_188 ();
 sg13g2_decap_8 FILLER_8_195 ();
 sg13g2_fill_2 FILLER_8_202 ();
 sg13g2_fill_1 FILLER_8_204 ();
 sg13g2_decap_4 FILLER_8_213 ();
 sg13g2_decap_8 FILLER_8_222 ();
 sg13g2_decap_8 FILLER_8_229 ();
 sg13g2_decap_8 FILLER_8_269 ();
 sg13g2_decap_4 FILLER_8_276 ();
 sg13g2_fill_1 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_298 ();
 sg13g2_decap_8 FILLER_8_305 ();
 sg13g2_decap_8 FILLER_8_312 ();
 sg13g2_decap_8 FILLER_8_319 ();
 sg13g2_decap_8 FILLER_8_326 ();
 sg13g2_decap_8 FILLER_8_333 ();
 sg13g2_decap_8 FILLER_8_340 ();
 sg13g2_decap_8 FILLER_8_347 ();
 sg13g2_decap_8 FILLER_8_354 ();
 sg13g2_decap_8 FILLER_8_361 ();
 sg13g2_decap_8 FILLER_8_368 ();
 sg13g2_decap_8 FILLER_8_375 ();
 sg13g2_decap_8 FILLER_8_382 ();
 sg13g2_decap_8 FILLER_8_389 ();
 sg13g2_decap_8 FILLER_8_396 ();
 sg13g2_decap_8 FILLER_8_403 ();
 sg13g2_decap_8 FILLER_8_410 ();
 sg13g2_decap_8 FILLER_8_417 ();
 sg13g2_decap_4 FILLER_8_424 ();
 sg13g2_fill_2 FILLER_8_428 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_fill_1 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_73 ();
 sg13g2_decap_8 FILLER_9_80 ();
 sg13g2_decap_4 FILLER_9_87 ();
 sg13g2_fill_1 FILLER_9_91 ();
 sg13g2_fill_1 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_136 ();
 sg13g2_decap_8 FILLER_9_143 ();
 sg13g2_decap_8 FILLER_9_150 ();
 sg13g2_decap_8 FILLER_9_157 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_decap_8 FILLER_9_191 ();
 sg13g2_decap_8 FILLER_9_198 ();
 sg13g2_decap_8 FILLER_9_205 ();
 sg13g2_decap_4 FILLER_9_212 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_fill_2 FILLER_9_245 ();
 sg13g2_decap_4 FILLER_9_251 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_fill_1 FILLER_9_280 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_fill_2 FILLER_9_427 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_fill_1 FILLER_10_64 ();
 sg13g2_decap_8 FILLER_10_70 ();
 sg13g2_decap_4 FILLER_10_77 ();
 sg13g2_fill_1 FILLER_10_81 ();
 sg13g2_fill_2 FILLER_10_87 ();
 sg13g2_fill_1 FILLER_10_89 ();
 sg13g2_fill_1 FILLER_10_102 ();
 sg13g2_fill_1 FILLER_10_113 ();
 sg13g2_decap_8 FILLER_10_118 ();
 sg13g2_decap_8 FILLER_10_125 ();
 sg13g2_decap_4 FILLER_10_132 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_4 FILLER_10_165 ();
 sg13g2_fill_1 FILLER_10_169 ();
 sg13g2_fill_2 FILLER_10_200 ();
 sg13g2_fill_1 FILLER_10_216 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_fill_2 FILLER_10_257 ();
 sg13g2_decap_8 FILLER_10_265 ();
 sg13g2_fill_2 FILLER_10_272 ();
 sg13g2_fill_1 FILLER_10_274 ();
 sg13g2_decap_8 FILLER_10_296 ();
 sg13g2_decap_4 FILLER_10_303 ();
 sg13g2_decap_8 FILLER_10_320 ();
 sg13g2_decap_8 FILLER_10_327 ();
 sg13g2_decap_8 FILLER_10_334 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_8 FILLER_10_404 ();
 sg13g2_decap_8 FILLER_10_411 ();
 sg13g2_decap_8 FILLER_10_418 ();
 sg13g2_decap_4 FILLER_10_425 ();
 sg13g2_fill_1 FILLER_10_429 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_fill_2 FILLER_11_7 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_fill_1 FILLER_11_37 ();
 sg13g2_decap_8 FILLER_11_41 ();
 sg13g2_fill_2 FILLER_11_48 ();
 sg13g2_fill_2 FILLER_11_53 ();
 sg13g2_fill_1 FILLER_11_55 ();
 sg13g2_fill_2 FILLER_11_61 ();
 sg13g2_fill_2 FILLER_11_67 ();
 sg13g2_fill_1 FILLER_11_69 ();
 sg13g2_fill_2 FILLER_11_78 ();
 sg13g2_fill_1 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_103 ();
 sg13g2_decap_8 FILLER_11_110 ();
 sg13g2_decap_8 FILLER_11_117 ();
 sg13g2_fill_1 FILLER_11_124 ();
 sg13g2_decap_4 FILLER_11_164 ();
 sg13g2_fill_1 FILLER_11_168 ();
 sg13g2_fill_2 FILLER_11_186 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_213 ();
 sg13g2_fill_1 FILLER_11_244 ();
 sg13g2_fill_2 FILLER_11_271 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_decap_8 FILLER_11_291 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_8 FILLER_11_403 ();
 sg13g2_decap_8 FILLER_11_410 ();
 sg13g2_decap_8 FILLER_11_417 ();
 sg13g2_decap_4 FILLER_11_424 ();
 sg13g2_fill_2 FILLER_11_428 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_fill_2 FILLER_12_14 ();
 sg13g2_decap_4 FILLER_12_47 ();
 sg13g2_fill_2 FILLER_12_51 ();
 sg13g2_fill_1 FILLER_12_84 ();
 sg13g2_decap_4 FILLER_12_100 ();
 sg13g2_fill_1 FILLER_12_109 ();
 sg13g2_fill_1 FILLER_12_114 ();
 sg13g2_fill_1 FILLER_12_126 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_decap_4 FILLER_12_145 ();
 sg13g2_decap_8 FILLER_12_152 ();
 sg13g2_decap_8 FILLER_12_159 ();
 sg13g2_decap_8 FILLER_12_166 ();
 sg13g2_fill_2 FILLER_12_181 ();
 sg13g2_fill_2 FILLER_12_195 ();
 sg13g2_fill_1 FILLER_12_205 ();
 sg13g2_fill_2 FILLER_12_267 ();
 sg13g2_fill_1 FILLER_12_269 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_decap_8 FILLER_12_406 ();
 sg13g2_decap_8 FILLER_12_413 ();
 sg13g2_decap_8 FILLER_12_420 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_4 FILLER_13_28 ();
 sg13g2_fill_1 FILLER_13_45 ();
 sg13g2_fill_1 FILLER_13_50 ();
 sg13g2_decap_8 FILLER_13_55 ();
 sg13g2_decap_8 FILLER_13_62 ();
 sg13g2_fill_1 FILLER_13_69 ();
 sg13g2_fill_2 FILLER_13_131 ();
 sg13g2_fill_1 FILLER_13_137 ();
 sg13g2_decap_8 FILLER_13_146 ();
 sg13g2_decap_8 FILLER_13_157 ();
 sg13g2_fill_2 FILLER_13_164 ();
 sg13g2_fill_1 FILLER_13_184 ();
 sg13g2_decap_8 FILLER_13_222 ();
 sg13g2_decap_8 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_236 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_4 FILLER_13_266 ();
 sg13g2_fill_2 FILLER_13_279 ();
 sg13g2_decap_8 FILLER_13_331 ();
 sg13g2_decap_8 FILLER_13_338 ();
 sg13g2_decap_8 FILLER_13_345 ();
 sg13g2_decap_8 FILLER_13_352 ();
 sg13g2_decap_8 FILLER_13_359 ();
 sg13g2_decap_8 FILLER_13_366 ();
 sg13g2_decap_8 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_380 ();
 sg13g2_decap_8 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_394 ();
 sg13g2_decap_8 FILLER_13_401 ();
 sg13g2_decap_8 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_13_415 ();
 sg13g2_decap_8 FILLER_13_422 ();
 sg13g2_fill_1 FILLER_13_429 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_2 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_52 ();
 sg13g2_decap_8 FILLER_14_59 ();
 sg13g2_decap_8 FILLER_14_66 ();
 sg13g2_decap_8 FILLER_14_73 ();
 sg13g2_decap_4 FILLER_14_80 ();
 sg13g2_fill_1 FILLER_14_84 ();
 sg13g2_fill_2 FILLER_14_101 ();
 sg13g2_fill_1 FILLER_14_115 ();
 sg13g2_fill_2 FILLER_14_127 ();
 sg13g2_fill_1 FILLER_14_134 ();
 sg13g2_fill_1 FILLER_14_139 ();
 sg13g2_fill_2 FILLER_14_144 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_fill_2 FILLER_14_187 ();
 sg13g2_decap_8 FILLER_14_193 ();
 sg13g2_decap_8 FILLER_14_200 ();
 sg13g2_decap_8 FILLER_14_207 ();
 sg13g2_fill_2 FILLER_14_214 ();
 sg13g2_fill_1 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_fill_2 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_decap_8 FILLER_14_298 ();
 sg13g2_decap_8 FILLER_14_305 ();
 sg13g2_decap_8 FILLER_14_312 ();
 sg13g2_decap_8 FILLER_14_319 ();
 sg13g2_decap_8 FILLER_14_326 ();
 sg13g2_decap_8 FILLER_14_333 ();
 sg13g2_decap_8 FILLER_14_340 ();
 sg13g2_decap_8 FILLER_14_347 ();
 sg13g2_decap_8 FILLER_14_354 ();
 sg13g2_decap_8 FILLER_14_361 ();
 sg13g2_decap_8 FILLER_14_368 ();
 sg13g2_decap_8 FILLER_14_375 ();
 sg13g2_decap_8 FILLER_14_382 ();
 sg13g2_decap_8 FILLER_14_389 ();
 sg13g2_decap_8 FILLER_14_396 ();
 sg13g2_decap_8 FILLER_14_403 ();
 sg13g2_decap_8 FILLER_14_410 ();
 sg13g2_decap_8 FILLER_14_417 ();
 sg13g2_decap_4 FILLER_14_424 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_8 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_28 ();
 sg13g2_decap_8 FILLER_15_59 ();
 sg13g2_decap_8 FILLER_15_66 ();
 sg13g2_decap_8 FILLER_15_73 ();
 sg13g2_decap_4 FILLER_15_80 ();
 sg13g2_fill_2 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_99 ();
 sg13g2_decap_4 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_123 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_decap_8 FILLER_15_204 ();
 sg13g2_decap_8 FILLER_15_211 ();
 sg13g2_decap_8 FILLER_15_218 ();
 sg13g2_decap_8 FILLER_15_225 ();
 sg13g2_decap_8 FILLER_15_232 ();
 sg13g2_decap_4 FILLER_15_239 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_decap_8 FILLER_15_248 ();
 sg13g2_decap_8 FILLER_15_255 ();
 sg13g2_fill_2 FILLER_15_262 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_4 FILLER_15_424 ();
 sg13g2_fill_2 FILLER_15_428 ();
 sg13g2_decap_4 FILLER_16_26 ();
 sg13g2_decap_8 FILLER_16_48 ();
 sg13g2_fill_2 FILLER_16_55 ();
 sg13g2_fill_2 FILLER_16_65 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_82 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_decap_8 FILLER_16_113 ();
 sg13g2_decap_8 FILLER_16_135 ();
 sg13g2_decap_8 FILLER_16_142 ();
 sg13g2_decap_8 FILLER_16_153 ();
 sg13g2_decap_4 FILLER_16_160 ();
 sg13g2_decap_8 FILLER_16_184 ();
 sg13g2_decap_8 FILLER_16_191 ();
 sg13g2_fill_2 FILLER_16_198 ();
 sg13g2_fill_2 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_233 ();
 sg13g2_fill_1 FILLER_16_235 ();
 sg13g2_decap_4 FILLER_16_244 ();
 sg13g2_decap_4 FILLER_16_251 ();
 sg13g2_decap_8 FILLER_16_279 ();
 sg13g2_decap_8 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_300 ();
 sg13g2_decap_8 FILLER_16_307 ();
 sg13g2_decap_8 FILLER_16_314 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_decap_8 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_335 ();
 sg13g2_decap_8 FILLER_16_342 ();
 sg13g2_decap_8 FILLER_16_349 ();
 sg13g2_decap_8 FILLER_16_356 ();
 sg13g2_decap_8 FILLER_16_363 ();
 sg13g2_decap_8 FILLER_16_370 ();
 sg13g2_decap_8 FILLER_16_377 ();
 sg13g2_decap_8 FILLER_16_384 ();
 sg13g2_decap_8 FILLER_16_391 ();
 sg13g2_decap_8 FILLER_16_398 ();
 sg13g2_decap_8 FILLER_16_405 ();
 sg13g2_decap_8 FILLER_16_412 ();
 sg13g2_decap_8 FILLER_16_419 ();
 sg13g2_decap_4 FILLER_16_426 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_fill_2 FILLER_17_21 ();
 sg13g2_fill_1 FILLER_17_23 ();
 sg13g2_decap_8 FILLER_17_75 ();
 sg13g2_decap_8 FILLER_17_82 ();
 sg13g2_decap_8 FILLER_17_89 ();
 sg13g2_decap_8 FILLER_17_96 ();
 sg13g2_decap_8 FILLER_17_103 ();
 sg13g2_decap_8 FILLER_17_110 ();
 sg13g2_decap_4 FILLER_17_117 ();
 sg13g2_fill_2 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_126 ();
 sg13g2_decap_8 FILLER_17_135 ();
 sg13g2_decap_8 FILLER_17_142 ();
 sg13g2_decap_8 FILLER_17_149 ();
 sg13g2_decap_8 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_163 ();
 sg13g2_fill_1 FILLER_17_165 ();
 sg13g2_fill_2 FILLER_17_169 ();
 sg13g2_fill_1 FILLER_17_181 ();
 sg13g2_decap_4 FILLER_17_190 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_fill_2 FILLER_17_205 ();
 sg13g2_fill_1 FILLER_17_215 ();
 sg13g2_fill_2 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_226 ();
 sg13g2_decap_4 FILLER_17_233 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_265 ();
 sg13g2_decap_4 FILLER_17_272 ();
 sg13g2_decap_8 FILLER_17_281 ();
 sg13g2_decap_8 FILLER_17_288 ();
 sg13g2_decap_8 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_302 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_decap_8 FILLER_17_316 ();
 sg13g2_decap_8 FILLER_17_323 ();
 sg13g2_decap_8 FILLER_17_330 ();
 sg13g2_decap_8 FILLER_17_337 ();
 sg13g2_decap_8 FILLER_17_344 ();
 sg13g2_decap_8 FILLER_17_351 ();
 sg13g2_decap_8 FILLER_17_358 ();
 sg13g2_decap_8 FILLER_17_365 ();
 sg13g2_decap_8 FILLER_17_372 ();
 sg13g2_decap_8 FILLER_17_379 ();
 sg13g2_decap_8 FILLER_17_386 ();
 sg13g2_decap_8 FILLER_17_393 ();
 sg13g2_decap_8 FILLER_17_400 ();
 sg13g2_decap_8 FILLER_17_407 ();
 sg13g2_decap_8 FILLER_17_414 ();
 sg13g2_decap_8 FILLER_17_421 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_fill_1 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_33 ();
 sg13g2_decap_4 FILLER_18_44 ();
 sg13g2_decap_4 FILLER_18_52 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_2 FILLER_18_65 ();
 sg13g2_fill_2 FILLER_18_71 ();
 sg13g2_decap_4 FILLER_18_77 ();
 sg13g2_decap_4 FILLER_18_85 ();
 sg13g2_fill_1 FILLER_18_113 ();
 sg13g2_fill_1 FILLER_18_118 ();
 sg13g2_fill_1 FILLER_18_123 ();
 sg13g2_fill_2 FILLER_18_136 ();
 sg13g2_fill_1 FILLER_18_138 ();
 sg13g2_decap_4 FILLER_18_143 ();
 sg13g2_fill_1 FILLER_18_147 ();
 sg13g2_fill_1 FILLER_18_179 ();
 sg13g2_decap_4 FILLER_18_183 ();
 sg13g2_decap_8 FILLER_18_205 ();
 sg13g2_decap_4 FILLER_18_212 ();
 sg13g2_fill_1 FILLER_18_216 ();
 sg13g2_decap_8 FILLER_18_225 ();
 sg13g2_decap_4 FILLER_18_232 ();
 sg13g2_fill_1 FILLER_18_236 ();
 sg13g2_decap_8 FILLER_18_246 ();
 sg13g2_fill_1 FILLER_18_253 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_fill_2 FILLER_18_287 ();
 sg13g2_fill_1 FILLER_18_297 ();
 sg13g2_decap_8 FILLER_18_306 ();
 sg13g2_decap_8 FILLER_18_313 ();
 sg13g2_decap_8 FILLER_18_320 ();
 sg13g2_decap_8 FILLER_18_327 ();
 sg13g2_decap_8 FILLER_18_334 ();
 sg13g2_decap_8 FILLER_18_341 ();
 sg13g2_decap_8 FILLER_18_348 ();
 sg13g2_decap_8 FILLER_18_355 ();
 sg13g2_decap_8 FILLER_18_362 ();
 sg13g2_decap_8 FILLER_18_369 ();
 sg13g2_decap_8 FILLER_18_376 ();
 sg13g2_decap_8 FILLER_18_383 ();
 sg13g2_decap_8 FILLER_18_390 ();
 sg13g2_decap_8 FILLER_18_397 ();
 sg13g2_decap_8 FILLER_18_404 ();
 sg13g2_decap_8 FILLER_18_411 ();
 sg13g2_decap_8 FILLER_18_418 ();
 sg13g2_decap_4 FILLER_18_425 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_18 ();
 sg13g2_fill_2 FILLER_19_24 ();
 sg13g2_fill_1 FILLER_19_26 ();
 sg13g2_fill_1 FILLER_19_45 ();
 sg13g2_decap_4 FILLER_19_49 ();
 sg13g2_fill_2 FILLER_19_53 ();
 sg13g2_decap_8 FILLER_19_59 ();
 sg13g2_decap_4 FILLER_19_66 ();
 sg13g2_fill_2 FILLER_19_79 ();
 sg13g2_fill_1 FILLER_19_81 ();
 sg13g2_fill_1 FILLER_19_94 ();
 sg13g2_fill_2 FILLER_19_121 ();
 sg13g2_fill_1 FILLER_19_123 ();
 sg13g2_fill_1 FILLER_19_165 ();
 sg13g2_fill_1 FILLER_19_205 ();
 sg13g2_fill_2 FILLER_19_214 ();
 sg13g2_decap_8 FILLER_19_220 ();
 sg13g2_fill_2 FILLER_19_227 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_fill_2 FILLER_19_266 ();
 sg13g2_fill_1 FILLER_19_268 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_4 FILLER_19_280 ();
 sg13g2_fill_1 FILLER_19_284 ();
 sg13g2_fill_2 FILLER_19_289 ();
 sg13g2_fill_1 FILLER_19_295 ();
 sg13g2_decap_8 FILLER_19_312 ();
 sg13g2_decap_8 FILLER_19_319 ();
 sg13g2_decap_8 FILLER_19_326 ();
 sg13g2_decap_8 FILLER_19_333 ();
 sg13g2_decap_8 FILLER_19_340 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_354 ();
 sg13g2_decap_8 FILLER_19_361 ();
 sg13g2_decap_8 FILLER_19_368 ();
 sg13g2_decap_8 FILLER_19_375 ();
 sg13g2_decap_8 FILLER_19_382 ();
 sg13g2_decap_8 FILLER_19_389 ();
 sg13g2_decap_8 FILLER_19_396 ();
 sg13g2_decap_8 FILLER_19_403 ();
 sg13g2_decap_8 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_417 ();
 sg13g2_decap_4 FILLER_19_424 ();
 sg13g2_fill_2 FILLER_19_428 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_8 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_14 ();
 sg13g2_decap_8 FILLER_20_21 ();
 sg13g2_decap_4 FILLER_20_43 ();
 sg13g2_fill_1 FILLER_20_47 ();
 sg13g2_decap_4 FILLER_20_61 ();
 sg13g2_fill_1 FILLER_20_65 ();
 sg13g2_fill_2 FILLER_20_109 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_fill_1 FILLER_20_125 ();
 sg13g2_decap_8 FILLER_20_129 ();
 sg13g2_fill_1 FILLER_20_136 ();
 sg13g2_decap_8 FILLER_20_142 ();
 sg13g2_decap_8 FILLER_20_149 ();
 sg13g2_fill_2 FILLER_20_156 ();
 sg13g2_fill_1 FILLER_20_158 ();
 sg13g2_decap_4 FILLER_20_167 ();
 sg13g2_decap_4 FILLER_20_175 ();
 sg13g2_fill_1 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_184 ();
 sg13g2_fill_1 FILLER_20_191 ();
 sg13g2_fill_2 FILLER_20_201 ();
 sg13g2_fill_1 FILLER_20_211 ();
 sg13g2_decap_8 FILLER_20_246 ();
 sg13g2_decap_8 FILLER_20_253 ();
 sg13g2_fill_2 FILLER_20_260 ();
 sg13g2_fill_1 FILLER_20_270 ();
 sg13g2_decap_4 FILLER_20_279 ();
 sg13g2_fill_2 FILLER_20_295 ();
 sg13g2_decap_8 FILLER_20_311 ();
 sg13g2_decap_8 FILLER_20_318 ();
 sg13g2_decap_8 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_332 ();
 sg13g2_decap_8 FILLER_20_339 ();
 sg13g2_decap_8 FILLER_20_346 ();
 sg13g2_decap_8 FILLER_20_353 ();
 sg13g2_decap_8 FILLER_20_360 ();
 sg13g2_decap_8 FILLER_20_367 ();
 sg13g2_decap_8 FILLER_20_374 ();
 sg13g2_decap_8 FILLER_20_381 ();
 sg13g2_decap_8 FILLER_20_388 ();
 sg13g2_decap_8 FILLER_20_395 ();
 sg13g2_decap_8 FILLER_20_402 ();
 sg13g2_decap_8 FILLER_20_409 ();
 sg13g2_decap_8 FILLER_20_416 ();
 sg13g2_decap_8 FILLER_20_423 ();
 sg13g2_decap_4 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_71 ();
 sg13g2_fill_2 FILLER_21_81 ();
 sg13g2_fill_1 FILLER_21_83 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_2 FILLER_21_95 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_decap_4 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_107 ();
 sg13g2_fill_2 FILLER_21_134 ();
 sg13g2_fill_1 FILLER_21_166 ();
 sg13g2_fill_2 FILLER_21_172 ();
 sg13g2_decap_4 FILLER_21_177 ();
 sg13g2_fill_2 FILLER_21_181 ();
 sg13g2_decap_4 FILLER_21_187 ();
 sg13g2_fill_1 FILLER_21_191 ();
 sg13g2_decap_8 FILLER_21_200 ();
 sg13g2_fill_1 FILLER_21_211 ();
 sg13g2_fill_1 FILLER_21_217 ();
 sg13g2_fill_2 FILLER_21_222 ();
 sg13g2_decap_8 FILLER_21_227 ();
 sg13g2_decap_4 FILLER_21_234 ();
 sg13g2_fill_1 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_243 ();
 sg13g2_fill_2 FILLER_21_250 ();
 sg13g2_fill_1 FILLER_21_252 ();
 sg13g2_decap_4 FILLER_21_263 ();
 sg13g2_fill_1 FILLER_21_267 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_4 FILLER_21_298 ();
 sg13g2_decap_8 FILLER_21_324 ();
 sg13g2_decap_8 FILLER_21_331 ();
 sg13g2_decap_8 FILLER_21_338 ();
 sg13g2_decap_8 FILLER_21_345 ();
 sg13g2_decap_8 FILLER_21_352 ();
 sg13g2_decap_8 FILLER_21_359 ();
 sg13g2_decap_8 FILLER_21_366 ();
 sg13g2_decap_8 FILLER_21_373 ();
 sg13g2_decap_8 FILLER_21_380 ();
 sg13g2_decap_8 FILLER_21_387 ();
 sg13g2_decap_8 FILLER_21_394 ();
 sg13g2_decap_8 FILLER_21_401 ();
 sg13g2_decap_8 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_decap_8 FILLER_21_422 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_decap_8 FILLER_22_28 ();
 sg13g2_decap_4 FILLER_22_35 ();
 sg13g2_decap_4 FILLER_22_42 ();
 sg13g2_decap_8 FILLER_22_64 ();
 sg13g2_decap_8 FILLER_22_71 ();
 sg13g2_fill_2 FILLER_22_78 ();
 sg13g2_fill_1 FILLER_22_80 ();
 sg13g2_decap_8 FILLER_22_111 ();
 sg13g2_decap_8 FILLER_22_118 ();
 sg13g2_decap_8 FILLER_22_125 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_199 ();
 sg13g2_decap_4 FILLER_22_206 ();
 sg13g2_fill_1 FILLER_22_210 ();
 sg13g2_decap_8 FILLER_22_219 ();
 sg13g2_decap_8 FILLER_22_229 ();
 sg13g2_decap_4 FILLER_22_236 ();
 sg13g2_decap_8 FILLER_22_244 ();
 sg13g2_decap_8 FILLER_22_251 ();
 sg13g2_fill_2 FILLER_22_258 ();
 sg13g2_decap_8 FILLER_22_265 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_291 ();
 sg13g2_fill_1 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_315 ();
 sg13g2_decap_8 FILLER_22_321 ();
 sg13g2_decap_8 FILLER_22_328 ();
 sg13g2_decap_8 FILLER_22_335 ();
 sg13g2_decap_8 FILLER_22_342 ();
 sg13g2_decap_8 FILLER_22_349 ();
 sg13g2_decap_8 FILLER_22_356 ();
 sg13g2_decap_8 FILLER_22_363 ();
 sg13g2_decap_8 FILLER_22_370 ();
 sg13g2_decap_8 FILLER_22_377 ();
 sg13g2_decap_8 FILLER_22_384 ();
 sg13g2_decap_8 FILLER_22_391 ();
 sg13g2_decap_8 FILLER_22_398 ();
 sg13g2_decap_8 FILLER_22_405 ();
 sg13g2_decap_8 FILLER_22_412 ();
 sg13g2_decap_8 FILLER_22_419 ();
 sg13g2_decap_4 FILLER_22_426 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_fill_2 FILLER_23_21 ();
 sg13g2_fill_1 FILLER_23_23 ();
 sg13g2_fill_2 FILLER_23_54 ();
 sg13g2_decap_8 FILLER_23_71 ();
 sg13g2_decap_8 FILLER_23_78 ();
 sg13g2_decap_4 FILLER_23_85 ();
 sg13g2_fill_2 FILLER_23_92 ();
 sg13g2_decap_8 FILLER_23_102 ();
 sg13g2_decap_8 FILLER_23_109 ();
 sg13g2_fill_2 FILLER_23_116 ();
 sg13g2_fill_1 FILLER_23_118 ();
 sg13g2_decap_8 FILLER_23_157 ();
 sg13g2_fill_2 FILLER_23_164 ();
 sg13g2_fill_1 FILLER_23_166 ();
 sg13g2_decap_4 FILLER_23_176 ();
 sg13g2_fill_1 FILLER_23_180 ();
 sg13g2_decap_4 FILLER_23_223 ();
 sg13g2_decap_4 FILLER_23_253 ();
 sg13g2_fill_1 FILLER_23_257 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_decap_4 FILLER_23_295 ();
 sg13g2_fill_1 FILLER_23_299 ();
 sg13g2_fill_1 FILLER_23_308 ();
 sg13g2_fill_1 FILLER_23_313 ();
 sg13g2_fill_1 FILLER_23_323 ();
 sg13g2_decap_8 FILLER_23_332 ();
 sg13g2_decap_8 FILLER_23_339 ();
 sg13g2_decap_8 FILLER_23_346 ();
 sg13g2_decap_8 FILLER_23_353 ();
 sg13g2_decap_8 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_367 ();
 sg13g2_decap_8 FILLER_23_374 ();
 sg13g2_decap_8 FILLER_23_381 ();
 sg13g2_decap_8 FILLER_23_388 ();
 sg13g2_decap_8 FILLER_23_395 ();
 sg13g2_decap_8 FILLER_23_402 ();
 sg13g2_decap_8 FILLER_23_409 ();
 sg13g2_decap_8 FILLER_23_416 ();
 sg13g2_decap_8 FILLER_23_423 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_fill_2 FILLER_24_14 ();
 sg13g2_fill_1 FILLER_24_16 ();
 sg13g2_fill_2 FILLER_24_107 ();
 sg13g2_decap_8 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_125 ();
 sg13g2_decap_4 FILLER_24_132 ();
 sg13g2_fill_1 FILLER_24_136 ();
 sg13g2_fill_2 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_175 ();
 sg13g2_fill_2 FILLER_24_194 ();
 sg13g2_fill_1 FILLER_24_196 ();
 sg13g2_fill_2 FILLER_24_213 ();
 sg13g2_fill_2 FILLER_24_218 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_fill_1 FILLER_24_247 ();
 sg13g2_decap_8 FILLER_24_253 ();
 sg13g2_decap_8 FILLER_24_296 ();
 sg13g2_decap_4 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_307 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_2 FILLER_24_321 ();
 sg13g2_fill_1 FILLER_24_327 ();
 sg13g2_decap_8 FILLER_24_332 ();
 sg13g2_decap_8 FILLER_24_339 ();
 sg13g2_decap_8 FILLER_24_346 ();
 sg13g2_decap_8 FILLER_24_353 ();
 sg13g2_decap_8 FILLER_24_360 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_24_409 ();
 sg13g2_decap_8 FILLER_24_416 ();
 sg13g2_decap_8 FILLER_24_423 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_4 FILLER_25_21 ();
 sg13g2_fill_1 FILLER_25_25 ();
 sg13g2_fill_1 FILLER_25_38 ();
 sg13g2_fill_2 FILLER_25_51 ();
 sg13g2_fill_1 FILLER_25_56 ();
 sg13g2_fill_1 FILLER_25_69 ();
 sg13g2_decap_8 FILLER_25_81 ();
 sg13g2_decap_8 FILLER_25_88 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_decap_8 FILLER_25_102 ();
 sg13g2_decap_4 FILLER_25_109 ();
 sg13g2_fill_1 FILLER_25_113 ();
 sg13g2_decap_4 FILLER_25_129 ();
 sg13g2_fill_2 FILLER_25_133 ();
 sg13g2_fill_1 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_156 ();
 sg13g2_decap_4 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_167 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_199 ();
 sg13g2_fill_2 FILLER_25_206 ();
 sg13g2_fill_2 FILLER_25_233 ();
 sg13g2_fill_2 FILLER_25_239 ();
 sg13g2_fill_1 FILLER_25_241 ();
 sg13g2_decap_8 FILLER_25_255 ();
 sg13g2_decap_8 FILLER_25_262 ();
 sg13g2_decap_4 FILLER_25_269 ();
 sg13g2_fill_1 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_284 ();
 sg13g2_decap_4 FILLER_25_316 ();
 sg13g2_fill_1 FILLER_25_320 ();
 sg13g2_fill_2 FILLER_25_324 ();
 sg13g2_fill_1 FILLER_25_326 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_decap_8 FILLER_25_347 ();
 sg13g2_decap_8 FILLER_25_354 ();
 sg13g2_decap_8 FILLER_25_361 ();
 sg13g2_decap_8 FILLER_25_368 ();
 sg13g2_decap_8 FILLER_25_375 ();
 sg13g2_decap_8 FILLER_25_382 ();
 sg13g2_decap_8 FILLER_25_389 ();
 sg13g2_decap_8 FILLER_25_396 ();
 sg13g2_decap_8 FILLER_25_403 ();
 sg13g2_decap_8 FILLER_25_410 ();
 sg13g2_decap_8 FILLER_25_417 ();
 sg13g2_decap_4 FILLER_25_424 ();
 sg13g2_fill_2 FILLER_25_428 ();
 sg13g2_fill_2 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_2 ();
 sg13g2_decap_8 FILLER_26_36 ();
 sg13g2_fill_1 FILLER_26_43 ();
 sg13g2_decap_4 FILLER_26_52 ();
 sg13g2_fill_2 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_fill_2 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_4 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_130 ();
 sg13g2_decap_8 FILLER_26_137 ();
 sg13g2_decap_8 FILLER_26_144 ();
 sg13g2_decap_4 FILLER_26_151 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_2 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_188 ();
 sg13g2_decap_4 FILLER_26_203 ();
 sg13g2_fill_2 FILLER_26_207 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_4 FILLER_26_245 ();
 sg13g2_decap_4 FILLER_26_254 ();
 sg13g2_fill_1 FILLER_26_258 ();
 sg13g2_fill_1 FILLER_26_267 ();
 sg13g2_fill_1 FILLER_26_272 ();
 sg13g2_fill_1 FILLER_26_276 ();
 sg13g2_fill_1 FILLER_26_281 ();
 sg13g2_decap_4 FILLER_26_287 ();
 sg13g2_fill_2 FILLER_26_291 ();
 sg13g2_fill_1 FILLER_26_297 ();
 sg13g2_fill_2 FILLER_26_312 ();
 sg13g2_fill_1 FILLER_26_314 ();
 sg13g2_decap_8 FILLER_26_319 ();
 sg13g2_fill_2 FILLER_26_326 ();
 sg13g2_decap_8 FILLER_26_341 ();
 sg13g2_decap_8 FILLER_26_348 ();
 sg13g2_decap_8 FILLER_26_355 ();
 sg13g2_decap_8 FILLER_26_362 ();
 sg13g2_decap_8 FILLER_26_369 ();
 sg13g2_decap_8 FILLER_26_376 ();
 sg13g2_decap_8 FILLER_26_383 ();
 sg13g2_decap_8 FILLER_26_390 ();
 sg13g2_decap_8 FILLER_26_397 ();
 sg13g2_decap_8 FILLER_26_404 ();
 sg13g2_decap_8 FILLER_26_411 ();
 sg13g2_decap_8 FILLER_26_418 ();
 sg13g2_decap_4 FILLER_26_425 ();
 sg13g2_fill_1 FILLER_26_429 ();
 sg13g2_decap_8 FILLER_27_0 ();
 sg13g2_decap_4 FILLER_27_7 ();
 sg13g2_decap_4 FILLER_27_15 ();
 sg13g2_fill_2 FILLER_27_23 ();
 sg13g2_fill_1 FILLER_27_25 ();
 sg13g2_decap_8 FILLER_27_39 ();
 sg13g2_decap_4 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_80 ();
 sg13g2_fill_2 FILLER_27_95 ();
 sg13g2_fill_2 FILLER_27_113 ();
 sg13g2_fill_1 FILLER_27_128 ();
 sg13g2_decap_8 FILLER_27_138 ();
 sg13g2_decap_8 FILLER_27_145 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_decap_8 FILLER_27_159 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_4 FILLER_27_228 ();
 sg13g2_fill_2 FILLER_27_232 ();
 sg13g2_decap_4 FILLER_27_239 ();
 sg13g2_fill_1 FILLER_27_243 ();
 sg13g2_fill_1 FILLER_27_282 ();
 sg13g2_decap_8 FILLER_27_301 ();
 sg13g2_decap_8 FILLER_27_308 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_1 FILLER_27_339 ();
 sg13g2_decap_8 FILLER_27_345 ();
 sg13g2_decap_8 FILLER_27_352 ();
 sg13g2_decap_8 FILLER_27_359 ();
 sg13g2_decap_8 FILLER_27_366 ();
 sg13g2_decap_8 FILLER_27_373 ();
 sg13g2_decap_8 FILLER_27_380 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_decap_8 FILLER_27_415 ();
 sg13g2_decap_8 FILLER_27_422 ();
 sg13g2_fill_1 FILLER_27_429 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_decap_4 FILLER_28_30 ();
 sg13g2_fill_2 FILLER_28_39 ();
 sg13g2_fill_1 FILLER_28_41 ();
 sg13g2_decap_8 FILLER_28_47 ();
 sg13g2_decap_8 FILLER_28_54 ();
 sg13g2_decap_8 FILLER_28_61 ();
 sg13g2_decap_4 FILLER_28_68 ();
 sg13g2_fill_1 FILLER_28_85 ();
 sg13g2_fill_2 FILLER_28_99 ();
 sg13g2_fill_1 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_130 ();
 sg13g2_decap_8 FILLER_28_143 ();
 sg13g2_decap_8 FILLER_28_150 ();
 sg13g2_fill_1 FILLER_28_157 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_fill_2 FILLER_28_175 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_192 ();
 sg13g2_fill_1 FILLER_28_196 ();
 sg13g2_fill_1 FILLER_28_207 ();
 sg13g2_fill_2 FILLER_28_213 ();
 sg13g2_fill_2 FILLER_28_241 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_283 ();
 sg13g2_decap_8 FILLER_28_292 ();
 sg13g2_decap_8 FILLER_28_299 ();
 sg13g2_fill_1 FILLER_28_306 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_fill_2 FILLER_28_322 ();
 sg13g2_fill_2 FILLER_28_345 ();
 sg13g2_decap_8 FILLER_28_360 ();
 sg13g2_decap_8 FILLER_28_367 ();
 sg13g2_decap_8 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_decap_8 FILLER_28_409 ();
 sg13g2_decap_8 FILLER_28_416 ();
 sg13g2_decap_8 FILLER_28_423 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_2 FILLER_29_7 ();
 sg13g2_decap_8 FILLER_29_43 ();
 sg13g2_fill_2 FILLER_29_50 ();
 sg13g2_fill_1 FILLER_29_52 ();
 sg13g2_decap_8 FILLER_29_58 ();
 sg13g2_decap_8 FILLER_29_65 ();
 sg13g2_decap_8 FILLER_29_72 ();
 sg13g2_decap_4 FILLER_29_79 ();
 sg13g2_fill_1 FILLER_29_83 ();
 sg13g2_decap_4 FILLER_29_89 ();
 sg13g2_fill_2 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_119 ();
 sg13g2_fill_1 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_130 ();
 sg13g2_fill_2 FILLER_29_140 ();
 sg13g2_decap_8 FILLER_29_155 ();
 sg13g2_decap_8 FILLER_29_162 ();
 sg13g2_decap_8 FILLER_29_169 ();
 sg13g2_decap_8 FILLER_29_176 ();
 sg13g2_decap_8 FILLER_29_183 ();
 sg13g2_decap_8 FILLER_29_190 ();
 sg13g2_fill_2 FILLER_29_201 ();
 sg13g2_fill_1 FILLER_29_203 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_fill_2 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_241 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_decap_8 FILLER_29_253 ();
 sg13g2_decap_8 FILLER_29_264 ();
 sg13g2_decap_8 FILLER_29_271 ();
 sg13g2_decap_4 FILLER_29_278 ();
 sg13g2_fill_1 FILLER_29_299 ();
 sg13g2_decap_4 FILLER_29_323 ();
 sg13g2_fill_2 FILLER_29_327 ();
 sg13g2_decap_8 FILLER_29_334 ();
 sg13g2_fill_2 FILLER_29_341 ();
 sg13g2_fill_1 FILLER_29_343 ();
 sg13g2_decap_8 FILLER_29_357 ();
 sg13g2_decap_8 FILLER_29_364 ();
 sg13g2_decap_8 FILLER_29_371 ();
 sg13g2_decap_8 FILLER_29_378 ();
 sg13g2_decap_8 FILLER_29_385 ();
 sg13g2_decap_8 FILLER_29_392 ();
 sg13g2_decap_8 FILLER_29_399 ();
 sg13g2_decap_8 FILLER_29_406 ();
 sg13g2_decap_8 FILLER_29_413 ();
 sg13g2_decap_8 FILLER_29_420 ();
 sg13g2_fill_2 FILLER_29_427 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_fill_1 FILLER_30_13 ();
 sg13g2_fill_2 FILLER_30_18 ();
 sg13g2_fill_1 FILLER_30_25 ();
 sg13g2_fill_2 FILLER_30_39 ();
 sg13g2_fill_1 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_52 ();
 sg13g2_decap_8 FILLER_30_74 ();
 sg13g2_decap_8 FILLER_30_81 ();
 sg13g2_decap_4 FILLER_30_95 ();
 sg13g2_fill_1 FILLER_30_99 ();
 sg13g2_fill_2 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_117 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_128 ();
 sg13g2_fill_1 FILLER_30_133 ();
 sg13g2_fill_2 FILLER_30_139 ();
 sg13g2_fill_2 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_146 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_fill_2 FILLER_30_157 ();
 sg13g2_fill_1 FILLER_30_159 ();
 sg13g2_decap_8 FILLER_30_164 ();
 sg13g2_decap_8 FILLER_30_171 ();
 sg13g2_decap_8 FILLER_30_178 ();
 sg13g2_fill_1 FILLER_30_185 ();
 sg13g2_decap_4 FILLER_30_189 ();
 sg13g2_fill_1 FILLER_30_193 ();
 sg13g2_fill_1 FILLER_30_201 ();
 sg13g2_decap_8 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_257 ();
 sg13g2_fill_1 FILLER_30_259 ();
 sg13g2_decap_4 FILLER_30_265 ();
 sg13g2_decap_8 FILLER_30_272 ();
 sg13g2_decap_8 FILLER_30_279 ();
 sg13g2_decap_8 FILLER_30_286 ();
 sg13g2_decap_8 FILLER_30_293 ();
 sg13g2_decap_4 FILLER_30_300 ();
 sg13g2_fill_1 FILLER_30_304 ();
 sg13g2_fill_1 FILLER_30_314 ();
 sg13g2_decap_8 FILLER_30_328 ();
 sg13g2_decap_8 FILLER_30_335 ();
 sg13g2_decap_4 FILLER_30_342 ();
 sg13g2_decap_8 FILLER_30_351 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_2 FILLER_31_36 ();
 sg13g2_decap_8 FILLER_31_41 ();
 sg13g2_fill_2 FILLER_31_48 ();
 sg13g2_fill_2 FILLER_31_57 ();
 sg13g2_fill_1 FILLER_31_68 ();
 sg13g2_decap_8 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_84 ();
 sg13g2_fill_2 FILLER_31_91 ();
 sg13g2_fill_1 FILLER_31_98 ();
 sg13g2_decap_4 FILLER_31_117 ();
 sg13g2_fill_1 FILLER_31_121 ();
 sg13g2_fill_2 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_146 ();
 sg13g2_fill_1 FILLER_31_158 ();
 sg13g2_fill_2 FILLER_31_165 ();
 sg13g2_fill_1 FILLER_31_171 ();
 sg13g2_fill_1 FILLER_31_206 ();
 sg13g2_fill_2 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_264 ();
 sg13g2_decap_8 FILLER_31_271 ();
 sg13g2_decap_8 FILLER_31_295 ();
 sg13g2_decap_8 FILLER_31_302 ();
 sg13g2_decap_8 FILLER_31_309 ();
 sg13g2_decap_4 FILLER_31_316 ();
 sg13g2_fill_1 FILLER_31_334 ();
 sg13g2_fill_2 FILLER_31_340 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_381 ();
 sg13g2_decap_8 FILLER_31_388 ();
 sg13g2_decap_8 FILLER_31_395 ();
 sg13g2_decap_8 FILLER_31_402 ();
 sg13g2_decap_8 FILLER_31_409 ();
 sg13g2_decap_8 FILLER_31_416 ();
 sg13g2_decap_8 FILLER_31_423 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_72 ();
 sg13g2_fill_2 FILLER_32_79 ();
 sg13g2_fill_1 FILLER_32_81 ();
 sg13g2_fill_2 FILLER_32_105 ();
 sg13g2_decap_4 FILLER_32_119 ();
 sg13g2_fill_2 FILLER_32_123 ();
 sg13g2_fill_1 FILLER_32_170 ();
 sg13g2_decap_8 FILLER_32_202 ();
 sg13g2_decap_8 FILLER_32_209 ();
 sg13g2_decap_4 FILLER_32_216 ();
 sg13g2_fill_2 FILLER_32_220 ();
 sg13g2_fill_2 FILLER_32_233 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_262 ();
 sg13g2_fill_2 FILLER_32_269 ();
 sg13g2_decap_8 FILLER_32_283 ();
 sg13g2_fill_1 FILLER_32_290 ();
 sg13g2_decap_8 FILLER_32_304 ();
 sg13g2_decap_4 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_decap_8 FILLER_32_356 ();
 sg13g2_fill_1 FILLER_32_363 ();
 sg13g2_decap_8 FILLER_32_381 ();
 sg13g2_decap_8 FILLER_32_388 ();
 sg13g2_decap_8 FILLER_32_395 ();
 sg13g2_decap_8 FILLER_32_402 ();
 sg13g2_decap_8 FILLER_32_409 ();
 sg13g2_decap_8 FILLER_32_416 ();
 sg13g2_decap_8 FILLER_32_423 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_29 ();
 sg13g2_decap_8 FILLER_33_36 ();
 sg13g2_fill_2 FILLER_33_43 ();
 sg13g2_fill_1 FILLER_33_45 ();
 sg13g2_fill_2 FILLER_33_50 ();
 sg13g2_fill_1 FILLER_33_52 ();
 sg13g2_fill_2 FILLER_33_58 ();
 sg13g2_decap_8 FILLER_33_67 ();
 sg13g2_decap_8 FILLER_33_74 ();
 sg13g2_decap_4 FILLER_33_81 ();
 sg13g2_fill_1 FILLER_33_85 ();
 sg13g2_decap_8 FILLER_33_89 ();
 sg13g2_decap_4 FILLER_33_96 ();
 sg13g2_fill_2 FILLER_33_100 ();
 sg13g2_decap_8 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_135 ();
 sg13g2_fill_2 FILLER_33_141 ();
 sg13g2_fill_2 FILLER_33_152 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_fill_1 FILLER_33_175 ();
 sg13g2_fill_2 FILLER_33_180 ();
 sg13g2_fill_1 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_263 ();
 sg13g2_fill_2 FILLER_33_270 ();
 sg13g2_fill_2 FILLER_33_276 ();
 sg13g2_fill_1 FILLER_33_278 ();
 sg13g2_decap_8 FILLER_33_283 ();
 sg13g2_decap_8 FILLER_33_290 ();
 sg13g2_fill_2 FILLER_33_297 ();
 sg13g2_decap_8 FILLER_33_303 ();
 sg13g2_decap_8 FILLER_33_310 ();
 sg13g2_decap_8 FILLER_33_317 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_326 ();
 sg13g2_fill_2 FILLER_33_331 ();
 sg13g2_decap_4 FILLER_33_357 ();
 sg13g2_fill_2 FILLER_33_366 ();
 sg13g2_decap_4 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_394 ();
 sg13g2_decap_8 FILLER_33_401 ();
 sg13g2_decap_8 FILLER_33_408 ();
 sg13g2_decap_8 FILLER_33_415 ();
 sg13g2_decap_8 FILLER_33_422 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_decap_8 FILLER_34_7 ();
 sg13g2_decap_4 FILLER_34_17 ();
 sg13g2_decap_8 FILLER_34_30 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_decap_8 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_77 ();
 sg13g2_fill_2 FILLER_34_90 ();
 sg13g2_decap_4 FILLER_34_95 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_115 ();
 sg13g2_fill_1 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_155 ();
 sg13g2_decap_8 FILLER_34_162 ();
 sg13g2_decap_8 FILLER_34_169 ();
 sg13g2_decap_8 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_8 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_197 ();
 sg13g2_fill_2 FILLER_34_213 ();
 sg13g2_fill_1 FILLER_34_219 ();
 sg13g2_fill_1 FILLER_34_225 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_fill_1 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_279 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_4 FILLER_34_291 ();
 sg13g2_decap_4 FILLER_34_300 ();
 sg13g2_fill_1 FILLER_34_317 ();
 sg13g2_fill_1 FILLER_34_358 ();
 sg13g2_fill_1 FILLER_34_363 ();
 sg13g2_fill_2 FILLER_34_373 ();
 sg13g2_fill_1 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_407 ();
 sg13g2_decap_8 FILLER_34_414 ();
 sg13g2_decap_8 FILLER_34_421 ();
 sg13g2_fill_2 FILLER_34_428 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_14 ();
 sg13g2_fill_2 FILLER_35_21 ();
 sg13g2_fill_2 FILLER_35_28 ();
 sg13g2_decap_4 FILLER_35_35 ();
 sg13g2_fill_1 FILLER_35_39 ();
 sg13g2_fill_2 FILLER_35_43 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_fill_2 FILLER_35_77 ();
 sg13g2_fill_1 FILLER_35_89 ();
 sg13g2_decap_4 FILLER_35_93 ();
 sg13g2_fill_2 FILLER_35_97 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_2 FILLER_35_125 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_fill_2 FILLER_35_147 ();
 sg13g2_fill_1 FILLER_35_149 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_decap_8 FILLER_35_169 ();
 sg13g2_decap_8 FILLER_35_176 ();
 sg13g2_fill_2 FILLER_35_183 ();
 sg13g2_fill_1 FILLER_35_185 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_232 ();
 sg13g2_decap_8 FILLER_35_239 ();
 sg13g2_decap_8 FILLER_35_246 ();
 sg13g2_decap_4 FILLER_35_253 ();
 sg13g2_decap_8 FILLER_35_265 ();
 sg13g2_decap_8 FILLER_35_272 ();
 sg13g2_fill_2 FILLER_35_279 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_4 FILLER_35_301 ();
 sg13g2_fill_2 FILLER_35_315 ();
 sg13g2_fill_1 FILLER_35_322 ();
 sg13g2_fill_2 FILLER_35_331 ();
 sg13g2_decap_8 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_371 ();
 sg13g2_fill_2 FILLER_35_386 ();
 sg13g2_decap_8 FILLER_35_401 ();
 sg13g2_decap_8 FILLER_35_408 ();
 sg13g2_decap_8 FILLER_35_415 ();
 sg13g2_decap_8 FILLER_35_422 ();
 sg13g2_fill_1 FILLER_35_429 ();
 sg13g2_decap_4 FILLER_36_52 ();
 sg13g2_fill_2 FILLER_36_56 ();
 sg13g2_decap_4 FILLER_36_66 ();
 sg13g2_fill_1 FILLER_36_70 ();
 sg13g2_fill_2 FILLER_36_87 ();
 sg13g2_decap_8 FILLER_36_94 ();
 sg13g2_fill_2 FILLER_36_101 ();
 sg13g2_fill_2 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_120 ();
 sg13g2_fill_1 FILLER_36_122 ();
 sg13g2_fill_2 FILLER_36_142 ();
 sg13g2_fill_1 FILLER_36_144 ();
 sg13g2_decap_4 FILLER_36_169 ();
 sg13g2_fill_1 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_1 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_215 ();
 sg13g2_decap_8 FILLER_36_222 ();
 sg13g2_decap_8 FILLER_36_229 ();
 sg13g2_decap_4 FILLER_36_236 ();
 sg13g2_decap_8 FILLER_36_244 ();
 sg13g2_decap_4 FILLER_36_251 ();
 sg13g2_fill_2 FILLER_36_255 ();
 sg13g2_decap_8 FILLER_36_278 ();
 sg13g2_decap_8 FILLER_36_285 ();
 sg13g2_fill_1 FILLER_36_292 ();
 sg13g2_fill_2 FILLER_36_309 ();
 sg13g2_fill_1 FILLER_36_311 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_1 FILLER_36_319 ();
 sg13g2_fill_1 FILLER_36_327 ();
 sg13g2_fill_2 FILLER_36_353 ();
 sg13g2_fill_1 FILLER_36_359 ();
 sg13g2_decap_8 FILLER_36_377 ();
 sg13g2_decap_8 FILLER_36_384 ();
 sg13g2_decap_8 FILLER_36_404 ();
 sg13g2_decap_8 FILLER_36_411 ();
 sg13g2_decap_8 FILLER_36_418 ();
 sg13g2_decap_4 FILLER_36_425 ();
 sg13g2_fill_1 FILLER_36_429 ();
 sg13g2_decap_4 FILLER_37_73 ();
 sg13g2_fill_1 FILLER_37_77 ();
 sg13g2_fill_2 FILLER_37_83 ();
 sg13g2_fill_1 FILLER_37_85 ();
 sg13g2_fill_1 FILLER_37_89 ();
 sg13g2_fill_2 FILLER_37_94 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_decap_8 FILLER_37_106 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_fill_2 FILLER_37_137 ();
 sg13g2_fill_1 FILLER_37_149 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_4 FILLER_37_179 ();
 sg13g2_fill_1 FILLER_37_183 ();
 sg13g2_fill_1 FILLER_37_202 ();
 sg13g2_decap_8 FILLER_37_215 ();
 sg13g2_decap_8 FILLER_37_222 ();
 sg13g2_fill_1 FILLER_37_229 ();
 sg13g2_fill_2 FILLER_37_237 ();
 sg13g2_decap_8 FILLER_37_275 ();
 sg13g2_decap_8 FILLER_37_282 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_fill_2 FILLER_37_338 ();
 sg13g2_fill_1 FILLER_37_340 ();
 sg13g2_fill_1 FILLER_37_349 ();
 sg13g2_fill_2 FILLER_37_356 ();
 sg13g2_fill_1 FILLER_37_376 ();
 sg13g2_fill_1 FILLER_37_381 ();
 sg13g2_fill_2 FILLER_37_387 ();
 sg13g2_fill_1 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_408 ();
 sg13g2_decap_8 FILLER_37_415 ();
 sg13g2_decap_8 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_decap_4 FILLER_38_18 ();
 sg13g2_decap_8 FILLER_38_30 ();
 sg13g2_fill_2 FILLER_38_37 ();
 sg13g2_fill_1 FILLER_38_39 ();
 sg13g2_fill_2 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_60 ();
 sg13g2_fill_1 FILLER_38_62 ();
 sg13g2_decap_8 FILLER_38_66 ();
 sg13g2_decap_4 FILLER_38_73 ();
 sg13g2_decap_4 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_93 ();
 sg13g2_fill_2 FILLER_38_97 ();
 sg13g2_decap_8 FILLER_38_107 ();
 sg13g2_decap_8 FILLER_38_114 ();
 sg13g2_decap_4 FILLER_38_121 ();
 sg13g2_fill_2 FILLER_38_125 ();
 sg13g2_decap_4 FILLER_38_149 ();
 sg13g2_fill_2 FILLER_38_157 ();
 sg13g2_fill_1 FILLER_38_163 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_4 FILLER_38_182 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_decap_8 FILLER_38_200 ();
 sg13g2_decap_8 FILLER_38_211 ();
 sg13g2_decap_4 FILLER_38_218 ();
 sg13g2_decap_8 FILLER_38_271 ();
 sg13g2_decap_8 FILLER_38_278 ();
 sg13g2_decap_4 FILLER_38_285 ();
 sg13g2_fill_1 FILLER_38_289 ();
 sg13g2_decap_8 FILLER_38_295 ();
 sg13g2_fill_2 FILLER_38_302 ();
 sg13g2_fill_1 FILLER_38_304 ();
 sg13g2_fill_1 FILLER_38_317 ();
 sg13g2_fill_2 FILLER_38_326 ();
 sg13g2_fill_1 FILLER_38_328 ();
 sg13g2_decap_8 FILLER_38_341 ();
 sg13g2_decap_4 FILLER_38_359 ();
 sg13g2_fill_1 FILLER_38_363 ();
 sg13g2_fill_1 FILLER_38_373 ();
 sg13g2_fill_1 FILLER_38_390 ();
 sg13g2_decap_8 FILLER_38_422 ();
 sg13g2_fill_1 FILLER_38_429 ();
 sg13g2_decap_8 FILLER_39_0 ();
 sg13g2_decap_8 FILLER_39_7 ();
 sg13g2_fill_2 FILLER_39_14 ();
 sg13g2_fill_2 FILLER_39_21 ();
 sg13g2_fill_1 FILLER_39_23 ();
 sg13g2_fill_2 FILLER_39_37 ();
 sg13g2_decap_8 FILLER_39_42 ();
 sg13g2_decap_8 FILLER_39_49 ();
 sg13g2_decap_8 FILLER_39_56 ();
 sg13g2_decap_8 FILLER_39_63 ();
 sg13g2_decap_8 FILLER_39_70 ();
 sg13g2_fill_1 FILLER_39_85 ();
 sg13g2_fill_2 FILLER_39_89 ();
 sg13g2_fill_1 FILLER_39_91 ();
 sg13g2_decap_4 FILLER_39_100 ();
 sg13g2_fill_1 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_128 ();
 sg13g2_fill_2 FILLER_39_161 ();
 sg13g2_fill_1 FILLER_39_163 ();
 sg13g2_decap_8 FILLER_39_167 ();
 sg13g2_decap_8 FILLER_39_174 ();
 sg13g2_decap_4 FILLER_39_181 ();
 sg13g2_fill_2 FILLER_39_231 ();
 sg13g2_fill_2 FILLER_39_261 ();
 sg13g2_fill_1 FILLER_39_271 ();
 sg13g2_fill_1 FILLER_39_275 ();
 sg13g2_fill_1 FILLER_39_281 ();
 sg13g2_fill_1 FILLER_39_295 ();
 sg13g2_decap_4 FILLER_39_301 ();
 sg13g2_fill_2 FILLER_39_305 ();
 sg13g2_fill_2 FILLER_39_322 ();
 sg13g2_fill_1 FILLER_39_329 ();
 sg13g2_fill_2 FILLER_39_341 ();
 sg13g2_fill_1 FILLER_39_343 ();
 sg13g2_decap_8 FILLER_39_352 ();
 sg13g2_decap_4 FILLER_39_359 ();
 sg13g2_fill_1 FILLER_39_372 ();
 sg13g2_fill_1 FILLER_39_377 ();
 sg13g2_decap_4 FILLER_39_389 ();
 sg13g2_fill_2 FILLER_39_393 ();
 sg13g2_fill_2 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_406 ();
 sg13g2_decap_8 FILLER_39_412 ();
 sg13g2_decap_8 FILLER_39_419 ();
 sg13g2_decap_4 FILLER_39_426 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_fill_2 FILLER_40_17 ();
 sg13g2_fill_1 FILLER_40_34 ();
 sg13g2_decap_4 FILLER_40_47 ();
 sg13g2_fill_2 FILLER_40_51 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_4 FILLER_40_63 ();
 sg13g2_fill_1 FILLER_40_67 ();
 sg13g2_fill_2 FILLER_40_83 ();
 sg13g2_fill_1 FILLER_40_89 ();
 sg13g2_fill_1 FILLER_40_129 ();
 sg13g2_fill_2 FILLER_40_153 ();
 sg13g2_fill_1 FILLER_40_159 ();
 sg13g2_fill_1 FILLER_40_165 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_1 FILLER_40_184 ();
 sg13g2_decap_4 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_207 ();
 sg13g2_decap_4 FILLER_40_214 ();
 sg13g2_fill_1 FILLER_40_218 ();
 sg13g2_fill_2 FILLER_40_224 ();
 sg13g2_fill_2 FILLER_40_231 ();
 sg13g2_fill_2 FILLER_40_242 ();
 sg13g2_fill_1 FILLER_40_244 ();
 sg13g2_decap_4 FILLER_40_249 ();
 sg13g2_fill_2 FILLER_40_256 ();
 sg13g2_fill_1 FILLER_40_258 ();
 sg13g2_decap_8 FILLER_40_270 ();
 sg13g2_decap_8 FILLER_40_277 ();
 sg13g2_decap_8 FILLER_40_284 ();
 sg13g2_decap_4 FILLER_40_291 ();
 sg13g2_fill_2 FILLER_40_299 ();
 sg13g2_fill_1 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_326 ();
 sg13g2_decap_8 FILLER_40_333 ();
 sg13g2_fill_2 FILLER_40_340 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_fill_1 FILLER_40_369 ();
 sg13g2_decap_4 FILLER_40_383 ();
 sg13g2_fill_2 FILLER_40_387 ();
 sg13g2_fill_1 FILLER_40_398 ();
 sg13g2_decap_8 FILLER_40_417 ();
 sg13g2_decap_4 FILLER_40_424 ();
 sg13g2_fill_2 FILLER_40_428 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_fill_2 FILLER_41_14 ();
 sg13g2_fill_1 FILLER_41_16 ();
 sg13g2_fill_2 FILLER_41_21 ();
 sg13g2_fill_1 FILLER_41_30 ();
 sg13g2_fill_2 FILLER_41_62 ();
 sg13g2_fill_1 FILLER_41_64 ();
 sg13g2_fill_1 FILLER_41_74 ();
 sg13g2_fill_1 FILLER_41_85 ();
 sg13g2_fill_2 FILLER_41_90 ();
 sg13g2_fill_1 FILLER_41_97 ();
 sg13g2_fill_1 FILLER_41_104 ();
 sg13g2_fill_1 FILLER_41_108 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_fill_2 FILLER_41_119 ();
 sg13g2_fill_1 FILLER_41_138 ();
 sg13g2_decap_8 FILLER_41_169 ();
 sg13g2_fill_2 FILLER_41_176 ();
 sg13g2_fill_2 FILLER_41_186 ();
 sg13g2_fill_1 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_199 ();
 sg13g2_decap_8 FILLER_41_206 ();
 sg13g2_decap_8 FILLER_41_213 ();
 sg13g2_fill_2 FILLER_41_220 ();
 sg13g2_fill_1 FILLER_41_222 ();
 sg13g2_decap_8 FILLER_41_228 ();
 sg13g2_decap_8 FILLER_41_235 ();
 sg13g2_decap_8 FILLER_41_242 ();
 sg13g2_fill_1 FILLER_41_254 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_4 FILLER_41_294 ();
 sg13g2_decap_4 FILLER_41_302 ();
 sg13g2_fill_2 FILLER_41_306 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_fill_1 FILLER_41_344 ();
 sg13g2_decap_8 FILLER_41_353 ();
 sg13g2_decap_4 FILLER_41_364 ();
 sg13g2_fill_2 FILLER_41_368 ();
 sg13g2_fill_2 FILLER_41_388 ();
 sg13g2_fill_1 FILLER_41_390 ();
 sg13g2_decap_4 FILLER_41_395 ();
 sg13g2_decap_8 FILLER_41_421 ();
 sg13g2_fill_2 FILLER_41_428 ();
 sg13g2_fill_1 FILLER_42_18 ();
 sg13g2_fill_2 FILLER_42_63 ();
 sg13g2_fill_1 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_76 ();
 sg13g2_fill_2 FILLER_42_104 ();
 sg13g2_fill_2 FILLER_42_118 ();
 sg13g2_fill_1 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_131 ();
 sg13g2_fill_1 FILLER_42_153 ();
 sg13g2_decap_8 FILLER_42_159 ();
 sg13g2_fill_2 FILLER_42_166 ();
 sg13g2_fill_2 FILLER_42_194 ();
 sg13g2_fill_2 FILLER_42_200 ();
 sg13g2_fill_1 FILLER_42_202 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_decap_8 FILLER_42_215 ();
 sg13g2_decap_8 FILLER_42_222 ();
 sg13g2_decap_4 FILLER_42_229 ();
 sg13g2_fill_2 FILLER_42_233 ();
 sg13g2_decap_4 FILLER_42_243 ();
 sg13g2_decap_8 FILLER_42_251 ();
 sg13g2_decap_8 FILLER_42_258 ();
 sg13g2_decap_8 FILLER_42_265 ();
 sg13g2_decap_8 FILLER_42_272 ();
 sg13g2_decap_4 FILLER_42_279 ();
 sg13g2_fill_1 FILLER_42_283 ();
 sg13g2_decap_4 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_297 ();
 sg13g2_fill_1 FILLER_42_306 ();
 sg13g2_decap_4 FILLER_42_321 ();
 sg13g2_fill_1 FILLER_42_325 ();
 sg13g2_fill_1 FILLER_42_330 ();
 sg13g2_fill_1 FILLER_42_368 ();
 sg13g2_fill_2 FILLER_42_378 ();
 sg13g2_decap_4 FILLER_42_389 ();
 sg13g2_decap_4 FILLER_42_398 ();
 sg13g2_decap_8 FILLER_42_412 ();
 sg13g2_decap_8 FILLER_42_419 ();
 sg13g2_decap_4 FILLER_42_426 ();
 sg13g2_fill_1 FILLER_43_0 ();
 sg13g2_fill_1 FILLER_43_27 ();
 sg13g2_fill_1 FILLER_43_33 ();
 sg13g2_fill_1 FILLER_43_39 ();
 sg13g2_decap_4 FILLER_43_44 ();
 sg13g2_fill_2 FILLER_43_55 ();
 sg13g2_fill_2 FILLER_43_61 ();
 sg13g2_decap_4 FILLER_43_68 ();
 sg13g2_decap_4 FILLER_43_77 ();
 sg13g2_decap_4 FILLER_43_88 ();
 sg13g2_fill_1 FILLER_43_92 ();
 sg13g2_fill_1 FILLER_43_97 ();
 sg13g2_decap_8 FILLER_43_110 ();
 sg13g2_fill_1 FILLER_43_121 ();
 sg13g2_decap_8 FILLER_43_157 ();
 sg13g2_decap_8 FILLER_43_164 ();
 sg13g2_decap_8 FILLER_43_171 ();
 sg13g2_decap_8 FILLER_43_178 ();
 sg13g2_decap_8 FILLER_43_185 ();
 sg13g2_fill_2 FILLER_43_192 ();
 sg13g2_decap_4 FILLER_43_202 ();
 sg13g2_decap_8 FILLER_43_219 ();
 sg13g2_decap_4 FILLER_43_256 ();
 sg13g2_fill_1 FILLER_43_260 ();
 sg13g2_fill_1 FILLER_43_269 ();
 sg13g2_decap_8 FILLER_43_279 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_fill_1 FILLER_43_296 ();
 sg13g2_fill_2 FILLER_43_307 ();
 sg13g2_fill_2 FILLER_43_313 ();
 sg13g2_fill_1 FILLER_43_315 ();
 sg13g2_fill_1 FILLER_43_342 ();
 sg13g2_fill_2 FILLER_43_353 ();
 sg13g2_fill_1 FILLER_43_355 ();
 sg13g2_fill_1 FILLER_43_406 ();
 sg13g2_decap_4 FILLER_43_424 ();
 sg13g2_fill_2 FILLER_43_428 ();
 sg13g2_fill_2 FILLER_44_35 ();
 sg13g2_decap_4 FILLER_44_41 ();
 sg13g2_fill_2 FILLER_44_45 ();
 sg13g2_decap_8 FILLER_44_63 ();
 sg13g2_decap_4 FILLER_44_70 ();
 sg13g2_decap_8 FILLER_44_80 ();
 sg13g2_decap_8 FILLER_44_87 ();
 sg13g2_fill_2 FILLER_44_94 ();
 sg13g2_fill_2 FILLER_44_115 ();
 sg13g2_fill_2 FILLER_44_128 ();
 sg13g2_fill_1 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_154 ();
 sg13g2_fill_2 FILLER_44_161 ();
 sg13g2_fill_1 FILLER_44_163 ();
 sg13g2_decap_8 FILLER_44_168 ();
 sg13g2_decap_8 FILLER_44_175 ();
 sg13g2_decap_8 FILLER_44_182 ();
 sg13g2_fill_1 FILLER_44_189 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_4 FILLER_44_210 ();
 sg13g2_fill_1 FILLER_44_214 ();
 sg13g2_fill_1 FILLER_44_240 ();
 sg13g2_fill_2 FILLER_44_249 ();
 sg13g2_fill_1 FILLER_44_251 ();
 sg13g2_decap_4 FILLER_44_256 ();
 sg13g2_fill_1 FILLER_44_268 ();
 sg13g2_decap_8 FILLER_44_279 ();
 sg13g2_decap_4 FILLER_44_286 ();
 sg13g2_fill_1 FILLER_44_290 ();
 sg13g2_decap_4 FILLER_44_295 ();
 sg13g2_fill_2 FILLER_44_299 ();
 sg13g2_fill_2 FILLER_44_306 ();
 sg13g2_fill_2 FILLER_44_320 ();
 sg13g2_fill_2 FILLER_44_346 ();
 sg13g2_fill_1 FILLER_44_348 ();
 sg13g2_fill_2 FILLER_44_354 ();
 sg13g2_fill_2 FILLER_44_360 ();
 sg13g2_fill_1 FILLER_44_376 ();
 sg13g2_fill_1 FILLER_44_382 ();
 sg13g2_fill_2 FILLER_44_386 ();
 sg13g2_fill_1 FILLER_44_392 ();
 sg13g2_fill_1 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_422 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_decap_4 FILLER_45_0 ();
 sg13g2_fill_2 FILLER_45_4 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_4 FILLER_45_35 ();
 sg13g2_decap_4 FILLER_45_47 ();
 sg13g2_fill_1 FILLER_45_51 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_4 FILLER_45_70 ();
 sg13g2_fill_1 FILLER_45_74 ();
 sg13g2_decap_4 FILLER_45_88 ();
 sg13g2_decap_4 FILLER_45_96 ();
 sg13g2_fill_1 FILLER_45_115 ();
 sg13g2_fill_1 FILLER_45_121 ();
 sg13g2_decap_4 FILLER_45_136 ();
 sg13g2_fill_2 FILLER_45_140 ();
 sg13g2_fill_2 FILLER_45_157 ();
 sg13g2_fill_1 FILLER_45_159 ();
 sg13g2_decap_4 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_180 ();
 sg13g2_decap_4 FILLER_45_187 ();
 sg13g2_decap_4 FILLER_45_196 ();
 sg13g2_fill_2 FILLER_45_200 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_209 ();
 sg13g2_fill_2 FILLER_45_246 ();
 sg13g2_fill_2 FILLER_45_260 ();
 sg13g2_decap_4 FILLER_45_266 ();
 sg13g2_fill_1 FILLER_45_270 ();
 sg13g2_decap_8 FILLER_45_276 ();
 sg13g2_decap_8 FILLER_45_283 ();
 sg13g2_fill_1 FILLER_45_290 ();
 sg13g2_fill_2 FILLER_45_303 ();
 sg13g2_fill_1 FILLER_45_305 ();
 sg13g2_fill_2 FILLER_45_312 ();
 sg13g2_decap_8 FILLER_45_319 ();
 sg13g2_fill_1 FILLER_45_335 ();
 sg13g2_fill_1 FILLER_45_340 ();
 sg13g2_decap_4 FILLER_45_351 ();
 sg13g2_fill_2 FILLER_45_359 ();
 sg13g2_decap_8 FILLER_45_365 ();
 sg13g2_decap_8 FILLER_45_372 ();
 sg13g2_fill_2 FILLER_45_379 ();
 sg13g2_fill_1 FILLER_45_381 ();
 sg13g2_fill_1 FILLER_45_387 ();
 sg13g2_fill_1 FILLER_45_392 ();
 sg13g2_fill_1 FILLER_45_401 ();
 sg13g2_fill_2 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_45_407 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_fill_2 FILLER_45_427 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_decap_4 FILLER_46_0 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_12 ();
 sg13g2_decap_8 FILLER_46_19 ();
 sg13g2_decap_4 FILLER_46_26 ();
 sg13g2_fill_1 FILLER_46_30 ();
 sg13g2_decap_8 FILLER_46_36 ();
 sg13g2_decap_8 FILLER_46_48 ();
 sg13g2_fill_2 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_63 ();
 sg13g2_fill_2 FILLER_46_69 ();
 sg13g2_fill_1 FILLER_46_71 ();
 sg13g2_fill_1 FILLER_46_82 ();
 sg13g2_fill_1 FILLER_46_88 ();
 sg13g2_fill_1 FILLER_46_93 ();
 sg13g2_fill_2 FILLER_46_99 ();
 sg13g2_fill_1 FILLER_46_108 ();
 sg13g2_fill_1 FILLER_46_120 ();
 sg13g2_fill_1 FILLER_46_125 ();
 sg13g2_decap_8 FILLER_46_134 ();
 sg13g2_decap_4 FILLER_46_146 ();
 sg13g2_fill_2 FILLER_46_155 ();
 sg13g2_fill_1 FILLER_46_178 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_fill_2 FILLER_46_198 ();
 sg13g2_fill_1 FILLER_46_204 ();
 sg13g2_fill_1 FILLER_46_236 ();
 sg13g2_decap_4 FILLER_46_247 ();
 sg13g2_fill_1 FILLER_46_262 ();
 sg13g2_decap_8 FILLER_46_289 ();
 sg13g2_fill_2 FILLER_46_296 ();
 sg13g2_fill_1 FILLER_46_298 ();
 sg13g2_fill_2 FILLER_46_308 ();
 sg13g2_fill_2 FILLER_46_318 ();
 sg13g2_fill_1 FILLER_46_320 ();
 sg13g2_fill_1 FILLER_46_338 ();
 sg13g2_fill_1 FILLER_46_342 ();
 sg13g2_decap_8 FILLER_46_348 ();
 sg13g2_decap_8 FILLER_46_355 ();
 sg13g2_decap_4 FILLER_46_374 ();
 sg13g2_fill_1 FILLER_46_378 ();
 sg13g2_fill_1 FILLER_46_383 ();
 sg13g2_fill_1 FILLER_46_392 ();
 sg13g2_fill_1 FILLER_46_397 ();
 sg13g2_fill_2 FILLER_46_412 ();
 sg13g2_decap_8 FILLER_46_418 ();
 sg13g2_decap_4 FILLER_46_425 ();
 sg13g2_fill_1 FILLER_46_429 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_4 FILLER_47_14 ();
 sg13g2_fill_1 FILLER_47_18 ();
 sg13g2_fill_2 FILLER_47_45 ();
 sg13g2_fill_1 FILLER_47_73 ();
 sg13g2_fill_2 FILLER_47_91 ();
 sg13g2_fill_2 FILLER_47_121 ();
 sg13g2_fill_1 FILLER_47_135 ();
 sg13g2_decap_4 FILLER_47_152 ();
 sg13g2_decap_4 FILLER_47_198 ();
 sg13g2_decap_8 FILLER_47_207 ();
 sg13g2_decap_8 FILLER_47_214 ();
 sg13g2_decap_8 FILLER_47_221 ();
 sg13g2_decap_8 FILLER_47_228 ();
 sg13g2_decap_8 FILLER_47_235 ();
 sg13g2_decap_8 FILLER_47_242 ();
 sg13g2_fill_1 FILLER_47_249 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_fill_2 FILLER_47_273 ();
 sg13g2_fill_1 FILLER_47_280 ();
 sg13g2_decap_4 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_293 ();
 sg13g2_decap_4 FILLER_47_299 ();
 sg13g2_decap_8 FILLER_47_307 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_1 FILLER_47_316 ();
 sg13g2_fill_2 FILLER_47_321 ();
 sg13g2_fill_1 FILLER_47_323 ();
 sg13g2_fill_1 FILLER_47_338 ();
 sg13g2_fill_1 FILLER_47_344 ();
 sg13g2_fill_1 FILLER_47_349 ();
 sg13g2_fill_1 FILLER_47_355 ();
 sg13g2_fill_1 FILLER_47_361 ();
 sg13g2_fill_2 FILLER_47_367 ();
 sg13g2_fill_2 FILLER_47_374 ();
 sg13g2_fill_1 FILLER_47_381 ();
 sg13g2_fill_2 FILLER_47_391 ();
 sg13g2_fill_1 FILLER_47_393 ();
 sg13g2_fill_1 FILLER_47_398 ();
 sg13g2_fill_2 FILLER_47_404 ();
 sg13g2_decap_8 FILLER_47_410 ();
 sg13g2_decap_8 FILLER_47_417 ();
 sg13g2_decap_4 FILLER_47_424 ();
 sg13g2_fill_2 FILLER_47_428 ();
 sg13g2_fill_1 FILLER_48_26 ();
 sg13g2_fill_1 FILLER_48_33 ();
 sg13g2_decap_4 FILLER_48_37 ();
 sg13g2_fill_1 FILLER_48_41 ();
 sg13g2_fill_2 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_55 ();
 sg13g2_fill_2 FILLER_48_62 ();
 sg13g2_fill_2 FILLER_48_69 ();
 sg13g2_fill_1 FILLER_48_71 ();
 sg13g2_decap_4 FILLER_48_106 ();
 sg13g2_fill_1 FILLER_48_110 ();
 sg13g2_fill_1 FILLER_48_116 ();
 sg13g2_decap_4 FILLER_48_121 ();
 sg13g2_decap_4 FILLER_48_133 ();
 sg13g2_decap_4 FILLER_48_142 ();
 sg13g2_fill_1 FILLER_48_146 ();
 sg13g2_fill_1 FILLER_48_173 ();
 sg13g2_fill_2 FILLER_48_179 ();
 sg13g2_fill_2 FILLER_48_185 ();
 sg13g2_fill_2 FILLER_48_195 ();
 sg13g2_fill_2 FILLER_48_200 ();
 sg13g2_fill_1 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_216 ();
 sg13g2_decap_8 FILLER_48_223 ();
 sg13g2_decap_8 FILLER_48_237 ();
 sg13g2_decap_8 FILLER_48_244 ();
 sg13g2_decap_8 FILLER_48_251 ();
 sg13g2_decap_8 FILLER_48_258 ();
 sg13g2_decap_8 FILLER_48_265 ();
 sg13g2_fill_1 FILLER_48_294 ();
 sg13g2_decap_4 FILLER_48_304 ();
 sg13g2_fill_2 FILLER_48_326 ();
 sg13g2_fill_2 FILLER_48_344 ();
 sg13g2_fill_2 FILLER_48_350 ();
 sg13g2_fill_2 FILLER_48_356 ();
 sg13g2_fill_2 FILLER_48_363 ();
 sg13g2_fill_1 FILLER_48_365 ();
 sg13g2_fill_1 FILLER_48_371 ();
 sg13g2_decap_4 FILLER_48_376 ();
 sg13g2_fill_2 FILLER_48_415 ();
 sg13g2_decap_8 FILLER_48_422 ();
 sg13g2_fill_1 FILLER_48_429 ();
 sg13g2_decap_8 FILLER_49_0 ();
 sg13g2_decap_4 FILLER_49_7 ();
 sg13g2_fill_1 FILLER_49_11 ();
 sg13g2_fill_2 FILLER_49_19 ();
 sg13g2_fill_2 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_35 ();
 sg13g2_fill_2 FILLER_49_51 ();
 sg13g2_fill_1 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_59 ();
 sg13g2_decap_8 FILLER_49_66 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_fill_2 FILLER_49_84 ();
 sg13g2_fill_1 FILLER_49_86 ();
 sg13g2_decap_4 FILLER_49_95 ();
 sg13g2_fill_2 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_106 ();
 sg13g2_decap_8 FILLER_49_111 ();
 sg13g2_fill_2 FILLER_49_118 ();
 sg13g2_decap_4 FILLER_49_124 ();
 sg13g2_decap_8 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_140 ();
 sg13g2_fill_2 FILLER_49_147 ();
 sg13g2_fill_2 FILLER_49_161 ();
 sg13g2_fill_1 FILLER_49_171 ();
 sg13g2_fill_2 FILLER_49_176 ();
 sg13g2_fill_1 FILLER_49_183 ();
 sg13g2_fill_1 FILLER_49_187 ();
 sg13g2_fill_1 FILLER_49_196 ();
 sg13g2_fill_1 FILLER_49_201 ();
 sg13g2_fill_2 FILLER_49_206 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_fill_1 FILLER_49_234 ();
 sg13g2_decap_8 FILLER_49_244 ();
 sg13g2_decap_8 FILLER_49_251 ();
 sg13g2_fill_2 FILLER_49_267 ();
 sg13g2_fill_1 FILLER_49_283 ();
 sg13g2_fill_2 FILLER_49_288 ();
 sg13g2_fill_2 FILLER_49_298 ();
 sg13g2_decap_4 FILLER_49_305 ();
 sg13g2_fill_1 FILLER_49_309 ();
 sg13g2_decap_8 FILLER_49_335 ();
 sg13g2_decap_8 FILLER_49_342 ();
 sg13g2_fill_1 FILLER_49_349 ();
 sg13g2_fill_2 FILLER_49_362 ();
 sg13g2_fill_1 FILLER_49_374 ();
 sg13g2_fill_2 FILLER_49_387 ();
 sg13g2_fill_2 FILLER_49_399 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_4 FILLER_49_424 ();
 sg13g2_fill_2 FILLER_49_428 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_4 FILLER_50_7 ();
 sg13g2_fill_2 FILLER_50_21 ();
 sg13g2_fill_1 FILLER_50_23 ();
 sg13g2_decap_4 FILLER_50_27 ();
 sg13g2_fill_1 FILLER_50_31 ();
 sg13g2_decap_8 FILLER_50_50 ();
 sg13g2_decap_8 FILLER_50_57 ();
 sg13g2_decap_8 FILLER_50_64 ();
 sg13g2_decap_8 FILLER_50_71 ();
 sg13g2_decap_8 FILLER_50_78 ();
 sg13g2_decap_4 FILLER_50_85 ();
 sg13g2_decap_8 FILLER_50_124 ();
 sg13g2_decap_8 FILLER_50_131 ();
 sg13g2_decap_8 FILLER_50_138 ();
 sg13g2_decap_4 FILLER_50_145 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_fill_1 FILLER_50_173 ();
 sg13g2_fill_1 FILLER_50_178 ();
 sg13g2_fill_1 FILLER_50_183 ();
 sg13g2_fill_1 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_194 ();
 sg13g2_decap_4 FILLER_50_206 ();
 sg13g2_fill_1 FILLER_50_221 ();
 sg13g2_fill_1 FILLER_50_226 ();
 sg13g2_fill_1 FILLER_50_231 ();
 sg13g2_fill_1 FILLER_50_238 ();
 sg13g2_decap_4 FILLER_50_243 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_fill_2 FILLER_50_283 ();
 sg13g2_decap_4 FILLER_50_291 ();
 sg13g2_fill_2 FILLER_50_295 ();
 sg13g2_decap_4 FILLER_50_304 ();
 sg13g2_fill_1 FILLER_50_308 ();
 sg13g2_fill_1 FILLER_50_313 ();
 sg13g2_decap_4 FILLER_50_318 ();
 sg13g2_fill_2 FILLER_50_327 ();
 sg13g2_fill_1 FILLER_50_329 ();
 sg13g2_fill_2 FILLER_50_334 ();
 sg13g2_decap_8 FILLER_50_347 ();
 sg13g2_decap_8 FILLER_50_375 ();
 sg13g2_fill_1 FILLER_50_382 ();
 sg13g2_fill_2 FILLER_50_396 ();
 sg13g2_fill_1 FILLER_50_398 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_fill_1 FILLER_50_413 ();
 sg13g2_decap_4 FILLER_50_426 ();
 sg13g2_fill_2 FILLER_51_0 ();
 sg13g2_fill_1 FILLER_51_26 ();
 sg13g2_fill_1 FILLER_51_40 ();
 sg13g2_decap_8 FILLER_51_67 ();
 sg13g2_fill_2 FILLER_51_74 ();
 sg13g2_decap_4 FILLER_51_86 ();
 sg13g2_decap_8 FILLER_51_94 ();
 sg13g2_fill_2 FILLER_51_106 ();
 sg13g2_decap_8 FILLER_51_116 ();
 sg13g2_decap_8 FILLER_51_123 ();
 sg13g2_decap_8 FILLER_51_130 ();
 sg13g2_fill_2 FILLER_51_137 ();
 sg13g2_fill_2 FILLER_51_143 ();
 sg13g2_decap_8 FILLER_51_174 ();
 sg13g2_fill_2 FILLER_51_181 ();
 sg13g2_fill_1 FILLER_51_183 ();
 sg13g2_fill_1 FILLER_51_195 ();
 sg13g2_fill_1 FILLER_51_212 ();
 sg13g2_decap_8 FILLER_51_218 ();
 sg13g2_fill_2 FILLER_51_225 ();
 sg13g2_fill_2 FILLER_51_240 ();
 sg13g2_fill_1 FILLER_51_242 ();
 sg13g2_decap_8 FILLER_51_246 ();
 sg13g2_decap_4 FILLER_51_253 ();
 sg13g2_fill_1 FILLER_51_262 ();
 sg13g2_fill_1 FILLER_51_267 ();
 sg13g2_decap_4 FILLER_51_273 ();
 sg13g2_fill_1 FILLER_51_277 ();
 sg13g2_decap_4 FILLER_51_282 ();
 sg13g2_decap_8 FILLER_51_290 ();
 sg13g2_decap_4 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_301 ();
 sg13g2_decap_4 FILLER_51_306 ();
 sg13g2_fill_2 FILLER_51_310 ();
 sg13g2_fill_2 FILLER_51_317 ();
 sg13g2_fill_1 FILLER_51_319 ();
 sg13g2_decap_4 FILLER_51_324 ();
 sg13g2_decap_8 FILLER_51_343 ();
 sg13g2_fill_2 FILLER_51_350 ();
 sg13g2_fill_2 FILLER_51_356 ();
 sg13g2_fill_2 FILLER_51_362 ();
 sg13g2_fill_1 FILLER_51_364 ();
 sg13g2_decap_4 FILLER_51_374 ();
 sg13g2_fill_1 FILLER_51_383 ();
 sg13g2_fill_2 FILLER_51_389 ();
 sg13g2_fill_1 FILLER_51_391 ();
 sg13g2_fill_1 FILLER_51_397 ();
 sg13g2_decap_8 FILLER_51_410 ();
 sg13g2_fill_1 FILLER_51_421 ();
 sg13g2_decap_4 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_52_8 ();
 sg13g2_fill_1 FILLER_52_18 ();
 sg13g2_fill_2 FILLER_52_34 ();
 sg13g2_decap_8 FILLER_52_60 ();
 sg13g2_fill_2 FILLER_52_67 ();
 sg13g2_decap_4 FILLER_52_95 ();
 sg13g2_fill_1 FILLER_52_99 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_fill_1 FILLER_52_133 ();
 sg13g2_fill_1 FILLER_52_152 ();
 sg13g2_fill_1 FILLER_52_161 ();
 sg13g2_fill_1 FILLER_52_167 ();
 sg13g2_fill_1 FILLER_52_176 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_4 FILLER_52_189 ();
 sg13g2_fill_1 FILLER_52_193 ();
 sg13g2_fill_2 FILLER_52_206 ();
 sg13g2_decap_8 FILLER_52_216 ();
 sg13g2_fill_1 FILLER_52_223 ();
 sg13g2_fill_1 FILLER_52_229 ();
 sg13g2_decap_8 FILLER_52_239 ();
 sg13g2_decap_8 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_300 ();
 sg13g2_fill_1 FILLER_52_302 ();
 sg13g2_decap_4 FILLER_52_323 ();
 sg13g2_fill_1 FILLER_52_336 ();
 sg13g2_fill_2 FILLER_52_346 ();
 sg13g2_fill_1 FILLER_52_348 ();
 sg13g2_decap_4 FILLER_52_357 ();
 sg13g2_fill_2 FILLER_52_361 ();
 sg13g2_fill_1 FILLER_52_367 ();
 sg13g2_fill_1 FILLER_52_378 ();
 sg13g2_decap_4 FILLER_52_383 ();
 sg13g2_fill_1 FILLER_52_396 ();
 sg13g2_decap_8 FILLER_52_408 ();
 sg13g2_fill_2 FILLER_52_415 ();
 sg13g2_decap_8 FILLER_52_421 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_2 FILLER_53_34 ();
 sg13g2_fill_1 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_90 ();
 sg13g2_fill_2 FILLER_53_97 ();
 sg13g2_fill_1 FILLER_53_99 ();
 sg13g2_fill_1 FILLER_53_109 ();
 sg13g2_fill_2 FILLER_53_115 ();
 sg13g2_fill_1 FILLER_53_117 ();
 sg13g2_decap_8 FILLER_53_123 ();
 sg13g2_decap_8 FILLER_53_130 ();
 sg13g2_fill_2 FILLER_53_137 ();
 sg13g2_fill_1 FILLER_53_139 ();
 sg13g2_fill_1 FILLER_53_163 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_4 FILLER_53_175 ();
 sg13g2_decap_4 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_4 FILLER_53_238 ();
 sg13g2_fill_2 FILLER_53_242 ();
 sg13g2_fill_1 FILLER_53_248 ();
 sg13g2_decap_4 FILLER_53_262 ();
 sg13g2_decap_4 FILLER_53_288 ();
 sg13g2_fill_2 FILLER_53_292 ();
 sg13g2_fill_1 FILLER_53_314 ();
 sg13g2_decap_8 FILLER_53_319 ();
 sg13g2_decap_4 FILLER_53_335 ();
 sg13g2_fill_2 FILLER_53_339 ();
 sg13g2_decap_8 FILLER_53_346 ();
 sg13g2_decap_8 FILLER_53_353 ();
 sg13g2_fill_2 FILLER_53_360 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_1 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_416 ();
 sg13g2_decap_8 FILLER_53_421 ();
 sg13g2_fill_2 FILLER_53_428 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_decap_8 FILLER_54_7 ();
 sg13g2_decap_4 FILLER_54_14 ();
 sg13g2_fill_1 FILLER_54_18 ();
 sg13g2_fill_1 FILLER_54_31 ();
 sg13g2_fill_1 FILLER_54_37 ();
 sg13g2_fill_1 FILLER_54_41 ();
 sg13g2_fill_2 FILLER_54_55 ();
 sg13g2_fill_1 FILLER_54_62 ();
 sg13g2_decap_8 FILLER_54_70 ();
 sg13g2_decap_4 FILLER_54_77 ();
 sg13g2_fill_2 FILLER_54_81 ();
 sg13g2_decap_8 FILLER_54_92 ();
 sg13g2_fill_1 FILLER_54_99 ();
 sg13g2_fill_2 FILLER_54_134 ();
 sg13g2_decap_8 FILLER_54_156 ();
 sg13g2_decap_8 FILLER_54_163 ();
 sg13g2_fill_2 FILLER_54_170 ();
 sg13g2_fill_1 FILLER_54_172 ();
 sg13g2_fill_2 FILLER_54_178 ();
 sg13g2_decap_8 FILLER_54_212 ();
 sg13g2_decap_8 FILLER_54_219 ();
 sg13g2_decap_4 FILLER_54_226 ();
 sg13g2_fill_1 FILLER_54_230 ();
 sg13g2_fill_1 FILLER_54_235 ();
 sg13g2_fill_2 FILLER_54_244 ();
 sg13g2_fill_1 FILLER_54_246 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_decap_4 FILLER_54_263 ();
 sg13g2_fill_2 FILLER_54_267 ();
 sg13g2_fill_1 FILLER_54_274 ();
 sg13g2_fill_2 FILLER_54_279 ();
 sg13g2_decap_8 FILLER_54_285 ();
 sg13g2_decap_4 FILLER_54_292 ();
 sg13g2_fill_2 FILLER_54_314 ();
 sg13g2_decap_8 FILLER_54_335 ();
 sg13g2_decap_4 FILLER_54_342 ();
 sg13g2_decap_8 FILLER_54_352 ();
 sg13g2_decap_8 FILLER_54_359 ();
 sg13g2_fill_1 FILLER_54_366 ();
 sg13g2_decap_4 FILLER_54_387 ();
 sg13g2_fill_2 FILLER_54_396 ();
 sg13g2_fill_1 FILLER_54_398 ();
 sg13g2_fill_2 FILLER_54_411 ();
 sg13g2_fill_1 FILLER_54_413 ();
 sg13g2_decap_8 FILLER_54_421 ();
 sg13g2_fill_2 FILLER_54_428 ();
 sg13g2_fill_2 FILLER_55_30 ();
 sg13g2_fill_2 FILLER_55_40 ();
 sg13g2_decap_4 FILLER_55_47 ();
 sg13g2_decap_4 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_65 ();
 sg13g2_decap_8 FILLER_55_72 ();
 sg13g2_fill_2 FILLER_55_79 ();
 sg13g2_fill_1 FILLER_55_81 ();
 sg13g2_fill_2 FILLER_55_91 ();
 sg13g2_fill_1 FILLER_55_93 ();
 sg13g2_fill_1 FILLER_55_98 ();
 sg13g2_fill_2 FILLER_55_104 ();
 sg13g2_fill_2 FILLER_55_110 ();
 sg13g2_fill_2 FILLER_55_116 ();
 sg13g2_fill_1 FILLER_55_118 ();
 sg13g2_decap_8 FILLER_55_124 ();
 sg13g2_decap_8 FILLER_55_131 ();
 sg13g2_decap_4 FILLER_55_138 ();
 sg13g2_fill_2 FILLER_55_142 ();
 sg13g2_decap_4 FILLER_55_149 ();
 sg13g2_decap_8 FILLER_55_157 ();
 sg13g2_decap_4 FILLER_55_164 ();
 sg13g2_fill_1 FILLER_55_168 ();
 sg13g2_fill_1 FILLER_55_174 ();
 sg13g2_fill_1 FILLER_55_182 ();
 sg13g2_fill_1 FILLER_55_186 ();
 sg13g2_decap_8 FILLER_55_191 ();
 sg13g2_decap_8 FILLER_55_198 ();
 sg13g2_decap_4 FILLER_55_205 ();
 sg13g2_fill_2 FILLER_55_209 ();
 sg13g2_fill_1 FILLER_55_216 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_decap_4 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_fill_1 FILLER_55_294 ();
 sg13g2_fill_2 FILLER_55_314 ();
 sg13g2_fill_1 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_fill_2 FILLER_55_338 ();
 sg13g2_fill_2 FILLER_55_344 ();
 sg13g2_decap_4 FILLER_55_355 ();
 sg13g2_fill_1 FILLER_55_359 ();
 sg13g2_decap_4 FILLER_55_363 ();
 sg13g2_fill_2 FILLER_55_392 ();
 sg13g2_fill_2 FILLER_55_399 ();
 sg13g2_fill_1 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_411 ();
 sg13g2_decap_8 FILLER_55_417 ();
 sg13g2_decap_4 FILLER_55_424 ();
 sg13g2_fill_2 FILLER_55_428 ();
 sg13g2_decap_8 FILLER_56_0 ();
 sg13g2_decap_8 FILLER_56_7 ();
 sg13g2_decap_8 FILLER_56_14 ();
 sg13g2_decap_8 FILLER_56_21 ();
 sg13g2_decap_8 FILLER_56_28 ();
 sg13g2_decap_4 FILLER_56_35 ();
 sg13g2_decap_4 FILLER_56_53 ();
 sg13g2_fill_1 FILLER_56_62 ();
 sg13g2_fill_1 FILLER_56_68 ();
 sg13g2_fill_2 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_128 ();
 sg13g2_decap_4 FILLER_56_135 ();
 sg13g2_fill_2 FILLER_56_139 ();
 sg13g2_fill_1 FILLER_56_170 ();
 sg13g2_decap_4 FILLER_56_220 ();
 sg13g2_fill_1 FILLER_56_224 ();
 sg13g2_fill_1 FILLER_56_243 ();
 sg13g2_fill_1 FILLER_56_249 ();
 sg13g2_fill_1 FILLER_56_254 ();
 sg13g2_fill_2 FILLER_56_264 ();
 sg13g2_fill_1 FILLER_56_266 ();
 sg13g2_fill_1 FILLER_56_271 ();
 sg13g2_fill_1 FILLER_56_276 ();
 sg13g2_decap_8 FILLER_56_281 ();
 sg13g2_decap_4 FILLER_56_288 ();
 sg13g2_fill_1 FILLER_56_292 ();
 sg13g2_decap_4 FILLER_56_302 ();
 sg13g2_decap_4 FILLER_56_311 ();
 sg13g2_decap_4 FILLER_56_319 ();
 sg13g2_fill_1 FILLER_56_333 ();
 sg13g2_fill_1 FILLER_56_340 ();
 sg13g2_fill_2 FILLER_56_350 ();
 sg13g2_fill_1 FILLER_56_360 ();
 sg13g2_fill_2 FILLER_56_368 ();
 sg13g2_fill_1 FILLER_56_370 ();
 sg13g2_decap_8 FILLER_56_379 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_decap_8 FILLER_56_421 ();
 sg13g2_fill_2 FILLER_56_428 ();
 sg13g2_decap_8 FILLER_57_26 ();
 sg13g2_decap_8 FILLER_57_33 ();
 sg13g2_decap_8 FILLER_57_40 ();
 sg13g2_decap_8 FILLER_57_47 ();
 sg13g2_decap_8 FILLER_57_54 ();
 sg13g2_decap_4 FILLER_57_61 ();
 sg13g2_decap_8 FILLER_57_73 ();
 sg13g2_fill_1 FILLER_57_80 ();
 sg13g2_decap_8 FILLER_57_107 ();
 sg13g2_decap_4 FILLER_57_114 ();
 sg13g2_decap_8 FILLER_57_127 ();
 sg13g2_decap_4 FILLER_57_134 ();
 sg13g2_fill_1 FILLER_57_138 ();
 sg13g2_decap_8 FILLER_57_157 ();
 sg13g2_fill_2 FILLER_57_164 ();
 sg13g2_fill_1 FILLER_57_169 ();
 sg13g2_decap_8 FILLER_57_191 ();
 sg13g2_decap_8 FILLER_57_198 ();
 sg13g2_decap_4 FILLER_57_205 ();
 sg13g2_fill_1 FILLER_57_209 ();
 sg13g2_decap_4 FILLER_57_226 ();
 sg13g2_fill_2 FILLER_57_237 ();
 sg13g2_fill_1 FILLER_57_243 ();
 sg13g2_fill_1 FILLER_57_248 ();
 sg13g2_decap_4 FILLER_57_253 ();
 sg13g2_fill_1 FILLER_57_257 ();
 sg13g2_decap_8 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_268 ();
 sg13g2_fill_2 FILLER_57_277 ();
 sg13g2_fill_2 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_307 ();
 sg13g2_decap_8 FILLER_57_323 ();
 sg13g2_decap_8 FILLER_57_330 ();
 sg13g2_fill_1 FILLER_57_341 ();
 sg13g2_fill_1 FILLER_57_346 ();
 sg13g2_fill_1 FILLER_57_351 ();
 sg13g2_fill_2 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_372 ();
 sg13g2_fill_2 FILLER_57_379 ();
 sg13g2_fill_1 FILLER_57_381 ();
 sg13g2_fill_1 FILLER_57_387 ();
 sg13g2_fill_1 FILLER_57_392 ();
 sg13g2_fill_1 FILLER_57_398 ();
 sg13g2_fill_1 FILLER_57_403 ();
 sg13g2_fill_1 FILLER_57_407 ();
 sg13g2_decap_8 FILLER_57_411 ();
 sg13g2_decap_8 FILLER_57_418 ();
 sg13g2_decap_4 FILLER_57_425 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_fill_2 FILLER_58_7 ();
 sg13g2_fill_1 FILLER_58_9 ();
 sg13g2_fill_1 FILLER_58_17 ();
 sg13g2_fill_1 FILLER_58_23 ();
 sg13g2_fill_1 FILLER_58_33 ();
 sg13g2_fill_2 FILLER_58_46 ();
 sg13g2_decap_8 FILLER_58_74 ();
 sg13g2_decap_8 FILLER_58_81 ();
 sg13g2_decap_8 FILLER_58_88 ();
 sg13g2_decap_4 FILLER_58_95 ();
 sg13g2_decap_8 FILLER_58_107 ();
 sg13g2_fill_2 FILLER_58_114 ();
 sg13g2_fill_1 FILLER_58_116 ();
 sg13g2_fill_2 FILLER_58_122 ();
 sg13g2_fill_2 FILLER_58_128 ();
 sg13g2_fill_1 FILLER_58_130 ();
 sg13g2_fill_1 FILLER_58_162 ();
 sg13g2_decap_4 FILLER_58_168 ();
 sg13g2_fill_2 FILLER_58_196 ();
 sg13g2_fill_2 FILLER_58_204 ();
 sg13g2_fill_1 FILLER_58_206 ();
 sg13g2_decap_8 FILLER_58_221 ();
 sg13g2_fill_2 FILLER_58_228 ();
 sg13g2_decap_4 FILLER_58_247 ();
 sg13g2_fill_1 FILLER_58_251 ();
 sg13g2_fill_1 FILLER_58_259 ();
 sg13g2_fill_2 FILLER_58_265 ();
 sg13g2_fill_1 FILLER_58_267 ();
 sg13g2_fill_1 FILLER_58_296 ();
 sg13g2_fill_2 FILLER_58_301 ();
 sg13g2_fill_1 FILLER_58_303 ();
 sg13g2_fill_2 FILLER_58_320 ();
 sg13g2_fill_1 FILLER_58_322 ();
 sg13g2_fill_2 FILLER_58_328 ();
 sg13g2_fill_1 FILLER_58_330 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_fill_1 FILLER_58_341 ();
 sg13g2_fill_1 FILLER_58_352 ();
 sg13g2_decap_8 FILLER_58_377 ();
 sg13g2_fill_2 FILLER_58_384 ();
 sg13g2_fill_1 FILLER_58_394 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_fill_2 FILLER_58_410 ();
 sg13g2_decap_8 FILLER_58_417 ();
 sg13g2_decap_4 FILLER_58_424 ();
 sg13g2_fill_2 FILLER_58_428 ();
 sg13g2_decap_8 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_7 ();
 sg13g2_fill_1 FILLER_59_17 ();
 sg13g2_decap_4 FILLER_59_23 ();
 sg13g2_fill_2 FILLER_59_68 ();
 sg13g2_decap_8 FILLER_59_75 ();
 sg13g2_decap_8 FILLER_59_82 ();
 sg13g2_decap_8 FILLER_59_89 ();
 sg13g2_decap_4 FILLER_59_106 ();
 sg13g2_fill_1 FILLER_59_110 ();
 sg13g2_fill_1 FILLER_59_116 ();
 sg13g2_decap_8 FILLER_59_148 ();
 sg13g2_decap_4 FILLER_59_155 ();
 sg13g2_fill_1 FILLER_59_159 ();
 sg13g2_fill_1 FILLER_59_174 ();
 sg13g2_fill_2 FILLER_59_188 ();
 sg13g2_fill_2 FILLER_59_199 ();
 sg13g2_decap_8 FILLER_59_210 ();
 sg13g2_decap_8 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_224 ();
 sg13g2_decap_4 FILLER_59_231 ();
 sg13g2_decap_4 FILLER_59_247 ();
 sg13g2_fill_1 FILLER_59_251 ();
 sg13g2_decap_4 FILLER_59_257 ();
 sg13g2_fill_1 FILLER_59_264 ();
 sg13g2_fill_1 FILLER_59_270 ();
 sg13g2_decap_4 FILLER_59_279 ();
 sg13g2_fill_2 FILLER_59_283 ();
 sg13g2_fill_1 FILLER_59_295 ();
 sg13g2_fill_1 FILLER_59_320 ();
 sg13g2_fill_1 FILLER_59_345 ();
 sg13g2_fill_1 FILLER_59_358 ();
 sg13g2_fill_2 FILLER_59_363 ();
 sg13g2_fill_1 FILLER_59_365 ();
 sg13g2_decap_8 FILLER_59_381 ();
 sg13g2_decap_4 FILLER_59_388 ();
 sg13g2_fill_1 FILLER_59_392 ();
 sg13g2_fill_1 FILLER_59_406 ();
 sg13g2_decap_8 FILLER_59_420 ();
 sg13g2_fill_2 FILLER_59_427 ();
 sg13g2_fill_1 FILLER_59_429 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_7 ();
 sg13g2_fill_1 FILLER_60_11 ();
 sg13g2_fill_1 FILLER_60_17 ();
 sg13g2_decap_8 FILLER_60_42 ();
 sg13g2_decap_8 FILLER_60_49 ();
 sg13g2_decap_8 FILLER_60_56 ();
 sg13g2_decap_8 FILLER_60_63 ();
 sg13g2_decap_4 FILLER_60_70 ();
 sg13g2_decap_8 FILLER_60_82 ();
 sg13g2_decap_8 FILLER_60_89 ();
 sg13g2_decap_4 FILLER_60_96 ();
 sg13g2_fill_1 FILLER_60_100 ();
 sg13g2_fill_2 FILLER_60_127 ();
 sg13g2_fill_1 FILLER_60_129 ();
 sg13g2_fill_2 FILLER_60_134 ();
 sg13g2_fill_1 FILLER_60_136 ();
 sg13g2_fill_2 FILLER_60_141 ();
 sg13g2_fill_1 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_150 ();
 sg13g2_fill_2 FILLER_60_161 ();
 sg13g2_fill_1 FILLER_60_163 ();
 sg13g2_decap_8 FILLER_60_168 ();
 sg13g2_fill_2 FILLER_60_175 ();
 sg13g2_fill_1 FILLER_60_177 ();
 sg13g2_fill_2 FILLER_60_191 ();
 sg13g2_fill_2 FILLER_60_198 ();
 sg13g2_decap_8 FILLER_60_210 ();
 sg13g2_decap_8 FILLER_60_217 ();
 sg13g2_decap_8 FILLER_60_224 ();
 sg13g2_fill_2 FILLER_60_231 ();
 sg13g2_fill_2 FILLER_60_239 ();
 sg13g2_fill_1 FILLER_60_241 ();
 sg13g2_fill_2 FILLER_60_247 ();
 sg13g2_fill_1 FILLER_60_249 ();
 sg13g2_decap_4 FILLER_60_266 ();
 sg13g2_fill_2 FILLER_60_270 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_283 ();
 sg13g2_fill_1 FILLER_60_301 ();
 sg13g2_fill_1 FILLER_60_323 ();
 sg13g2_fill_1 FILLER_60_329 ();
 sg13g2_decap_4 FILLER_60_339 ();
 sg13g2_fill_2 FILLER_60_343 ();
 sg13g2_decap_4 FILLER_60_349 ();
 sg13g2_fill_1 FILLER_60_353 ();
 sg13g2_fill_2 FILLER_60_378 ();
 sg13g2_fill_1 FILLER_60_380 ();
 sg13g2_fill_1 FILLER_60_390 ();
 sg13g2_fill_1 FILLER_60_395 ();
 sg13g2_fill_2 FILLER_60_404 ();
 sg13g2_fill_1 FILLER_60_406 ();
 sg13g2_fill_1 FILLER_60_412 ();
 sg13g2_decap_8 FILLER_60_417 ();
 sg13g2_decap_4 FILLER_60_424 ();
 sg13g2_fill_2 FILLER_60_428 ();
 sg13g2_fill_2 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_26 ();
 sg13g2_decap_4 FILLER_61_57 ();
 sg13g2_fill_2 FILLER_61_61 ();
 sg13g2_fill_2 FILLER_61_71 ();
 sg13g2_fill_1 FILLER_61_73 ();
 sg13g2_fill_2 FILLER_61_89 ();
 sg13g2_fill_2 FILLER_61_96 ();
 sg13g2_decap_8 FILLER_61_106 ();
 sg13g2_decap_8 FILLER_61_113 ();
 sg13g2_decap_8 FILLER_61_120 ();
 sg13g2_decap_8 FILLER_61_127 ();
 sg13g2_decap_8 FILLER_61_134 ();
 sg13g2_fill_1 FILLER_61_141 ();
 sg13g2_decap_4 FILLER_61_168 ();
 sg13g2_fill_2 FILLER_61_180 ();
 sg13g2_fill_1 FILLER_61_182 ();
 sg13g2_decap_4 FILLER_61_195 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_decap_4 FILLER_61_214 ();
 sg13g2_fill_2 FILLER_61_218 ();
 sg13g2_decap_8 FILLER_61_246 ();
 sg13g2_fill_2 FILLER_61_253 ();
 sg13g2_decap_8 FILLER_61_269 ();
 sg13g2_decap_4 FILLER_61_276 ();
 sg13g2_fill_1 FILLER_61_280 ();
 sg13g2_fill_1 FILLER_61_285 ();
 sg13g2_decap_8 FILLER_61_301 ();
 sg13g2_decap_8 FILLER_61_308 ();
 sg13g2_fill_2 FILLER_61_315 ();
 sg13g2_fill_2 FILLER_61_321 ();
 sg13g2_fill_1 FILLER_61_323 ();
 sg13g2_decap_4 FILLER_61_330 ();
 sg13g2_fill_1 FILLER_61_334 ();
 sg13g2_decap_4 FILLER_61_340 ();
 sg13g2_fill_1 FILLER_61_344 ();
 sg13g2_decap_8 FILLER_61_352 ();
 sg13g2_decap_4 FILLER_61_363 ();
 sg13g2_fill_1 FILLER_61_367 ();
 sg13g2_fill_2 FILLER_61_378 ();
 sg13g2_decap_4 FILLER_61_388 ();
 sg13g2_fill_1 FILLER_61_395 ();
 sg13g2_decap_8 FILLER_61_416 ();
 sg13g2_decap_8 FILLER_61_423 ();
 sg13g2_decap_4 FILLER_62_0 ();
 sg13g2_fill_1 FILLER_62_4 ();
 sg13g2_fill_1 FILLER_62_18 ();
 sg13g2_fill_1 FILLER_62_27 ();
 sg13g2_fill_2 FILLER_62_32 ();
 sg13g2_fill_1 FILLER_62_34 ();
 sg13g2_decap_8 FILLER_62_38 ();
 sg13g2_fill_1 FILLER_62_45 ();
 sg13g2_fill_1 FILLER_62_59 ();
 sg13g2_decap_4 FILLER_62_65 ();
 sg13g2_fill_1 FILLER_62_77 ();
 sg13g2_fill_2 FILLER_62_93 ();
 sg13g2_decap_8 FILLER_62_108 ();
 sg13g2_decap_8 FILLER_62_115 ();
 sg13g2_decap_8 FILLER_62_122 ();
 sg13g2_decap_8 FILLER_62_129 ();
 sg13g2_decap_4 FILLER_62_136 ();
 sg13g2_fill_1 FILLER_62_140 ();
 sg13g2_fill_1 FILLER_62_146 ();
 sg13g2_fill_1 FILLER_62_151 ();
 sg13g2_decap_8 FILLER_62_155 ();
 sg13g2_decap_8 FILLER_62_162 ();
 sg13g2_fill_2 FILLER_62_177 ();
 sg13g2_decap_8 FILLER_62_187 ();
 sg13g2_fill_2 FILLER_62_205 ();
 sg13g2_decap_4 FILLER_62_217 ();
 sg13g2_fill_2 FILLER_62_221 ();
 sg13g2_fill_1 FILLER_62_241 ();
 sg13g2_decap_8 FILLER_62_247 ();
 sg13g2_decap_4 FILLER_62_254 ();
 sg13g2_decap_8 FILLER_62_262 ();
 sg13g2_decap_4 FILLER_62_269 ();
 sg13g2_decap_8 FILLER_62_278 ();
 sg13g2_fill_2 FILLER_62_285 ();
 sg13g2_fill_1 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_296 ();
 sg13g2_decap_8 FILLER_62_312 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_decap_8 FILLER_62_348 ();
 sg13g2_fill_2 FILLER_62_355 ();
 sg13g2_fill_1 FILLER_62_357 ();
 sg13g2_fill_1 FILLER_62_363 ();
 sg13g2_decap_8 FILLER_62_368 ();
 sg13g2_decap_8 FILLER_62_375 ();
 sg13g2_fill_2 FILLER_62_388 ();
 sg13g2_fill_1 FILLER_62_390 ();
 sg13g2_fill_1 FILLER_62_405 ();
 sg13g2_decap_4 FILLER_62_410 ();
 sg13g2_decap_8 FILLER_62_419 ();
 sg13g2_decap_4 FILLER_62_426 ();
 sg13g2_decap_4 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_4 ();
 sg13g2_decap_8 FILLER_63_24 ();
 sg13g2_decap_8 FILLER_63_31 ();
 sg13g2_decap_4 FILLER_63_38 ();
 sg13g2_fill_2 FILLER_63_52 ();
 sg13g2_fill_1 FILLER_63_54 ();
 sg13g2_decap_8 FILLER_63_65 ();
 sg13g2_fill_1 FILLER_63_72 ();
 sg13g2_fill_1 FILLER_63_78 ();
 sg13g2_fill_1 FILLER_63_87 ();
 sg13g2_decap_8 FILLER_63_92 ();
 sg13g2_fill_1 FILLER_63_99 ();
 sg13g2_decap_8 FILLER_63_113 ();
 sg13g2_decap_4 FILLER_63_120 ();
 sg13g2_fill_2 FILLER_63_124 ();
 sg13g2_decap_4 FILLER_63_164 ();
 sg13g2_fill_1 FILLER_63_198 ();
 sg13g2_fill_2 FILLER_63_207 ();
 sg13g2_fill_1 FILLER_63_209 ();
 sg13g2_fill_2 FILLER_63_218 ();
 sg13g2_fill_1 FILLER_63_220 ();
 sg13g2_decap_4 FILLER_63_251 ();
 sg13g2_fill_1 FILLER_63_255 ();
 sg13g2_decap_8 FILLER_63_275 ();
 sg13g2_decap_4 FILLER_63_282 ();
 sg13g2_decap_4 FILLER_63_290 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_fill_2 FILLER_63_300 ();
 sg13g2_fill_1 FILLER_63_302 ();
 sg13g2_decap_4 FILLER_63_312 ();
 sg13g2_fill_2 FILLER_63_316 ();
 sg13g2_fill_2 FILLER_63_321 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_fill_1 FILLER_63_355 ();
 sg13g2_decap_4 FILLER_63_371 ();
 sg13g2_fill_1 FILLER_63_375 ();
 sg13g2_fill_1 FILLER_63_381 ();
 sg13g2_fill_2 FILLER_63_389 ();
 sg13g2_fill_2 FILLER_63_405 ();
 sg13g2_fill_1 FILLER_63_407 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_fill_2 FILLER_63_427 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_2 ();
 sg13g2_fill_1 FILLER_64_29 ();
 sg13g2_fill_2 FILLER_64_35 ();
 sg13g2_fill_2 FILLER_64_45 ();
 sg13g2_fill_2 FILLER_64_51 ();
 sg13g2_fill_1 FILLER_64_53 ();
 sg13g2_decap_8 FILLER_64_59 ();
 sg13g2_decap_8 FILLER_64_66 ();
 sg13g2_fill_2 FILLER_64_73 ();
 sg13g2_fill_1 FILLER_64_75 ();
 sg13g2_fill_1 FILLER_64_87 ();
 sg13g2_decap_4 FILLER_64_105 ();
 sg13g2_fill_2 FILLER_64_109 ();
 sg13g2_decap_8 FILLER_64_119 ();
 sg13g2_decap_8 FILLER_64_126 ();
 sg13g2_fill_1 FILLER_64_133 ();
 sg13g2_decap_4 FILLER_64_138 ();
 sg13g2_fill_2 FILLER_64_142 ();
 sg13g2_fill_2 FILLER_64_162 ();
 sg13g2_decap_4 FILLER_64_168 ();
 sg13g2_fill_2 FILLER_64_172 ();
 sg13g2_decap_4 FILLER_64_178 ();
 sg13g2_decap_4 FILLER_64_190 ();
 sg13g2_fill_1 FILLER_64_207 ();
 sg13g2_decap_8 FILLER_64_212 ();
 sg13g2_decap_8 FILLER_64_219 ();
 sg13g2_decap_4 FILLER_64_226 ();
 sg13g2_decap_8 FILLER_64_235 ();
 sg13g2_decap_4 FILLER_64_242 ();
 sg13g2_fill_1 FILLER_64_246 ();
 sg13g2_decap_4 FILLER_64_251 ();
 sg13g2_decap_4 FILLER_64_260 ();
 sg13g2_fill_2 FILLER_64_268 ();
 sg13g2_fill_2 FILLER_64_299 ();
 sg13g2_fill_1 FILLER_64_301 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_fill_1 FILLER_64_314 ();
 sg13g2_decap_8 FILLER_64_324 ();
 sg13g2_decap_4 FILLER_64_331 ();
 sg13g2_decap_8 FILLER_64_344 ();
 sg13g2_fill_1 FILLER_64_351 ();
 sg13g2_decap_8 FILLER_64_374 ();
 sg13g2_decap_4 FILLER_64_392 ();
 sg13g2_fill_2 FILLER_64_396 ();
 sg13g2_fill_2 FILLER_64_409 ();
 sg13g2_decap_4 FILLER_64_424 ();
 sg13g2_fill_2 FILLER_64_428 ();
 sg13g2_decap_4 FILLER_65_44 ();
 sg13g2_fill_1 FILLER_65_48 ();
 sg13g2_decap_4 FILLER_65_54 ();
 sg13g2_fill_1 FILLER_65_62 ();
 sg13g2_fill_2 FILLER_65_67 ();
 sg13g2_decap_8 FILLER_65_73 ();
 sg13g2_fill_2 FILLER_65_80 ();
 sg13g2_fill_1 FILLER_65_82 ();
 sg13g2_fill_2 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_101 ();
 sg13g2_fill_2 FILLER_65_108 ();
 sg13g2_fill_2 FILLER_65_113 ();
 sg13g2_fill_1 FILLER_65_115 ();
 sg13g2_decap_8 FILLER_65_124 ();
 sg13g2_decap_8 FILLER_65_131 ();
 sg13g2_decap_4 FILLER_65_138 ();
 sg13g2_decap_4 FILLER_65_155 ();
 sg13g2_fill_1 FILLER_65_185 ();
 sg13g2_decap_8 FILLER_65_198 ();
 sg13g2_decap_8 FILLER_65_205 ();
 sg13g2_decap_4 FILLER_65_212 ();
 sg13g2_decap_8 FILLER_65_221 ();
 sg13g2_fill_1 FILLER_65_228 ();
 sg13g2_decap_8 FILLER_65_234 ();
 sg13g2_decap_8 FILLER_65_241 ();
 sg13g2_decap_8 FILLER_65_248 ();
 sg13g2_fill_2 FILLER_65_255 ();
 sg13g2_fill_2 FILLER_65_277 ();
 sg13g2_fill_2 FILLER_65_283 ();
 sg13g2_decap_8 FILLER_65_303 ();
 sg13g2_fill_2 FILLER_65_310 ();
 sg13g2_decap_8 FILLER_65_317 ();
 sg13g2_decap_8 FILLER_65_324 ();
 sg13g2_decap_4 FILLER_65_331 ();
 sg13g2_fill_1 FILLER_65_352 ();
 sg13g2_fill_1 FILLER_65_366 ();
 sg13g2_fill_2 FILLER_65_382 ();
 sg13g2_decap_4 FILLER_65_424 ();
 sg13g2_fill_2 FILLER_65_428 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_4 FILLER_66_7 ();
 sg13g2_decap_8 FILLER_66_15 ();
 sg13g2_decap_4 FILLER_66_22 ();
 sg13g2_fill_1 FILLER_66_30 ();
 sg13g2_decap_4 FILLER_66_41 ();
 sg13g2_fill_2 FILLER_66_57 ();
 sg13g2_fill_1 FILLER_66_59 ();
 sg13g2_decap_4 FILLER_66_64 ();
 sg13g2_fill_1 FILLER_66_78 ();
 sg13g2_fill_1 FILLER_66_83 ();
 sg13g2_fill_2 FILLER_66_92 ();
 sg13g2_fill_2 FILLER_66_97 ();
 sg13g2_fill_2 FILLER_66_103 ();
 sg13g2_fill_2 FILLER_66_110 ();
 sg13g2_decap_8 FILLER_66_142 ();
 sg13g2_decap_8 FILLER_66_154 ();
 sg13g2_decap_4 FILLER_66_161 ();
 sg13g2_fill_2 FILLER_66_165 ();
 sg13g2_decap_8 FILLER_66_171 ();
 sg13g2_decap_8 FILLER_66_178 ();
 sg13g2_fill_1 FILLER_66_185 ();
 sg13g2_decap_8 FILLER_66_190 ();
 sg13g2_decap_8 FILLER_66_202 ();
 sg13g2_decap_4 FILLER_66_209 ();
 sg13g2_decap_8 FILLER_66_226 ();
 sg13g2_decap_8 FILLER_66_233 ();
 sg13g2_decap_8 FILLER_66_240 ();
 sg13g2_decap_8 FILLER_66_247 ();
 sg13g2_decap_8 FILLER_66_254 ();
 sg13g2_fill_1 FILLER_66_261 ();
 sg13g2_fill_1 FILLER_66_281 ();
 sg13g2_decap_8 FILLER_66_306 ();
 sg13g2_fill_1 FILLER_66_313 ();
 sg13g2_decap_4 FILLER_66_319 ();
 sg13g2_decap_4 FILLER_66_333 ();
 sg13g2_fill_2 FILLER_66_347 ();
 sg13g2_decap_8 FILLER_66_377 ();
 sg13g2_decap_4 FILLER_66_384 ();
 sg13g2_fill_2 FILLER_66_393 ();
 sg13g2_decap_8 FILLER_66_414 ();
 sg13g2_decap_8 FILLER_66_421 ();
 sg13g2_fill_2 FILLER_66_428 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_2 FILLER_67_14 ();
 sg13g2_decap_8 FILLER_67_21 ();
 sg13g2_decap_4 FILLER_67_28 ();
 sg13g2_fill_2 FILLER_67_37 ();
 sg13g2_fill_1 FILLER_67_39 ();
 sg13g2_decap_4 FILLER_67_48 ();
 sg13g2_fill_2 FILLER_67_65 ();
 sg13g2_fill_1 FILLER_67_79 ();
 sg13g2_fill_2 FILLER_67_93 ();
 sg13g2_fill_2 FILLER_67_98 ();
 sg13g2_fill_2 FILLER_67_115 ();
 sg13g2_fill_1 FILLER_67_117 ();
 sg13g2_fill_2 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_137 ();
 sg13g2_fill_2 FILLER_67_144 ();
 sg13g2_fill_1 FILLER_67_177 ();
 sg13g2_fill_2 FILLER_67_202 ();
 sg13g2_decap_4 FILLER_67_207 ();
 sg13g2_fill_2 FILLER_67_211 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_fill_2 FILLER_67_252 ();
 sg13g2_fill_1 FILLER_67_267 ();
 sg13g2_decap_8 FILLER_67_272 ();
 sg13g2_decap_4 FILLER_67_279 ();
 sg13g2_fill_1 FILLER_67_283 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_decap_8 FILLER_67_320 ();
 sg13g2_decap_8 FILLER_67_331 ();
 sg13g2_decap_8 FILLER_67_338 ();
 sg13g2_decap_4 FILLER_67_345 ();
 sg13g2_decap_4 FILLER_67_377 ();
 sg13g2_fill_1 FILLER_67_381 ();
 sg13g2_fill_1 FILLER_67_401 ();
 sg13g2_decap_8 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_67_414 ();
 sg13g2_decap_8 FILLER_67_421 ();
 sg13g2_fill_2 FILLER_67_428 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_11 ();
 sg13g2_decap_4 FILLER_68_18 ();
 sg13g2_fill_1 FILLER_68_22 ();
 sg13g2_fill_2 FILLER_68_27 ();
 sg13g2_decap_4 FILLER_68_45 ();
 sg13g2_fill_2 FILLER_68_66 ();
 sg13g2_fill_1 FILLER_68_68 ();
 sg13g2_decap_4 FILLER_68_77 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_94 ();
 sg13g2_fill_1 FILLER_68_100 ();
 sg13g2_fill_2 FILLER_68_118 ();
 sg13g2_decap_8 FILLER_68_140 ();
 sg13g2_fill_2 FILLER_68_177 ();
 sg13g2_fill_1 FILLER_68_190 ();
 sg13g2_decap_8 FILLER_68_209 ();
 sg13g2_decap_4 FILLER_68_216 ();
 sg13g2_fill_2 FILLER_68_229 ();
 sg13g2_fill_1 FILLER_68_231 ();
 sg13g2_decap_4 FILLER_68_236 ();
 sg13g2_fill_1 FILLER_68_240 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_fill_1 FILLER_68_248 ();
 sg13g2_fill_1 FILLER_68_265 ();
 sg13g2_fill_1 FILLER_68_270 ();
 sg13g2_fill_1 FILLER_68_275 ();
 sg13g2_fill_2 FILLER_68_282 ();
 sg13g2_fill_2 FILLER_68_288 ();
 sg13g2_fill_1 FILLER_68_297 ();
 sg13g2_fill_1 FILLER_68_303 ();
 sg13g2_decap_4 FILLER_68_317 ();
 sg13g2_fill_2 FILLER_68_325 ();
 sg13g2_fill_2 FILLER_68_342 ();
 sg13g2_fill_1 FILLER_68_344 ();
 sg13g2_fill_1 FILLER_68_356 ();
 sg13g2_fill_2 FILLER_68_361 ();
 sg13g2_fill_1 FILLER_68_363 ();
 sg13g2_fill_2 FILLER_68_374 ();
 sg13g2_decap_8 FILLER_68_380 ();
 sg13g2_fill_1 FILLER_68_391 ();
 sg13g2_fill_2 FILLER_68_396 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_4 FILLER_68_424 ();
 sg13g2_fill_2 FILLER_68_428 ();
 sg13g2_fill_2 FILLER_69_30 ();
 sg13g2_fill_1 FILLER_69_40 ();
 sg13g2_decap_8 FILLER_69_57 ();
 sg13g2_fill_1 FILLER_69_82 ();
 sg13g2_fill_1 FILLER_69_88 ();
 sg13g2_decap_8 FILLER_69_141 ();
 sg13g2_decap_4 FILLER_69_148 ();
 sg13g2_decap_4 FILLER_69_156 ();
 sg13g2_decap_4 FILLER_69_164 ();
 sg13g2_fill_2 FILLER_69_173 ();
 sg13g2_fill_1 FILLER_69_175 ();
 sg13g2_decap_4 FILLER_69_187 ();
 sg13g2_fill_1 FILLER_69_191 ();
 sg13g2_fill_1 FILLER_69_213 ();
 sg13g2_decap_8 FILLER_69_217 ();
 sg13g2_decap_8 FILLER_69_224 ();
 sg13g2_decap_8 FILLER_69_231 ();
 sg13g2_decap_8 FILLER_69_238 ();
 sg13g2_decap_8 FILLER_69_245 ();
 sg13g2_decap_8 FILLER_69_252 ();
 sg13g2_fill_1 FILLER_69_300 ();
 sg13g2_fill_2 FILLER_69_309 ();
 sg13g2_fill_1 FILLER_69_316 ();
 sg13g2_fill_1 FILLER_69_321 ();
 sg13g2_fill_2 FILLER_69_339 ();
 sg13g2_fill_1 FILLER_69_341 ();
 sg13g2_decap_8 FILLER_69_353 ();
 sg13g2_fill_2 FILLER_69_360 ();
 sg13g2_fill_1 FILLER_69_368 ();
 sg13g2_decap_4 FILLER_69_373 ();
 sg13g2_decap_8 FILLER_69_385 ();
 sg13g2_fill_2 FILLER_69_397 ();
 sg13g2_fill_1 FILLER_69_399 ();
 sg13g2_decap_8 FILLER_69_405 ();
 sg13g2_decap_8 FILLER_69_412 ();
 sg13g2_decap_8 FILLER_69_419 ();
 sg13g2_decap_4 FILLER_69_426 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_4 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_25 ();
 sg13g2_fill_2 FILLER_70_46 ();
 sg13g2_decap_8 FILLER_70_53 ();
 sg13g2_fill_2 FILLER_70_60 ();
 sg13g2_fill_1 FILLER_70_62 ();
 sg13g2_fill_2 FILLER_70_68 ();
 sg13g2_decap_4 FILLER_70_73 ();
 sg13g2_fill_1 FILLER_70_77 ();
 sg13g2_fill_2 FILLER_70_86 ();
 sg13g2_fill_1 FILLER_70_88 ();
 sg13g2_decap_4 FILLER_70_100 ();
 sg13g2_decap_4 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_fill_2 FILLER_70_189 ();
 sg13g2_fill_1 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_230 ();
 sg13g2_decap_8 FILLER_70_237 ();
 sg13g2_decap_8 FILLER_70_244 ();
 sg13g2_decap_4 FILLER_70_251 ();
 sg13g2_fill_2 FILLER_70_255 ();
 sg13g2_decap_8 FILLER_70_260 ();
 sg13g2_fill_2 FILLER_70_267 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_2 FILLER_70_302 ();
 sg13g2_fill_2 FILLER_70_308 ();
 sg13g2_fill_1 FILLER_70_310 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_4 FILLER_70_329 ();
 sg13g2_fill_1 FILLER_70_333 ();
 sg13g2_fill_2 FILLER_70_337 ();
 sg13g2_fill_1 FILLER_70_344 ();
 sg13g2_fill_2 FILLER_70_357 ();
 sg13g2_fill_1 FILLER_70_359 ();
 sg13g2_decap_4 FILLER_70_373 ();
 sg13g2_fill_1 FILLER_70_377 ();
 sg13g2_decap_8 FILLER_70_383 ();
 sg13g2_decap_8 FILLER_70_390 ();
 sg13g2_decap_4 FILLER_70_397 ();
 sg13g2_decap_8 FILLER_70_417 ();
 sg13g2_decap_4 FILLER_70_424 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_decap_4 FILLER_71_42 ();
 sg13g2_fill_2 FILLER_71_46 ();
 sg13g2_decap_8 FILLER_71_67 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_decap_8 FILLER_71_81 ();
 sg13g2_fill_1 FILLER_71_88 ();
 sg13g2_decap_8 FILLER_71_92 ();
 sg13g2_decap_8 FILLER_71_99 ();
 sg13g2_fill_2 FILLER_71_106 ();
 sg13g2_decap_4 FILLER_71_124 ();
 sg13g2_fill_1 FILLER_71_128 ();
 sg13g2_fill_1 FILLER_71_159 ();
 sg13g2_decap_8 FILLER_71_165 ();
 sg13g2_decap_4 FILLER_71_172 ();
 sg13g2_fill_1 FILLER_71_176 ();
 sg13g2_fill_1 FILLER_71_189 ();
 sg13g2_fill_1 FILLER_71_207 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_decap_8 FILLER_71_238 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_decap_8 FILLER_71_256 ();
 sg13g2_decap_4 FILLER_71_263 ();
 sg13g2_fill_1 FILLER_71_267 ();
 sg13g2_fill_1 FILLER_71_279 ();
 sg13g2_decap_4 FILLER_71_285 ();
 sg13g2_decap_8 FILLER_71_293 ();
 sg13g2_fill_2 FILLER_71_300 ();
 sg13g2_fill_1 FILLER_71_302 ();
 sg13g2_decap_8 FILLER_71_311 ();
 sg13g2_decap_8 FILLER_71_318 ();
 sg13g2_decap_4 FILLER_71_325 ();
 sg13g2_fill_1 FILLER_71_333 ();
 sg13g2_fill_2 FILLER_71_338 ();
 sg13g2_fill_1 FILLER_71_340 ();
 sg13g2_decap_4 FILLER_71_349 ();
 sg13g2_fill_2 FILLER_71_365 ();
 sg13g2_fill_2 FILLER_71_376 ();
 sg13g2_fill_2 FILLER_71_400 ();
 sg13g2_fill_1 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_71_413 ();
 sg13g2_decap_8 FILLER_71_420 ();
 sg13g2_fill_2 FILLER_71_427 ();
 sg13g2_fill_1 FILLER_71_429 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_11 ();
 sg13g2_decap_4 FILLER_72_18 ();
 sg13g2_fill_1 FILLER_72_34 ();
 sg13g2_decap_4 FILLER_72_87 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_decap_4 FILLER_72_102 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_fill_2 FILLER_72_122 ();
 sg13g2_fill_1 FILLER_72_131 ();
 sg13g2_fill_2 FILLER_72_136 ();
 sg13g2_fill_1 FILLER_72_138 ();
 sg13g2_decap_4 FILLER_72_173 ();
 sg13g2_fill_1 FILLER_72_200 ();
 sg13g2_fill_1 FILLER_72_206 ();
 sg13g2_fill_1 FILLER_72_211 ();
 sg13g2_fill_1 FILLER_72_246 ();
 sg13g2_fill_2 FILLER_72_264 ();
 sg13g2_fill_2 FILLER_72_282 ();
 sg13g2_fill_2 FILLER_72_297 ();
 sg13g2_fill_1 FILLER_72_310 ();
 sg13g2_decap_4 FILLER_72_315 ();
 sg13g2_fill_1 FILLER_72_319 ();
 sg13g2_decap_4 FILLER_72_325 ();
 sg13g2_fill_1 FILLER_72_329 ();
 sg13g2_decap_4 FILLER_72_334 ();
 sg13g2_fill_1 FILLER_72_338 ();
 sg13g2_fill_1 FILLER_72_344 ();
 sg13g2_decap_8 FILLER_72_349 ();
 sg13g2_decap_4 FILLER_72_356 ();
 sg13g2_fill_1 FILLER_72_380 ();
 sg13g2_fill_1 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_391 ();
 sg13g2_decap_8 FILLER_72_415 ();
 sg13g2_decap_8 FILLER_72_422 ();
 sg13g2_fill_1 FILLER_72_429 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_fill_2 FILLER_73_7 ();
 sg13g2_fill_1 FILLER_73_9 ();
 sg13g2_fill_1 FILLER_73_47 ();
 sg13g2_fill_1 FILLER_73_70 ();
 sg13g2_fill_1 FILLER_73_97 ();
 sg13g2_fill_1 FILLER_73_124 ();
 sg13g2_decap_8 FILLER_73_129 ();
 sg13g2_fill_1 FILLER_73_136 ();
 sg13g2_decap_4 FILLER_73_145 ();
 sg13g2_fill_1 FILLER_73_149 ();
 sg13g2_decap_8 FILLER_73_158 ();
 sg13g2_decap_8 FILLER_73_165 ();
 sg13g2_decap_4 FILLER_73_172 ();
 sg13g2_fill_1 FILLER_73_176 ();
 sg13g2_fill_1 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_196 ();
 sg13g2_fill_2 FILLER_73_202 ();
 sg13g2_decap_4 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_241 ();
 sg13g2_decap_8 FILLER_73_247 ();
 sg13g2_decap_8 FILLER_73_254 ();
 sg13g2_decap_4 FILLER_73_261 ();
 sg13g2_fill_1 FILLER_73_265 ();
 sg13g2_decap_4 FILLER_73_276 ();
 sg13g2_fill_2 FILLER_73_285 ();
 sg13g2_fill_2 FILLER_73_309 ();
 sg13g2_fill_1 FILLER_73_315 ();
 sg13g2_fill_1 FILLER_73_321 ();
 sg13g2_decap_8 FILLER_73_326 ();
 sg13g2_fill_2 FILLER_73_333 ();
 sg13g2_fill_1 FILLER_73_335 ();
 sg13g2_fill_2 FILLER_73_345 ();
 sg13g2_fill_1 FILLER_73_347 ();
 sg13g2_fill_1 FILLER_73_353 ();
 sg13g2_fill_2 FILLER_73_371 ();
 sg13g2_decap_4 FILLER_73_379 ();
 sg13g2_fill_2 FILLER_73_383 ();
 sg13g2_fill_1 FILLER_73_390 ();
 sg13g2_fill_1 FILLER_73_396 ();
 sg13g2_decap_8 FILLER_73_402 ();
 sg13g2_decap_8 FILLER_73_413 ();
 sg13g2_decap_8 FILLER_73_420 ();
 sg13g2_fill_2 FILLER_73_427 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_fill_2 FILLER_74_0 ();
 sg13g2_fill_1 FILLER_74_32 ();
 sg13g2_fill_2 FILLER_74_67 ();
 sg13g2_decap_4 FILLER_74_73 ();
 sg13g2_fill_1 FILLER_74_77 ();
 sg13g2_decap_8 FILLER_74_82 ();
 sg13g2_fill_1 FILLER_74_89 ();
 sg13g2_decap_4 FILLER_74_94 ();
 sg13g2_decap_4 FILLER_74_103 ();
 sg13g2_decap_8 FILLER_74_111 ();
 sg13g2_fill_2 FILLER_74_118 ();
 sg13g2_fill_1 FILLER_74_120 ();
 sg13g2_decap_8 FILLER_74_124 ();
 sg13g2_decap_8 FILLER_74_131 ();
 sg13g2_fill_2 FILLER_74_138 ();
 sg13g2_fill_1 FILLER_74_140 ();
 sg13g2_decap_8 FILLER_74_145 ();
 sg13g2_decap_8 FILLER_74_152 ();
 sg13g2_decap_8 FILLER_74_159 ();
 sg13g2_decap_8 FILLER_74_166 ();
 sg13g2_fill_2 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_175 ();
 sg13g2_decap_4 FILLER_74_180 ();
 sg13g2_decap_8 FILLER_74_188 ();
 sg13g2_fill_2 FILLER_74_195 ();
 sg13g2_decap_8 FILLER_74_200 ();
 sg13g2_decap_8 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_214 ();
 sg13g2_decap_8 FILLER_74_219 ();
 sg13g2_decap_8 FILLER_74_226 ();
 sg13g2_decap_8 FILLER_74_233 ();
 sg13g2_decap_8 FILLER_74_240 ();
 sg13g2_decap_8 FILLER_74_247 ();
 sg13g2_decap_8 FILLER_74_254 ();
 sg13g2_decap_4 FILLER_74_261 ();
 sg13g2_fill_1 FILLER_74_265 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_1 FILLER_74_276 ();
 sg13g2_decap_4 FILLER_74_292 ();
 sg13g2_fill_1 FILLER_74_296 ();
 sg13g2_decap_4 FILLER_74_311 ();
 sg13g2_decap_4 FILLER_74_319 ();
 sg13g2_decap_4 FILLER_74_329 ();
 sg13g2_fill_1 FILLER_74_333 ();
 sg13g2_decap_8 FILLER_74_347 ();
 sg13g2_decap_4 FILLER_74_358 ();
 sg13g2_fill_2 FILLER_74_367 ();
 sg13g2_fill_1 FILLER_74_369 ();
 sg13g2_fill_2 FILLER_74_378 ();
 sg13g2_fill_1 FILLER_74_380 ();
 sg13g2_fill_2 FILLER_74_386 ();
 sg13g2_fill_1 FILLER_74_388 ();
 sg13g2_fill_2 FILLER_74_398 ();
 sg13g2_decap_8 FILLER_74_404 ();
 sg13g2_decap_8 FILLER_74_411 ();
 sg13g2_decap_8 FILLER_74_418 ();
 sg13g2_decap_4 FILLER_74_425 ();
 sg13g2_fill_1 FILLER_74_429 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_4 FILLER_75_14 ();
 sg13g2_decap_4 FILLER_75_42 ();
 sg13g2_decap_4 FILLER_75_50 ();
 sg13g2_fill_1 FILLER_75_54 ();
 sg13g2_decap_8 FILLER_75_62 ();
 sg13g2_decap_8 FILLER_75_69 ();
 sg13g2_decap_8 FILLER_75_76 ();
 sg13g2_decap_8 FILLER_75_83 ();
 sg13g2_decap_4 FILLER_75_90 ();
 sg13g2_fill_1 FILLER_75_94 ();
 sg13g2_fill_2 FILLER_75_104 ();
 sg13g2_fill_1 FILLER_75_106 ();
 sg13g2_fill_1 FILLER_75_126 ();
 sg13g2_fill_2 FILLER_75_131 ();
 sg13g2_fill_2 FILLER_75_137 ();
 sg13g2_fill_1 FILLER_75_142 ();
 sg13g2_decap_8 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_176 ();
 sg13g2_fill_2 FILLER_75_182 ();
 sg13g2_fill_1 FILLER_75_184 ();
 sg13g2_fill_2 FILLER_75_201 ();
 sg13g2_decap_8 FILLER_75_247 ();
 sg13g2_decap_8 FILLER_75_254 ();
 sg13g2_decap_8 FILLER_75_261 ();
 sg13g2_fill_1 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_285 ();
 sg13g2_decap_8 FILLER_75_299 ();
 sg13g2_decap_8 FILLER_75_306 ();
 sg13g2_decap_4 FILLER_75_313 ();
 sg13g2_fill_1 FILLER_75_317 ();
 sg13g2_decap_8 FILLER_75_327 ();
 sg13g2_fill_2 FILLER_75_334 ();
 sg13g2_decap_4 FILLER_75_348 ();
 sg13g2_decap_4 FILLER_75_380 ();
 sg13g2_fill_1 FILLER_75_392 ();
 sg13g2_fill_2 FILLER_75_398 ();
 sg13g2_decap_8 FILLER_75_408 ();
 sg13g2_decap_8 FILLER_75_415 ();
 sg13g2_decap_8 FILLER_75_422 ();
 sg13g2_fill_1 FILLER_75_429 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_4 FILLER_76_28 ();
 sg13g2_fill_1 FILLER_76_32 ();
 sg13g2_decap_8 FILLER_76_46 ();
 sg13g2_decap_8 FILLER_76_61 ();
 sg13g2_decap_4 FILLER_76_68 ();
 sg13g2_fill_1 FILLER_76_79 ();
 sg13g2_fill_1 FILLER_76_84 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_fill_1 FILLER_76_91 ();
 sg13g2_decap_8 FILLER_76_152 ();
 sg13g2_decap_8 FILLER_76_159 ();
 sg13g2_decap_8 FILLER_76_166 ();
 sg13g2_fill_2 FILLER_76_173 ();
 sg13g2_fill_1 FILLER_76_186 ();
 sg13g2_fill_1 FILLER_76_191 ();
 sg13g2_fill_2 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_221 ();
 sg13g2_fill_2 FILLER_76_228 ();
 sg13g2_decap_8 FILLER_76_245 ();
 sg13g2_decap_8 FILLER_76_252 ();
 sg13g2_decap_8 FILLER_76_259 ();
 sg13g2_fill_1 FILLER_76_278 ();
 sg13g2_decap_4 FILLER_76_283 ();
 sg13g2_fill_2 FILLER_76_307 ();
 sg13g2_fill_1 FILLER_76_309 ();
 sg13g2_fill_2 FILLER_76_320 ();
 sg13g2_fill_2 FILLER_76_326 ();
 sg13g2_fill_1 FILLER_76_328 ();
 sg13g2_fill_2 FILLER_76_333 ();
 sg13g2_fill_1 FILLER_76_335 ();
 sg13g2_fill_1 FILLER_76_358 ();
 sg13g2_fill_2 FILLER_76_364 ();
 sg13g2_fill_1 FILLER_76_371 ();
 sg13g2_fill_2 FILLER_76_383 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_decap_8 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_76_415 ();
 sg13g2_decap_8 FILLER_76_422 ();
 sg13g2_fill_1 FILLER_76_429 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_4 FILLER_77_21 ();
 sg13g2_fill_2 FILLER_77_56 ();
 sg13g2_fill_1 FILLER_77_58 ();
 sg13g2_fill_2 FILLER_77_109 ();
 sg13g2_fill_1 FILLER_77_111 ();
 sg13g2_fill_1 FILLER_77_116 ();
 sg13g2_fill_2 FILLER_77_147 ();
 sg13g2_fill_1 FILLER_77_149 ();
 sg13g2_decap_8 FILLER_77_166 ();
 sg13g2_fill_2 FILLER_77_173 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_fill_2 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_182 ();
 sg13g2_fill_2 FILLER_77_188 ();
 sg13g2_fill_1 FILLER_77_190 ();
 sg13g2_fill_2 FILLER_77_195 ();
 sg13g2_fill_1 FILLER_77_197 ();
 sg13g2_fill_2 FILLER_77_205 ();
 sg13g2_decap_4 FILLER_77_212 ();
 sg13g2_decap_4 FILLER_77_221 ();
 sg13g2_fill_1 FILLER_77_225 ();
 sg13g2_decap_8 FILLER_77_256 ();
 sg13g2_decap_8 FILLER_77_263 ();
 sg13g2_decap_4 FILLER_77_279 ();
 sg13g2_fill_2 FILLER_77_283 ();
 sg13g2_fill_1 FILLER_77_289 ();
 sg13g2_fill_2 FILLER_77_307 ();
 sg13g2_fill_2 FILLER_77_313 ();
 sg13g2_fill_1 FILLER_77_315 ();
 sg13g2_fill_2 FILLER_77_320 ();
 sg13g2_fill_2 FILLER_77_331 ();
 sg13g2_fill_1 FILLER_77_333 ();
 sg13g2_fill_1 FILLER_77_353 ();
 sg13g2_fill_2 FILLER_77_359 ();
 sg13g2_fill_2 FILLER_77_371 ();
 sg13g2_fill_1 FILLER_77_373 ();
 sg13g2_decap_4 FILLER_77_379 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_fill_2 FILLER_77_427 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_4 FILLER_78_28 ();
 sg13g2_fill_2 FILLER_78_89 ();
 sg13g2_fill_1 FILLER_78_91 ();
 sg13g2_fill_1 FILLER_78_104 ();
 sg13g2_fill_1 FILLER_78_110 ();
 sg13g2_fill_1 FILLER_78_136 ();
 sg13g2_fill_1 FILLER_78_153 ();
 sg13g2_fill_2 FILLER_78_180 ();
 sg13g2_fill_2 FILLER_78_186 ();
 sg13g2_decap_4 FILLER_78_192 ();
 sg13g2_fill_2 FILLER_78_196 ();
 sg13g2_decap_8 FILLER_78_202 ();
 sg13g2_fill_1 FILLER_78_209 ();
 sg13g2_fill_1 FILLER_78_236 ();
 sg13g2_fill_1 FILLER_78_241 ();
 sg13g2_fill_2 FILLER_78_268 ();
 sg13g2_fill_2 FILLER_78_274 ();
 sg13g2_fill_2 FILLER_78_283 ();
 sg13g2_fill_2 FILLER_78_308 ();
 sg13g2_fill_1 FILLER_78_323 ();
 sg13g2_fill_1 FILLER_78_329 ();
 sg13g2_fill_1 FILLER_78_334 ();
 sg13g2_fill_1 FILLER_78_339 ();
 sg13g2_fill_2 FILLER_78_344 ();
 sg13g2_fill_2 FILLER_78_350 ();
 sg13g2_fill_1 FILLER_78_362 ();
 sg13g2_fill_2 FILLER_78_367 ();
 sg13g2_fill_1 FILLER_78_378 ();
 sg13g2_decap_8 FILLER_78_393 ();
 sg13g2_decap_8 FILLER_78_400 ();
 sg13g2_decap_8 FILLER_78_407 ();
 sg13g2_decap_8 FILLER_78_414 ();
 sg13g2_decap_8 FILLER_78_421 ();
 sg13g2_fill_2 FILLER_78_428 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_4 FILLER_79_42 ();
 sg13g2_fill_2 FILLER_79_46 ();
 sg13g2_decap_4 FILLER_79_69 ();
 sg13g2_fill_2 FILLER_79_73 ();
 sg13g2_decap_4 FILLER_79_88 ();
 sg13g2_decap_8 FILLER_79_96 ();
 sg13g2_decap_8 FILLER_79_103 ();
 sg13g2_decap_8 FILLER_79_110 ();
 sg13g2_decap_4 FILLER_79_117 ();
 sg13g2_fill_1 FILLER_79_125 ();
 sg13g2_fill_1 FILLER_79_130 ();
 sg13g2_decap_4 FILLER_79_136 ();
 sg13g2_fill_2 FILLER_79_140 ();
 sg13g2_fill_2 FILLER_79_146 ();
 sg13g2_fill_2 FILLER_79_152 ();
 sg13g2_fill_1 FILLER_79_154 ();
 sg13g2_fill_2 FILLER_79_159 ();
 sg13g2_fill_1 FILLER_79_161 ();
 sg13g2_decap_8 FILLER_79_166 ();
 sg13g2_fill_2 FILLER_79_203 ();
 sg13g2_decap_4 FILLER_79_274 ();
 sg13g2_fill_1 FILLER_79_278 ();
 sg13g2_decap_8 FILLER_79_284 ();
 sg13g2_decap_8 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_306 ();
 sg13g2_decap_4 FILLER_79_313 ();
 sg13g2_fill_2 FILLER_79_329 ();
 sg13g2_fill_1 FILLER_79_331 ();
 sg13g2_decap_4 FILLER_79_348 ();
 sg13g2_fill_2 FILLER_79_352 ();
 sg13g2_decap_8 FILLER_79_358 ();
 sg13g2_decap_8 FILLER_79_365 ();
 sg13g2_decap_8 FILLER_79_372 ();
 sg13g2_decap_8 FILLER_79_379 ();
 sg13g2_decap_8 FILLER_79_386 ();
 sg13g2_decap_8 FILLER_79_393 ();
 sg13g2_decap_8 FILLER_79_400 ();
 sg13g2_decap_8 FILLER_79_407 ();
 sg13g2_decap_8 FILLER_79_414 ();
 sg13g2_decap_8 FILLER_79_421 ();
 sg13g2_fill_2 FILLER_79_428 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_fill_2 FILLER_80_70 ();
 sg13g2_fill_1 FILLER_80_72 ();
 sg13g2_fill_2 FILLER_80_81 ();
 sg13g2_fill_1 FILLER_80_83 ();
 sg13g2_fill_2 FILLER_80_116 ();
 sg13g2_fill_2 FILLER_80_122 ();
 sg13g2_fill_2 FILLER_80_128 ();
 sg13g2_decap_4 FILLER_80_134 ();
 sg13g2_fill_1 FILLER_80_138 ();
 sg13g2_fill_1 FILLER_80_143 ();
 sg13g2_fill_2 FILLER_80_156 ();
 sg13g2_fill_1 FILLER_80_162 ();
 sg13g2_decap_4 FILLER_80_167 ();
 sg13g2_fill_2 FILLER_80_183 ();
 sg13g2_decap_4 FILLER_80_189 ();
 sg13g2_fill_2 FILLER_80_231 ();
 sg13g2_fill_1 FILLER_80_233 ();
 sg13g2_fill_1 FILLER_80_238 ();
 sg13g2_fill_1 FILLER_80_247 ();
 sg13g2_decap_4 FILLER_80_252 ();
 sg13g2_fill_2 FILLER_80_260 ();
 sg13g2_fill_1 FILLER_80_262 ();
 sg13g2_decap_8 FILLER_80_267 ();
 sg13g2_decap_8 FILLER_80_274 ();
 sg13g2_decap_8 FILLER_80_281 ();
 sg13g2_decap_8 FILLER_80_288 ();
 sg13g2_decap_8 FILLER_80_295 ();
 sg13g2_decap_8 FILLER_80_302 ();
 sg13g2_decap_8 FILLER_80_309 ();
 sg13g2_decap_8 FILLER_80_316 ();
 sg13g2_decap_8 FILLER_80_323 ();
 sg13g2_decap_8 FILLER_80_330 ();
 sg13g2_decap_8 FILLER_80_337 ();
 sg13g2_decap_8 FILLER_80_344 ();
 sg13g2_decap_8 FILLER_80_351 ();
 sg13g2_decap_4 FILLER_80_358 ();
 sg13g2_fill_1 FILLER_80_362 ();
 sg13g2_decap_8 FILLER_80_367 ();
 sg13g2_decap_8 FILLER_80_374 ();
 sg13g2_decap_8 FILLER_80_381 ();
 sg13g2_decap_8 FILLER_80_388 ();
 sg13g2_decap_8 FILLER_80_395 ();
 sg13g2_decap_8 FILLER_80_402 ();
 sg13g2_decap_8 FILLER_80_409 ();
 sg13g2_decap_8 FILLER_80_416 ();
 sg13g2_decap_8 FILLER_80_423 ();
endmodule
