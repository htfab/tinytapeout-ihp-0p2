module tt_um_rejunity_vga_test01 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire clknet_0_clk;
 wire \center_x[0] ;
 wire \center_x[1] ;
 wire \center_x[2] ;
 wire \center_x[3] ;
 wire \center_x[4] ;
 wire \center_x[5] ;
 wire \center_y[0] ;
 wire \envelopeA[0] ;
 wire \frame_counter[7] ;
 wire \frame_counter[8] ;
 wire \frame_counter[9] ;
 wire frame_counter_frac;
 wire hsync;
 wire \hvsync_gen.hpos[0] ;
 wire \hvsync_gen.hpos[1] ;
 wire \hvsync_gen.hpos[2] ;
 wire \hvsync_gen.hpos[3] ;
 wire \hvsync_gen.hpos[4] ;
 wire \hvsync_gen.hpos[5] ;
 wire \hvsync_gen.hpos[6] ;
 wire \hvsync_gen.hpos[7] ;
 wire \hvsync_gen.hpos[8] ;
 wire \hvsync_gen.hpos[9] ;
 wire \hvsync_gen.vpos[0] ;
 wire \hvsync_gen.vpos[1] ;
 wire \hvsync_gen.vpos[2] ;
 wire \hvsync_gen.vpos[3] ;
 wire \hvsync_gen.vpos[4] ;
 wire \hvsync_gen.vpos[5] ;
 wire \hvsync_gen.vpos[6] ;
 wire \hvsync_gen.vpos[7] ;
 wire \hvsync_gen.vpos[8] ;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire noise;
 wire \noise_counter[0] ;
 wire \noise_counter[1] ;
 wire \noise_counter[2] ;
 wire note;
 wire note2;
 wire \note2_counter[0] ;
 wire \note2_counter[1] ;
 wire \note2_counter[2] ;
 wire \note2_counter[3] ;
 wire \note2_counter[4] ;
 wire \note2_counter[5] ;
 wire \note2_counter[6] ;
 wire \note2_counter[7] ;
 wire \note2_counter[8] ;
 wire \note2_freq[0] ;
 wire \note2_freq[1] ;
 wire \note2_freq[3] ;
 wire \note2_freq[4] ;
 wire \note2_freq[5] ;
 wire \note2_freq[6] ;
 wire \note2_freq[7] ;
 wire \note2_freq[8] ;
 wire \note_counter[0] ;
 wire \note_counter[1] ;
 wire \note_counter[2] ;
 wire \note_counter[3] ;
 wire \note_counter[4] ;
 wire \note_counter[5] ;
 wire \note_counter[6] ;
 wire \note_counter[7] ;
 wire \note_freq[0] ;
 wire \note_freq[1] ;
 wire \note_freq[2] ;
 wire \note_freq[4] ;
 wire \note_freq[5] ;
 wire \note_freq[6] ;
 wire \note_freq[7] ;
 wire \r1[0] ;
 wire \r1[10] ;
 wire \r1[11] ;
 wire \r1[12] ;
 wire \r1[13] ;
 wire \r1[14] ;
 wire \r1[15] ;
 wire \r1[16] ;
 wire \r1[17] ;
 wire \r1[1] ;
 wire \r1[2] ;
 wire \r1[3] ;
 wire \r1[4] ;
 wire \r1[5] ;
 wire \r1[6] ;
 wire \r1[7] ;
 wire \r1[8] ;
 wire \r1[9] ;
 wire \r2[0] ;
 wire \r2[10] ;
 wire \r2[11] ;
 wire \r2[12] ;
 wire \r2[13] ;
 wire \r2[14] ;
 wire \r2[15] ;
 wire \r2[16] ;
 wire \r2[17] ;
 wire \r2[18] ;
 wire \r2[1] ;
 wire \r2[2] ;
 wire \r2[3] ;
 wire \r2[4] ;
 wire \r2[5] ;
 wire \r2[6] ;
 wire \r2[7] ;
 wire \r2[8] ;
 wire \r2[9] ;
 wire \title_r[0] ;
 wire \title_r[10] ;
 wire \title_r[11] ;
 wire \title_r[12] ;
 wire \title_r[13] ;
 wire \title_r[1] ;
 wire \title_r[2] ;
 wire \title_r[3] ;
 wire \title_r[4] ;
 wire \title_r[5] ;
 wire \title_r[6] ;
 wire \title_r[7] ;
 wire \title_r[8] ;
 wire \title_r[9] ;
 wire \title_r_pixels_in_scanline[0] ;
 wire \title_r_pixels_in_scanline[1] ;
 wire \title_r_pixels_in_scanline[2] ;
 wire \title_r_pixels_in_scanline[3] ;
 wire \title_r_pixels_in_scanline[4] ;
 wire \title_r_pixels_in_scanline[5] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_dfrbp_1 \AUDIO_OUT[0]$_SDFF_PN0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net131),
    .D(_00064_),
    .Q_N(_05689_),
    .Q(net8));
 sg13g2_dfrbp_1 \VIDEO_OUT[0]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net132),
    .D(_00065_),
    .Q_N(_05688_),
    .Q(net9));
 sg13g2_dfrbp_1 \VIDEO_OUT[1]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net133),
    .D(_00066_),
    .Q_N(_05687_),
    .Q(net10));
 sg13g2_dfrbp_1 \VIDEO_OUT[2]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net134),
    .D(_00067_),
    .Q_N(_05686_),
    .Q(net11));
 sg13g2_dfrbp_1 \VIDEO_OUT[3]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net135),
    .D(_00068_),
    .Q_N(_05685_),
    .Q(net12));
 sg13g2_dfrbp_1 \VIDEO_OUT[4]$_SDFF_PN0_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net136),
    .D(_00069_),
    .Q_N(_05684_),
    .Q(net13));
 sg13g2_dfrbp_1 \VIDEO_OUT[5]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net137),
    .D(_00070_),
    .Q_N(_05683_),
    .Q(net14));
 sg13g2_dfrbp_1 \VIDEO_OUT[6]$_SDFF_PN0_  (.CLK(clknet_5_31__leaf_clk),
    .RESET_B(net138),
    .D(_00071_),
    .Q_N(_05682_),
    .Q(net15));
 sg13g2_dfrbp_1 \VIDEO_OUT[7]$_SDFF_PN0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net139),
    .D(_00072_),
    .Q_N(_05681_),
    .Q(net16));
 sg13g2_buf_1 _05702_ (.A(\hvsync_gen.vpos[8] ),
    .X(_02389_));
 sg13g2_buf_2 _05703_ (.A(\hvsync_gen.vpos[6] ),
    .X(_02400_));
 sg13g2_buf_2 _05704_ (.A(\hvsync_gen.vpos[7] ),
    .X(_02411_));
 sg13g2_and3_1 _05705_ (.X(_02422_),
    .A(_02389_),
    .B(_02400_),
    .C(_02411_));
 sg13g2_inv_1 _05706_ (.Y(_02433_),
    .A(_02422_));
 sg13g2_buf_2 _05707_ (.A(\hvsync_gen.vpos[4] ),
    .X(_02444_));
 sg13g2_inv_1 _05708_ (.Y(_02455_),
    .A(_02444_));
 sg13g2_buf_1 _05709_ (.A(\hvsync_gen.vpos[3] ),
    .X(_02466_));
 sg13g2_buf_1 _05710_ (.A(\hvsync_gen.vpos[1] ),
    .X(_02477_));
 sg13g2_nand3_1 _05711_ (.B(net129),
    .C(net128),
    .A(_02455_),
    .Y(_02488_));
 sg13g2_buf_2 _05712_ (.A(\hvsync_gen.vpos[0] ),
    .X(_02499_));
 sg13g2_buf_1 _05713_ (.A(\hvsync_gen.vpos[2] ),
    .X(_02510_));
 sg13g2_nand2b_1 _05714_ (.Y(_02521_),
    .B(net127),
    .A_N(_02499_));
 sg13g2_nand2_1 _05715_ (.Y(_02532_),
    .A(net129),
    .B(net127));
 sg13g2_inv_2 _05716_ (.Y(_02543_),
    .A(\hvsync_gen.vpos[9] ));
 sg13g2_buf_2 _05717_ (.A(\hvsync_gen.vpos[5] ),
    .X(_02554_));
 sg13g2_nand4_1 _05718_ (.B(_02532_),
    .C(_02543_),
    .A(_02521_),
    .Y(_02565_),
    .D(_02554_));
 sg13g2_nor3_1 _05719_ (.A(_02433_),
    .B(_02488_),
    .C(_02565_),
    .Y(_00011_));
 sg13g2_buf_1 _05720_ (.A(\hvsync_gen.hpos[7] ),
    .X(_02586_));
 sg13g2_buf_1 _05721_ (.A(\hvsync_gen.hpos[6] ),
    .X(_02597_));
 sg13g2_buf_1 _05722_ (.A(_02597_),
    .X(_02608_));
 sg13g2_nand2_1 _05723_ (.Y(_02619_),
    .A(net126),
    .B(net116));
 sg13g2_inv_1 _05724_ (.Y(_02630_),
    .A(_02619_));
 sg13g2_buf_1 _05725_ (.A(\hvsync_gen.hpos[8] ),
    .X(_02641_));
 sg13g2_buf_1 _05726_ (.A(\hvsync_gen.hpos[9] ),
    .X(_02652_));
 sg13g2_inv_1 _05727_ (.Y(_02663_),
    .A(_02652_));
 sg13g2_nor2_2 _05728_ (.A(net125),
    .B(_02663_),
    .Y(_02674_));
 sg13g2_nand2_1 _05729_ (.Y(_02685_),
    .A(_02652_),
    .B(net125));
 sg13g2_inv_1 _05730_ (.Y(_02696_),
    .A(_02685_));
 sg13g2_a21oi_1 _05731_ (.A1(_02630_),
    .A2(_02674_),
    .Y(_02707_),
    .B1(_02696_));
 sg13g2_buf_1 _05732_ (.A(\hvsync_gen.hpos[4] ),
    .X(_02718_));
 sg13g2_inv_1 _05733_ (.Y(_02729_),
    .A(_02718_));
 sg13g2_buf_2 _05734_ (.A(\hvsync_gen.hpos[5] ),
    .X(_02740_));
 sg13g2_inv_2 _05735_ (.Y(_02751_),
    .A(_02740_));
 sg13g2_nand2_1 _05736_ (.Y(_02762_),
    .A(net115),
    .B(_02751_));
 sg13g2_inv_2 _05737_ (.Y(_02773_),
    .A(net126));
 sg13g2_nor2_1 _05738_ (.A(_02597_),
    .B(_02773_),
    .Y(_02784_));
 sg13g2_nand3_1 _05739_ (.B(_02762_),
    .C(_02784_),
    .A(_02674_),
    .Y(_02795_));
 sg13g2_buf_1 _05740_ (.A(_00017_),
    .X(_02806_));
 sg13g2_inv_1 _05741_ (.Y(_02817_),
    .A(_02806_));
 sg13g2_buf_1 _05742_ (.A(_02718_),
    .X(_02828_));
 sg13g2_buf_1 _05743_ (.A(_02740_),
    .X(_02839_));
 sg13g2_nand3_1 _05744_ (.B(net114),
    .C(_02839_),
    .A(_02630_),
    .Y(_02850_));
 sg13g2_nand2_1 _05745_ (.Y(_02861_),
    .A(_02850_),
    .B(_02674_));
 sg13g2_a22oi_1 _05746_ (.Y(_00010_),
    .B1(_02817_),
    .B2(_02861_),
    .A2(_02795_),
    .A1(_02707_));
 sg13g2_buf_8 _05747_ (.A(rst_n),
    .X(_02882_));
 sg13g2_inv_1 _05748_ (.Y(_02893_),
    .A(net130));
 sg13g2_buf_1 _05749_ (.A(_00033_),
    .X(_02904_));
 sg13g2_inv_1 _05750_ (.Y(_02915_),
    .A(_02904_));
 sg13g2_buf_1 _05751_ (.A(\hvsync_gen.hpos[0] ),
    .X(_02926_));
 sg13g2_buf_1 _05752_ (.A(\hvsync_gen.hpos[1] ),
    .X(_02937_));
 sg13g2_nor2_1 _05753_ (.A(net124),
    .B(net123),
    .Y(_02948_));
 sg13g2_buf_1 _05754_ (.A(\hvsync_gen.hpos[2] ),
    .X(_02959_));
 sg13g2_inv_2 _05755_ (.Y(_02970_),
    .A(net122));
 sg13g2_buf_1 _05756_ (.A(\hvsync_gen.hpos[3] ),
    .X(_02981_));
 sg13g2_inv_1 _05757_ (.Y(_02992_),
    .A(_02981_));
 sg13g2_nand3_1 _05758_ (.B(_02970_),
    .C(_02992_),
    .A(_02948_),
    .Y(_03003_));
 sg13g2_nor2_1 _05759_ (.A(_02652_),
    .B(net125),
    .Y(_03014_));
 sg13g2_inv_1 _05760_ (.Y(_03025_),
    .A(_03014_));
 sg13g2_nor4_1 _05761_ (.A(net126),
    .B(net116),
    .C(_02762_),
    .D(_03025_),
    .Y(_03036_));
 sg13g2_nor2b_1 _05762_ (.A(_03003_),
    .B_N(_03036_),
    .Y(_03047_));
 sg13g2_buf_1 _05763_ (.A(_03047_),
    .X(_03058_));
 sg13g2_inv_1 _05764_ (.Y(_03069_),
    .A(_02389_));
 sg13g2_nand2_1 _05765_ (.Y(_03080_),
    .A(_03069_),
    .B(_02543_));
 sg13g2_nor2_1 _05766_ (.A(net128),
    .B(_02499_),
    .Y(_03091_));
 sg13g2_inv_1 _05767_ (.Y(_03102_),
    .A(_03091_));
 sg13g2_nor3_1 _05768_ (.A(net129),
    .B(net127),
    .C(_03102_),
    .Y(_03113_));
 sg13g2_inv_1 _05769_ (.Y(_03124_),
    .A(_03113_));
 sg13g2_nor3_1 _05770_ (.A(_02400_),
    .B(_02554_),
    .C(_02444_),
    .Y(_03135_));
 sg13g2_inv_1 _05771_ (.Y(_03146_),
    .A(_03135_));
 sg13g2_nor2_1 _05772_ (.A(_02411_),
    .B(_03146_),
    .Y(_03157_));
 sg13g2_inv_1 _05773_ (.Y(_03168_),
    .A(_03157_));
 sg13g2_nor3_2 _05774_ (.A(_03080_),
    .B(_03124_),
    .C(_03168_),
    .Y(_03179_));
 sg13g2_nand2_1 _05775_ (.Y(_03190_),
    .A(_03058_),
    .B(_03179_));
 sg13g2_buf_2 _05776_ (.A(_03190_),
    .X(_03201_));
 sg13g2_buf_8 _05777_ (.A(\center_x[2] ),
    .X(_03212_));
 sg13g2_inv_4 _05778_ (.A(_03212_),
    .Y(_03223_));
 sg13g2_buf_8 _05779_ (.A(\center_x[0] ),
    .X(_03234_));
 sg13g2_buf_1 _05780_ (.A(net121),
    .X(_03245_));
 sg13g2_buf_1 _05781_ (.A(net110),
    .X(_03256_));
 sg13g2_buf_8 _05782_ (.A(\center_x[1] ),
    .X(_03267_));
 sg13g2_buf_8 _05783_ (.A(net120),
    .X(_03278_));
 sg13g2_buf_8 _05784_ (.A(\center_y[0] ),
    .X(_03289_));
 sg13g2_buf_1 _05785_ (.A(_03289_),
    .X(_03300_));
 sg13g2_buf_1 _05786_ (.A(frame_counter_frac),
    .X(_03311_));
 sg13g2_nand4_1 _05787_ (.B(net109),
    .C(net108),
    .A(net98),
    .Y(_03322_),
    .D(_03311_));
 sg13g2_nor2_2 _05788_ (.A(net111),
    .B(_03322_),
    .Y(_03333_));
 sg13g2_inv_1 _05789_ (.Y(_03344_),
    .A(_03333_));
 sg13g2_inv_2 _05790_ (.Y(_03355_),
    .A(_03201_));
 sg13g2_o21ai_1 _05791_ (.B1(_03355_),
    .Y(_03366_),
    .A1(_02904_),
    .A2(_03344_));
 sg13g2_a21oi_1 _05792_ (.A1(_02904_),
    .A2(_03344_),
    .Y(_03377_),
    .B1(_03366_));
 sg13g2_a21oi_1 _05793_ (.A1(_02915_),
    .A2(_03201_),
    .Y(_03388_),
    .B1(_03377_));
 sg13g2_nor2_1 _05794_ (.A(_02893_),
    .B(_03388_),
    .Y(_03399_));
 sg13g2_buf_2 _05795_ (.A(_00029_),
    .X(_03410_));
 sg13g2_inv_4 _05796_ (.A(_03410_),
    .Y(_03421_));
 sg13g2_buf_8 _05797_ (.A(\center_x[3] ),
    .X(_03432_));
 sg13g2_buf_8 _05798_ (.A(net119),
    .X(_03443_));
 sg13g2_nand2_1 _05799_ (.Y(_03454_),
    .A(_03333_),
    .B(net106));
 sg13g2_o21ai_1 _05800_ (.B1(_03355_),
    .Y(_03465_),
    .A1(_03410_),
    .A2(_03454_));
 sg13g2_a21oi_1 _05801_ (.A1(_03410_),
    .A2(_03454_),
    .Y(_03476_),
    .B1(_03465_));
 sg13g2_a21oi_1 _05802_ (.A1(net107),
    .A2(_03201_),
    .Y(_03487_),
    .B1(_03476_));
 sg13g2_nor2_1 _05803_ (.A(_02893_),
    .B(_03487_),
    .Y(_03498_));
 sg13g2_buf_2 _05804_ (.A(_03498_),
    .X(_03509_));
 sg13g2_buf_1 _05805_ (.A(_02893_),
    .X(_03520_));
 sg13g2_buf_8 _05806_ (.A(_00035_),
    .X(_03531_));
 sg13g2_inv_2 _05807_ (.Y(_03542_),
    .A(_03531_));
 sg13g2_buf_1 _05808_ (.A(_03201_),
    .X(_03553_));
 sg13g2_xnor2_1 _05809_ (.Y(_03564_),
    .A(_03531_),
    .B(_03322_));
 sg13g2_nor2_1 _05810_ (.A(_03564_),
    .B(_03201_),
    .Y(_03575_));
 sg13g2_a21oi_2 _05811_ (.B1(_03575_),
    .Y(_03586_),
    .A2(net47),
    .A1(_03542_));
 sg13g2_nor2_1 _05812_ (.A(net105),
    .B(_03586_),
    .Y(_03597_));
 sg13g2_inv_1 _05813_ (.Y(_03608_),
    .A(_03597_));
 sg13g2_o21ai_1 _05814_ (.B1(_03608_),
    .Y(_00006_),
    .A1(_03399_),
    .A2(_03509_));
 sg13g2_buf_8 _05815_ (.A(_00027_),
    .X(_03629_));
 sg13g2_inv_4 _05816_ (.A(_03629_),
    .Y(_03640_));
 sg13g2_buf_8 _05817_ (.A(\center_x[4] ),
    .X(_03651_));
 sg13g2_nand2_1 _05818_ (.Y(_03662_),
    .A(_03651_),
    .B(net119));
 sg13g2_xnor2_1 _05819_ (.Y(_03673_),
    .A(_03629_),
    .B(_03662_));
 sg13g2_buf_8 _05820_ (.A(_03673_),
    .X(_03684_));
 sg13g2_nor2_1 _05821_ (.A(_03640_),
    .B(_03333_),
    .Y(_03695_));
 sg13g2_a21oi_1 _05822_ (.A1(_03333_),
    .A2(net78),
    .Y(_03706_),
    .B1(_03695_));
 sg13g2_nand2_1 _05823_ (.Y(_03717_),
    .A(_03355_),
    .B(_03706_));
 sg13g2_inv_1 _05824_ (.Y(_03728_),
    .A(_03717_));
 sg13g2_a21oi_1 _05825_ (.A1(_03640_),
    .A2(_03201_),
    .Y(_03739_),
    .B1(_03728_));
 sg13g2_nor2_1 _05826_ (.A(_02893_),
    .B(_03739_),
    .Y(_03750_));
 sg13g2_inv_1 _05827_ (.Y(_03761_),
    .A(_03750_));
 sg13g2_nor2_1 _05828_ (.A(_03487_),
    .B(_03761_),
    .Y(_03772_));
 sg13g2_o21ai_1 _05829_ (.B1(_03586_),
    .Y(_00005_),
    .A1(_03399_),
    .A2(_03772_));
 sg13g2_inv_1 _05830_ (.Y(_03793_),
    .A(_03388_));
 sg13g2_inv_1 _05831_ (.Y(_00002_),
    .A(_03509_));
 sg13g2_nor3_1 _05832_ (.A(_03793_),
    .B(_03750_),
    .C(_00002_),
    .Y(_03814_));
 sg13g2_nor2_1 _05833_ (.A(_03608_),
    .B(_03814_),
    .Y(_03825_));
 sg13g2_a21oi_1 _05834_ (.A1(_03586_),
    .A2(_03814_),
    .Y(_00007_),
    .B1(_03825_));
 sg13g2_nor2_1 _05835_ (.A(_03597_),
    .B(_03399_),
    .Y(_03846_));
 sg13g2_nand2_1 _05836_ (.Y(_03857_),
    .A(_03772_),
    .B(_03586_));
 sg13g2_inv_1 _05837_ (.Y(_03868_),
    .A(_03857_));
 sg13g2_nor2_1 _05838_ (.A(_03846_),
    .B(_03868_),
    .Y(_00008_));
 sg13g2_inv_1 _05839_ (.Y(_00009_),
    .A(_00008_));
 sg13g2_buf_1 _05840_ (.A(_00026_),
    .X(_03899_));
 sg13g2_inv_2 _05841_ (.Y(_03910_),
    .A(\center_x[3] ));
 sg13g2_buf_8 _05842_ (.A(_03910_),
    .X(_03921_));
 sg13g2_buf_1 _05843_ (.A(\center_x[5] ),
    .X(_03932_));
 sg13g2_nand2_1 _05844_ (.Y(_03943_),
    .A(_03651_),
    .B(_03932_));
 sg13g2_nor2_1 _05845_ (.A(net104),
    .B(_03943_),
    .Y(_03954_));
 sg13g2_buf_8 _05846_ (.A(_03954_),
    .X(_03965_));
 sg13g2_buf_8 _05847_ (.A(_03965_),
    .X(_03976_));
 sg13g2_nand2_1 _05848_ (.Y(_03987_),
    .A(_03333_),
    .B(_03976_));
 sg13g2_a21oi_1 _05849_ (.A1(_03899_),
    .A2(_03987_),
    .Y(_03998_),
    .B1(_03201_));
 sg13g2_o21ai_1 _05850_ (.B1(_03998_),
    .Y(_04009_),
    .A1(_03899_),
    .A2(_03987_));
 sg13g2_o21ai_1 _05851_ (.B1(_04009_),
    .Y(_04020_),
    .A1(_03899_),
    .A2(_03355_));
 sg13g2_nand2_2 _05852_ (.Y(_04031_),
    .A(_04020_),
    .B(net130));
 sg13g2_nor2_1 _05853_ (.A(_03761_),
    .B(_04031_),
    .Y(_04042_));
 sg13g2_nor2_1 _05854_ (.A(_03761_),
    .B(_03509_),
    .Y(_04053_));
 sg13g2_a22oi_1 _05855_ (.Y(_00000_),
    .B1(_04031_),
    .B2(_04053_),
    .A2(_03509_),
    .A1(_04042_));
 sg13g2_nor2_1 _05856_ (.A(_03509_),
    .B(_04042_),
    .Y(_00001_));
 sg13g2_nand2_1 _05857_ (.Y(_00120_),
    .A(_04042_),
    .B(_03509_));
 sg13g2_nand2b_1 _05858_ (.Y(_00003_),
    .B(_00120_),
    .A_N(_00001_));
 sg13g2_a21oi_1 _05859_ (.A1(_03509_),
    .A2(_04031_),
    .Y(_00004_),
    .B1(_03761_));
 sg13g2_inv_1 _05860_ (.Y(_04114_),
    .A(_00061_));
 sg13g2_nand2_1 _05861_ (.Y(_04125_),
    .A(net124),
    .B(net123));
 sg13g2_nor2_1 _05862_ (.A(_02970_),
    .B(_04125_),
    .Y(_04136_));
 sg13g2_buf_1 _05863_ (.A(_02981_),
    .X(_04147_));
 sg13g2_nand2_1 _05864_ (.Y(_04158_),
    .A(_04136_),
    .B(net103));
 sg13g2_nor2_1 _05865_ (.A(net115),
    .B(_04158_),
    .Y(_04169_));
 sg13g2_nor2_1 _05866_ (.A(net126),
    .B(net116),
    .Y(_04180_));
 sg13g2_nand4_1 _05867_ (.B(_02751_),
    .C(_02696_),
    .A(_04169_),
    .Y(_04191_),
    .D(_04180_));
 sg13g2_nor4_1 _05868_ (.A(_02389_),
    .B(_02543_),
    .C(_02532_),
    .D(_03102_),
    .Y(_04202_));
 sg13g2_a21oi_1 _05869_ (.A1(_04202_),
    .A2(_03157_),
    .Y(_04213_),
    .B1(_02893_));
 sg13g2_nand2b_1 _05870_ (.Y(_04224_),
    .B(_04213_),
    .A_N(_04191_));
 sg13g2_nand2_1 _05871_ (.Y(_04235_),
    .A(_04191_),
    .B(net130));
 sg13g2_buf_1 _05872_ (.A(_04235_),
    .X(_04245_));
 sg13g2_inv_2 _05873_ (.Y(_04256_),
    .A(_04245_));
 sg13g2_nand2_1 _05874_ (.Y(_04266_),
    .A(_04256_),
    .B(_02499_));
 sg13g2_o21ai_1 _05875_ (.B1(_04266_),
    .Y(_00094_),
    .A1(_04114_),
    .A2(_04224_));
 sg13g2_nor2_1 _05876_ (.A(_04213_),
    .B(_04256_),
    .Y(_04286_));
 sg13g2_buf_2 _05877_ (.A(_04286_),
    .X(_04295_));
 sg13g2_nand2_2 _05878_ (.Y(_04305_),
    .A(net128),
    .B(_02499_));
 sg13g2_nor2_1 _05879_ (.A(_04305_),
    .B(_04256_),
    .Y(_04313_));
 sg13g2_a21oi_1 _05880_ (.A1(_04245_),
    .A2(_02499_),
    .Y(_04320_),
    .B1(net128));
 sg13g2_nor3_1 _05881_ (.A(_04295_),
    .B(_04313_),
    .C(_04320_),
    .Y(_00095_));
 sg13g2_inv_1 _05882_ (.Y(_04335_),
    .A(net127));
 sg13g2_xnor2_1 _05883_ (.Y(_04346_),
    .A(_04335_),
    .B(_04305_));
 sg13g2_nand2_1 _05884_ (.Y(_04357_),
    .A(_04256_),
    .B(net127));
 sg13g2_o21ai_1 _05885_ (.B1(_04357_),
    .Y(_00096_),
    .A1(_04346_),
    .A2(_04224_));
 sg13g2_inv_1 _05886_ (.Y(_04374_),
    .A(_02466_));
 sg13g2_buf_1 _05887_ (.A(_04245_),
    .X(_04385_));
 sg13g2_nor2_1 _05888_ (.A(_02532_),
    .B(_04305_),
    .Y(_04395_));
 sg13g2_inv_1 _05889_ (.Y(_04406_),
    .A(_04395_));
 sg13g2_o21ai_1 _05890_ (.B1(_04374_),
    .Y(_04417_),
    .A1(_04335_),
    .A2(_04305_));
 sg13g2_nand4_1 _05891_ (.B(_04213_),
    .C(_04406_),
    .A(net46),
    .Y(_04428_),
    .D(_04417_));
 sg13g2_o21ai_1 _05892_ (.B1(_04428_),
    .Y(_00097_),
    .A1(_04374_),
    .A2(_04385_));
 sg13g2_a21oi_1 _05893_ (.A1(_04245_),
    .A2(_04395_),
    .Y(_04447_),
    .B1(_02444_));
 sg13g2_nor3_1 _05894_ (.A(_02455_),
    .B(_04406_),
    .C(_04256_),
    .Y(_04456_));
 sg13g2_nor3_1 _05895_ (.A(_04295_),
    .B(_04447_),
    .C(_04456_),
    .Y(_00098_));
 sg13g2_nand2_1 _05896_ (.Y(_04472_),
    .A(_02554_),
    .B(_02444_));
 sg13g2_nor3_1 _05897_ (.A(_04406_),
    .B(_04472_),
    .C(_04256_),
    .Y(_04480_));
 sg13g2_nor2_1 _05898_ (.A(_02554_),
    .B(_04456_),
    .Y(_04488_));
 sg13g2_nor3_1 _05899_ (.A(_04295_),
    .B(_04480_),
    .C(_04488_),
    .Y(_00099_));
 sg13g2_inv_1 _05900_ (.Y(_04503_),
    .A(_02400_));
 sg13g2_buf_1 _05901_ (.A(_04503_),
    .X(_04514_));
 sg13g2_nor3_1 _05902_ (.A(net97),
    .B(_02532_),
    .C(_04472_),
    .Y(_04525_));
 sg13g2_and2_1 _05903_ (.A(_04313_),
    .B(_04525_),
    .X(_04536_));
 sg13g2_buf_1 _05904_ (.A(_04536_),
    .X(_04547_));
 sg13g2_nor2_1 _05905_ (.A(_02400_),
    .B(_04480_),
    .Y(_04558_));
 sg13g2_nor3_1 _05906_ (.A(_04295_),
    .B(_04547_),
    .C(_04558_),
    .Y(_00100_));
 sg13g2_nor2_1 _05907_ (.A(_02411_),
    .B(_04547_),
    .Y(_04578_));
 sg13g2_nand2_1 _05908_ (.Y(_04589_),
    .A(_04547_),
    .B(_02411_));
 sg13g2_inv_1 _05909_ (.Y(_04600_),
    .A(_04589_));
 sg13g2_nor3_1 _05910_ (.A(_04295_),
    .B(_04578_),
    .C(_04600_),
    .Y(_00101_));
 sg13g2_nor2_1 _05911_ (.A(_03069_),
    .B(_04589_),
    .Y(_04621_));
 sg13g2_nor2_1 _05912_ (.A(_02389_),
    .B(_04600_),
    .Y(_04632_));
 sg13g2_nor3_1 _05913_ (.A(_04295_),
    .B(_04621_),
    .C(_04632_),
    .Y(_00102_));
 sg13g2_nor4_1 _05914_ (.A(_02543_),
    .B(_04472_),
    .C(_04406_),
    .D(_02433_),
    .Y(_04653_));
 sg13g2_inv_1 _05915_ (.Y(_04664_),
    .A(_04621_));
 sg13g2_a221oi_1 _05916_ (.B2(_02543_),
    .C1(_04295_),
    .B1(_04664_),
    .A1(net46),
    .Y(_00103_),
    .A2(_04653_));
 sg13g2_buf_1 _05917_ (.A(\title_r_pixels_in_scanline[0] ),
    .X(_04684_));
 sg13g2_inv_1 _05918_ (.Y(_04694_),
    .A(_04684_));
 sg13g2_inv_1 _05919_ (.Y(_04705_),
    .A(_02784_));
 sg13g2_inv_1 _05920_ (.Y(_04715_),
    .A(net124));
 sg13g2_nand3_1 _05921_ (.B(_04715_),
    .C(net115),
    .A(_02674_),
    .Y(_04725_));
 sg13g2_nor4_2 _05922_ (.A(net122),
    .B(net123),
    .C(net103),
    .Y(_04736_),
    .D(_02740_));
 sg13g2_inv_1 _05923_ (.Y(_04746_),
    .A(_04736_));
 sg13g2_nor3_1 _05924_ (.A(_04705_),
    .B(_04725_),
    .C(_04746_),
    .Y(_04756_));
 sg13g2_buf_2 _05925_ (.A(_04756_),
    .X(_04767_));
 sg13g2_inv_1 _05926_ (.Y(_04777_),
    .A(_04767_));
 sg13g2_nor2_1 _05927_ (.A(net126),
    .B(net125),
    .Y(_04787_));
 sg13g2_nor2_1 _05928_ (.A(_02806_),
    .B(_04787_),
    .Y(_04797_));
 sg13g2_inv_1 _05929_ (.Y(_04807_),
    .A(_02554_));
 sg13g2_nor2_1 _05930_ (.A(_04807_),
    .B(_02433_),
    .Y(_04816_));
 sg13g2_nor3_1 _05931_ (.A(\hvsync_gen.vpos[9] ),
    .B(_04797_),
    .C(_04816_),
    .Y(_04826_));
 sg13g2_buf_8 _05932_ (.A(_04826_),
    .X(_04836_));
 sg13g2_inv_2 _05933_ (.Y(_04846_),
    .A(_04836_));
 sg13g2_nand3_1 _05934_ (.B(_03135_),
    .C(_03113_),
    .A(_04846_),
    .Y(_04856_));
 sg13g2_inv_1 _05935_ (.Y(_04866_),
    .A(_04856_));
 sg13g2_nor2_1 _05936_ (.A(_02893_),
    .B(_04866_),
    .Y(_04877_));
 sg13g2_inv_1 _05937_ (.Y(_04888_),
    .A(_04877_));
 sg13g2_nor2_2 _05938_ (.A(_04777_),
    .B(_04888_),
    .Y(_04898_));
 sg13g2_buf_2 _05939_ (.A(\title_r[6] ),
    .X(_04909_));
 sg13g2_buf_2 _05940_ (.A(\title_r[5] ),
    .X(_04920_));
 sg13g2_buf_2 _05941_ (.A(\title_r[4] ),
    .X(_04931_));
 sg13g2_nor3_1 _05942_ (.A(_04909_),
    .B(_04920_),
    .C(_04931_),
    .Y(_04942_));
 sg13g2_buf_2 _05943_ (.A(\title_r[8] ),
    .X(_04953_));
 sg13g2_inv_1 _05944_ (.Y(_04964_),
    .A(_04953_));
 sg13g2_buf_1 _05945_ (.A(\title_r[7] ),
    .X(_04975_));
 sg13g2_inv_1 _05946_ (.Y(_04985_),
    .A(_04975_));
 sg13g2_nand3_1 _05947_ (.B(_04964_),
    .C(_04985_),
    .A(_04942_),
    .Y(_04996_));
 sg13g2_buf_2 _05948_ (.A(\title_r[11] ),
    .X(_05007_));
 sg13g2_buf_2 _05949_ (.A(\title_r[10] ),
    .X(_05017_));
 sg13g2_buf_2 _05950_ (.A(\title_r[9] ),
    .X(_05028_));
 sg13g2_nand4_1 _05951_ (.B(_05007_),
    .C(_05017_),
    .A(_04996_),
    .Y(_05038_),
    .D(_05028_));
 sg13g2_buf_1 _05952_ (.A(\title_r[12] ),
    .X(_05049_));
 sg13g2_inv_1 _05953_ (.Y(_05059_),
    .A(_05049_));
 sg13g2_buf_1 _05954_ (.A(\title_r[13] ),
    .X(_05069_));
 sg13g2_a21o_1 _05955_ (.A2(_05059_),
    .A1(_05038_),
    .B1(_05069_),
    .X(_05080_));
 sg13g2_nor2_1 _05956_ (.A(_02619_),
    .B(_04725_),
    .Y(_05090_));
 sg13g2_a21oi_1 _05957_ (.A1(_05090_),
    .A2(_04736_),
    .Y(_05101_),
    .B1(_02707_));
 sg13g2_inv_1 _05958_ (.Y(_05111_),
    .A(_04797_));
 sg13g2_nor2_1 _05959_ (.A(_05111_),
    .B(_04767_),
    .Y(_05122_));
 sg13g2_inv_1 _05960_ (.Y(_05132_),
    .A(_05122_));
 sg13g2_nor2_1 _05961_ (.A(_02696_),
    .B(_05132_),
    .Y(_05142_));
 sg13g2_nand4_1 _05962_ (.B(_05080_),
    .C(_05101_),
    .A(_04877_),
    .Y(_05152_),
    .D(_05142_));
 sg13g2_nand2b_1 _05963_ (.Y(_05162_),
    .B(_05152_),
    .A_N(_04898_));
 sg13g2_buf_1 _05964_ (.A(_04777_),
    .X(_05172_));
 sg13g2_nand3_1 _05965_ (.B(_00063_),
    .C(_05172_),
    .A(_05162_),
    .Y(_05182_));
 sg13g2_o21ai_1 _05966_ (.B1(_05182_),
    .Y(_00183_),
    .A1(_04694_),
    .A2(_05162_));
 sg13g2_buf_1 _05967_ (.A(\title_r_pixels_in_scanline[1] ),
    .X(_05201_));
 sg13g2_a21oi_1 _05968_ (.A1(_05162_),
    .A2(_04684_),
    .Y(_05211_),
    .B1(_05201_));
 sg13g2_nand3_1 _05969_ (.B(_05201_),
    .C(_04684_),
    .A(_05162_),
    .Y(_05221_));
 sg13g2_inv_1 _05970_ (.Y(_05231_),
    .A(_05221_));
 sg13g2_nor3_1 _05971_ (.A(_04898_),
    .B(_05211_),
    .C(_05231_),
    .Y(_00184_));
 sg13g2_inv_1 _05972_ (.Y(_05236_),
    .A(\title_r_pixels_in_scanline[2] ));
 sg13g2_nor2_1 _05973_ (.A(_05236_),
    .B(_05221_),
    .Y(_05237_));
 sg13g2_nor2_1 _05974_ (.A(\title_r_pixels_in_scanline[2] ),
    .B(_05231_),
    .Y(_05238_));
 sg13g2_nor3_1 _05975_ (.A(_04898_),
    .B(_05237_),
    .C(_05238_),
    .Y(_00185_));
 sg13g2_buf_1 _05976_ (.A(\title_r_pixels_in_scanline[3] ),
    .X(_05239_));
 sg13g2_nor2_1 _05977_ (.A(_05239_),
    .B(_05237_),
    .Y(_05240_));
 sg13g2_nand2_1 _05978_ (.Y(_05241_),
    .A(_05237_),
    .B(_05239_));
 sg13g2_inv_1 _05979_ (.Y(_05242_),
    .A(_05241_));
 sg13g2_nor3_1 _05980_ (.A(_04898_),
    .B(_05240_),
    .C(_05242_),
    .Y(_00186_));
 sg13g2_buf_1 _05981_ (.A(\title_r_pixels_in_scanline[4] ),
    .X(_05243_));
 sg13g2_inv_1 _05982_ (.Y(_05244_),
    .A(_05243_));
 sg13g2_nor2_1 _05983_ (.A(_05244_),
    .B(_05241_),
    .Y(_05245_));
 sg13g2_nor2_1 _05984_ (.A(_05243_),
    .B(_05242_),
    .Y(_05246_));
 sg13g2_nor3_1 _05985_ (.A(_04898_),
    .B(_05245_),
    .C(_05246_),
    .Y(_00187_));
 sg13g2_buf_1 _05986_ (.A(\title_r_pixels_in_scanline[5] ),
    .X(_05247_));
 sg13g2_nor2_1 _05987_ (.A(_05247_),
    .B(_05245_),
    .Y(_05248_));
 sg13g2_a21oi_1 _05988_ (.A1(_05245_),
    .A2(_05247_),
    .Y(_05249_),
    .B1(_04898_));
 sg13g2_nor2b_1 _05989_ (.A(_05248_),
    .B_N(_05249_),
    .Y(_00188_));
 sg13g2_nor2b_1 _05990_ (.A(net46),
    .B_N(_00060_),
    .Y(_00084_));
 sg13g2_inv_1 _05991_ (.Y(_05250_),
    .A(_04125_));
 sg13g2_nor3_1 _05992_ (.A(_02948_),
    .B(_05250_),
    .C(net46),
    .Y(_00085_));
 sg13g2_nor2_1 _05993_ (.A(net122),
    .B(_05250_),
    .Y(_05251_));
 sg13g2_nor3_1 _05994_ (.A(_04136_),
    .B(_05251_),
    .C(net46),
    .Y(_00086_));
 sg13g2_buf_1 _05995_ (.A(net105),
    .X(_05252_));
 sg13g2_nor2_1 _05996_ (.A(net103),
    .B(_04136_),
    .Y(_05253_));
 sg13g2_inv_1 _05997_ (.Y(_05254_),
    .A(_04158_));
 sg13g2_nor3_1 _05998_ (.A(_05252_),
    .B(_05253_),
    .C(_05254_),
    .Y(_00087_));
 sg13g2_nor2_1 _05999_ (.A(net114),
    .B(_05254_),
    .Y(_05255_));
 sg13g2_nor3_1 _06000_ (.A(_05252_),
    .B(_04169_),
    .C(_05255_),
    .Y(_00088_));
 sg13g2_nor2_1 _06001_ (.A(_02839_),
    .B(_04169_),
    .Y(_05256_));
 sg13g2_nand2_1 _06002_ (.Y(_05257_),
    .A(_04169_),
    .B(net113));
 sg13g2_inv_1 _06003_ (.Y(_05258_),
    .A(_05257_));
 sg13g2_nor3_1 _06004_ (.A(_05256_),
    .B(_05258_),
    .C(net46),
    .Y(_00089_));
 sg13g2_buf_1 _06005_ (.A(_02608_),
    .X(_05259_));
 sg13g2_nor2_1 _06006_ (.A(net95),
    .B(_05258_),
    .Y(_05260_));
 sg13g2_inv_1 _06007_ (.Y(_05261_),
    .A(net116));
 sg13g2_buf_1 _06008_ (.A(_05261_),
    .X(_05262_));
 sg13g2_nor2_1 _06009_ (.A(net77),
    .B(_05257_),
    .Y(_05263_));
 sg13g2_nor3_1 _06010_ (.A(_05260_),
    .B(_05263_),
    .C(_04385_),
    .Y(_00090_));
 sg13g2_nor2_1 _06011_ (.A(net126),
    .B(_05263_),
    .Y(_05264_));
 sg13g2_nor2_1 _06012_ (.A(_04158_),
    .B(_02850_),
    .Y(_05265_));
 sg13g2_nor3_1 _06013_ (.A(_05264_),
    .B(_05265_),
    .C(net46),
    .Y(_00091_));
 sg13g2_nand2_1 _06014_ (.Y(_05266_),
    .A(_05265_),
    .B(_02641_));
 sg13g2_inv_1 _06015_ (.Y(_05267_),
    .A(_05266_));
 sg13g2_nor2_1 _06016_ (.A(_02641_),
    .B(_05265_),
    .Y(_05268_));
 sg13g2_nor3_1 _06017_ (.A(_05267_),
    .B(_05268_),
    .C(net46),
    .Y(_00092_));
 sg13g2_o21ai_1 _06018_ (.B1(_04256_),
    .Y(_05269_),
    .A1(_02663_),
    .A2(_05266_));
 sg13g2_a21oi_1 _06019_ (.A1(_02663_),
    .A2(_05266_),
    .Y(_00093_),
    .B1(_05269_));
 sg13g2_nand2_1 _06020_ (.Y(_00121_),
    .A(_04053_),
    .B(_04031_));
 sg13g2_inv_1 _06021_ (.Y(_05270_),
    .A(\title_r[0] ));
 sg13g2_nor2_1 _06022_ (.A(_04767_),
    .B(_05142_),
    .Y(_05271_));
 sg13g2_buf_1 _06023_ (.A(_05271_),
    .X(_05272_));
 sg13g2_buf_1 _06024_ (.A(_05272_),
    .X(_05273_));
 sg13g2_buf_1 _06025_ (.A(_04877_),
    .X(_05274_));
 sg13g2_o21ai_1 _06026_ (.B1(net37),
    .Y(_05275_),
    .A1(_00062_),
    .A2(net31));
 sg13g2_a21oi_1 _06027_ (.A1(_05270_),
    .A2(net31),
    .Y(_00169_),
    .B1(_05275_));
 sg13g2_xnor2_1 _06028_ (.Y(_05276_),
    .A(net95),
    .B(_05017_));
 sg13g2_nor2_1 _06029_ (.A(net114),
    .B(_04920_),
    .Y(_05277_));
 sg13g2_nor2_1 _06030_ (.A(net103),
    .B(_04931_),
    .Y(_05278_));
 sg13g2_buf_1 _06031_ (.A(\title_r[2] ),
    .X(_05279_));
 sg13g2_xor2_1 _06032_ (.B(_05279_),
    .A(net123),
    .X(_05280_));
 sg13g2_inv_1 _06033_ (.Y(_05281_),
    .A(_05280_));
 sg13g2_buf_1 _06034_ (.A(\title_r[1] ),
    .X(_05282_));
 sg13g2_xor2_1 _06035_ (.B(_05282_),
    .A(net124),
    .X(_05283_));
 sg13g2_inv_1 _06036_ (.Y(_05284_),
    .A(_05283_));
 sg13g2_nor2_1 _06037_ (.A(_05270_),
    .B(_05284_),
    .Y(_05285_));
 sg13g2_a21oi_1 _06038_ (.A1(net124),
    .A2(_05282_),
    .Y(_05286_),
    .B1(_05285_));
 sg13g2_nor2_1 _06039_ (.A(_05281_),
    .B(_05286_),
    .Y(_05287_));
 sg13g2_inv_1 _06040_ (.Y(_05288_),
    .A(_05287_));
 sg13g2_nand2_1 _06041_ (.Y(_05289_),
    .A(net123),
    .B(_05279_));
 sg13g2_nand2_1 _06042_ (.Y(_05290_),
    .A(_05288_),
    .B(_05289_));
 sg13g2_inv_1 _06043_ (.Y(_05291_),
    .A(_05290_));
 sg13g2_buf_1 _06044_ (.A(\title_r[3] ),
    .X(_05292_));
 sg13g2_nand2_1 _06045_ (.Y(_05293_),
    .A(net122),
    .B(_05292_));
 sg13g2_nor2_1 _06046_ (.A(net122),
    .B(_05292_),
    .Y(_05294_));
 sg13g2_a21oi_1 _06047_ (.A1(_05291_),
    .A2(_05293_),
    .Y(_05295_),
    .B1(_05294_));
 sg13g2_inv_1 _06048_ (.Y(_05296_),
    .A(_05295_));
 sg13g2_nand2_1 _06049_ (.Y(_05297_),
    .A(net103),
    .B(_04931_));
 sg13g2_o21ai_1 _06050_ (.B1(_05297_),
    .Y(_05298_),
    .A1(_05278_),
    .A2(_05296_));
 sg13g2_inv_1 _06051_ (.Y(_05299_),
    .A(_05298_));
 sg13g2_nand2_1 _06052_ (.Y(_05300_),
    .A(_02828_),
    .B(_04920_));
 sg13g2_o21ai_1 _06053_ (.B1(_05300_),
    .Y(_05301_),
    .A1(_05277_),
    .A2(_05299_));
 sg13g2_nor2_1 _06054_ (.A(_02740_),
    .B(_04909_),
    .Y(_05302_));
 sg13g2_nand2_1 _06055_ (.Y(_05303_),
    .A(_02740_),
    .B(_04909_));
 sg13g2_inv_1 _06056_ (.Y(_05304_),
    .A(_05303_));
 sg13g2_nor2_1 _06057_ (.A(_05302_),
    .B(_05304_),
    .Y(_05305_));
 sg13g2_nand2_1 _06058_ (.Y(_05306_),
    .A(_05301_),
    .B(_05305_));
 sg13g2_nor2_1 _06059_ (.A(net116),
    .B(_04985_),
    .Y(_05307_));
 sg13g2_nor2_1 _06060_ (.A(_05307_),
    .B(_05304_),
    .Y(_05308_));
 sg13g2_nor2_1 _06061_ (.A(_04975_),
    .B(_05261_),
    .Y(_05309_));
 sg13g2_a21oi_1 _06062_ (.A1(_05306_),
    .A2(_05308_),
    .Y(_05310_),
    .B1(_05309_));
 sg13g2_xnor2_1 _06063_ (.Y(_05311_),
    .A(net116),
    .B(_04953_));
 sg13g2_inv_1 _06064_ (.Y(_05312_),
    .A(_05311_));
 sg13g2_xnor2_1 _06065_ (.Y(_05313_),
    .A(_05259_),
    .B(_05028_));
 sg13g2_nor2b_1 _06066_ (.A(_05312_),
    .B_N(_05313_),
    .Y(_05314_));
 sg13g2_nor2_1 _06067_ (.A(net116),
    .B(_04964_),
    .Y(_05315_));
 sg13g2_a221oi_1 _06068_ (.B2(_05314_),
    .C1(_05315_),
    .B1(_05310_),
    .A1(net77),
    .Y(_05316_),
    .A2(_05028_));
 sg13g2_xnor2_1 _06069_ (.Y(_05317_),
    .A(_05276_),
    .B(_05316_));
 sg13g2_a21oi_1 _06070_ (.A1(_05317_),
    .A2(net52),
    .Y(_05318_),
    .B1(net31));
 sg13g2_nor2_1 _06071_ (.A(_04975_),
    .B(net97),
    .Y(_05319_));
 sg13g2_nor2_1 _06072_ (.A(_04953_),
    .B(_04503_),
    .Y(_05320_));
 sg13g2_inv_1 _06073_ (.Y(_05321_),
    .A(_05320_));
 sg13g2_nand2_1 _06074_ (.Y(_05322_),
    .A(_04514_),
    .B(_04953_));
 sg13g2_a21oi_1 _06075_ (.A1(_05321_),
    .A2(_05322_),
    .Y(_05323_),
    .B1(_05319_));
 sg13g2_a21oi_1 _06076_ (.A1(_04953_),
    .A2(_05319_),
    .Y(_05324_),
    .B1(_05323_));
 sg13g2_inv_1 _06077_ (.Y(_05325_),
    .A(_05324_));
 sg13g2_nand2_1 _06078_ (.Y(_05326_),
    .A(_04920_),
    .B(_02444_));
 sg13g2_xor2_1 _06079_ (.B(_02554_),
    .A(_04909_),
    .X(_05327_));
 sg13g2_xnor2_1 _06080_ (.Y(_05328_),
    .A(_05326_),
    .B(_05327_));
 sg13g2_inv_1 _06081_ (.Y(_05329_),
    .A(_05328_));
 sg13g2_nand2_1 _06082_ (.Y(_05330_),
    .A(_04931_),
    .B(net129));
 sg13g2_xor2_1 _06083_ (.B(_02444_),
    .A(_04920_),
    .X(_05331_));
 sg13g2_nor2b_1 _06084_ (.A(_05330_),
    .B_N(_05331_),
    .Y(_05332_));
 sg13g2_xnor2_1 _06085_ (.Y(_05333_),
    .A(_05330_),
    .B(_05331_));
 sg13g2_inv_1 _06086_ (.Y(_05334_),
    .A(_05333_));
 sg13g2_nand2_1 _06087_ (.Y(_05335_),
    .A(_05292_),
    .B(_02510_));
 sg13g2_xor2_1 _06088_ (.B(net129),
    .A(_04931_),
    .X(_05336_));
 sg13g2_nor2b_1 _06089_ (.A(_05335_),
    .B_N(_05336_),
    .Y(_05337_));
 sg13g2_xnor2_1 _06090_ (.Y(_05338_),
    .A(_05335_),
    .B(_05336_));
 sg13g2_inv_1 _06091_ (.Y(_05339_),
    .A(_05338_));
 sg13g2_nand2_1 _06092_ (.Y(_05340_),
    .A(_05279_),
    .B(net128));
 sg13g2_xor2_1 _06093_ (.B(_02510_),
    .A(_05292_),
    .X(_05341_));
 sg13g2_nor2b_1 _06094_ (.A(_05340_),
    .B_N(_05341_),
    .Y(_05342_));
 sg13g2_xnor2_1 _06095_ (.Y(_05343_),
    .A(_05340_),
    .B(_05341_));
 sg13g2_inv_1 _06096_ (.Y(_05344_),
    .A(_05343_));
 sg13g2_xor2_1 _06097_ (.B(_02499_),
    .A(_05282_),
    .X(_05345_));
 sg13g2_inv_1 _06098_ (.Y(_05346_),
    .A(_05345_));
 sg13g2_nand2_1 _06099_ (.Y(_05347_),
    .A(_05282_),
    .B(_02499_));
 sg13g2_o21ai_1 _06100_ (.B1(_05347_),
    .Y(_05348_),
    .A1(_05270_),
    .A2(_05346_));
 sg13g2_xor2_1 _06101_ (.B(net128),
    .A(_05279_),
    .X(_05349_));
 sg13g2_nand2_1 _06102_ (.Y(_05350_),
    .A(_05348_),
    .B(_05349_));
 sg13g2_nor2_1 _06103_ (.A(_05344_),
    .B(_05350_),
    .Y(_05351_));
 sg13g2_nor2_1 _06104_ (.A(_05342_),
    .B(_05351_),
    .Y(_05352_));
 sg13g2_nor2_1 _06105_ (.A(_05339_),
    .B(_05352_),
    .Y(_05353_));
 sg13g2_nor2_1 _06106_ (.A(_05337_),
    .B(_05353_),
    .Y(_05354_));
 sg13g2_nor2_1 _06107_ (.A(_05334_),
    .B(_05354_),
    .Y(_05355_));
 sg13g2_nor2_1 _06108_ (.A(_05332_),
    .B(_05355_),
    .Y(_05356_));
 sg13g2_nand2_1 _06109_ (.Y(_05357_),
    .A(_04909_),
    .B(_02554_));
 sg13g2_xnor2_1 _06110_ (.Y(_05358_),
    .A(_04975_),
    .B(_02400_));
 sg13g2_nor2_1 _06111_ (.A(_05357_),
    .B(_05358_),
    .Y(_05359_));
 sg13g2_nor2b_1 _06112_ (.A(_05326_),
    .B_N(_05327_),
    .Y(_05360_));
 sg13g2_nor2_1 _06113_ (.A(_05359_),
    .B(_05360_),
    .Y(_05361_));
 sg13g2_o21ai_1 _06114_ (.B1(_05361_),
    .Y(_05362_),
    .A1(_05329_),
    .A2(_05356_));
 sg13g2_nand2_1 _06115_ (.Y(_05363_),
    .A(_05358_),
    .B(_05357_));
 sg13g2_nand2_1 _06116_ (.Y(_05364_),
    .A(_05362_),
    .B(_05363_));
 sg13g2_nor2_1 _06117_ (.A(_05325_),
    .B(_05364_),
    .Y(_05365_));
 sg13g2_nor2_1 _06118_ (.A(_05028_),
    .B(net97),
    .Y(_05366_));
 sg13g2_inv_1 _06119_ (.Y(_05367_),
    .A(_05366_));
 sg13g2_nand2_1 _06120_ (.Y(_05368_),
    .A(net97),
    .B(_05028_));
 sg13g2_a21oi_1 _06121_ (.A1(_05367_),
    .A2(_05368_),
    .Y(_05369_),
    .B1(_05320_));
 sg13g2_a21oi_2 _06122_ (.B1(_05369_),
    .Y(_05370_),
    .A2(_05320_),
    .A1(_05028_));
 sg13g2_nand2_1 _06123_ (.Y(_05371_),
    .A(_05365_),
    .B(_05370_));
 sg13g2_a21oi_1 _06124_ (.A1(_05370_),
    .A2(_05323_),
    .Y(_05372_),
    .B1(_05369_));
 sg13g2_nor2_1 _06125_ (.A(_05017_),
    .B(net97),
    .Y(_05373_));
 sg13g2_inv_1 _06126_ (.Y(_05374_),
    .A(_05373_));
 sg13g2_nand2_1 _06127_ (.Y(_05375_),
    .A(net97),
    .B(_05017_));
 sg13g2_a21oi_1 _06128_ (.A1(_05374_),
    .A2(_05375_),
    .Y(_05376_),
    .B1(_05366_));
 sg13g2_a21oi_1 _06129_ (.A1(_05017_),
    .A2(_05366_),
    .Y(_05377_),
    .B1(_05376_));
 sg13g2_inv_1 _06130_ (.Y(_05378_),
    .A(_05377_));
 sg13g2_a21o_1 _06131_ (.A2(_05372_),
    .A1(_05371_),
    .B1(_05378_),
    .X(_05379_));
 sg13g2_buf_1 _06132_ (.A(_04767_),
    .X(_05380_));
 sg13g2_nand3_1 _06133_ (.B(_05372_),
    .C(_05378_),
    .A(_05371_),
    .Y(_05381_));
 sg13g2_nand3_1 _06134_ (.B(net58),
    .C(_05381_),
    .A(_05379_),
    .Y(_05382_));
 sg13g2_inv_1 _06135_ (.Y(_05383_),
    .A(_05272_));
 sg13g2_buf_1 _06136_ (.A(_05383_),
    .X(_05384_));
 sg13g2_o21ai_1 _06137_ (.B1(net37),
    .Y(_05385_),
    .A1(_05017_),
    .A2(net28));
 sg13g2_a21oi_1 _06138_ (.A1(_05318_),
    .A2(_05382_),
    .Y(_00170_),
    .B1(_05385_));
 sg13g2_inv_1 _06139_ (.Y(_05386_),
    .A(_05007_));
 sg13g2_xnor2_1 _06140_ (.Y(_05387_),
    .A(net95),
    .B(_05007_));
 sg13g2_inv_1 _06141_ (.Y(_05388_),
    .A(_05276_));
 sg13g2_inv_1 _06142_ (.Y(_05389_),
    .A(_05302_));
 sg13g2_a21oi_1 _06143_ (.A1(_05301_),
    .A2(_05389_),
    .Y(_05390_),
    .B1(_05304_));
 sg13g2_inv_1 _06144_ (.Y(_05391_),
    .A(_05390_));
 sg13g2_nor2_1 _06145_ (.A(_05309_),
    .B(_05307_),
    .Y(_05392_));
 sg13g2_nand2_1 _06146_ (.Y(_05393_),
    .A(_05391_),
    .B(_05392_));
 sg13g2_nor2_1 _06147_ (.A(_05315_),
    .B(_05307_),
    .Y(_05394_));
 sg13g2_o21ai_1 _06148_ (.B1(_05394_),
    .Y(_05395_),
    .A1(_05312_),
    .A2(_05393_));
 sg13g2_nand2_1 _06149_ (.Y(_05396_),
    .A(_05395_),
    .B(_05313_));
 sg13g2_o21ai_1 _06150_ (.B1(net77),
    .Y(_05397_),
    .A1(_05017_),
    .A2(_05028_));
 sg13g2_o21ai_1 _06151_ (.B1(_05397_),
    .Y(_05398_),
    .A1(_05388_),
    .A2(_05396_));
 sg13g2_nor2_1 _06152_ (.A(_05387_),
    .B(_05398_),
    .Y(_05399_));
 sg13g2_nand2_1 _06153_ (.Y(_05400_),
    .A(_05398_),
    .B(_05387_));
 sg13g2_nand3b_1 _06154_ (.B(net52),
    .C(_05400_),
    .Y(_05401_),
    .A_N(_05399_));
 sg13g2_nor2_1 _06155_ (.A(_05386_),
    .B(_05374_),
    .Y(_05402_));
 sg13g2_xnor2_1 _06156_ (.Y(_05403_),
    .A(_05007_),
    .B(_02400_));
 sg13g2_nor2_1 _06157_ (.A(_05373_),
    .B(_05403_),
    .Y(_05404_));
 sg13g2_nor2_1 _06158_ (.A(_05402_),
    .B(_05404_),
    .Y(_05405_));
 sg13g2_inv_1 _06159_ (.Y(_05406_),
    .A(_05355_));
 sg13g2_a21oi_1 _06160_ (.A1(_05332_),
    .A2(_05327_),
    .Y(_05407_),
    .B1(_05360_));
 sg13g2_o21ai_1 _06161_ (.B1(_05407_),
    .Y(_05408_),
    .A1(_05329_),
    .A2(_05406_));
 sg13g2_inv_1 _06162_ (.Y(_05409_),
    .A(_05359_));
 sg13g2_nand2_1 _06163_ (.Y(_05410_),
    .A(_05409_),
    .B(_05363_));
 sg13g2_nor2_1 _06164_ (.A(_05410_),
    .B(_05325_),
    .Y(_05411_));
 sg13g2_a221oi_1 _06165_ (.B2(_05411_),
    .C1(_05323_),
    .B1(_05408_),
    .A1(_05324_),
    .Y(_05412_),
    .A2(_05359_));
 sg13g2_inv_1 _06166_ (.Y(_05413_),
    .A(_05412_));
 sg13g2_nand3_1 _06167_ (.B(_05370_),
    .C(_05377_),
    .A(_05413_),
    .Y(_05414_));
 sg13g2_a21oi_1 _06168_ (.A1(_05377_),
    .A2(_05369_),
    .Y(_05415_),
    .B1(_05376_));
 sg13g2_nand2_1 _06169_ (.Y(_05416_),
    .A(_05414_),
    .B(_05415_));
 sg13g2_nor2_1 _06170_ (.A(_05405_),
    .B(_05416_),
    .Y(_05417_));
 sg13g2_nor2_1 _06171_ (.A(_04777_),
    .B(_05417_),
    .Y(_05418_));
 sg13g2_nand2_1 _06172_ (.Y(_05419_),
    .A(_05416_),
    .B(_05405_));
 sg13g2_a21oi_1 _06173_ (.A1(_05418_),
    .A2(_05419_),
    .Y(_05420_),
    .B1(_05272_));
 sg13g2_a221oi_1 _06174_ (.B2(_05420_),
    .C1(_04888_),
    .B1(_05401_),
    .A1(_05386_),
    .Y(_00171_),
    .A2(net31));
 sg13g2_xnor2_1 _06175_ (.Y(_05421_),
    .A(net95),
    .B(_05049_));
 sg13g2_inv_1 _06176_ (.Y(_05422_),
    .A(_05421_));
 sg13g2_nand2_1 _06177_ (.Y(_05423_),
    .A(_05276_),
    .B(_05387_));
 sg13g2_o21ai_1 _06178_ (.B1(net77),
    .Y(_05424_),
    .A1(_05007_),
    .A2(_05017_));
 sg13g2_o21ai_1 _06179_ (.B1(_05424_),
    .Y(_05425_),
    .A1(_05423_),
    .A2(_05316_));
 sg13g2_xnor2_1 _06180_ (.Y(_05426_),
    .A(_05422_),
    .B(_05425_));
 sg13g2_a21oi_1 _06181_ (.A1(_05405_),
    .A2(_05376_),
    .Y(_05427_),
    .B1(_05404_));
 sg13g2_o21ai_1 _06182_ (.B1(_05427_),
    .Y(_05428_),
    .A1(_05402_),
    .A2(_05379_));
 sg13g2_nand2_1 _06183_ (.Y(_05429_),
    .A(_05049_),
    .B(_02400_));
 sg13g2_nor2_1 _06184_ (.A(_05007_),
    .B(_05429_),
    .Y(_05430_));
 sg13g2_a21oi_1 _06185_ (.A1(_05059_),
    .A2(_05007_),
    .Y(_05431_),
    .B1(net97));
 sg13g2_a21oi_1 _06186_ (.A1(_05059_),
    .A2(net97),
    .Y(_05432_),
    .B1(_05431_));
 sg13g2_nor2_1 _06187_ (.A(_05430_),
    .B(_05432_),
    .Y(_05433_));
 sg13g2_o21ai_1 _06188_ (.B1(_04767_),
    .Y(_05434_),
    .A1(_05433_),
    .A2(_05428_));
 sg13g2_a21oi_1 _06189_ (.A1(_05428_),
    .A2(_05433_),
    .Y(_05435_),
    .B1(_05434_));
 sg13g2_a21oi_1 _06190_ (.A1(_05426_),
    .A2(net52),
    .Y(_05436_),
    .B1(_05435_));
 sg13g2_o21ai_1 _06191_ (.B1(net37),
    .Y(_05437_),
    .A1(_05049_),
    .A2(net28));
 sg13g2_a21oi_1 _06192_ (.A1(_05436_),
    .A2(net28),
    .Y(_00172_),
    .B1(_05437_));
 sg13g2_nor2_1 _06193_ (.A(_05284_),
    .B(_04767_),
    .Y(_05438_));
 sg13g2_a21oi_1 _06194_ (.A1(net58),
    .A2(_05345_),
    .Y(_05439_),
    .B1(_05438_));
 sg13g2_xnor2_1 _06195_ (.Y(_05440_),
    .A(_00062_),
    .B(_05439_));
 sg13g2_o21ai_1 _06196_ (.B1(net37),
    .Y(_05441_),
    .A1(_05282_),
    .A2(net28));
 sg13g2_a21oi_1 _06197_ (.A1(_05440_),
    .A2(net28),
    .Y(_00174_),
    .B1(_05441_));
 sg13g2_nor2_1 _06198_ (.A(_05349_),
    .B(_05348_),
    .Y(_05442_));
 sg13g2_nor2_1 _06199_ (.A(_05442_),
    .B(net52),
    .Y(_05443_));
 sg13g2_a21oi_1 _06200_ (.A1(_05286_),
    .A2(_05281_),
    .Y(_05444_),
    .B1(net58));
 sg13g2_a22oi_1 _06201_ (.Y(_05445_),
    .B1(_05288_),
    .B2(_05444_),
    .A2(_05350_),
    .A1(_05443_));
 sg13g2_o21ai_1 _06202_ (.B1(net37),
    .Y(_05446_),
    .A1(_05279_),
    .A2(net28));
 sg13g2_a21oi_1 _06203_ (.A1(net28),
    .A2(_05445_),
    .Y(_00175_),
    .B1(_05446_));
 sg13g2_inv_1 _06204_ (.Y(_05447_),
    .A(_05292_));
 sg13g2_xnor2_1 _06205_ (.Y(_05448_),
    .A(_05344_),
    .B(_05350_));
 sg13g2_nor2b_1 _06206_ (.A(_05294_),
    .B_N(_05293_),
    .Y(_05449_));
 sg13g2_xnor2_1 _06207_ (.Y(_05450_),
    .A(_05449_),
    .B(_05290_));
 sg13g2_a21o_1 _06208_ (.A2(_05142_),
    .A1(_05450_),
    .B1(_04888_),
    .X(_05451_));
 sg13g2_a221oi_1 _06209_ (.B2(_05448_),
    .C1(_05451_),
    .B1(net58),
    .A1(_05447_),
    .Y(_00176_),
    .A2(net31));
 sg13g2_nor2b_1 _06210_ (.A(_05278_),
    .B_N(_05297_),
    .Y(_05452_));
 sg13g2_xor2_1 _06211_ (.B(_05295_),
    .A(_05452_),
    .X(_05453_));
 sg13g2_a21oi_1 _06212_ (.A1(_05453_),
    .A2(_05172_),
    .Y(_05454_),
    .B1(_05273_));
 sg13g2_nand2_1 _06213_ (.Y(_05455_),
    .A(_05352_),
    .B(_05339_));
 sg13g2_nand3b_1 _06214_ (.B(net58),
    .C(_05455_),
    .Y(_05456_),
    .A_N(_05353_));
 sg13g2_o21ai_1 _06215_ (.B1(net37),
    .Y(_05457_),
    .A1(_04931_),
    .A2(_05384_));
 sg13g2_a21oi_1 _06216_ (.A1(_05454_),
    .A2(_05456_),
    .Y(_00177_),
    .B1(_05457_));
 sg13g2_nor2b_1 _06217_ (.A(_05277_),
    .B_N(_05300_),
    .Y(_05458_));
 sg13g2_xor2_1 _06218_ (.B(_05298_),
    .A(_05458_),
    .X(_05459_));
 sg13g2_a21oi_1 _06219_ (.A1(_05459_),
    .A2(net52),
    .Y(_05460_),
    .B1(net31));
 sg13g2_nand2_1 _06220_ (.Y(_05461_),
    .A(_05354_),
    .B(_05334_));
 sg13g2_nand3_1 _06221_ (.B(net58),
    .C(_05461_),
    .A(_05406_),
    .Y(_05462_));
 sg13g2_o21ai_1 _06222_ (.B1(_05274_),
    .Y(_05463_),
    .A1(_04920_),
    .A2(_05383_));
 sg13g2_a21oi_1 _06223_ (.A1(_05460_),
    .A2(_05462_),
    .Y(_00178_),
    .B1(_05463_));
 sg13g2_xnor2_1 _06224_ (.Y(_05464_),
    .A(_05329_),
    .B(_05356_));
 sg13g2_xnor2_1 _06225_ (.Y(_05465_),
    .A(_05305_),
    .B(_05301_));
 sg13g2_o21ai_1 _06226_ (.B1(net37),
    .Y(_05466_),
    .A1(_04909_),
    .A2(_05383_));
 sg13g2_a221oi_1 _06227_ (.B2(_05142_),
    .C1(_05466_),
    .B1(_05465_),
    .A1(_05380_),
    .Y(_00179_),
    .A2(_05464_));
 sg13g2_nand2b_1 _06228_ (.Y(_05467_),
    .B(_05390_),
    .A_N(_05392_));
 sg13g2_nand3_1 _06229_ (.B(net52),
    .C(_05467_),
    .A(_05393_),
    .Y(_05468_));
 sg13g2_xnor2_1 _06230_ (.Y(_05469_),
    .A(_05410_),
    .B(_05408_));
 sg13g2_a21oi_1 _06231_ (.A1(_05469_),
    .A2(_05380_),
    .Y(_05470_),
    .B1(_05272_));
 sg13g2_a221oi_1 _06232_ (.B2(_05470_),
    .C1(_04888_),
    .B1(_05468_),
    .A1(_04985_),
    .Y(_00180_),
    .A2(_05273_));
 sg13g2_inv_1 _06233_ (.Y(_05471_),
    .A(_05365_));
 sg13g2_a21oi_1 _06234_ (.A1(_05364_),
    .A2(_05325_),
    .Y(_05472_),
    .B1(_04777_));
 sg13g2_xnor2_1 _06235_ (.Y(_05473_),
    .A(_05312_),
    .B(_05310_));
 sg13g2_a22oi_1 _06236_ (.Y(_05474_),
    .B1(net52),
    .B2(_05473_),
    .A2(_05472_),
    .A1(_05471_));
 sg13g2_o21ai_1 _06237_ (.B1(_05274_),
    .Y(_05475_),
    .A1(_04953_),
    .A2(_05383_));
 sg13g2_a21oi_1 _06238_ (.A1(_05474_),
    .A2(_05384_),
    .Y(_00181_),
    .B1(_05475_));
 sg13g2_a21oi_1 _06239_ (.A1(_05395_),
    .A2(_05313_),
    .Y(_05476_),
    .B1(net58));
 sg13g2_o21ai_1 _06240_ (.B1(_05476_),
    .Y(_05477_),
    .A1(_05313_),
    .A2(_05395_));
 sg13g2_a21oi_1 _06241_ (.A1(_05413_),
    .A2(_05370_),
    .Y(_05478_),
    .B1(net52));
 sg13g2_nand2b_1 _06242_ (.Y(_05479_),
    .B(_05412_),
    .A_N(_05370_));
 sg13g2_a21oi_1 _06243_ (.A1(_05478_),
    .A2(_05479_),
    .Y(_05480_),
    .B1(net31));
 sg13g2_o21ai_1 _06244_ (.B1(net37),
    .Y(_05481_),
    .A1(_05028_),
    .A2(_05383_));
 sg13g2_a21oi_1 _06245_ (.A1(_05477_),
    .A2(_05480_),
    .Y(_00182_),
    .B1(_05481_));
 sg13g2_buf_1 _06246_ (.A(net105),
    .X(_05482_));
 sg13g2_buf_1 _06247_ (.A(_03212_),
    .X(_05483_));
 sg13g2_buf_1 _06248_ (.A(_05483_),
    .X(_05484_));
 sg13g2_inv_4 _06249_ (.A(net121),
    .Y(_05485_));
 sg13g2_buf_8 _06250_ (.A(_05485_),
    .X(_05486_));
 sg13g2_nand2_1 _06251_ (.Y(_05487_),
    .A(net115),
    .B(net92));
 sg13g2_o21ai_1 _06252_ (.B1(_05487_),
    .Y(_05488_),
    .A1(net113),
    .A2(net109));
 sg13g2_inv_1 _06253_ (.Y(_05489_),
    .A(_03311_));
 sg13g2_inv_2 _06254_ (.Y(_05490_),
    .A(net108));
 sg13g2_a22oi_1 _06255_ (.Y(_05491_),
    .B1(net112),
    .B2(_05490_),
    .A2(_05489_),
    .A1(_02970_));
 sg13g2_a221oi_1 _06256_ (.B2(net108),
    .C1(_05491_),
    .B1(net103),
    .A1(net114),
    .Y(_05492_),
    .A2(net98));
 sg13g2_inv_2 _06257_ (.Y(_05493_),
    .A(net120));
 sg13g2_buf_8 _06258_ (.A(_05493_),
    .X(_05494_));
 sg13g2_buf_8 _06259_ (.A(net91),
    .X(_05495_));
 sg13g2_nand2_1 _06260_ (.Y(_05496_),
    .A(net95),
    .B(net93));
 sg13g2_o21ai_1 _06261_ (.B1(_05496_),
    .Y(_05497_),
    .A1(_02751_),
    .A2(net76));
 sg13g2_inv_1 _06262_ (.Y(_05498_),
    .A(_05497_));
 sg13g2_o21ai_1 _06263_ (.B1(_05498_),
    .Y(_05499_),
    .A1(_05488_),
    .A2(_05492_));
 sg13g2_o21ai_1 _06264_ (.B1(_05499_),
    .Y(_05500_),
    .A1(_05259_),
    .A2(net93));
 sg13g2_nor2_1 _06265_ (.A(net126),
    .B(_03025_),
    .Y(_05501_));
 sg13g2_nor2_1 _06266_ (.A(\hvsync_gen.vpos[9] ),
    .B(_03069_),
    .Y(_05502_));
 sg13g2_inv_1 _06267_ (.Y(_05503_),
    .A(_05502_));
 sg13g2_nor2_1 _06268_ (.A(_02411_),
    .B(_05503_),
    .Y(_05504_));
 sg13g2_nand2_1 _06269_ (.Y(_05505_),
    .A(_05504_),
    .B(_03135_));
 sg13g2_o21ai_1 _06270_ (.B1(_03080_),
    .Y(_05506_),
    .A1(_04417_),
    .A2(_05505_));
 sg13g2_inv_1 _06271_ (.Y(_05507_),
    .A(net128));
 sg13g2_or4_1 _06272_ (.A(net129),
    .B(_05507_),
    .C(_02521_),
    .D(_05505_),
    .X(_05508_));
 sg13g2_nand4_1 _06273_ (.B(_05501_),
    .C(_05506_),
    .A(_05500_),
    .Y(_05509_),
    .D(_05508_));
 sg13g2_nand2_1 _06274_ (.Y(_05510_),
    .A(net103),
    .B(_03311_));
 sg13g2_o21ai_1 _06275_ (.B1(_05510_),
    .Y(_05511_),
    .A1(net115),
    .A2(_05490_));
 sg13g2_buf_1 _06276_ (.A(_00024_),
    .X(_05512_));
 sg13g2_inv_1 _06277_ (.Y(_05513_),
    .A(_05512_));
 sg13g2_o21ai_1 _06278_ (.B1(_05513_),
    .Y(_05514_),
    .A1(net77),
    .A2(net76));
 sg13g2_nand2_1 _06279_ (.Y(_05515_),
    .A(net113),
    .B(net98));
 sg13g2_nand3b_1 _06280_ (.B(_02948_),
    .C(_05515_),
    .Y(_05516_),
    .A_N(_05514_));
 sg13g2_o21ai_1 _06281_ (.B1(_02773_),
    .Y(_05517_),
    .A1(_05511_),
    .A2(_05516_));
 sg13g2_nand2_1 _06282_ (.Y(_05518_),
    .A(net77),
    .B(net76));
 sg13g2_a21oi_1 _06283_ (.A1(net112),
    .A2(_05489_),
    .Y(_05519_),
    .B1(_00034_));
 sg13g2_a22oi_1 _06284_ (.Y(_05520_),
    .B1(_02751_),
    .B2(net92),
    .A2(_05490_),
    .A1(net115));
 sg13g2_o21ai_1 _06285_ (.B1(_05520_),
    .Y(_05521_),
    .A1(_05519_),
    .A2(_05511_));
 sg13g2_nand3b_1 _06286_ (.B(_05521_),
    .C(_05515_),
    .Y(_05522_),
    .A_N(_05514_));
 sg13g2_nand3_1 _06287_ (.B(_05518_),
    .C(_05522_),
    .A(_05517_),
    .Y(_05523_));
 sg13g2_inv_1 _06288_ (.Y(_05524_),
    .A(noise));
 sg13g2_nor2_1 _06289_ (.A(net102),
    .B(net104),
    .Y(_05525_));
 sg13g2_inv_1 _06290_ (.Y(_05526_),
    .A(_05525_));
 sg13g2_nor3_1 _06291_ (.A(_05524_),
    .B(_03025_),
    .C(_05526_),
    .Y(_05527_));
 sg13g2_buf_8 _06292_ (.A(\frame_counter[8] ),
    .X(_05528_));
 sg13g2_buf_8 _06293_ (.A(\frame_counter[7] ),
    .X(_05529_));
 sg13g2_inv_2 _06294_ (.Y(_05530_),
    .A(_00036_));
 sg13g2_nor2_1 _06295_ (.A(_05529_),
    .B(_05530_),
    .Y(_05531_));
 sg13g2_inv_1 _06296_ (.Y(_05532_),
    .A(_05531_));
 sg13g2_nor2_2 _06297_ (.A(_05528_),
    .B(_05532_),
    .Y(_05533_));
 sg13g2_nor2_1 _06298_ (.A(_05501_),
    .B(_05533_),
    .Y(_05534_));
 sg13g2_nand3_1 _06299_ (.B(_05527_),
    .C(_05534_),
    .A(_05523_),
    .Y(_05535_));
 sg13g2_a22oi_1 _06300_ (.Y(_05536_),
    .B1(_05262_),
    .B2(net92),
    .A2(_05490_),
    .A1(_02751_));
 sg13g2_o21ai_1 _06301_ (.B1(net114),
    .Y(_05537_),
    .A1(_04147_),
    .A2(_03311_));
 sg13g2_nand2_1 _06302_ (.Y(_05538_),
    .A(net113),
    .B(net108));
 sg13g2_nand3_1 _06303_ (.B(_05510_),
    .C(_05538_),
    .A(_05537_),
    .Y(_05539_));
 sg13g2_a22oi_1 _06304_ (.Y(_05540_),
    .B1(_05536_),
    .B2(_05539_),
    .A2(net98),
    .A1(net95));
 sg13g2_a21o_1 _06305_ (.A2(net76),
    .A1(_02773_),
    .B1(_05540_),
    .X(_05541_));
 sg13g2_inv_2 _06306_ (.Y(_05542_),
    .A(_05528_));
 sg13g2_inv_2 _06307_ (.Y(_05543_),
    .A(\frame_counter[9] ));
 sg13g2_o21ai_1 _06308_ (.B1(_05543_),
    .Y(_05544_),
    .A1(_03899_),
    .A2(_05542_));
 sg13g2_nand2_1 _06309_ (.Y(_05545_),
    .A(_02586_),
    .B(net109));
 sg13g2_inv_1 _06310_ (.Y(_05546_),
    .A(net125));
 sg13g2_inv_1 _06311_ (.Y(_05547_),
    .A(note));
 sg13g2_nor3_1 _06312_ (.A(_02652_),
    .B(_05546_),
    .C(_05547_),
    .Y(_05548_));
 sg13g2_nand4_1 _06313_ (.B(_05544_),
    .C(_05545_),
    .A(_05541_),
    .Y(_05549_),
    .D(_05548_));
 sg13g2_nand2_1 _06314_ (.Y(_05550_),
    .A(_04736_),
    .B(_04180_));
 sg13g2_o21ai_1 _06315_ (.B1(_02806_),
    .Y(_05551_),
    .A1(_04725_),
    .A2(_05550_));
 sg13g2_inv_1 _06316_ (.Y(_05552_),
    .A(_00021_));
 sg13g2_nand2_1 _06317_ (.Y(_05553_),
    .A(net77),
    .B(_05552_));
 sg13g2_nand2_1 _06318_ (.Y(_05554_),
    .A(_02751_),
    .B(net77));
 sg13g2_nand3_1 _06319_ (.B(_05554_),
    .C(_05512_),
    .A(_05553_),
    .Y(_05555_));
 sg13g2_nand3_1 _06320_ (.B(_02773_),
    .C(_05525_),
    .A(_05555_),
    .Y(_05556_));
 sg13g2_a21o_1 _06321_ (.A2(_05513_),
    .A1(_05553_),
    .B1(_05525_),
    .X(_05557_));
 sg13g2_nand3_1 _06322_ (.B(_02674_),
    .C(_05557_),
    .A(_05556_),
    .Y(_05558_));
 sg13g2_nand4_1 _06323_ (.B(_05558_),
    .C(note2),
    .A(_05551_),
    .Y(_05559_),
    .D(_02685_));
 sg13g2_nand4_1 _06324_ (.B(_05535_),
    .C(_05549_),
    .A(_05509_),
    .Y(_05560_),
    .D(_05559_));
 sg13g2_nor2b_1 _06325_ (.A(_05482_),
    .B_N(_05560_),
    .Y(_00064_));
 sg13g2_buf_8 _06326_ (.A(_00037_),
    .X(_05561_));
 sg13g2_inv_2 _06327_ (.Y(_05562_),
    .A(_05561_));
 sg13g2_nor3_1 _06328_ (.A(net121),
    .B(net120),
    .C(_05562_),
    .Y(_05563_));
 sg13g2_xnor2_1 _06329_ (.Y(_05564_),
    .A(_03212_),
    .B(_05563_));
 sg13g2_buf_1 _06330_ (.A(_05564_),
    .X(_05565_));
 sg13g2_inv_2 _06331_ (.Y(_05566_),
    .A(net71));
 sg13g2_buf_8 _06332_ (.A(_05566_),
    .X(_05567_));
 sg13g2_buf_2 _06333_ (.A(_00056_),
    .X(_05568_));
 sg13g2_buf_8 _06334_ (.A(\r1[1] ),
    .X(_05569_));
 sg13g2_xnor2_1 _06335_ (.Y(_05570_),
    .A(_03289_),
    .B(_05569_));
 sg13g2_xor2_1 _06336_ (.B(_05570_),
    .A(_00057_),
    .X(_05571_));
 sg13g2_xnor2_1 _06337_ (.Y(_05572_),
    .A(_05568_),
    .B(_05571_));
 sg13g2_buf_2 _06338_ (.A(\r2[1] ),
    .X(_05573_));
 sg13g2_buf_2 _06339_ (.A(\r1[0] ),
    .X(_05574_));
 sg13g2_nor2_1 _06340_ (.A(_05573_),
    .B(_05574_),
    .Y(_05575_));
 sg13g2_nand2_1 _06341_ (.Y(_05576_),
    .A(_05572_),
    .B(_05575_));
 sg13g2_xor2_1 _06342_ (.B(_05574_),
    .A(_05573_),
    .X(_05577_));
 sg13g2_inv_1 _06343_ (.Y(_05578_),
    .A(_05577_));
 sg13g2_nor2_1 _06344_ (.A(_05485_),
    .B(_05578_),
    .Y(_05579_));
 sg13g2_inv_2 _06345_ (.Y(_05580_),
    .A(_05579_));
 sg13g2_nor2_1 _06346_ (.A(_05575_),
    .B(_05572_),
    .Y(_05581_));
 sg13g2_a21oi_2 _06347_ (.B1(_05581_),
    .Y(_05582_),
    .A2(_05580_),
    .A1(_05576_));
 sg13g2_buf_1 _06348_ (.A(\r2[2] ),
    .X(_05583_));
 sg13g2_inv_1 _06349_ (.Y(_05584_),
    .A(_05583_));
 sg13g2_nand2_1 _06350_ (.Y(_05585_),
    .A(_05571_),
    .B(_05568_));
 sg13g2_o21ai_1 _06351_ (.B1(_05585_),
    .Y(_05586_),
    .A1(_05584_),
    .A2(_05570_));
 sg13g2_buf_8 _06352_ (.A(\r1[2] ),
    .X(_05587_));
 sg13g2_xor2_1 _06353_ (.B(_05587_),
    .A(net121),
    .X(_05588_));
 sg13g2_inv_8 _06354_ (.Y(_05589_),
    .A(_05569_));
 sg13g2_nand2_2 _06355_ (.Y(_05590_),
    .A(_05589_),
    .B(_03289_));
 sg13g2_inv_1 _06356_ (.Y(_05591_),
    .A(_05590_));
 sg13g2_nand2_1 _06357_ (.Y(_05592_),
    .A(_05588_),
    .B(_05591_));
 sg13g2_xnor2_1 _06358_ (.Y(_05593_),
    .A(\center_x[0] ),
    .B(_05587_));
 sg13g2_nand2_1 _06359_ (.Y(_05594_),
    .A(_05593_),
    .B(_05590_));
 sg13g2_nand2_1 _06360_ (.Y(_05595_),
    .A(_05592_),
    .B(_05594_));
 sg13g2_buf_1 _06361_ (.A(\r2[3] ),
    .X(_05596_));
 sg13g2_nand2_1 _06362_ (.Y(_05597_),
    .A(_05595_),
    .B(_05596_));
 sg13g2_inv_1 _06363_ (.Y(_05598_),
    .A(_05596_));
 sg13g2_nand3_1 _06364_ (.B(_05594_),
    .C(_05598_),
    .A(_05592_),
    .Y(_05599_));
 sg13g2_nand2_1 _06365_ (.Y(_05600_),
    .A(_05597_),
    .B(_05599_));
 sg13g2_nand2_1 _06366_ (.Y(_05601_),
    .A(_05600_),
    .B(_03531_));
 sg13g2_nand3_1 _06367_ (.B(_05599_),
    .C(_03542_),
    .A(_05597_),
    .Y(_05602_));
 sg13g2_nand2_1 _06368_ (.Y(_05603_),
    .A(_05601_),
    .B(_05602_));
 sg13g2_nand2b_1 _06369_ (.Y(_05604_),
    .B(_05603_),
    .A_N(_05586_));
 sg13g2_nand3_1 _06370_ (.B(_05586_),
    .C(_05602_),
    .A(_05601_),
    .Y(_05605_));
 sg13g2_buf_2 _06371_ (.A(_05605_),
    .X(_05606_));
 sg13g2_nand2_1 _06372_ (.Y(_05607_),
    .A(_05604_),
    .B(_05606_));
 sg13g2_nor2_1 _06373_ (.A(_05582_),
    .B(_05607_),
    .Y(_05608_));
 sg13g2_inv_1 _06374_ (.Y(_05609_),
    .A(_05608_));
 sg13g2_nand2_1 _06375_ (.Y(_05610_),
    .A(_05607_),
    .B(_05582_));
 sg13g2_nand2_1 _06376_ (.Y(_05611_),
    .A(_05609_),
    .B(_05610_));
 sg13g2_buf_1 _06377_ (.A(_05611_),
    .X(_05612_));
 sg13g2_nor2_1 _06378_ (.A(_05580_),
    .B(_05572_),
    .Y(_05613_));
 sg13g2_nor2b_1 _06379_ (.A(_05581_),
    .B_N(_05576_),
    .Y(_05614_));
 sg13g2_nor2b_1 _06380_ (.A(_05579_),
    .B_N(_05614_),
    .Y(_05615_));
 sg13g2_nor2_1 _06381_ (.A(_05613_),
    .B(_05615_),
    .Y(_05616_));
 sg13g2_nor3_1 _06382_ (.A(net121),
    .B(net120),
    .C(_03289_),
    .Y(_00189_));
 sg13g2_nand2_1 _06383_ (.Y(_00190_),
    .A(_00189_),
    .B(_03223_));
 sg13g2_xnor2_1 _06384_ (.Y(_00191_),
    .A(_03921_),
    .B(_00190_));
 sg13g2_buf_2 _06385_ (.A(_00191_),
    .X(_00192_));
 sg13g2_buf_8 _06386_ (.A(_00192_),
    .X(_00193_));
 sg13g2_nand2_1 _06387_ (.Y(_00194_),
    .A(_05616_),
    .B(net65));
 sg13g2_o21ai_1 _06388_ (.B1(_00194_),
    .Y(_00195_),
    .A1(net57),
    .A2(_05612_));
 sg13g2_xnor2_1 _06389_ (.Y(_00196_),
    .A(_05485_),
    .B(_05577_));
 sg13g2_buf_1 _06390_ (.A(_00196_),
    .X(_00197_));
 sg13g2_inv_8 _06391_ (.Y(_00198_),
    .A(_03651_));
 sg13g2_nand2_2 _06392_ (.Y(_00199_),
    .A(_00198_),
    .B(net104));
 sg13g2_nand2_1 _06393_ (.Y(_00200_),
    .A(_00199_),
    .B(_03662_));
 sg13g2_buf_8 _06394_ (.A(_00200_),
    .X(_00201_));
 sg13g2_inv_4 _06395_ (.A(net70),
    .Y(_00202_));
 sg13g2_inv_1 _06396_ (.Y(_00203_),
    .A(_05563_));
 sg13g2_nor2_1 _06397_ (.A(_05483_),
    .B(_00203_),
    .Y(_00204_));
 sg13g2_nor2_1 _06398_ (.A(_03651_),
    .B(_00204_),
    .Y(_00205_));
 sg13g2_a21oi_1 _06399_ (.A1(_00202_),
    .A2(_00204_),
    .Y(_00206_),
    .B1(_00205_));
 sg13g2_buf_1 _06400_ (.A(_00206_),
    .X(_00207_));
 sg13g2_nor2_1 _06401_ (.A(_00197_),
    .B(net51),
    .Y(_00208_));
 sg13g2_inv_2 _06402_ (.Y(_00209_),
    .A(_05616_));
 sg13g2_nor2_1 _06403_ (.A(net57),
    .B(_00209_),
    .Y(_00210_));
 sg13g2_inv_1 _06404_ (.Y(_00211_),
    .A(_00210_));
 sg13g2_inv_1 _06405_ (.Y(_00212_),
    .A(_05612_));
 sg13g2_nand2_1 _06406_ (.Y(_00213_),
    .A(_00212_),
    .B(_00192_));
 sg13g2_nor2_1 _06407_ (.A(_00211_),
    .B(_00213_),
    .Y(_00214_));
 sg13g2_a21oi_1 _06408_ (.A1(_00195_),
    .A2(_00208_),
    .Y(_00215_),
    .B1(_00214_));
 sg13g2_buf_1 _06409_ (.A(_00012_),
    .X(_00216_));
 sg13g2_buf_1 _06410_ (.A(\r2[0] ),
    .X(_00217_));
 sg13g2_xnor2_1 _06411_ (.Y(_00218_),
    .A(net121),
    .B(_00217_));
 sg13g2_xnor2_1 _06412_ (.Y(_00219_),
    .A(_00216_),
    .B(_00218_));
 sg13g2_buf_1 _06413_ (.A(_00219_),
    .X(_00220_));
 sg13g2_nor2_1 _06414_ (.A(_00199_),
    .B(_00190_),
    .Y(_00221_));
 sg13g2_xnor2_1 _06415_ (.Y(_00222_),
    .A(net118),
    .B(_00221_));
 sg13g2_buf_1 _06416_ (.A(_00222_),
    .X(_00223_));
 sg13g2_inv_1 _06417_ (.Y(_00224_),
    .A(_00223_));
 sg13g2_nor2_1 _06418_ (.A(_00220_),
    .B(_00224_),
    .Y(_00225_));
 sg13g2_nor2_1 _06419_ (.A(_03651_),
    .B(\center_x[5] ),
    .Y(_00226_));
 sg13g2_nand2_1 _06420_ (.Y(_00227_),
    .A(_00226_),
    .B(_03921_));
 sg13g2_buf_8 _06421_ (.A(_00227_),
    .X(_00228_));
 sg13g2_inv_1 _06422_ (.Y(_00229_),
    .A(_00204_));
 sg13g2_nor2_1 _06423_ (.A(_00228_),
    .B(_00229_),
    .Y(_00230_));
 sg13g2_buf_1 _06424_ (.A(_00230_),
    .X(_00231_));
 sg13g2_inv_1 _06425_ (.Y(_00232_),
    .A(net50));
 sg13g2_nor2_1 _06426_ (.A(_00197_),
    .B(net45),
    .Y(_00233_));
 sg13g2_nand2_1 _06427_ (.Y(_00234_),
    .A(_00225_),
    .B(_00233_));
 sg13g2_inv_1 _06428_ (.Y(_00235_),
    .A(_00234_));
 sg13g2_inv_1 _06429_ (.Y(_00236_),
    .A(_00220_));
 sg13g2_nor2_1 _06430_ (.A(_00197_),
    .B(_00224_),
    .Y(_00237_));
 sg13g2_a21oi_1 _06431_ (.A1(net50),
    .A2(_00236_),
    .Y(_00238_),
    .B1(_00237_));
 sg13g2_nor2_1 _06432_ (.A(_00235_),
    .B(_00238_),
    .Y(_00239_));
 sg13g2_nor2b_1 _06433_ (.A(_00215_),
    .B_N(_00239_),
    .Y(_00240_));
 sg13g2_buf_1 _06434_ (.A(_00240_),
    .X(_00241_));
 sg13g2_nor2_1 _06435_ (.A(_00224_),
    .B(_00209_),
    .Y(_00242_));
 sg13g2_nor2_1 _06436_ (.A(_00233_),
    .B(_00242_),
    .Y(_00243_));
 sg13g2_nor2_1 _06437_ (.A(net45),
    .B(_00209_),
    .Y(_00244_));
 sg13g2_nand2_1 _06438_ (.Y(_00245_),
    .A(_00244_),
    .B(_00237_));
 sg13g2_inv_1 _06439_ (.Y(_00246_),
    .A(_00245_));
 sg13g2_nor2_1 _06440_ (.A(_00243_),
    .B(_00246_),
    .Y(_00247_));
 sg13g2_inv_1 _06441_ (.Y(_00248_),
    .A(_05604_));
 sg13g2_a21oi_2 _06442_ (.B1(_00248_),
    .Y(_00249_),
    .A2(_05606_),
    .A1(_05582_));
 sg13g2_buf_8 _06443_ (.A(\r1[3] ),
    .X(_00250_));
 sg13g2_xnor2_1 _06444_ (.Y(_00251_),
    .A(net120),
    .B(_00250_));
 sg13g2_inv_2 _06445_ (.Y(_00252_),
    .A(_00251_));
 sg13g2_inv_8 _06446_ (.Y(_00253_),
    .A(_05587_));
 sg13g2_nand2_1 _06447_ (.Y(_00254_),
    .A(_00253_),
    .B(net121));
 sg13g2_nor2_1 _06448_ (.A(net121),
    .B(_00253_),
    .Y(_00255_));
 sg13g2_a21oi_2 _06449_ (.B1(_00255_),
    .Y(_00256_),
    .A2(_00254_),
    .A1(_05590_));
 sg13g2_xnor2_1 _06450_ (.Y(_00257_),
    .A(_00252_),
    .B(_00256_));
 sg13g2_buf_2 _06451_ (.A(\r2[4] ),
    .X(_00258_));
 sg13g2_nand2_1 _06452_ (.Y(_00259_),
    .A(_00257_),
    .B(_00258_));
 sg13g2_xnor2_1 _06453_ (.Y(_00260_),
    .A(_00251_),
    .B(_00256_));
 sg13g2_inv_1 _06454_ (.Y(_00261_),
    .A(_00258_));
 sg13g2_nand2_1 _06455_ (.Y(_00262_),
    .A(_00260_),
    .B(_00261_));
 sg13g2_nand2_1 _06456_ (.Y(_00263_),
    .A(_00259_),
    .B(_00262_));
 sg13g2_nand2_1 _06457_ (.Y(_00264_),
    .A(_00263_),
    .B(_02904_));
 sg13g2_nand3_1 _06458_ (.B(_00262_),
    .C(_02915_),
    .A(_00259_),
    .Y(_00265_));
 sg13g2_nand2_1 _06459_ (.Y(_00266_),
    .A(_00264_),
    .B(_00265_));
 sg13g2_nor2_1 _06460_ (.A(_00055_),
    .B(_05595_),
    .Y(_00267_));
 sg13g2_nand2b_1 _06461_ (.Y(_00268_),
    .B(_05601_),
    .A_N(_00267_));
 sg13g2_nand2_1 _06462_ (.Y(_00269_),
    .A(_00266_),
    .B(_00268_));
 sg13g2_a21oi_1 _06463_ (.A1(_05600_),
    .A2(_03531_),
    .Y(_00270_),
    .B1(_00267_));
 sg13g2_nand3_1 _06464_ (.B(_00265_),
    .C(_00270_),
    .A(_00264_),
    .Y(_00271_));
 sg13g2_nand2_2 _06465_ (.Y(_00272_),
    .A(_00269_),
    .B(_00271_));
 sg13g2_xnor2_1 _06466_ (.Y(_00273_),
    .A(_00249_),
    .B(_00272_));
 sg13g2_buf_2 _06467_ (.A(_00273_),
    .X(_00274_));
 sg13g2_nor2_1 _06468_ (.A(_05566_),
    .B(_00274_),
    .Y(_00275_));
 sg13g2_inv_1 _06469_ (.Y(_00276_),
    .A(_00275_));
 sg13g2_nand2_1 _06470_ (.Y(_00277_),
    .A(_00276_),
    .B(_00213_));
 sg13g2_nor2_1 _06471_ (.A(net51),
    .B(_00209_),
    .Y(_00278_));
 sg13g2_nor2_1 _06472_ (.A(_00213_),
    .B(_00276_),
    .Y(_00279_));
 sg13g2_a21oi_1 _06473_ (.A1(_00277_),
    .A2(_00278_),
    .Y(_00280_),
    .B1(_00279_));
 sg13g2_xnor2_1 _06474_ (.Y(_00281_),
    .A(_00247_),
    .B(_00280_));
 sg13g2_xnor2_1 _06475_ (.Y(_00282_),
    .A(_00234_),
    .B(_00281_));
 sg13g2_nor2_1 _06476_ (.A(net51),
    .B(_05612_),
    .Y(_00283_));
 sg13g2_nand2b_1 _06477_ (.Y(_00284_),
    .B(_00260_),
    .A_N(_00054_));
 sg13g2_nand2_1 _06478_ (.Y(_00285_),
    .A(_00264_),
    .B(_00284_));
 sg13g2_inv_8 _06479_ (.Y(_00286_),
    .A(_00250_));
 sg13g2_nor2_1 _06480_ (.A(net120),
    .B(_00286_),
    .Y(_00287_));
 sg13g2_nor2_1 _06481_ (.A(_00255_),
    .B(_00287_),
    .Y(_00288_));
 sg13g2_nand2_1 _06482_ (.Y(_00289_),
    .A(_05594_),
    .B(_00288_));
 sg13g2_nand2_1 _06483_ (.Y(_00290_),
    .A(_00286_),
    .B(net120));
 sg13g2_nand2_1 _06484_ (.Y(_00291_),
    .A(_00289_),
    .B(_00290_));
 sg13g2_buf_2 _06485_ (.A(\r1[4] ),
    .X(_00292_));
 sg13g2_xnor2_1 _06486_ (.Y(_00293_),
    .A(_03212_),
    .B(_00292_));
 sg13g2_nand2_1 _06487_ (.Y(_00294_),
    .A(_00291_),
    .B(_00293_));
 sg13g2_xor2_1 _06488_ (.B(_00292_),
    .A(_03212_),
    .X(_00295_));
 sg13g2_nand3_1 _06489_ (.B(_00295_),
    .C(_00290_),
    .A(_00289_),
    .Y(_00296_));
 sg13g2_nand2_1 _06490_ (.Y(_00297_),
    .A(_00294_),
    .B(_00296_));
 sg13g2_buf_1 _06491_ (.A(\r2[5] ),
    .X(_00298_));
 sg13g2_inv_1 _06492_ (.Y(_00299_),
    .A(_00298_));
 sg13g2_nand2_1 _06493_ (.Y(_00300_),
    .A(_00297_),
    .B(_00299_));
 sg13g2_nand3_1 _06494_ (.B(_00296_),
    .C(_00298_),
    .A(_00294_),
    .Y(_00301_));
 sg13g2_nand2_1 _06495_ (.Y(_00302_),
    .A(_00300_),
    .B(_00301_));
 sg13g2_nand2_1 _06496_ (.Y(_00303_),
    .A(_00302_),
    .B(_03410_));
 sg13g2_nand3_1 _06497_ (.B(_00301_),
    .C(net107),
    .A(_00300_),
    .Y(_00304_));
 sg13g2_nand2_1 _06498_ (.Y(_00305_),
    .A(_00303_),
    .B(_00304_));
 sg13g2_nand2b_1 _06499_ (.Y(_00306_),
    .B(_00305_),
    .A_N(_00285_));
 sg13g2_buf_1 _06500_ (.A(_00306_),
    .X(_00307_));
 sg13g2_nand3_1 _06501_ (.B(_00304_),
    .C(_00285_),
    .A(_00303_),
    .Y(_00308_));
 sg13g2_buf_1 _06502_ (.A(_00308_),
    .X(_00309_));
 sg13g2_nand2_1 _06503_ (.Y(_00310_),
    .A(_00307_),
    .B(_00309_));
 sg13g2_nand3_1 _06504_ (.B(_00265_),
    .C(_00268_),
    .A(_00264_),
    .Y(_00311_));
 sg13g2_nand2_1 _06505_ (.Y(_00312_),
    .A(_00311_),
    .B(_05606_));
 sg13g2_nand2_1 _06506_ (.Y(_00313_),
    .A(_00266_),
    .B(_00270_));
 sg13g2_nand2_1 _06507_ (.Y(_00314_),
    .A(_00312_),
    .B(_00313_));
 sg13g2_nand2_1 _06508_ (.Y(_00315_),
    .A(_00272_),
    .B(_05608_));
 sg13g2_nand3_1 _06509_ (.B(_00314_),
    .C(_00315_),
    .A(_00310_),
    .Y(_00316_));
 sg13g2_nand2_1 _06510_ (.Y(_00317_),
    .A(_00315_),
    .B(_00314_));
 sg13g2_inv_1 _06511_ (.Y(_00318_),
    .A(_00310_));
 sg13g2_nand2_1 _06512_ (.Y(_00319_),
    .A(_00317_),
    .B(_00318_));
 sg13g2_nand2_1 _06513_ (.Y(_00320_),
    .A(_00316_),
    .B(_00319_));
 sg13g2_buf_2 _06514_ (.A(_00320_),
    .X(_00321_));
 sg13g2_inv_1 _06515_ (.Y(_00322_),
    .A(_00321_));
 sg13g2_nand2_1 _06516_ (.Y(_00323_),
    .A(_00322_),
    .B(net65));
 sg13g2_nor2_1 _06517_ (.A(_00276_),
    .B(_00323_),
    .Y(_00324_));
 sg13g2_inv_4 _06518_ (.A(_00192_),
    .Y(_00325_));
 sg13g2_nor2_1 _06519_ (.A(_05566_),
    .B(_00321_),
    .Y(_00326_));
 sg13g2_inv_1 _06520_ (.Y(_00327_),
    .A(_00326_));
 sg13g2_o21ai_1 _06521_ (.B1(_00327_),
    .Y(_00328_),
    .A1(net63),
    .A2(_00274_));
 sg13g2_nand2b_1 _06522_ (.Y(_00329_),
    .B(_00328_),
    .A_N(_00324_));
 sg13g2_xnor2_1 _06523_ (.Y(_00330_),
    .A(_00283_),
    .B(_00329_));
 sg13g2_nor2_1 _06524_ (.A(_03234_),
    .B(_03289_),
    .Y(_00331_));
 sg13g2_xnor2_1 _06525_ (.Y(_00332_),
    .A(net120),
    .B(_00331_));
 sg13g2_inv_4 _06526_ (.A(_00332_),
    .Y(_00333_));
 sg13g2_nand2_1 _06527_ (.Y(_00334_),
    .A(_00272_),
    .B(_00249_));
 sg13g2_nand3_1 _06528_ (.B(_00311_),
    .C(_00309_),
    .A(_00334_),
    .Y(_00335_));
 sg13g2_nand2_1 _06529_ (.Y(_00336_),
    .A(_00335_),
    .B(_00307_));
 sg13g2_nand2b_1 _06530_ (.Y(_00337_),
    .B(_00297_),
    .A_N(_00053_));
 sg13g2_nand2_1 _06531_ (.Y(_00338_),
    .A(_00303_),
    .B(_00337_));
 sg13g2_nand2_1 _06532_ (.Y(_00339_),
    .A(_00293_),
    .B(_00251_));
 sg13g2_inv_2 _06533_ (.Y(_00340_),
    .A(_00292_));
 sg13g2_nand2_1 _06534_ (.Y(_00341_),
    .A(_00340_),
    .B(_03212_));
 sg13g2_nor2_1 _06535_ (.A(_03212_),
    .B(_00340_),
    .Y(_00342_));
 sg13g2_a21oi_1 _06536_ (.A1(_00287_),
    .A2(_00341_),
    .Y(_00343_),
    .B1(_00342_));
 sg13g2_o21ai_1 _06537_ (.B1(_00343_),
    .Y(_00344_),
    .A1(_00339_),
    .A2(_00256_));
 sg13g2_buf_1 _06538_ (.A(_00344_),
    .X(_00345_));
 sg13g2_buf_8 _06539_ (.A(\r1[5] ),
    .X(_00346_));
 sg13g2_xor2_1 _06540_ (.B(_00346_),
    .A(net119),
    .X(_00347_));
 sg13g2_nand2_1 _06541_ (.Y(_00348_),
    .A(_00345_),
    .B(_00347_));
 sg13g2_nor2_1 _06542_ (.A(_00339_),
    .B(_00256_),
    .Y(_00349_));
 sg13g2_nor2b_1 _06543_ (.A(_00349_),
    .B_N(_00343_),
    .Y(_00350_));
 sg13g2_xnor2_1 _06544_ (.Y(_00351_),
    .A(net119),
    .B(_00346_));
 sg13g2_nand2_1 _06545_ (.Y(_00352_),
    .A(_00350_),
    .B(_00351_));
 sg13g2_nand2_1 _06546_ (.Y(_00353_),
    .A(_00348_),
    .B(_00352_));
 sg13g2_buf_2 _06547_ (.A(\r2[6] ),
    .X(_00354_));
 sg13g2_nand2_1 _06548_ (.Y(_00355_),
    .A(_00353_),
    .B(_00354_));
 sg13g2_inv_1 _06549_ (.Y(_00356_),
    .A(_00354_));
 sg13g2_nand3_1 _06550_ (.B(_00352_),
    .C(_00356_),
    .A(_00348_),
    .Y(_00357_));
 sg13g2_nand2_1 _06551_ (.Y(_00358_),
    .A(_00355_),
    .B(_00357_));
 sg13g2_nand2_1 _06552_ (.Y(_00359_),
    .A(_00358_),
    .B(_03629_));
 sg13g2_nand3_1 _06553_ (.B(_00357_),
    .C(_03640_),
    .A(_00355_),
    .Y(_00360_));
 sg13g2_nand3_1 _06554_ (.B(_00359_),
    .C(_00360_),
    .A(_00338_),
    .Y(_00361_));
 sg13g2_nand2_1 _06555_ (.Y(_00362_),
    .A(_00359_),
    .B(_00360_));
 sg13g2_nand2b_1 _06556_ (.Y(_00363_),
    .B(_00362_),
    .A_N(_00338_));
 sg13g2_nand2_1 _06557_ (.Y(_00364_),
    .A(_00361_),
    .B(_00363_));
 sg13g2_nand2_1 _06558_ (.Y(_00365_),
    .A(_00336_),
    .B(_00364_));
 sg13g2_xnor2_1 _06559_ (.Y(_00366_),
    .A(_00338_),
    .B(_00362_));
 sg13g2_nand3_1 _06560_ (.B(_00366_),
    .C(_00307_),
    .A(_00335_),
    .Y(_00367_));
 sg13g2_nand2_1 _06561_ (.Y(_00368_),
    .A(_00365_),
    .B(_00367_));
 sg13g2_buf_2 _06562_ (.A(_00368_),
    .X(_00369_));
 sg13g2_nor2_1 _06563_ (.A(net75),
    .B(_00369_),
    .Y(_00370_));
 sg13g2_nand2_1 _06564_ (.Y(_00371_),
    .A(_00347_),
    .B(_00342_));
 sg13g2_nand2_1 _06565_ (.Y(_00372_),
    .A(net119),
    .B(_00346_));
 sg13g2_nand2_1 _06566_ (.Y(_00373_),
    .A(_00371_),
    .B(_00372_));
 sg13g2_nand2_1 _06567_ (.Y(_00374_),
    .A(_00347_),
    .B(_00293_));
 sg13g2_a21oi_1 _06568_ (.A1(_00255_),
    .A2(_00290_),
    .Y(_00375_),
    .B1(_00287_));
 sg13g2_nor2_1 _06569_ (.A(_00374_),
    .B(_00375_),
    .Y(_00376_));
 sg13g2_nor2_1 _06570_ (.A(_00373_),
    .B(_00376_),
    .Y(_00377_));
 sg13g2_nor2_1 _06571_ (.A(_05588_),
    .B(_00252_),
    .Y(_00378_));
 sg13g2_nor2_1 _06572_ (.A(_00351_),
    .B(_00295_),
    .Y(_00379_));
 sg13g2_nand3_1 _06573_ (.B(_00379_),
    .C(_05590_),
    .A(_00378_),
    .Y(_00380_));
 sg13g2_nand2_1 _06574_ (.Y(_00381_),
    .A(_00377_),
    .B(_00380_));
 sg13g2_buf_8 _06575_ (.A(\r1[6] ),
    .X(_00382_));
 sg13g2_inv_2 _06576_ (.Y(_00383_),
    .A(_00382_));
 sg13g2_nand2_1 _06577_ (.Y(_00384_),
    .A(_00200_),
    .B(_00383_));
 sg13g2_nand3_1 _06578_ (.B(_00382_),
    .C(_03662_),
    .A(_00199_),
    .Y(_00385_));
 sg13g2_nand2_1 _06579_ (.Y(_00386_),
    .A(_00384_),
    .B(_00385_));
 sg13g2_nand2_1 _06580_ (.Y(_00387_),
    .A(_00381_),
    .B(_00386_));
 sg13g2_xnor2_1 _06581_ (.Y(_00388_),
    .A(_00382_),
    .B(net70));
 sg13g2_nand3_1 _06582_ (.B(_00380_),
    .C(_00388_),
    .A(_00377_),
    .Y(_00389_));
 sg13g2_buf_1 _06583_ (.A(_00389_),
    .X(_00390_));
 sg13g2_nand2_1 _06584_ (.Y(_00391_),
    .A(_00387_),
    .B(_00390_));
 sg13g2_inv_1 _06585_ (.Y(_00392_),
    .A(_00051_));
 sg13g2_nand2_1 _06586_ (.Y(_00393_),
    .A(_00391_),
    .B(_00392_));
 sg13g2_nand3_1 _06587_ (.B(_00390_),
    .C(_00051_),
    .A(_00387_),
    .Y(_00394_));
 sg13g2_nand2_1 _06588_ (.Y(_00395_),
    .A(_00393_),
    .B(_00394_));
 sg13g2_inv_1 _06589_ (.Y(_00396_),
    .A(_00052_));
 sg13g2_nand3_1 _06590_ (.B(_00352_),
    .C(_00396_),
    .A(_00348_),
    .Y(_00397_));
 sg13g2_nand2_1 _06591_ (.Y(_00398_),
    .A(_00359_),
    .B(_00397_));
 sg13g2_nand2b_1 _06592_ (.Y(_00399_),
    .B(_00398_),
    .A_N(_00395_));
 sg13g2_nand3_1 _06593_ (.B(_00395_),
    .C(_00397_),
    .A(_00359_),
    .Y(_00400_));
 sg13g2_nand2_1 _06594_ (.Y(_00401_),
    .A(_00399_),
    .B(_00400_));
 sg13g2_nand3_1 _06595_ (.B(_00317_),
    .C(_00318_),
    .A(_00366_),
    .Y(_00402_));
 sg13g2_nand2_1 _06596_ (.Y(_00403_),
    .A(_00361_),
    .B(_00309_));
 sg13g2_nand2_1 _06597_ (.Y(_00404_),
    .A(_00403_),
    .B(_00363_));
 sg13g2_nand2_1 _06598_ (.Y(_00405_),
    .A(_00402_),
    .B(_00404_));
 sg13g2_xnor2_1 _06599_ (.Y(_00406_),
    .A(_00401_),
    .B(_00405_));
 sg13g2_buf_2 _06600_ (.A(_00406_),
    .X(_00407_));
 sg13g2_nand2_1 _06601_ (.Y(_00408_),
    .A(_03234_),
    .B(_03289_));
 sg13g2_nor2b_1 _06602_ (.A(_00331_),
    .B_N(_00408_),
    .Y(_00409_));
 sg13g2_buf_1 _06603_ (.A(_00409_),
    .X(_00410_));
 sg13g2_nand2_1 _06604_ (.Y(_00411_),
    .A(_00407_),
    .B(_00410_));
 sg13g2_buf_8 _06605_ (.A(_05561_),
    .X(_00412_));
 sg13g2_nor2_1 _06606_ (.A(_00401_),
    .B(_00364_),
    .Y(_00413_));
 sg13g2_inv_1 _06607_ (.Y(_00414_),
    .A(_00311_));
 sg13g2_inv_1 _06608_ (.Y(_00415_),
    .A(_00309_));
 sg13g2_a21oi_1 _06609_ (.A1(_00307_),
    .A2(_00414_),
    .Y(_00416_),
    .B1(_00415_));
 sg13g2_inv_1 _06610_ (.Y(_00417_),
    .A(_00416_));
 sg13g2_nor2b_1 _06611_ (.A(_00398_),
    .B_N(_00395_),
    .Y(_00418_));
 sg13g2_o21ai_1 _06612_ (.B1(_00399_),
    .Y(_00419_),
    .A1(_00418_),
    .A2(_00361_));
 sg13g2_a21oi_1 _06613_ (.A1(_00413_),
    .A2(_00417_),
    .Y(_00420_),
    .B1(_00419_));
 sg13g2_inv_1 _06614_ (.Y(_00421_),
    .A(_00272_));
 sg13g2_nor2_1 _06615_ (.A(_00421_),
    .B(_00310_),
    .Y(_00422_));
 sg13g2_nand3_1 _06616_ (.B(_00249_),
    .C(_00422_),
    .A(_00413_),
    .Y(_00423_));
 sg13g2_nand2_1 _06617_ (.Y(_00424_),
    .A(_00420_),
    .B(_00423_));
 sg13g2_nand2_1 _06618_ (.Y(_00425_),
    .A(_00199_),
    .B(_03629_));
 sg13g2_nor2_1 _06619_ (.A(_03651_),
    .B(net119),
    .Y(_00426_));
 sg13g2_nand2_1 _06620_ (.Y(_00427_),
    .A(_00426_),
    .B(_03640_));
 sg13g2_nand3_1 _06621_ (.B(_00044_),
    .C(_00427_),
    .A(_00425_),
    .Y(_00428_));
 sg13g2_nand2_1 _06622_ (.Y(_00429_),
    .A(_00199_),
    .B(_03640_));
 sg13g2_inv_1 _06623_ (.Y(_00430_),
    .A(_00044_));
 sg13g2_nand2_1 _06624_ (.Y(_00431_),
    .A(_00426_),
    .B(_03629_));
 sg13g2_buf_8 _06625_ (.A(_00431_),
    .X(_00432_));
 sg13g2_nand3_1 _06626_ (.B(_00430_),
    .C(net74),
    .A(_00429_),
    .Y(_00433_));
 sg13g2_nand2_1 _06627_ (.Y(_00434_),
    .A(_00428_),
    .B(_00433_));
 sg13g2_buf_8 _06628_ (.A(_00434_),
    .X(_00435_));
 sg13g2_nor2_1 _06629_ (.A(_00351_),
    .B(_00386_),
    .Y(_00436_));
 sg13g2_nand2_1 _06630_ (.Y(_00437_),
    .A(_00345_),
    .B(_00436_));
 sg13g2_nor2_1 _06631_ (.A(_00043_),
    .B(net70),
    .Y(_00438_));
 sg13g2_inv_1 _06632_ (.Y(_00439_),
    .A(_00372_));
 sg13g2_nand3_1 _06633_ (.B(_00385_),
    .C(_00439_),
    .A(_00384_),
    .Y(_00440_));
 sg13g2_nand2b_2 _06634_ (.Y(_00441_),
    .B(_00440_),
    .A_N(_00438_));
 sg13g2_inv_4 _06635_ (.A(_00441_),
    .Y(_00442_));
 sg13g2_nand2_1 _06636_ (.Y(_00443_),
    .A(_00437_),
    .B(_00442_));
 sg13g2_nand2b_1 _06637_ (.Y(_00444_),
    .B(_00443_),
    .A_N(_00435_));
 sg13g2_nand3_1 _06638_ (.B(_00442_),
    .C(_00435_),
    .A(_00437_),
    .Y(_00445_));
 sg13g2_nand2_1 _06639_ (.Y(_00446_),
    .A(_00444_),
    .B(_00445_));
 sg13g2_buf_1 _06640_ (.A(\r2[8] ),
    .X(_00447_));
 sg13g2_nand2_1 _06641_ (.Y(_00448_),
    .A(_00446_),
    .B(_00447_));
 sg13g2_inv_1 _06642_ (.Y(_00449_),
    .A(_00447_));
 sg13g2_nand3_1 _06643_ (.B(_00445_),
    .C(_00449_),
    .A(_00444_),
    .Y(_00450_));
 sg13g2_inv_1 _06644_ (.Y(_00451_),
    .A(\r2[7] ));
 sg13g2_a21oi_2 _06645_ (.B1(_00451_),
    .Y(_00452_),
    .A2(_00390_),
    .A1(_00387_));
 sg13g2_a21oi_1 _06646_ (.A1(_00448_),
    .A2(_00450_),
    .Y(_00453_),
    .B1(_00452_));
 sg13g2_nand3_1 _06647_ (.B(_00450_),
    .C(_00452_),
    .A(_00448_),
    .Y(_00454_));
 sg13g2_inv_1 _06648_ (.Y(_00455_),
    .A(_00454_));
 sg13g2_nor2_1 _06649_ (.A(_00453_),
    .B(_00455_),
    .Y(_00456_));
 sg13g2_nand2_1 _06650_ (.Y(_00457_),
    .A(_00424_),
    .B(_00456_));
 sg13g2_nand2_1 _06651_ (.Y(_00458_),
    .A(_00448_),
    .B(_00450_));
 sg13g2_xor2_1 _06652_ (.B(_00458_),
    .A(_00452_),
    .X(_00459_));
 sg13g2_nand3_1 _06653_ (.B(_00423_),
    .C(_00459_),
    .A(_00420_),
    .Y(_00460_));
 sg13g2_nand2_1 _06654_ (.Y(_00461_),
    .A(_00457_),
    .B(_00460_));
 sg13g2_buf_8 _06655_ (.A(_00461_),
    .X(_00462_));
 sg13g2_nor2_1 _06656_ (.A(net101),
    .B(_00462_),
    .Y(_00463_));
 sg13g2_nand2b_1 _06657_ (.Y(_00464_),
    .B(_00463_),
    .A_N(_00411_));
 sg13g2_nand3_1 _06658_ (.B(_00460_),
    .C(_05562_),
    .A(_00457_),
    .Y(_00465_));
 sg13g2_nand2_1 _06659_ (.Y(_00466_),
    .A(_00465_),
    .B(_00411_));
 sg13g2_nand2_1 _06660_ (.Y(_00467_),
    .A(_00464_),
    .B(_00466_));
 sg13g2_nand2b_1 _06661_ (.Y(_00468_),
    .B(_00467_),
    .A_N(_00370_));
 sg13g2_nand3_1 _06662_ (.B(_00466_),
    .C(_00370_),
    .A(_00464_),
    .Y(_00469_));
 sg13g2_nand2_1 _06663_ (.Y(_00470_),
    .A(_00468_),
    .B(_00469_));
 sg13g2_nand2_1 _06664_ (.Y(_00471_),
    .A(_00407_),
    .B(_05562_));
 sg13g2_inv_1 _06665_ (.Y(_00472_),
    .A(_00369_));
 sg13g2_nand2_1 _06666_ (.Y(_00473_),
    .A(_00472_),
    .B(_00410_));
 sg13g2_nand2_1 _06667_ (.Y(_00474_),
    .A(_00471_),
    .B(_00473_));
 sg13g2_nor2_1 _06668_ (.A(net75),
    .B(_00321_),
    .Y(_00475_));
 sg13g2_nor2_1 _06669_ (.A(_05561_),
    .B(_00369_),
    .Y(_00476_));
 sg13g2_inv_1 _06670_ (.Y(_00477_),
    .A(_00476_));
 sg13g2_nor2_1 _06671_ (.A(_00477_),
    .B(_00411_),
    .Y(_00478_));
 sg13g2_a21oi_1 _06672_ (.A1(_00474_),
    .A2(_00475_),
    .Y(_00479_),
    .B1(_00478_));
 sg13g2_nand2_1 _06673_ (.Y(_00480_),
    .A(_00470_),
    .B(_00479_));
 sg13g2_inv_1 _06674_ (.Y(_00481_),
    .A(_00479_));
 sg13g2_nand3_1 _06675_ (.B(_00469_),
    .C(_00481_),
    .A(_00468_),
    .Y(_00482_));
 sg13g2_nand2_1 _06676_ (.Y(_00483_),
    .A(_00480_),
    .B(_00482_));
 sg13g2_nand2b_1 _06677_ (.Y(_00484_),
    .B(_00483_),
    .A_N(_00330_));
 sg13g2_nand3_1 _06678_ (.B(_00482_),
    .C(_00330_),
    .A(_00480_),
    .Y(_00485_));
 sg13g2_nand2_1 _06679_ (.Y(_00486_),
    .A(_00484_),
    .B(_00485_));
 sg13g2_nand3b_1 _06680_ (.B(_00475_),
    .C(_00474_),
    .Y(_00487_),
    .A_N(_00478_));
 sg13g2_xnor2_1 _06681_ (.Y(_00488_),
    .A(_00473_),
    .B(_00471_));
 sg13g2_nand2b_1 _06682_ (.Y(_00489_),
    .B(_00488_),
    .A_N(_00475_));
 sg13g2_nand2_1 _06683_ (.Y(_00490_),
    .A(_00487_),
    .B(_00489_));
 sg13g2_nand2_1 _06684_ (.Y(_00491_),
    .A(_00322_),
    .B(_00410_));
 sg13g2_nand2_1 _06685_ (.Y(_00492_),
    .A(_00477_),
    .B(_00491_));
 sg13g2_nor2_1 _06686_ (.A(net75),
    .B(_00274_),
    .Y(_00493_));
 sg13g2_nor2_1 _06687_ (.A(_05561_),
    .B(_00321_),
    .Y(_00494_));
 sg13g2_inv_1 _06688_ (.Y(_00495_),
    .A(_00494_));
 sg13g2_nor2_1 _06689_ (.A(_00495_),
    .B(_00473_),
    .Y(_00496_));
 sg13g2_a21oi_1 _06690_ (.A1(_00492_),
    .A2(_00493_),
    .Y(_00497_),
    .B1(_00496_));
 sg13g2_nand2_1 _06691_ (.Y(_00498_),
    .A(_00490_),
    .B(_00497_));
 sg13g2_nand2b_1 _06692_ (.Y(_00499_),
    .B(_00277_),
    .A_N(_00279_));
 sg13g2_xnor2_1 _06693_ (.Y(_00500_),
    .A(_00278_),
    .B(_00499_));
 sg13g2_inv_1 _06694_ (.Y(_00501_),
    .A(_00497_));
 sg13g2_nand3_1 _06695_ (.B(_00489_),
    .C(_00501_),
    .A(_00487_),
    .Y(_00502_));
 sg13g2_inv_1 _06696_ (.Y(_00503_),
    .A(_00502_));
 sg13g2_a21oi_1 _06697_ (.A1(_00498_),
    .A2(_00500_),
    .Y(_00504_),
    .B1(_00503_));
 sg13g2_nand2_1 _06698_ (.Y(_00505_),
    .A(_00486_),
    .B(_00504_));
 sg13g2_inv_1 _06699_ (.Y(_00506_),
    .A(_00504_));
 sg13g2_nand3_1 _06700_ (.B(_00485_),
    .C(_00506_),
    .A(_00484_),
    .Y(_00507_));
 sg13g2_nand2_1 _06701_ (.Y(_00508_),
    .A(_00505_),
    .B(_00507_));
 sg13g2_nand2b_1 _06702_ (.Y(_00509_),
    .B(_00508_),
    .A_N(_00282_));
 sg13g2_nand3_1 _06703_ (.B(_00507_),
    .C(_00282_),
    .A(_00505_),
    .Y(_00510_));
 sg13g2_nand2_1 _06704_ (.Y(_00511_),
    .A(_00509_),
    .B(_00510_));
 sg13g2_nand2_1 _06705_ (.Y(_00512_),
    .A(_00498_),
    .B(_00502_));
 sg13g2_nand2b_1 _06706_ (.Y(_00513_),
    .B(_00512_),
    .A_N(_00500_));
 sg13g2_nand3_1 _06707_ (.B(_00502_),
    .C(_00500_),
    .A(_00498_),
    .Y(_00514_));
 sg13g2_nand2_1 _06708_ (.Y(_00515_),
    .A(_00513_),
    .B(_00514_));
 sg13g2_xor2_1 _06709_ (.B(_00476_),
    .A(_00491_),
    .X(_00516_));
 sg13g2_xor2_1 _06710_ (.B(_00516_),
    .A(_00493_),
    .X(_00517_));
 sg13g2_inv_2 _06711_ (.Y(_00518_),
    .A(_00410_));
 sg13g2_nor2_1 _06712_ (.A(_00518_),
    .B(_00274_),
    .Y(_00519_));
 sg13g2_inv_1 _06713_ (.Y(_00520_),
    .A(_00519_));
 sg13g2_nand2_1 _06714_ (.Y(_00521_),
    .A(_00495_),
    .B(_00520_));
 sg13g2_nor2_1 _06715_ (.A(net75),
    .B(_05612_),
    .Y(_00522_));
 sg13g2_nor2_1 _06716_ (.A(_00520_),
    .B(_00495_),
    .Y(_00523_));
 sg13g2_a21oi_2 _06717_ (.B1(_00523_),
    .Y(_00524_),
    .A2(_00522_),
    .A1(_00521_));
 sg13g2_nand2_1 _06718_ (.Y(_00525_),
    .A(_00517_),
    .B(_00524_));
 sg13g2_o21ai_1 _06719_ (.B1(_00195_),
    .Y(_00526_),
    .A1(_00213_),
    .A2(_00211_));
 sg13g2_xnor2_1 _06720_ (.Y(_00527_),
    .A(_00208_),
    .B(_00526_));
 sg13g2_nor2_1 _06721_ (.A(_00524_),
    .B(_00517_),
    .Y(_00528_));
 sg13g2_a21oi_1 _06722_ (.A1(_00525_),
    .A2(_00527_),
    .Y(_00529_),
    .B1(_00528_));
 sg13g2_nand2_1 _06723_ (.Y(_00530_),
    .A(_00515_),
    .B(_00529_));
 sg13g2_xnor2_1 _06724_ (.Y(_00531_),
    .A(_00239_),
    .B(_00215_));
 sg13g2_inv_1 _06725_ (.Y(_00532_),
    .A(_00529_));
 sg13g2_nand3_1 _06726_ (.B(_00514_),
    .C(_00532_),
    .A(_00513_),
    .Y(_00533_));
 sg13g2_inv_1 _06727_ (.Y(_00534_),
    .A(_00533_));
 sg13g2_a21oi_1 _06728_ (.A1(_00530_),
    .A2(_00531_),
    .Y(_00535_),
    .B1(_00534_));
 sg13g2_nand2_1 _06729_ (.Y(_00536_),
    .A(_00511_),
    .B(_00535_));
 sg13g2_inv_1 _06730_ (.Y(_00537_),
    .A(_00535_));
 sg13g2_nand3_1 _06731_ (.B(_00510_),
    .C(_00537_),
    .A(_00509_),
    .Y(_00538_));
 sg13g2_nand2_1 _06732_ (.Y(_00539_),
    .A(_00536_),
    .B(_00538_));
 sg13g2_nand2b_1 _06733_ (.Y(_00540_),
    .B(_00539_),
    .A_N(_00241_));
 sg13g2_nand3_1 _06734_ (.B(_00538_),
    .C(_00241_),
    .A(_00536_),
    .Y(_00541_));
 sg13g2_nand2_1 _06735_ (.Y(_00542_),
    .A(_00540_),
    .B(_00541_));
 sg13g2_nand2_1 _06736_ (.Y(_00543_),
    .A(_00530_),
    .B(_00533_));
 sg13g2_nand2b_1 _06737_ (.Y(_00544_),
    .B(_00543_),
    .A_N(_00531_));
 sg13g2_nand3_1 _06738_ (.B(_00533_),
    .C(_00531_),
    .A(_00530_),
    .Y(_00545_));
 sg13g2_nand2_1 _06739_ (.Y(_00546_),
    .A(_00544_),
    .B(_00545_));
 sg13g2_xnor2_1 _06740_ (.Y(_00547_),
    .A(_00524_),
    .B(_00517_));
 sg13g2_xor2_1 _06741_ (.B(_00547_),
    .A(_00527_),
    .X(_00548_));
 sg13g2_nor2b_1 _06742_ (.A(_00523_),
    .B_N(_00521_),
    .Y(_00549_));
 sg13g2_xnor2_1 _06743_ (.Y(_00550_),
    .A(_00522_),
    .B(_00549_));
 sg13g2_buf_8 _06744_ (.A(_00518_),
    .X(_00551_));
 sg13g2_nor2_1 _06745_ (.A(net62),
    .B(_05612_),
    .Y(_00552_));
 sg13g2_inv_1 _06746_ (.Y(_00553_),
    .A(_00552_));
 sg13g2_o21ai_1 _06747_ (.B1(_00553_),
    .Y(_00554_),
    .A1(net101),
    .A2(_00274_));
 sg13g2_buf_1 _06748_ (.A(_00333_),
    .X(_00555_));
 sg13g2_nor2_1 _06749_ (.A(net69),
    .B(_00209_),
    .Y(_00556_));
 sg13g2_nand2_1 _06750_ (.Y(_00557_),
    .A(_00212_),
    .B(_05562_));
 sg13g2_nor2_1 _06751_ (.A(_00557_),
    .B(_00520_),
    .Y(_00558_));
 sg13g2_a21oi_1 _06752_ (.A1(_00554_),
    .A2(_00556_),
    .Y(_00559_),
    .B1(_00558_));
 sg13g2_nand2_1 _06753_ (.Y(_00560_),
    .A(_00550_),
    .B(_00559_));
 sg13g2_nor2_1 _06754_ (.A(_00220_),
    .B(net51),
    .Y(_00561_));
 sg13g2_nor2_1 _06755_ (.A(_00197_),
    .B(net63),
    .Y(_00562_));
 sg13g2_inv_1 _06756_ (.Y(_00563_),
    .A(_00562_));
 sg13g2_nor2_1 _06757_ (.A(_00563_),
    .B(_00211_),
    .Y(_00564_));
 sg13g2_nand2_1 _06758_ (.Y(_00565_),
    .A(_00211_),
    .B(_00563_));
 sg13g2_nand2b_1 _06759_ (.Y(_00566_),
    .B(_00565_),
    .A_N(_00564_));
 sg13g2_xnor2_1 _06760_ (.Y(_00567_),
    .A(_00561_),
    .B(_00566_));
 sg13g2_nor2_1 _06761_ (.A(_00559_),
    .B(_00550_),
    .Y(_00568_));
 sg13g2_a21oi_1 _06762_ (.A1(_00560_),
    .A2(_00567_),
    .Y(_00569_),
    .B1(_00568_));
 sg13g2_nand2_1 _06763_ (.Y(_00570_),
    .A(_00548_),
    .B(_00569_));
 sg13g2_a21oi_1 _06764_ (.A1(_00565_),
    .A2(_00561_),
    .Y(_00571_),
    .B1(_00564_));
 sg13g2_xnor2_1 _06765_ (.Y(_00572_),
    .A(_00225_),
    .B(_00571_));
 sg13g2_nor2_1 _06766_ (.A(_00569_),
    .B(_00548_),
    .Y(_00573_));
 sg13g2_a21oi_1 _06767_ (.A1(_00570_),
    .A2(_00572_),
    .Y(_00574_),
    .B1(_00573_));
 sg13g2_nand2_1 _06768_ (.Y(_00575_),
    .A(_00546_),
    .B(_00574_));
 sg13g2_nor2b_1 _06769_ (.A(_00571_),
    .B_N(_00225_),
    .Y(_00576_));
 sg13g2_inv_1 _06770_ (.Y(_00577_),
    .A(_00574_));
 sg13g2_nand3_1 _06771_ (.B(_00577_),
    .C(_00545_),
    .A(_00544_),
    .Y(_00578_));
 sg13g2_inv_1 _06772_ (.Y(_00579_),
    .A(_00578_));
 sg13g2_a21oi_1 _06773_ (.A1(_00575_),
    .A2(_00576_),
    .Y(_00580_),
    .B1(_00579_));
 sg13g2_nand2_1 _06774_ (.Y(_00581_),
    .A(_00542_),
    .B(_00580_));
 sg13g2_inv_1 _06775_ (.Y(_00582_),
    .A(_00580_));
 sg13g2_nand3_1 _06776_ (.B(_00541_),
    .C(_00582_),
    .A(_00540_),
    .Y(_00583_));
 sg13g2_inv_1 _06777_ (.Y(_00584_),
    .A(_00576_));
 sg13g2_nand2_1 _06778_ (.Y(_00585_),
    .A(_00575_),
    .B(_00578_));
 sg13g2_nor2_1 _06779_ (.A(_00584_),
    .B(_00585_),
    .Y(_00586_));
 sg13g2_nand2_1 _06780_ (.Y(_00587_),
    .A(_00585_),
    .B(_00584_));
 sg13g2_nor2b_1 _06781_ (.A(_00558_),
    .B_N(_00554_),
    .Y(_00588_));
 sg13g2_xnor2_1 _06782_ (.Y(_00589_),
    .A(_00556_),
    .B(_00588_));
 sg13g2_o21ai_1 _06783_ (.B1(_00557_),
    .Y(_00590_),
    .A1(net62),
    .A2(_00209_));
 sg13g2_nor2_1 _06784_ (.A(net75),
    .B(_00197_),
    .Y(_00591_));
 sg13g2_nor2_1 _06785_ (.A(_05561_),
    .B(_00209_),
    .Y(_00592_));
 sg13g2_inv_1 _06786_ (.Y(_00593_),
    .A(_00592_));
 sg13g2_nor2_1 _06787_ (.A(_00593_),
    .B(_00553_),
    .Y(_00594_));
 sg13g2_a21oi_2 _06788_ (.B1(_00594_),
    .Y(_00595_),
    .A2(_00591_),
    .A1(_00590_));
 sg13g2_nand2_1 _06789_ (.Y(_00596_),
    .A(_00589_),
    .B(_00595_));
 sg13g2_inv_1 _06790_ (.Y(_00597_),
    .A(_00197_));
 sg13g2_a22oi_1 _06791_ (.Y(_00598_),
    .B1(_00236_),
    .B2(net65),
    .A2(net71),
    .A1(_00597_));
 sg13g2_nor2_1 _06792_ (.A(_00220_),
    .B(net57),
    .Y(_00599_));
 sg13g2_inv_1 _06793_ (.Y(_00600_),
    .A(_00599_));
 sg13g2_nor2_1 _06794_ (.A(_00600_),
    .B(_00563_),
    .Y(_00601_));
 sg13g2_nor2_1 _06795_ (.A(_00598_),
    .B(_00601_),
    .Y(_00602_));
 sg13g2_nor2_1 _06796_ (.A(_00595_),
    .B(_00589_),
    .Y(_00603_));
 sg13g2_a21oi_1 _06797_ (.A1(_00596_),
    .A2(_00602_),
    .Y(_00604_),
    .B1(_00603_));
 sg13g2_nor2b_1 _06798_ (.A(_00568_),
    .B_N(_00560_),
    .Y(_00605_));
 sg13g2_xnor2_1 _06799_ (.Y(_00606_),
    .A(_00567_),
    .B(_00605_));
 sg13g2_nor2_1 _06800_ (.A(_00604_),
    .B(_00606_),
    .Y(_00607_));
 sg13g2_nand2_1 _06801_ (.Y(_00608_),
    .A(_00606_),
    .B(_00604_));
 sg13g2_nand2b_1 _06802_ (.Y(_00609_),
    .B(_00608_),
    .A_N(_00607_));
 sg13g2_buf_1 _06803_ (.A(_00410_),
    .X(_00610_));
 sg13g2_nand2_1 _06804_ (.Y(_00611_),
    .A(_00597_),
    .B(net68));
 sg13g2_nand2_1 _06805_ (.Y(_00612_),
    .A(_00593_),
    .B(_00611_));
 sg13g2_nor2_1 _06806_ (.A(net75),
    .B(_00220_),
    .Y(_00613_));
 sg13g2_nor2_1 _06807_ (.A(_00611_),
    .B(_00593_),
    .Y(_00614_));
 sg13g2_a21oi_1 _06808_ (.A1(_00612_),
    .A2(_00613_),
    .Y(_00615_),
    .B1(_00614_));
 sg13g2_nand2b_1 _06809_ (.Y(_00616_),
    .B(_00590_),
    .A_N(_00594_));
 sg13g2_xor2_1 _06810_ (.B(_00616_),
    .A(_00591_),
    .X(_00617_));
 sg13g2_xnor2_1 _06811_ (.Y(_00618_),
    .A(_00615_),
    .B(_00617_));
 sg13g2_nand2b_1 _06812_ (.Y(_00619_),
    .B(_00599_),
    .A_N(_00618_));
 sg13g2_nand2_1 _06813_ (.Y(_00620_),
    .A(_00618_),
    .B(_00600_));
 sg13g2_nor2b_1 _06814_ (.A(_00614_),
    .B_N(_00612_),
    .Y(_00621_));
 sg13g2_xnor2_1 _06815_ (.Y(_00622_),
    .A(_00613_),
    .B(_00621_));
 sg13g2_nor4_1 _06816_ (.A(net101),
    .B(_00220_),
    .C(_00611_),
    .D(_00622_),
    .Y(_00623_));
 sg13g2_nand3_1 _06817_ (.B(_00620_),
    .C(_00623_),
    .A(_00619_),
    .Y(_00624_));
 sg13g2_xnor2_1 _06818_ (.Y(_00625_),
    .A(_00595_),
    .B(_00589_));
 sg13g2_xor2_1 _06819_ (.B(_00625_),
    .A(_00602_),
    .X(_00626_));
 sg13g2_nand2_1 _06820_ (.Y(_00627_),
    .A(_00624_),
    .B(_00626_));
 sg13g2_nor2_1 _06821_ (.A(_00615_),
    .B(_00617_),
    .Y(_00628_));
 sg13g2_nor2b_1 _06822_ (.A(_00628_),
    .B_N(_00619_),
    .Y(_00629_));
 sg13g2_inv_1 _06823_ (.Y(_00630_),
    .A(_00629_));
 sg13g2_nor2_1 _06824_ (.A(_00626_),
    .B(_00624_),
    .Y(_00631_));
 sg13g2_a21oi_1 _06825_ (.A1(_00627_),
    .A2(_00630_),
    .Y(_00632_),
    .B1(_00631_));
 sg13g2_nand2_1 _06826_ (.Y(_00633_),
    .A(_00609_),
    .B(_00632_));
 sg13g2_nand2_1 _06827_ (.Y(_00634_),
    .A(_00633_),
    .B(_00601_));
 sg13g2_inv_1 _06828_ (.Y(_00635_),
    .A(_00632_));
 sg13g2_a21oi_1 _06829_ (.A1(_00635_),
    .A2(_00608_),
    .Y(_00636_),
    .B1(_00607_));
 sg13g2_nand2_1 _06830_ (.Y(_00637_),
    .A(_00634_),
    .B(_00636_));
 sg13g2_nand2b_1 _06831_ (.Y(_00638_),
    .B(_00570_),
    .A_N(_00573_));
 sg13g2_xnor2_1 _06832_ (.Y(_00639_),
    .A(_00572_),
    .B(_00638_));
 sg13g2_nand2_1 _06833_ (.Y(_00640_),
    .A(_00637_),
    .B(_00639_));
 sg13g2_nand2b_1 _06834_ (.Y(_00641_),
    .B(_00609_),
    .A_N(_00601_));
 sg13g2_nand3_1 _06835_ (.B(_00607_),
    .C(_00635_),
    .A(_00641_),
    .Y(_00642_));
 sg13g2_nand2_1 _06836_ (.Y(_00643_),
    .A(_00640_),
    .B(_00642_));
 sg13g2_nand2_1 _06837_ (.Y(_00644_),
    .A(_00587_),
    .B(_00643_));
 sg13g2_nor2_1 _06838_ (.A(_00586_),
    .B(_00644_),
    .Y(_00645_));
 sg13g2_nand3_1 _06839_ (.B(_00583_),
    .C(_00645_),
    .A(_00581_),
    .Y(_00646_));
 sg13g2_inv_1 _06840_ (.Y(_00647_),
    .A(_00538_));
 sg13g2_a21oi_2 _06841_ (.B1(_00647_),
    .Y(_00648_),
    .A2(_00241_),
    .A1(_00536_));
 sg13g2_buf_1 _06842_ (.A(_00224_),
    .X(_00649_));
 sg13g2_nor2_1 _06843_ (.A(net49),
    .B(_05612_),
    .Y(_00650_));
 sg13g2_xnor2_1 _06844_ (.Y(_00651_),
    .A(_00244_),
    .B(_00650_));
 sg13g2_a21oi_1 _06845_ (.A1(_00328_),
    .A2(_00283_),
    .Y(_00652_),
    .B1(_00324_));
 sg13g2_xnor2_1 _06846_ (.Y(_00653_),
    .A(_00651_),
    .B(_00652_));
 sg13g2_xnor2_1 _06847_ (.Y(_00654_),
    .A(_00246_),
    .B(_00653_));
 sg13g2_nor2_1 _06848_ (.A(net51),
    .B(_00274_),
    .Y(_00655_));
 sg13g2_nand2_1 _06849_ (.Y(_00656_),
    .A(_00472_),
    .B(net65));
 sg13g2_nor2_1 _06850_ (.A(_00327_),
    .B(_00656_),
    .Y(_00657_));
 sg13g2_nor2_1 _06851_ (.A(net57),
    .B(_00369_),
    .Y(_00658_));
 sg13g2_inv_1 _06852_ (.Y(_00659_),
    .A(_00658_));
 sg13g2_nand2_1 _06853_ (.Y(_00660_),
    .A(_00659_),
    .B(_00323_));
 sg13g2_nand2b_1 _06854_ (.Y(_00661_),
    .B(_00660_),
    .A_N(_00657_));
 sg13g2_xnor2_1 _06855_ (.Y(_00662_),
    .A(_00655_),
    .B(_00661_));
 sg13g2_inv_1 _06856_ (.Y(_00663_),
    .A(_00464_));
 sg13g2_a21oi_1 _06857_ (.A1(_00466_),
    .A2(_00370_),
    .Y(_00664_),
    .B1(_00663_));
 sg13g2_nor2_1 _06858_ (.A(_00386_),
    .B(_00435_),
    .Y(_00665_));
 sg13g2_nand2_1 _06859_ (.Y(_00666_),
    .A(_00381_),
    .B(_00665_));
 sg13g2_nor2b_1 _06860_ (.A(_00435_),
    .B_N(_00438_),
    .Y(_00667_));
 sg13g2_buf_8 _06861_ (.A(\r1[7] ),
    .X(_00668_));
 sg13g2_nand3_1 _06862_ (.B(_00668_),
    .C(net74),
    .A(_00429_),
    .Y(_00669_));
 sg13g2_nor2b_1 _06863_ (.A(_00667_),
    .B_N(_00669_),
    .Y(_00670_));
 sg13g2_nand2_1 _06864_ (.Y(_00671_),
    .A(_00666_),
    .B(_00670_));
 sg13g2_buf_1 _06865_ (.A(\r1[8] ),
    .X(_00672_));
 sg13g2_xnor2_1 _06866_ (.Y(_00673_),
    .A(_00672_),
    .B(_00228_));
 sg13g2_buf_2 _06867_ (.A(_00673_),
    .X(_00674_));
 sg13g2_inv_1 _06868_ (.Y(_00675_),
    .A(_00674_));
 sg13g2_nand2_1 _06869_ (.Y(_00676_),
    .A(_00671_),
    .B(_00675_));
 sg13g2_nand3_1 _06870_ (.B(_00670_),
    .C(_00674_),
    .A(_00666_),
    .Y(_00677_));
 sg13g2_buf_8 _06871_ (.A(\r2[9] ),
    .X(_00678_));
 sg13g2_nand3_1 _06872_ (.B(_00677_),
    .C(_00678_),
    .A(_00676_),
    .Y(_00679_));
 sg13g2_buf_1 _06873_ (.A(_00679_),
    .X(_00680_));
 sg13g2_nand2_1 _06874_ (.Y(_00681_),
    .A(_00671_),
    .B(_00674_));
 sg13g2_nand3_1 _06875_ (.B(_00670_),
    .C(_00675_),
    .A(_00666_),
    .Y(_00682_));
 sg13g2_inv_1 _06876_ (.Y(_00683_),
    .A(_00678_));
 sg13g2_nand3_1 _06877_ (.B(_00682_),
    .C(_00683_),
    .A(_00681_),
    .Y(_00684_));
 sg13g2_nand2_1 _06878_ (.Y(_00685_),
    .A(_00680_),
    .B(_00684_));
 sg13g2_nand2_1 _06879_ (.Y(_00686_),
    .A(_00446_),
    .B(_00050_));
 sg13g2_inv_1 _06880_ (.Y(_00687_),
    .A(_00686_));
 sg13g2_nand2_1 _06881_ (.Y(_00688_),
    .A(_00685_),
    .B(_00687_));
 sg13g2_nand3_1 _06882_ (.B(_00684_),
    .C(_00686_),
    .A(_00680_),
    .Y(_00689_));
 sg13g2_nand2_1 _06883_ (.Y(_00690_),
    .A(_00688_),
    .B(_00689_));
 sg13g2_buf_2 _06884_ (.A(_00690_),
    .X(_00691_));
 sg13g2_xnor2_1 _06885_ (.Y(_00692_),
    .A(_00395_),
    .B(_00398_));
 sg13g2_nand2_1 _06886_ (.Y(_00693_),
    .A(_00456_),
    .B(_00692_));
 sg13g2_inv_1 _06887_ (.Y(_00694_),
    .A(_00693_));
 sg13g2_nand2_1 _06888_ (.Y(_00695_),
    .A(_00405_),
    .B(_00694_));
 sg13g2_nand2_1 _06889_ (.Y(_00696_),
    .A(_00399_),
    .B(_00454_));
 sg13g2_nand2b_1 _06890_ (.Y(_00697_),
    .B(_00696_),
    .A_N(_00453_));
 sg13g2_nand2_1 _06891_ (.Y(_00698_),
    .A(_00695_),
    .B(_00697_));
 sg13g2_nand2b_1 _06892_ (.Y(_00699_),
    .B(_00698_),
    .A_N(_00691_));
 sg13g2_nand3_1 _06893_ (.B(_00691_),
    .C(_00697_),
    .A(_00695_),
    .Y(_00700_));
 sg13g2_nand2_1 _06894_ (.Y(_00701_),
    .A(_00699_),
    .B(_00700_));
 sg13g2_buf_8 _06895_ (.A(_00701_),
    .X(_00702_));
 sg13g2_nor2_1 _06896_ (.A(_00518_),
    .B(_00702_),
    .Y(_00703_));
 sg13g2_nand2_1 _06897_ (.Y(_00704_),
    .A(_00703_),
    .B(_00463_));
 sg13g2_nand3_1 _06898_ (.B(_00700_),
    .C(_05562_),
    .A(_00699_),
    .Y(_00705_));
 sg13g2_inv_2 _06899_ (.Y(_00706_),
    .A(_00462_));
 sg13g2_nand2_1 _06900_ (.Y(_00707_),
    .A(_00706_),
    .B(net68));
 sg13g2_nand2_1 _06901_ (.Y(_00708_),
    .A(_00705_),
    .B(_00707_));
 sg13g2_nand2_1 _06902_ (.Y(_00709_),
    .A(_00704_),
    .B(_00708_));
 sg13g2_inv_1 _06903_ (.Y(_00710_),
    .A(_00407_));
 sg13g2_nor2_1 _06904_ (.A(net75),
    .B(_00710_),
    .Y(_00711_));
 sg13g2_nand2_1 _06905_ (.Y(_00712_),
    .A(_00709_),
    .B(_00711_));
 sg13g2_inv_1 _06906_ (.Y(_00713_),
    .A(_00711_));
 sg13g2_nand3_1 _06907_ (.B(_00708_),
    .C(_00713_),
    .A(_00704_),
    .Y(_00714_));
 sg13g2_nand2_1 _06908_ (.Y(_00715_),
    .A(_00712_),
    .B(_00714_));
 sg13g2_nand2b_1 _06909_ (.Y(_00716_),
    .B(_00715_),
    .A_N(_00664_));
 sg13g2_nand3_1 _06910_ (.B(_00714_),
    .C(_00664_),
    .A(_00712_),
    .Y(_00717_));
 sg13g2_nand2_1 _06911_ (.Y(_00718_),
    .A(_00716_),
    .B(_00717_));
 sg13g2_nand2b_1 _06912_ (.Y(_00719_),
    .B(_00718_),
    .A_N(_00662_));
 sg13g2_nand3_1 _06913_ (.B(_00717_),
    .C(_00662_),
    .A(_00716_),
    .Y(_00720_));
 sg13g2_nand2_1 _06914_ (.Y(_00721_),
    .A(_00719_),
    .B(_00720_));
 sg13g2_inv_1 _06915_ (.Y(_00722_),
    .A(_00482_));
 sg13g2_a21oi_1 _06916_ (.A1(_00480_),
    .A2(_00330_),
    .Y(_00723_),
    .B1(_00722_));
 sg13g2_nand2_1 _06917_ (.Y(_00724_),
    .A(_00721_),
    .B(_00723_));
 sg13g2_inv_1 _06918_ (.Y(_00725_),
    .A(_00723_));
 sg13g2_nand3_1 _06919_ (.B(_00720_),
    .C(_00725_),
    .A(_00719_),
    .Y(_00726_));
 sg13g2_nand2_1 _06920_ (.Y(_00727_),
    .A(_00724_),
    .B(_00726_));
 sg13g2_nand2b_1 _06921_ (.Y(_00728_),
    .B(_00727_),
    .A_N(_00654_));
 sg13g2_nand3_1 _06922_ (.B(_00726_),
    .C(_00654_),
    .A(_00724_),
    .Y(_00729_));
 sg13g2_nand2_1 _06923_ (.Y(_00730_),
    .A(_00728_),
    .B(_00729_));
 sg13g2_inv_1 _06924_ (.Y(_00731_),
    .A(_00507_));
 sg13g2_a21oi_1 _06925_ (.A1(_00505_),
    .A2(_00282_),
    .Y(_00732_),
    .B1(_00731_));
 sg13g2_nand2_1 _06926_ (.Y(_00733_),
    .A(_00730_),
    .B(_00732_));
 sg13g2_inv_1 _06927_ (.Y(_00734_),
    .A(_00732_));
 sg13g2_nand3_1 _06928_ (.B(_00729_),
    .C(_00734_),
    .A(_00728_),
    .Y(_00735_));
 sg13g2_nand2_1 _06929_ (.Y(_00736_),
    .A(_00733_),
    .B(_00735_));
 sg13g2_nor2b_1 _06930_ (.A(_00280_),
    .B_N(_00247_),
    .Y(_00737_));
 sg13g2_a21oi_1 _06931_ (.A1(_00281_),
    .A2(_00235_),
    .Y(_00738_),
    .B1(_00737_));
 sg13g2_nand2_1 _06932_ (.Y(_00739_),
    .A(_00736_),
    .B(_00738_));
 sg13g2_inv_1 _06933_ (.Y(_00740_),
    .A(_00738_));
 sg13g2_nand3_1 _06934_ (.B(_00735_),
    .C(_00740_),
    .A(_00733_),
    .Y(_00741_));
 sg13g2_nand2_1 _06935_ (.Y(_00742_),
    .A(_00739_),
    .B(_00741_));
 sg13g2_nor2_1 _06936_ (.A(_00648_),
    .B(_00742_),
    .Y(_00743_));
 sg13g2_nor2b_1 _06937_ (.A(_00743_),
    .B_N(_00583_),
    .Y(_00744_));
 sg13g2_nand2_1 _06938_ (.Y(_00745_),
    .A(_00742_),
    .B(_00648_));
 sg13g2_inv_1 _06939_ (.Y(_00746_),
    .A(_00745_));
 sg13g2_a21oi_1 _06940_ (.A1(_00646_),
    .A2(_00744_),
    .Y(_00747_),
    .B1(_00746_));
 sg13g2_nand2_1 _06941_ (.Y(_00748_),
    .A(_00212_),
    .B(net50));
 sg13g2_nor2b_1 _06942_ (.A(_00748_),
    .B_N(_00242_),
    .Y(_00749_));
 sg13g2_nor2_1 _06943_ (.A(net49),
    .B(_00274_),
    .Y(_00750_));
 sg13g2_xor2_1 _06944_ (.B(_00750_),
    .A(_00748_),
    .X(_00751_));
 sg13g2_a21oi_1 _06945_ (.A1(_00660_),
    .A2(_00655_),
    .Y(_00752_),
    .B1(_00657_));
 sg13g2_xnor2_1 _06946_ (.Y(_00753_),
    .A(_00751_),
    .B(_00752_));
 sg13g2_xnor2_1 _06947_ (.Y(_00754_),
    .A(_00749_),
    .B(_00753_));
 sg13g2_inv_1 _06948_ (.Y(_00755_),
    .A(_00704_));
 sg13g2_a21oi_1 _06949_ (.A1(_00708_),
    .A2(_00711_),
    .Y(_00756_),
    .B1(_00755_));
 sg13g2_nor2_2 _06950_ (.A(_00459_),
    .B(_00691_),
    .Y(_00757_));
 sg13g2_nand2_1 _06951_ (.Y(_00758_),
    .A(_00757_),
    .B(_00419_));
 sg13g2_nand2_1 _06952_ (.Y(_00759_),
    .A(_00689_),
    .B(_00454_));
 sg13g2_nand2_1 _06953_ (.Y(_00760_),
    .A(_00759_),
    .B(_00688_));
 sg13g2_nand2_1 _06954_ (.Y(_00761_),
    .A(_00758_),
    .B(_00760_));
 sg13g2_inv_1 _06955_ (.Y(_00762_),
    .A(_05606_));
 sg13g2_a21oi_1 _06956_ (.A1(_05604_),
    .A2(_05581_),
    .Y(_00763_),
    .B1(_00762_));
 sg13g2_inv_1 _06957_ (.Y(_00764_),
    .A(_00763_));
 sg13g2_a21oi_1 _06958_ (.A1(_00422_),
    .A2(_00764_),
    .Y(_00765_),
    .B1(_00417_));
 sg13g2_nand2_1 _06959_ (.Y(_00766_),
    .A(_00757_),
    .B(_00413_));
 sg13g2_nor2_1 _06960_ (.A(_00765_),
    .B(_00766_),
    .Y(_00767_));
 sg13g2_nor2_1 _06961_ (.A(_00761_),
    .B(_00767_),
    .Y(_00768_));
 sg13g2_inv_1 _06962_ (.Y(_00769_),
    .A(_05607_));
 sg13g2_nand2_1 _06963_ (.Y(_00770_),
    .A(_00769_),
    .B(_05614_));
 sg13g2_nor3_1 _06964_ (.A(_00770_),
    .B(_00421_),
    .C(_00310_),
    .Y(_00771_));
 sg13g2_nand4_1 _06965_ (.B(_00771_),
    .C(_00413_),
    .A(_00757_),
    .Y(_00772_),
    .D(_05580_));
 sg13g2_nand2_1 _06966_ (.Y(_00773_),
    .A(_00768_),
    .B(_00772_));
 sg13g2_nor2_2 _06967_ (.A(_00674_),
    .B(_00435_),
    .Y(_00774_));
 sg13g2_nor2_1 _06968_ (.A(_00669_),
    .B(_00674_),
    .Y(_00775_));
 sg13g2_inv_1 _06969_ (.Y(_00776_),
    .A(_00042_));
 sg13g2_nand2_1 _06970_ (.Y(_00777_),
    .A(_00228_),
    .B(_00776_));
 sg13g2_nor2b_1 _06971_ (.A(_00775_),
    .B_N(_00777_),
    .Y(_00778_));
 sg13g2_inv_1 _06972_ (.Y(_00779_),
    .A(_00778_));
 sg13g2_a21oi_1 _06973_ (.A1(_00774_),
    .A2(_00441_),
    .Y(_00780_),
    .B1(_00779_));
 sg13g2_nand3_1 _06974_ (.B(_00436_),
    .C(_00345_),
    .A(_00774_),
    .Y(_00781_));
 sg13g2_nand2_1 _06975_ (.Y(_00782_),
    .A(_00780_),
    .B(_00781_));
 sg13g2_nand2_1 _06976_ (.Y(_00783_),
    .A(net74),
    .B(_00040_));
 sg13g2_inv_1 _06977_ (.Y(_00784_),
    .A(_00040_));
 sg13g2_nand3_1 _06978_ (.B(_03629_),
    .C(_00784_),
    .A(_00426_),
    .Y(_00785_));
 sg13g2_buf_2 _06979_ (.A(_00785_),
    .X(_00786_));
 sg13g2_nand2_2 _06980_ (.Y(_00787_),
    .A(_00783_),
    .B(_00786_));
 sg13g2_inv_1 _06981_ (.Y(_00788_),
    .A(_00787_));
 sg13g2_nand2_1 _06982_ (.Y(_00789_),
    .A(_00782_),
    .B(_00788_));
 sg13g2_nand3_1 _06983_ (.B(_00781_),
    .C(_00787_),
    .A(_00780_),
    .Y(_00790_));
 sg13g2_nand2_1 _06984_ (.Y(_00791_),
    .A(_00789_),
    .B(_00790_));
 sg13g2_buf_1 _06985_ (.A(\r2[10] ),
    .X(_00792_));
 sg13g2_inv_1 _06986_ (.Y(_00793_),
    .A(_00792_));
 sg13g2_nand2_1 _06987_ (.Y(_00794_),
    .A(_00791_),
    .B(_00793_));
 sg13g2_nand3_1 _06988_ (.B(_00790_),
    .C(_00792_),
    .A(_00789_),
    .Y(_00795_));
 sg13g2_nand2_1 _06989_ (.Y(_00796_),
    .A(_00794_),
    .B(_00795_));
 sg13g2_nand2b_1 _06990_ (.Y(_00797_),
    .B(_00796_),
    .A_N(_00680_));
 sg13g2_nand3_1 _06991_ (.B(_00795_),
    .C(_00680_),
    .A(_00794_),
    .Y(_00798_));
 sg13g2_nand2_1 _06992_ (.Y(_00799_),
    .A(_00797_),
    .B(_00798_));
 sg13g2_buf_8 _06993_ (.A(_00799_),
    .X(_00800_));
 sg13g2_inv_1 _06994_ (.Y(_00801_),
    .A(_00800_));
 sg13g2_nand2_1 _06995_ (.Y(_00802_),
    .A(_00773_),
    .B(_00801_));
 sg13g2_nand3_1 _06996_ (.B(_00800_),
    .C(_00772_),
    .A(_00768_),
    .Y(_00803_));
 sg13g2_buf_8 _06997_ (.A(_00803_),
    .X(_00804_));
 sg13g2_nand2_2 _06998_ (.Y(_00805_),
    .A(_00802_),
    .B(_00804_));
 sg13g2_nor2_1 _06999_ (.A(net101),
    .B(_00805_),
    .Y(_00806_));
 sg13g2_nand2_1 _07000_ (.Y(_00807_),
    .A(_00806_),
    .B(_00703_));
 sg13g2_nand3_1 _07001_ (.B(_00804_),
    .C(_05562_),
    .A(_00802_),
    .Y(_00808_));
 sg13g2_inv_1 _07002_ (.Y(_00809_),
    .A(_00703_));
 sg13g2_nand2_1 _07003_ (.Y(_00810_),
    .A(_00808_),
    .B(_00809_));
 sg13g2_nand2_1 _07004_ (.Y(_00811_),
    .A(_00807_),
    .B(_00810_));
 sg13g2_nor2_1 _07005_ (.A(_00333_),
    .B(_00462_),
    .Y(_00812_));
 sg13g2_nand2_1 _07006_ (.Y(_00813_),
    .A(_00811_),
    .B(_00812_));
 sg13g2_inv_1 _07007_ (.Y(_00814_),
    .A(_00812_));
 sg13g2_nand3_1 _07008_ (.B(_00810_),
    .C(_00814_),
    .A(_00807_),
    .Y(_00815_));
 sg13g2_nand2_1 _07009_ (.Y(_00816_),
    .A(_00813_),
    .B(_00815_));
 sg13g2_nand2b_1 _07010_ (.Y(_00817_),
    .B(_00816_),
    .A_N(_00756_));
 sg13g2_nand3_1 _07011_ (.B(_00815_),
    .C(_00756_),
    .A(_00813_),
    .Y(_00818_));
 sg13g2_buf_1 _07012_ (.A(_00818_),
    .X(_00819_));
 sg13g2_nand2_1 _07013_ (.Y(_00820_),
    .A(_00817_),
    .B(_00819_));
 sg13g2_nor2_1 _07014_ (.A(_00207_),
    .B(_00321_),
    .Y(_00821_));
 sg13g2_nand2_1 _07015_ (.Y(_00822_),
    .A(_00407_),
    .B(net65));
 sg13g2_nand2_1 _07016_ (.Y(_00823_),
    .A(_00407_),
    .B(net71));
 sg13g2_nand2_1 _07017_ (.Y(_00824_),
    .A(_00823_),
    .B(_00656_));
 sg13g2_o21ai_1 _07018_ (.B1(_00824_),
    .Y(_00825_),
    .A1(_00822_),
    .A2(_00659_));
 sg13g2_xnor2_1 _07019_ (.Y(_00826_),
    .A(_00821_),
    .B(_00825_));
 sg13g2_inv_1 _07020_ (.Y(_00827_),
    .A(_00826_));
 sg13g2_nand2_1 _07021_ (.Y(_00828_),
    .A(_00820_),
    .B(_00827_));
 sg13g2_nand3_1 _07022_ (.B(_00819_),
    .C(_00826_),
    .A(_00817_),
    .Y(_00829_));
 sg13g2_inv_1 _07023_ (.Y(_00830_),
    .A(_00716_));
 sg13g2_a21oi_1 _07024_ (.A1(_00717_),
    .A2(_00662_),
    .Y(_00831_),
    .B1(_00830_));
 sg13g2_inv_1 _07025_ (.Y(_00832_),
    .A(_00831_));
 sg13g2_nand3_1 _07026_ (.B(_00829_),
    .C(_00832_),
    .A(_00828_),
    .Y(_00833_));
 sg13g2_nand2_1 _07027_ (.Y(_00834_),
    .A(_00820_),
    .B(_00826_));
 sg13g2_nand3_1 _07028_ (.B(_00819_),
    .C(_00827_),
    .A(_00817_),
    .Y(_00835_));
 sg13g2_nand3_1 _07029_ (.B(_00835_),
    .C(_00831_),
    .A(_00834_),
    .Y(_00836_));
 sg13g2_nand2_1 _07030_ (.Y(_00837_),
    .A(_00833_),
    .B(_00836_));
 sg13g2_nand2b_1 _07031_ (.Y(_00838_),
    .B(_00837_),
    .A_N(_00754_));
 sg13g2_nand3_1 _07032_ (.B(_00836_),
    .C(_00754_),
    .A(_00833_),
    .Y(_00839_));
 sg13g2_nand2_1 _07033_ (.Y(_00840_),
    .A(_00838_),
    .B(_00839_));
 sg13g2_inv_1 _07034_ (.Y(_00841_),
    .A(_00726_));
 sg13g2_a21oi_1 _07035_ (.A1(_00724_),
    .A2(_00654_),
    .Y(_00842_),
    .B1(_00841_));
 sg13g2_nand2_1 _07036_ (.Y(_00843_),
    .A(_00840_),
    .B(_00842_));
 sg13g2_inv_1 _07037_ (.Y(_00844_),
    .A(_00842_));
 sg13g2_nand3_1 _07038_ (.B(_00839_),
    .C(_00844_),
    .A(_00838_),
    .Y(_00845_));
 sg13g2_nand2_1 _07039_ (.Y(_00846_),
    .A(_00843_),
    .B(_00845_));
 sg13g2_nor2_1 _07040_ (.A(_00651_),
    .B(_00652_),
    .Y(_00847_));
 sg13g2_nor2_1 _07041_ (.A(_00245_),
    .B(_00653_),
    .Y(_00848_));
 sg13g2_nor2_1 _07042_ (.A(_00847_),
    .B(_00848_),
    .Y(_00849_));
 sg13g2_nand2_1 _07043_ (.Y(_00850_),
    .A(_00846_),
    .B(_00849_));
 sg13g2_inv_1 _07044_ (.Y(_00851_),
    .A(_00849_));
 sg13g2_nand3_1 _07045_ (.B(_00845_),
    .C(_00851_),
    .A(_00843_),
    .Y(_00852_));
 sg13g2_nand2_1 _07046_ (.Y(_00853_),
    .A(_00850_),
    .B(_00852_));
 sg13g2_inv_1 _07047_ (.Y(_00854_),
    .A(_00735_));
 sg13g2_a21oi_1 _07048_ (.A1(_00733_),
    .A2(_00740_),
    .Y(_00855_),
    .B1(_00854_));
 sg13g2_nand2_1 _07049_ (.Y(_00856_),
    .A(_00853_),
    .B(_00855_));
 sg13g2_inv_1 _07050_ (.Y(_00857_),
    .A(_00855_));
 sg13g2_nand3_1 _07051_ (.B(_00852_),
    .C(_00857_),
    .A(_00850_),
    .Y(_00858_));
 sg13g2_nand2_1 _07052_ (.Y(_00859_),
    .A(_00856_),
    .B(_00858_));
 sg13g2_inv_1 _07053_ (.Y(_00860_),
    .A(_00845_));
 sg13g2_a21oi_1 _07054_ (.A1(_00843_),
    .A2(_00851_),
    .Y(_00861_),
    .B1(_00860_));
 sg13g2_inv_1 _07055_ (.Y(_00862_),
    .A(_00861_));
 sg13g2_a21oi_1 _07056_ (.A1(_00834_),
    .A2(_00835_),
    .Y(_00863_),
    .B1(_00831_));
 sg13g2_a21oi_1 _07057_ (.A1(_00836_),
    .A2(_00754_),
    .Y(_00864_),
    .B1(_00863_));
 sg13g2_a21oi_1 _07058_ (.A1(_00813_),
    .A2(_00815_),
    .Y(_00865_),
    .B1(_00756_));
 sg13g2_a21oi_1 _07059_ (.A1(_00819_),
    .A2(_00826_),
    .Y(_00866_),
    .B1(_00865_));
 sg13g2_nand3_1 _07060_ (.B(_00804_),
    .C(net68),
    .A(_00802_),
    .Y(_00867_));
 sg13g2_nor2_1 _07061_ (.A(_00705_),
    .B(_00867_),
    .Y(_00868_));
 sg13g2_a21oi_1 _07062_ (.A1(_00810_),
    .A2(_00812_),
    .Y(_00869_),
    .B1(_00868_));
 sg13g2_nor2_1 _07063_ (.A(_00787_),
    .B(_00674_),
    .Y(_00870_));
 sg13g2_nand2_1 _07064_ (.Y(_00871_),
    .A(_00671_),
    .B(_00870_));
 sg13g2_o21ai_1 _07065_ (.B1(_00786_),
    .Y(_00872_),
    .A1(_00777_),
    .A2(_00787_));
 sg13g2_buf_1 _07066_ (.A(_00872_),
    .X(_00873_));
 sg13g2_inv_1 _07067_ (.Y(_00874_),
    .A(_00873_));
 sg13g2_nand2_1 _07068_ (.Y(_00875_),
    .A(_00871_),
    .B(_00874_));
 sg13g2_buf_1 _07069_ (.A(_00041_),
    .X(_00876_));
 sg13g2_inv_1 _07070_ (.Y(_00877_),
    .A(_00876_));
 sg13g2_nand2_1 _07071_ (.Y(_00878_),
    .A(_00875_),
    .B(_00877_));
 sg13g2_nand3_1 _07072_ (.B(_00876_),
    .C(_00874_),
    .A(_00871_),
    .Y(_00879_));
 sg13g2_buf_1 _07073_ (.A(\r2[11] ),
    .X(_00880_));
 sg13g2_inv_2 _07074_ (.Y(_00881_),
    .A(_00880_));
 sg13g2_nand3_1 _07075_ (.B(_00879_),
    .C(_00881_),
    .A(_00878_),
    .Y(_00882_));
 sg13g2_buf_1 _07076_ (.A(_00882_),
    .X(_00883_));
 sg13g2_nand2_1 _07077_ (.Y(_00884_),
    .A(_00875_),
    .B(_00876_));
 sg13g2_nand3_1 _07078_ (.B(_00877_),
    .C(_00874_),
    .A(_00871_),
    .Y(_00885_));
 sg13g2_nand3_1 _07079_ (.B(_00885_),
    .C(_00880_),
    .A(_00884_),
    .Y(_00886_));
 sg13g2_nand2_1 _07080_ (.Y(_00887_),
    .A(_00883_),
    .B(_00886_));
 sg13g2_nand2_1 _07081_ (.Y(_00888_),
    .A(_00887_),
    .B(_00794_));
 sg13g2_inv_1 _07082_ (.Y(_00889_),
    .A(_00794_));
 sg13g2_nand3_1 _07083_ (.B(_00886_),
    .C(_00889_),
    .A(_00883_),
    .Y(_00890_));
 sg13g2_nand2_2 _07084_ (.Y(_00891_),
    .A(_00888_),
    .B(_00890_));
 sg13g2_nand2_1 _07085_ (.Y(_00892_),
    .A(_00797_),
    .B(_00689_));
 sg13g2_nand2_1 _07086_ (.Y(_00893_),
    .A(_00892_),
    .B(_00798_));
 sg13g2_inv_1 _07087_ (.Y(_00894_),
    .A(_00893_));
 sg13g2_nor3_1 _07088_ (.A(_00691_),
    .B(_00697_),
    .C(_00800_),
    .Y(_00895_));
 sg13g2_nor2_1 _07089_ (.A(_00894_),
    .B(_00895_),
    .Y(_00896_));
 sg13g2_nor3_1 _07090_ (.A(_00691_),
    .B(_00693_),
    .C(_00800_),
    .Y(_00897_));
 sg13g2_nand2_1 _07091_ (.Y(_00898_),
    .A(_00897_),
    .B(_00405_));
 sg13g2_nand2_1 _07092_ (.Y(_00899_),
    .A(_00896_),
    .B(_00898_));
 sg13g2_nand2b_1 _07093_ (.Y(_00900_),
    .B(_00899_),
    .A_N(_00891_));
 sg13g2_nand3_1 _07094_ (.B(_00898_),
    .C(_00891_),
    .A(_00896_),
    .Y(_00901_));
 sg13g2_nand2_1 _07095_ (.Y(_00902_),
    .A(_00900_),
    .B(_00901_));
 sg13g2_buf_8 _07096_ (.A(_00902_),
    .X(_00903_));
 sg13g2_nor2_1 _07097_ (.A(net62),
    .B(_00903_),
    .Y(_00904_));
 sg13g2_nand2_1 _07098_ (.Y(_00905_),
    .A(_00806_),
    .B(_00904_));
 sg13g2_nand3_1 _07099_ (.B(_00901_),
    .C(_05562_),
    .A(_00900_),
    .Y(_00906_));
 sg13g2_nand2_1 _07100_ (.Y(_00907_),
    .A(_00867_),
    .B(_00906_));
 sg13g2_nand2_1 _07101_ (.Y(_00908_),
    .A(_00905_),
    .B(_00907_));
 sg13g2_nor2_1 _07102_ (.A(net75),
    .B(_00702_),
    .Y(_00909_));
 sg13g2_nand2_1 _07103_ (.Y(_00910_),
    .A(_00908_),
    .B(_00909_));
 sg13g2_inv_1 _07104_ (.Y(_00911_),
    .A(_00909_));
 sg13g2_nand3_1 _07105_ (.B(_00907_),
    .C(_00911_),
    .A(_00905_),
    .Y(_00912_));
 sg13g2_nand2_1 _07106_ (.Y(_00913_),
    .A(_00910_),
    .B(_00912_));
 sg13g2_nand2b_1 _07107_ (.Y(_00914_),
    .B(_00913_),
    .A_N(_00869_));
 sg13g2_nand3_1 _07108_ (.B(_00869_),
    .C(_00912_),
    .A(_00910_),
    .Y(_00915_));
 sg13g2_nand2_1 _07109_ (.Y(_00916_),
    .A(_00914_),
    .B(_00915_));
 sg13g2_nor2_1 _07110_ (.A(_00207_),
    .B(_00369_),
    .Y(_00917_));
 sg13g2_nand2_1 _07111_ (.Y(_00918_),
    .A(_00706_),
    .B(net65));
 sg13g2_nor2_1 _07112_ (.A(_00823_),
    .B(_00918_),
    .Y(_00919_));
 sg13g2_nor2_1 _07113_ (.A(net57),
    .B(_00462_),
    .Y(_00920_));
 sg13g2_inv_1 _07114_ (.Y(_00921_),
    .A(_00920_));
 sg13g2_nand2_1 _07115_ (.Y(_00922_),
    .A(_00921_),
    .B(_00822_));
 sg13g2_nand2b_1 _07116_ (.Y(_00923_),
    .B(_00922_),
    .A_N(_00919_));
 sg13g2_xor2_1 _07117_ (.B(_00923_),
    .A(_00917_),
    .X(_00924_));
 sg13g2_inv_1 _07118_ (.Y(_00925_),
    .A(_00924_));
 sg13g2_nand2_1 _07119_ (.Y(_00926_),
    .A(_00916_),
    .B(_00925_));
 sg13g2_nand3_1 _07120_ (.B(_00915_),
    .C(_00924_),
    .A(_00914_),
    .Y(_00927_));
 sg13g2_nand2_1 _07121_ (.Y(_00928_),
    .A(_00926_),
    .B(_00927_));
 sg13g2_nand2b_1 _07122_ (.Y(_00929_),
    .B(_00928_),
    .A_N(_00866_));
 sg13g2_nand3_1 _07123_ (.B(_00927_),
    .C(_00866_),
    .A(_00926_),
    .Y(_00930_));
 sg13g2_nand2_1 _07124_ (.Y(_00931_),
    .A(_00929_),
    .B(_00930_));
 sg13g2_inv_1 _07125_ (.Y(_00932_),
    .A(_00650_));
 sg13g2_nor2_1 _07126_ (.A(net45),
    .B(_00274_),
    .Y(_00933_));
 sg13g2_inv_1 _07127_ (.Y(_00934_),
    .A(_00933_));
 sg13g2_nor2_1 _07128_ (.A(_00932_),
    .B(_00934_),
    .Y(_00935_));
 sg13g2_inv_1 _07129_ (.Y(_00936_),
    .A(_00935_));
 sg13g2_nor2_1 _07130_ (.A(net49),
    .B(_00321_),
    .Y(_00937_));
 sg13g2_xnor2_1 _07131_ (.Y(_00938_),
    .A(_00934_),
    .B(_00937_));
 sg13g2_nor2_1 _07132_ (.A(_00659_),
    .B(_00822_),
    .Y(_00939_));
 sg13g2_a21oi_1 _07133_ (.A1(_00824_),
    .A2(_00821_),
    .Y(_00940_),
    .B1(_00939_));
 sg13g2_xnor2_1 _07134_ (.Y(_00941_),
    .A(_00938_),
    .B(_00940_));
 sg13g2_xnor2_1 _07135_ (.Y(_00942_),
    .A(_00936_),
    .B(_00941_));
 sg13g2_nand2_1 _07136_ (.Y(_00943_),
    .A(_00931_),
    .B(_00942_));
 sg13g2_inv_1 _07137_ (.Y(_00944_),
    .A(_00942_));
 sg13g2_nand3_1 _07138_ (.B(_00930_),
    .C(_00944_),
    .A(_00929_),
    .Y(_00945_));
 sg13g2_nand2_1 _07139_ (.Y(_00946_),
    .A(_00943_),
    .B(_00945_));
 sg13g2_nand2b_1 _07140_ (.Y(_00947_),
    .B(_00946_),
    .A_N(_00864_));
 sg13g2_nand3_1 _07141_ (.B(_00945_),
    .C(_00864_),
    .A(_00943_),
    .Y(_00948_));
 sg13g2_nor2_1 _07142_ (.A(_00751_),
    .B(_00752_),
    .Y(_00949_));
 sg13g2_nand2b_1 _07143_ (.Y(_00950_),
    .B(_00749_),
    .A_N(_00753_));
 sg13g2_nor2b_1 _07144_ (.A(_00949_),
    .B_N(_00950_),
    .Y(_00951_));
 sg13g2_inv_1 _07145_ (.Y(_00952_),
    .A(_00951_));
 sg13g2_nand3_1 _07146_ (.B(_00948_),
    .C(_00952_),
    .A(_00947_),
    .Y(_00953_));
 sg13g2_nand2_1 _07147_ (.Y(_00954_),
    .A(_00947_),
    .B(_00948_));
 sg13g2_nand2_1 _07148_ (.Y(_00955_),
    .A(_00954_),
    .B(_00951_));
 sg13g2_nand3_1 _07149_ (.B(_00953_),
    .C(_00955_),
    .A(_00862_),
    .Y(_00956_));
 sg13g2_buf_1 _07150_ (.A(_00956_),
    .X(_00957_));
 sg13g2_nand2_1 _07151_ (.Y(_00958_),
    .A(_00955_),
    .B(_00953_));
 sg13g2_nand2_1 _07152_ (.Y(_00959_),
    .A(_00958_),
    .B(_00861_));
 sg13g2_nand2_1 _07153_ (.Y(_00960_),
    .A(_00957_),
    .B(_00959_));
 sg13g2_nor2_1 _07154_ (.A(_00859_),
    .B(_00960_),
    .Y(_00961_));
 sg13g2_nand2_1 _07155_ (.Y(_00962_),
    .A(_00747_),
    .B(_00961_));
 sg13g2_inv_1 _07156_ (.Y(_00963_),
    .A(_00858_));
 sg13g2_inv_1 _07157_ (.Y(_00964_),
    .A(_00957_));
 sg13g2_o21ai_1 _07158_ (.B1(_00959_),
    .Y(_00965_),
    .A1(_00963_),
    .A2(_00964_));
 sg13g2_nand2_1 _07159_ (.Y(_00966_),
    .A(_00962_),
    .B(_00965_));
 sg13g2_inv_1 _07160_ (.Y(_00967_),
    .A(_00947_));
 sg13g2_a21oi_1 _07161_ (.A1(_00948_),
    .A2(_00952_),
    .Y(_00968_),
    .B1(_00967_));
 sg13g2_inv_1 _07162_ (.Y(_00969_),
    .A(_00929_));
 sg13g2_a21oi_1 _07163_ (.A1(_00930_),
    .A2(_00942_),
    .Y(_00970_),
    .B1(_00969_));
 sg13g2_inv_1 _07164_ (.Y(_00971_),
    .A(_00914_));
 sg13g2_a21oi_1 _07165_ (.A1(_00915_),
    .A2(_00925_),
    .Y(_00972_),
    .B1(_00971_));
 sg13g2_a22oi_1 _07166_ (.Y(_00973_),
    .B1(_00909_),
    .B2(_00907_),
    .A2(_00806_),
    .A1(_00904_));
 sg13g2_nand3_1 _07167_ (.B(_00786_),
    .C(_00876_),
    .A(_00783_),
    .Y(_00974_));
 sg13g2_buf_2 _07168_ (.A(_00974_),
    .X(_00975_));
 sg13g2_inv_1 _07169_ (.Y(_00976_),
    .A(_00975_));
 sg13g2_nand3_1 _07170_ (.B(_00976_),
    .C(_00774_),
    .A(_00443_),
    .Y(_00977_));
 sg13g2_inv_1 _07171_ (.Y(_00978_),
    .A(\r1[10] ));
 sg13g2_nand2_1 _07172_ (.Y(_00979_),
    .A(_00786_),
    .B(_00978_));
 sg13g2_nor2_1 _07173_ (.A(_00975_),
    .B(_00778_),
    .Y(_00980_));
 sg13g2_nor2_1 _07174_ (.A(_00979_),
    .B(_00980_),
    .Y(_00981_));
 sg13g2_nand2_1 _07175_ (.Y(_00982_),
    .A(_00977_),
    .B(_00981_));
 sg13g2_inv_1 _07176_ (.Y(_00983_),
    .A(_00049_));
 sg13g2_nand2_1 _07177_ (.Y(_00984_),
    .A(_00982_),
    .B(_00983_));
 sg13g2_nand3_1 _07178_ (.B(_00049_),
    .C(_00981_),
    .A(_00977_),
    .Y(_00985_));
 sg13g2_inv_1 _07179_ (.Y(_00986_),
    .A(\r2[12] ));
 sg13g2_nand3_1 _07180_ (.B(_00985_),
    .C(_00986_),
    .A(_00984_),
    .Y(_00987_));
 sg13g2_buf_8 _07181_ (.A(_00987_),
    .X(_00988_));
 sg13g2_nand2_1 _07182_ (.Y(_00989_),
    .A(_00982_),
    .B(_00049_));
 sg13g2_nand3_1 _07183_ (.B(_00983_),
    .C(_00981_),
    .A(_00977_),
    .Y(_00990_));
 sg13g2_nand3_1 _07184_ (.B(_00990_),
    .C(\r2[12] ),
    .A(_00989_),
    .Y(_00991_));
 sg13g2_nand2_1 _07185_ (.Y(_00992_),
    .A(_00988_),
    .B(_00991_));
 sg13g2_nand2_1 _07186_ (.Y(_00993_),
    .A(_00992_),
    .B(_00883_));
 sg13g2_a21oi_1 _07187_ (.A1(_00884_),
    .A2(_00885_),
    .Y(_00994_),
    .B1(_00880_));
 sg13g2_nand3_1 _07188_ (.B(_00988_),
    .C(_00991_),
    .A(_00994_),
    .Y(_00995_));
 sg13g2_nand2_2 _07189_ (.Y(_00996_),
    .A(_00993_),
    .B(_00995_));
 sg13g2_nor2_1 _07190_ (.A(_00800_),
    .B(_00891_),
    .Y(_00997_));
 sg13g2_nand3_1 _07191_ (.B(_00997_),
    .C(_00757_),
    .A(_00424_),
    .Y(_00998_));
 sg13g2_inv_1 _07192_ (.Y(_00999_),
    .A(_00890_));
 sg13g2_a21oi_1 _07193_ (.A1(_00888_),
    .A2(_00797_),
    .Y(_01000_),
    .B1(_00999_));
 sg13g2_nor3_1 _07194_ (.A(_00800_),
    .B(_00760_),
    .C(_00891_),
    .Y(_01001_));
 sg13g2_nor2_1 _07195_ (.A(_01000_),
    .B(_01001_),
    .Y(_01002_));
 sg13g2_nand2_1 _07196_ (.Y(_01003_),
    .A(_00998_),
    .B(_01002_));
 sg13g2_xor2_1 _07197_ (.B(_01003_),
    .A(_00996_),
    .X(_01004_));
 sg13g2_buf_2 _07198_ (.A(_01004_),
    .X(_01005_));
 sg13g2_nor2_1 _07199_ (.A(net101),
    .B(_01005_),
    .Y(_01006_));
 sg13g2_nand2_1 _07200_ (.Y(_01007_),
    .A(_01006_),
    .B(_00904_));
 sg13g2_xnor2_1 _07201_ (.Y(_01008_),
    .A(_00996_),
    .B(_01003_));
 sg13g2_buf_8 _07202_ (.A(_05562_),
    .X(_01009_));
 sg13g2_nand2_1 _07203_ (.Y(_01010_),
    .A(_01008_),
    .B(net90));
 sg13g2_nand2b_1 _07204_ (.Y(_01011_),
    .B(_01010_),
    .A_N(_00904_));
 sg13g2_nand2_1 _07205_ (.Y(_01012_),
    .A(_01007_),
    .B(_01011_));
 sg13g2_nor2_1 _07206_ (.A(net69),
    .B(_00805_),
    .Y(_01013_));
 sg13g2_nand2_1 _07207_ (.Y(_01014_),
    .A(_01012_),
    .B(_01013_));
 sg13g2_inv_1 _07208_ (.Y(_01015_),
    .A(_01013_));
 sg13g2_nand3_1 _07209_ (.B(_01011_),
    .C(_01015_),
    .A(_01007_),
    .Y(_01016_));
 sg13g2_nand2_1 _07210_ (.Y(_01017_),
    .A(_01014_),
    .B(_01016_));
 sg13g2_nand2b_1 _07211_ (.Y(_01018_),
    .B(_01017_),
    .A_N(_00973_));
 sg13g2_nand3_1 _07212_ (.B(_01016_),
    .C(_00973_),
    .A(_01014_),
    .Y(_01019_));
 sg13g2_nand2_1 _07213_ (.Y(_01020_),
    .A(_01018_),
    .B(_01019_));
 sg13g2_nor2_1 _07214_ (.A(net51),
    .B(_00710_),
    .Y(_01021_));
 sg13g2_nor2_1 _07215_ (.A(net63),
    .B(_00702_),
    .Y(_01022_));
 sg13g2_inv_1 _07216_ (.Y(_01023_),
    .A(_01022_));
 sg13g2_o21ai_1 _07217_ (.B1(_00918_),
    .Y(_01024_),
    .A1(net57),
    .A2(_00702_));
 sg13g2_o21ai_1 _07218_ (.B1(_01024_),
    .Y(_01025_),
    .A1(_01023_),
    .A2(_00921_));
 sg13g2_xnor2_1 _07219_ (.Y(_01026_),
    .A(_01021_),
    .B(_01025_));
 sg13g2_nand2_1 _07220_ (.Y(_01027_),
    .A(_01020_),
    .B(_01026_));
 sg13g2_inv_1 _07221_ (.Y(_01028_),
    .A(_01026_));
 sg13g2_nand3_1 _07222_ (.B(_01019_),
    .C(_01028_),
    .A(_01018_),
    .Y(_01029_));
 sg13g2_nand2_1 _07223_ (.Y(_01030_),
    .A(_01027_),
    .B(_01029_));
 sg13g2_nand2b_1 _07224_ (.Y(_01031_),
    .B(_01030_),
    .A_N(_00972_));
 sg13g2_nand3_1 _07225_ (.B(_01029_),
    .C(_00972_),
    .A(_01027_),
    .Y(_01032_));
 sg13g2_nand2_1 _07226_ (.Y(_01033_),
    .A(_01031_),
    .B(_01032_));
 sg13g2_inv_1 _07227_ (.Y(_01034_),
    .A(_00750_));
 sg13g2_nor2_1 _07228_ (.A(net45),
    .B(_00321_),
    .Y(_01035_));
 sg13g2_inv_1 _07229_ (.Y(_01036_),
    .A(_01035_));
 sg13g2_nor2_1 _07230_ (.A(_01034_),
    .B(_01036_),
    .Y(_01037_));
 sg13g2_inv_1 _07231_ (.Y(_01038_),
    .A(_01037_));
 sg13g2_nor2_1 _07232_ (.A(net49),
    .B(_00369_),
    .Y(_01039_));
 sg13g2_xnor2_1 _07233_ (.Y(_01040_),
    .A(_01036_),
    .B(_01039_));
 sg13g2_a21oi_1 _07234_ (.A1(_00922_),
    .A2(_00917_),
    .Y(_01041_),
    .B1(_00919_));
 sg13g2_xnor2_1 _07235_ (.Y(_01042_),
    .A(_01040_),
    .B(_01041_));
 sg13g2_xnor2_1 _07236_ (.Y(_01043_),
    .A(_01038_),
    .B(_01042_));
 sg13g2_nand2_1 _07237_ (.Y(_01044_),
    .A(_01033_),
    .B(_01043_));
 sg13g2_inv_1 _07238_ (.Y(_01045_),
    .A(_01043_));
 sg13g2_nand3_1 _07239_ (.B(_01032_),
    .C(_01045_),
    .A(_01031_),
    .Y(_01046_));
 sg13g2_nand2_1 _07240_ (.Y(_01047_),
    .A(_01044_),
    .B(_01046_));
 sg13g2_nand2b_1 _07241_ (.Y(_01048_),
    .B(_01047_),
    .A_N(_00970_));
 sg13g2_nand3_1 _07242_ (.B(_01046_),
    .C(_00970_),
    .A(_01044_),
    .Y(_01049_));
 sg13g2_nand2_1 _07243_ (.Y(_01050_),
    .A(_01048_),
    .B(_01049_));
 sg13g2_nor2b_1 _07244_ (.A(_00940_),
    .B_N(_00938_),
    .Y(_01051_));
 sg13g2_a21oi_1 _07245_ (.A1(_00941_),
    .A2(_00935_),
    .Y(_01052_),
    .B1(_01051_));
 sg13g2_nand2_1 _07246_ (.Y(_01053_),
    .A(_01050_),
    .B(_01052_));
 sg13g2_inv_1 _07247_ (.Y(_01054_),
    .A(_01052_));
 sg13g2_nand3_1 _07248_ (.B(_01049_),
    .C(_01054_),
    .A(_01048_),
    .Y(_01055_));
 sg13g2_nand3b_1 _07249_ (.B(_01053_),
    .C(_01055_),
    .Y(_01056_),
    .A_N(_00968_));
 sg13g2_buf_1 _07250_ (.A(_01056_),
    .X(_01057_));
 sg13g2_nand2_1 _07251_ (.Y(_01058_),
    .A(_01053_),
    .B(_01055_));
 sg13g2_nand2_1 _07252_ (.Y(_01059_),
    .A(_01058_),
    .B(_00968_));
 sg13g2_nand2_1 _07253_ (.Y(_01060_),
    .A(_01057_),
    .B(_01059_));
 sg13g2_inv_1 _07254_ (.Y(_01061_),
    .A(_01048_));
 sg13g2_a21oi_1 _07255_ (.A1(_01049_),
    .A2(_01054_),
    .Y(_01062_),
    .B1(_01061_));
 sg13g2_inv_1 _07256_ (.Y(_01063_),
    .A(_01031_));
 sg13g2_a21oi_1 _07257_ (.A1(_01032_),
    .A2(_01043_),
    .Y(_01064_),
    .B1(_01063_));
 sg13g2_inv_1 _07258_ (.Y(_01065_),
    .A(_01018_));
 sg13g2_a21oi_1 _07259_ (.A1(_01019_),
    .A2(_01026_),
    .Y(_01066_),
    .B1(_01065_));
 sg13g2_inv_1 _07260_ (.Y(_01067_),
    .A(_01007_));
 sg13g2_a21oi_1 _07261_ (.A1(_01011_),
    .A2(_01013_),
    .Y(_01068_),
    .B1(_01067_));
 sg13g2_nor2_1 _07262_ (.A(net69),
    .B(_00903_),
    .Y(_01069_));
 sg13g2_buf_1 _07263_ (.A(\r1[11] ),
    .X(_01070_));
 sg13g2_nor2_1 _07264_ (.A(_01070_),
    .B(\r1[10] ),
    .Y(_01071_));
 sg13g2_inv_1 _07265_ (.Y(_01072_),
    .A(_01071_));
 sg13g2_nor3_1 _07266_ (.A(_01072_),
    .B(_00787_),
    .C(_00674_),
    .Y(_01073_));
 sg13g2_nand2_1 _07267_ (.Y(_01074_),
    .A(_00671_),
    .B(_01073_));
 sg13g2_nor2_1 _07268_ (.A(_01072_),
    .B(_00873_),
    .Y(_01075_));
 sg13g2_nand2_1 _07269_ (.Y(_01076_),
    .A(_01074_),
    .B(_01075_));
 sg13g2_inv_1 _07270_ (.Y(_01077_),
    .A(_00048_));
 sg13g2_nand2_1 _07271_ (.Y(_01078_),
    .A(_01076_),
    .B(_01077_));
 sg13g2_nand3_1 _07272_ (.B(_00048_),
    .C(_01075_),
    .A(_01074_),
    .Y(_01079_));
 sg13g2_nand2_1 _07273_ (.Y(_01080_),
    .A(_01078_),
    .B(_01079_));
 sg13g2_buf_2 _07274_ (.A(\r2[13] ),
    .X(_01081_));
 sg13g2_nand2_1 _07275_ (.Y(_01082_),
    .A(_01080_),
    .B(_01081_));
 sg13g2_inv_1 _07276_ (.Y(_01083_),
    .A(_01081_));
 sg13g2_nand3_1 _07277_ (.B(_01079_),
    .C(_01083_),
    .A(_01078_),
    .Y(_01084_));
 sg13g2_buf_2 _07278_ (.A(_01084_),
    .X(_01085_));
 sg13g2_nand2_1 _07279_ (.Y(_01086_),
    .A(_01082_),
    .B(_01085_));
 sg13g2_xnor2_1 _07280_ (.Y(_01087_),
    .A(_00988_),
    .B(_01086_));
 sg13g2_buf_1 _07281_ (.A(_01087_),
    .X(_01088_));
 sg13g2_nor2_1 _07282_ (.A(_00891_),
    .B(_00996_),
    .Y(_01089_));
 sg13g2_nor2_1 _07283_ (.A(_00691_),
    .B(_00800_),
    .Y(_01090_));
 sg13g2_nand3_1 _07284_ (.B(_01089_),
    .C(_01090_),
    .A(_00698_),
    .Y(_01091_));
 sg13g2_nor2_1 _07285_ (.A(_00883_),
    .B(_00992_),
    .Y(_01092_));
 sg13g2_o21ai_1 _07286_ (.B1(_00993_),
    .Y(_01093_),
    .A1(_00888_),
    .A2(_01092_));
 sg13g2_a21oi_1 _07287_ (.A1(_01089_),
    .A2(_00894_),
    .Y(_01094_),
    .B1(_01093_));
 sg13g2_nand2_1 _07288_ (.Y(_01095_),
    .A(_01091_),
    .B(_01094_));
 sg13g2_nand2b_1 _07289_ (.Y(_01096_),
    .B(_01095_),
    .A_N(_01088_));
 sg13g2_nand3_1 _07290_ (.B(_01088_),
    .C(_01094_),
    .A(_01091_),
    .Y(_01097_));
 sg13g2_nand2_1 _07291_ (.Y(_01098_),
    .A(_01096_),
    .B(_01097_));
 sg13g2_buf_8 _07292_ (.A(_01098_),
    .X(_01099_));
 sg13g2_nor2_1 _07293_ (.A(net62),
    .B(_01099_),
    .Y(_01100_));
 sg13g2_nand2_1 _07294_ (.Y(_01101_),
    .A(_01100_),
    .B(_01006_));
 sg13g2_nand3_1 _07295_ (.B(_01097_),
    .C(net90),
    .A(_01096_),
    .Y(_01102_));
 sg13g2_nand2_1 _07296_ (.Y(_01103_),
    .A(_01008_),
    .B(_00610_));
 sg13g2_nand2_1 _07297_ (.Y(_01104_),
    .A(_01102_),
    .B(_01103_));
 sg13g2_nand3b_1 _07298_ (.B(_01101_),
    .C(_01104_),
    .Y(_01105_),
    .A_N(_01069_));
 sg13g2_nand2_1 _07299_ (.Y(_01106_),
    .A(_01101_),
    .B(_01104_));
 sg13g2_nand2_1 _07300_ (.Y(_01107_),
    .A(_01106_),
    .B(_01069_));
 sg13g2_nand2_1 _07301_ (.Y(_01108_),
    .A(_01105_),
    .B(_01107_));
 sg13g2_nand2b_1 _07302_ (.Y(_01109_),
    .B(_01108_),
    .A_N(_01068_));
 sg13g2_nand3_1 _07303_ (.B(_01107_),
    .C(_01068_),
    .A(_01105_),
    .Y(_01110_));
 sg13g2_nand2_1 _07304_ (.Y(_01111_),
    .A(_01109_),
    .B(_01110_));
 sg13g2_buf_1 _07305_ (.A(net51),
    .X(_01112_));
 sg13g2_nor2_1 _07306_ (.A(net44),
    .B(_00462_),
    .Y(_01113_));
 sg13g2_nor2_1 _07307_ (.A(net57),
    .B(_00805_),
    .Y(_01114_));
 sg13g2_xnor2_1 _07308_ (.Y(_01115_),
    .A(_01023_),
    .B(_01114_));
 sg13g2_xor2_1 _07309_ (.B(_01115_),
    .A(_01113_),
    .X(_01116_));
 sg13g2_nand2_1 _07310_ (.Y(_01117_),
    .A(_01111_),
    .B(_01116_));
 sg13g2_inv_1 _07311_ (.Y(_01118_),
    .A(_01116_));
 sg13g2_nand3_1 _07312_ (.B(_01110_),
    .C(_01118_),
    .A(_01109_),
    .Y(_01119_));
 sg13g2_nand2_1 _07313_ (.Y(_01120_),
    .A(_01117_),
    .B(_01119_));
 sg13g2_nand2b_1 _07314_ (.Y(_01121_),
    .B(_01120_),
    .A_N(_01066_));
 sg13g2_nand3_1 _07315_ (.B(_01119_),
    .C(_01066_),
    .A(_01117_),
    .Y(_01122_));
 sg13g2_nand2_1 _07316_ (.Y(_01123_),
    .A(_01121_),
    .B(_01122_));
 sg13g2_inv_1 _07317_ (.Y(_01124_),
    .A(_00937_));
 sg13g2_nor2_1 _07318_ (.A(net45),
    .B(_00369_),
    .Y(_01125_));
 sg13g2_inv_1 _07319_ (.Y(_01126_),
    .A(_01125_));
 sg13g2_nor2_1 _07320_ (.A(_01124_),
    .B(_01126_),
    .Y(_01127_));
 sg13g2_inv_1 _07321_ (.Y(_01128_),
    .A(_01127_));
 sg13g2_nand2_1 _07322_ (.Y(_01129_),
    .A(_00407_),
    .B(_00223_));
 sg13g2_xnor2_1 _07323_ (.Y(_01130_),
    .A(_01125_),
    .B(_01129_));
 sg13g2_a22oi_1 _07324_ (.Y(_01131_),
    .B1(_01021_),
    .B2(_01024_),
    .A2(_00920_),
    .A1(_01022_));
 sg13g2_xnor2_1 _07325_ (.Y(_01132_),
    .A(_01130_),
    .B(_01131_));
 sg13g2_xnor2_1 _07326_ (.Y(_01133_),
    .A(_01128_),
    .B(_01132_));
 sg13g2_nand2_1 _07327_ (.Y(_01134_),
    .A(_01123_),
    .B(_01133_));
 sg13g2_inv_1 _07328_ (.Y(_01135_),
    .A(_01133_));
 sg13g2_nand3_1 _07329_ (.B(_01122_),
    .C(_01135_),
    .A(_01121_),
    .Y(_01136_));
 sg13g2_nand2_1 _07330_ (.Y(_01137_),
    .A(_01134_),
    .B(_01136_));
 sg13g2_nand2b_1 _07331_ (.Y(_01138_),
    .B(_01137_),
    .A_N(_01064_));
 sg13g2_nand3_1 _07332_ (.B(_01136_),
    .C(_01064_),
    .A(_01134_),
    .Y(_01139_));
 sg13g2_nand2_1 _07333_ (.Y(_01140_),
    .A(_01138_),
    .B(_01139_));
 sg13g2_nor2b_1 _07334_ (.A(_01041_),
    .B_N(_01040_),
    .Y(_01141_));
 sg13g2_a21oi_1 _07335_ (.A1(_01042_),
    .A2(_01037_),
    .Y(_01142_),
    .B1(_01141_));
 sg13g2_nand2_1 _07336_ (.Y(_01143_),
    .A(_01140_),
    .B(_01142_));
 sg13g2_inv_1 _07337_ (.Y(_01144_),
    .A(_01142_));
 sg13g2_nand3_1 _07338_ (.B(_01139_),
    .C(_01144_),
    .A(_01138_),
    .Y(_01145_));
 sg13g2_nand3b_1 _07339_ (.B(_01143_),
    .C(_01145_),
    .Y(_01146_),
    .A_N(_01062_));
 sg13g2_buf_1 _07340_ (.A(_01146_),
    .X(_01147_));
 sg13g2_nand2_1 _07341_ (.Y(_01148_),
    .A(_01143_),
    .B(_01145_));
 sg13g2_nand2_1 _07342_ (.Y(_01149_),
    .A(_01148_),
    .B(_01062_));
 sg13g2_nand2_1 _07343_ (.Y(_01150_),
    .A(_01147_),
    .B(_01149_));
 sg13g2_nor2_1 _07344_ (.A(_01060_),
    .B(_01150_),
    .Y(_01151_));
 sg13g2_nand2_1 _07345_ (.Y(_01152_),
    .A(_00966_),
    .B(_01151_));
 sg13g2_nand2_1 _07346_ (.Y(_01153_),
    .A(_01147_),
    .B(_01057_));
 sg13g2_nand2_1 _07347_ (.Y(_01154_),
    .A(_01153_),
    .B(_01149_));
 sg13g2_nand2_1 _07348_ (.Y(_01155_),
    .A(_01152_),
    .B(_01154_));
 sg13g2_inv_1 _07349_ (.Y(_01156_),
    .A(_01138_));
 sg13g2_a21oi_1 _07350_ (.A1(_01139_),
    .A2(_01144_),
    .Y(_01157_),
    .B1(_01156_));
 sg13g2_inv_1 _07351_ (.Y(_01158_),
    .A(_01157_));
 sg13g2_a21oi_1 _07352_ (.A1(_01117_),
    .A2(_01119_),
    .Y(_01159_),
    .B1(_01066_));
 sg13g2_a21oi_1 _07353_ (.A1(_01122_),
    .A2(_01133_),
    .Y(_01160_),
    .B1(_01159_));
 sg13g2_inv_1 _07354_ (.Y(_01161_),
    .A(_01109_));
 sg13g2_a21oi_1 _07355_ (.A1(_01110_),
    .A2(_01116_),
    .Y(_01162_),
    .B1(_01161_));
 sg13g2_a22oi_1 _07356_ (.Y(_01163_),
    .B1(_01069_),
    .B2(_01104_),
    .A2(_01006_),
    .A1(_01100_));
 sg13g2_nand2_1 _07357_ (.Y(_01164_),
    .A(_01086_),
    .B(_00988_));
 sg13g2_nor2_1 _07358_ (.A(_00988_),
    .B(_01086_),
    .Y(_01165_));
 sg13g2_a21oi_1 _07359_ (.A1(_00993_),
    .A2(_01164_),
    .Y(_01166_),
    .B1(_01165_));
 sg13g2_nor2_1 _07360_ (.A(_00996_),
    .B(_01088_),
    .Y(_01167_));
 sg13g2_nand2_1 _07361_ (.Y(_01168_),
    .A(_01167_),
    .B(_01000_));
 sg13g2_nand2b_1 _07362_ (.Y(_01169_),
    .B(_01168_),
    .A_N(_01166_));
 sg13g2_nand2_1 _07363_ (.Y(_01170_),
    .A(_01167_),
    .B(_00997_));
 sg13g2_nor2b_1 _07364_ (.A(_01170_),
    .B_N(_00761_),
    .Y(_01171_));
 sg13g2_nor2_1 _07365_ (.A(_01169_),
    .B(_01171_),
    .Y(_01172_));
 sg13g2_nor2_1 _07366_ (.A(_00766_),
    .B(_01170_),
    .Y(_01173_));
 sg13g2_nand2b_1 _07367_ (.Y(_01174_),
    .B(_01173_),
    .A_N(_00336_));
 sg13g2_nand2_1 _07368_ (.Y(_01175_),
    .A(_01172_),
    .B(_01174_));
 sg13g2_inv_4 _07369_ (.A(_01085_),
    .Y(_01176_));
 sg13g2_nand2_1 _07370_ (.Y(_01177_),
    .A(_00774_),
    .B(_00441_));
 sg13g2_nand2_1 _07371_ (.Y(_01178_),
    .A(_01177_),
    .B(_00778_));
 sg13g2_buf_1 _07372_ (.A(\r1[12] ),
    .X(_01179_));
 sg13g2_nor2_1 _07373_ (.A(_01070_),
    .B(_01179_),
    .Y(_01180_));
 sg13g2_inv_1 _07374_ (.Y(_01181_),
    .A(_01180_));
 sg13g2_nor2_1 _07375_ (.A(_01181_),
    .B(_00975_),
    .Y(_01182_));
 sg13g2_nand2_1 _07376_ (.Y(_01183_),
    .A(_01178_),
    .B(_01182_));
 sg13g2_nand4_1 _07377_ (.B(_01182_),
    .C(_00345_),
    .A(_00774_),
    .Y(_01184_),
    .D(_00436_));
 sg13g2_nor2_1 _07378_ (.A(_01181_),
    .B(_00979_),
    .Y(_01185_));
 sg13g2_nand3_1 _07379_ (.B(_01184_),
    .C(_01185_),
    .A(_01183_),
    .Y(_01186_));
 sg13g2_buf_1 _07380_ (.A(_00047_),
    .X(_01187_));
 sg13g2_nand2_1 _07381_ (.Y(_01188_),
    .A(_01186_),
    .B(_01187_));
 sg13g2_inv_1 _07382_ (.Y(_01189_),
    .A(_01187_));
 sg13g2_nand4_1 _07383_ (.B(_01184_),
    .C(_01189_),
    .A(_01183_),
    .Y(_01190_),
    .D(_01185_));
 sg13g2_nand2_1 _07384_ (.Y(_01191_),
    .A(_01188_),
    .B(_01190_));
 sg13g2_buf_1 _07385_ (.A(\r2[14] ),
    .X(_01192_));
 sg13g2_inv_1 _07386_ (.Y(_01193_),
    .A(_01192_));
 sg13g2_nand2_1 _07387_ (.Y(_01194_),
    .A(_01191_),
    .B(_01193_));
 sg13g2_nand3_1 _07388_ (.B(_01190_),
    .C(_01192_),
    .A(_01188_),
    .Y(_01195_));
 sg13g2_nand2_1 _07389_ (.Y(_01196_),
    .A(_01194_),
    .B(_01195_));
 sg13g2_xnor2_1 _07390_ (.Y(_01197_),
    .A(_01176_),
    .B(_01196_));
 sg13g2_nand2_1 _07391_ (.Y(_01198_),
    .A(_01175_),
    .B(_01197_));
 sg13g2_nand2_1 _07392_ (.Y(_01199_),
    .A(_01196_),
    .B(_01085_));
 sg13g2_nand3_1 _07393_ (.B(_01195_),
    .C(_01176_),
    .A(_01194_),
    .Y(_01200_));
 sg13g2_nand2_1 _07394_ (.Y(_01201_),
    .A(_01199_),
    .B(_01200_));
 sg13g2_nand3_1 _07395_ (.B(_01174_),
    .C(_01201_),
    .A(_01172_),
    .Y(_01202_));
 sg13g2_nand2_1 _07396_ (.Y(_01203_),
    .A(_01198_),
    .B(_01202_));
 sg13g2_buf_8 _07397_ (.A(_01203_),
    .X(_01204_));
 sg13g2_nor2_1 _07398_ (.A(net62),
    .B(_01204_),
    .Y(_01205_));
 sg13g2_nand2b_1 _07399_ (.Y(_01206_),
    .B(_01205_),
    .A_N(_01102_));
 sg13g2_nand3_1 _07400_ (.B(_01202_),
    .C(net90),
    .A(_01198_),
    .Y(_01207_));
 sg13g2_xnor2_1 _07401_ (.Y(_01208_),
    .A(_01088_),
    .B(_01095_));
 sg13g2_nand2_1 _07402_ (.Y(_01209_),
    .A(_01208_),
    .B(net68));
 sg13g2_nand2_1 _07403_ (.Y(_01210_),
    .A(_01207_),
    .B(_01209_));
 sg13g2_nand2_1 _07404_ (.Y(_01211_),
    .A(_01206_),
    .B(_01210_));
 sg13g2_nor2_1 _07405_ (.A(net69),
    .B(_01005_),
    .Y(_01212_));
 sg13g2_nand2_1 _07406_ (.Y(_01213_),
    .A(_01211_),
    .B(_01212_));
 sg13g2_inv_1 _07407_ (.Y(_01214_),
    .A(_01212_));
 sg13g2_nand3_1 _07408_ (.B(_01210_),
    .C(_01214_),
    .A(_01206_),
    .Y(_01215_));
 sg13g2_nand2_1 _07409_ (.Y(_01216_),
    .A(_01213_),
    .B(_01215_));
 sg13g2_nand2b_1 _07410_ (.Y(_01217_),
    .B(_01216_),
    .A_N(_01163_));
 sg13g2_nand3_1 _07411_ (.B(_01215_),
    .C(_01163_),
    .A(_01213_),
    .Y(_01218_));
 sg13g2_buf_1 _07412_ (.A(_01218_),
    .X(_01219_));
 sg13g2_nand2_1 _07413_ (.Y(_01220_),
    .A(_01217_),
    .B(_01219_));
 sg13g2_nor2_1 _07414_ (.A(net44),
    .B(_00702_),
    .Y(_01221_));
 sg13g2_nor2_1 _07415_ (.A(net63),
    .B(_00903_),
    .Y(_01222_));
 sg13g2_inv_1 _07416_ (.Y(_01223_),
    .A(_01222_));
 sg13g2_inv_2 _07417_ (.Y(_01224_),
    .A(_01114_));
 sg13g2_nor2_1 _07418_ (.A(_01223_),
    .B(_01224_),
    .Y(_01225_));
 sg13g2_inv_1 _07419_ (.Y(_01226_),
    .A(_00903_));
 sg13g2_nand2_1 _07420_ (.Y(_01227_),
    .A(_01226_),
    .B(net71));
 sg13g2_o21ai_1 _07421_ (.B1(_01227_),
    .Y(_01228_),
    .A1(net63),
    .A2(_00805_));
 sg13g2_nand2b_1 _07422_ (.Y(_01229_),
    .B(_01228_),
    .A_N(_01225_));
 sg13g2_xnor2_1 _07423_ (.Y(_01230_),
    .A(_01221_),
    .B(_01229_));
 sg13g2_nand2_1 _07424_ (.Y(_01231_),
    .A(_01220_),
    .B(_01230_));
 sg13g2_inv_1 _07425_ (.Y(_01232_),
    .A(_01230_));
 sg13g2_nand3_1 _07426_ (.B(_01219_),
    .C(_01232_),
    .A(_01217_),
    .Y(_01233_));
 sg13g2_nand2_1 _07427_ (.Y(_01234_),
    .A(_01231_),
    .B(_01233_));
 sg13g2_nand2b_1 _07428_ (.Y(_01235_),
    .B(_01234_),
    .A_N(_01162_));
 sg13g2_nand3_1 _07429_ (.B(_01233_),
    .C(_01162_),
    .A(_01231_),
    .Y(_01236_));
 sg13g2_buf_1 _07430_ (.A(_01236_),
    .X(_01237_));
 sg13g2_nand2_1 _07431_ (.Y(_01238_),
    .A(_01235_),
    .B(_01237_));
 sg13g2_nor2_1 _07432_ (.A(_01126_),
    .B(_01129_),
    .Y(_01239_));
 sg13g2_nand2_1 _07433_ (.Y(_01240_),
    .A(_00407_),
    .B(net50));
 sg13g2_nor2_1 _07434_ (.A(net49),
    .B(_00462_),
    .Y(_01241_));
 sg13g2_xnor2_1 _07435_ (.Y(_01242_),
    .A(_01240_),
    .B(_01241_));
 sg13g2_nor2_1 _07436_ (.A(_01023_),
    .B(_01224_),
    .Y(_01243_));
 sg13g2_a21oi_1 _07437_ (.A1(_01115_),
    .A2(_01113_),
    .Y(_01244_),
    .B1(_01243_));
 sg13g2_xnor2_1 _07438_ (.Y(_01245_),
    .A(_01242_),
    .B(_01244_));
 sg13g2_xor2_1 _07439_ (.B(_01245_),
    .A(_01239_),
    .X(_01246_));
 sg13g2_nand2_1 _07440_ (.Y(_01247_),
    .A(_01238_),
    .B(_01246_));
 sg13g2_inv_1 _07441_ (.Y(_01248_),
    .A(_01246_));
 sg13g2_nand3_1 _07442_ (.B(_01237_),
    .C(_01248_),
    .A(_01235_),
    .Y(_01249_));
 sg13g2_nand2_1 _07443_ (.Y(_01250_),
    .A(_01247_),
    .B(_01249_));
 sg13g2_nand2b_1 _07444_ (.Y(_01251_),
    .B(_01250_),
    .A_N(_01160_));
 sg13g2_nand3_1 _07445_ (.B(_01249_),
    .C(_01160_),
    .A(_01247_),
    .Y(_01252_));
 sg13g2_nand2_1 _07446_ (.Y(_01253_),
    .A(_01251_),
    .B(_01252_));
 sg13g2_nor2b_1 _07447_ (.A(_01131_),
    .B_N(_01130_),
    .Y(_01254_));
 sg13g2_a21oi_1 _07448_ (.A1(_01132_),
    .A2(_01127_),
    .Y(_01255_),
    .B1(_01254_));
 sg13g2_nand2_1 _07449_ (.Y(_01256_),
    .A(_01253_),
    .B(_01255_));
 sg13g2_inv_1 _07450_ (.Y(_01257_),
    .A(_01255_));
 sg13g2_nand3_1 _07451_ (.B(_01252_),
    .C(_01257_),
    .A(_01251_),
    .Y(_01258_));
 sg13g2_nand2_1 _07452_ (.Y(_01259_),
    .A(_01256_),
    .B(_01258_));
 sg13g2_xnor2_1 _07453_ (.Y(_01260_),
    .A(_01158_),
    .B(_01259_));
 sg13g2_inv_1 _07454_ (.Y(_01261_),
    .A(_01260_));
 sg13g2_inv_1 _07455_ (.Y(_01262_),
    .A(_01251_));
 sg13g2_a21oi_1 _07456_ (.A1(_01252_),
    .A2(_01257_),
    .Y(_01263_),
    .B1(_01262_));
 sg13g2_inv_2 _07457_ (.Y(_01264_),
    .A(_01263_));
 sg13g2_a21oi_1 _07458_ (.A1(_01231_),
    .A2(_01233_),
    .Y(_01265_),
    .B1(_01162_));
 sg13g2_a21oi_1 _07459_ (.A1(_01237_),
    .A2(_01246_),
    .Y(_01266_),
    .B1(_01265_));
 sg13g2_a21oi_1 _07460_ (.A1(_01213_),
    .A2(_01215_),
    .Y(_01267_),
    .B1(_01163_));
 sg13g2_a21oi_2 _07461_ (.B1(_01267_),
    .Y(_01268_),
    .A2(_01230_),
    .A1(_01219_));
 sg13g2_nand3_1 _07462_ (.B(_01202_),
    .C(net68),
    .A(_01198_),
    .Y(_01269_));
 sg13g2_nor2_1 _07463_ (.A(_01102_),
    .B(_01269_),
    .Y(_01270_));
 sg13g2_a21oi_2 _07464_ (.B1(_01270_),
    .Y(_01271_),
    .A2(_01212_),
    .A1(_01210_));
 sg13g2_nor2_1 _07465_ (.A(net69),
    .B(_01099_),
    .Y(_01272_));
 sg13g2_nor2_1 _07466_ (.A(_01088_),
    .B(_01201_),
    .Y(_01273_));
 sg13g2_nand3_1 _07467_ (.B(_01089_),
    .C(_01273_),
    .A(_00899_),
    .Y(_01274_));
 sg13g2_nand2_1 _07468_ (.Y(_01275_),
    .A(_01273_),
    .B(_01093_));
 sg13g2_inv_1 _07469_ (.Y(_01276_),
    .A(_01164_));
 sg13g2_inv_1 _07470_ (.Y(_01277_),
    .A(_01199_));
 sg13g2_a21oi_1 _07471_ (.A1(_01200_),
    .A2(_01276_),
    .Y(_01278_),
    .B1(_01277_));
 sg13g2_nand2_1 _07472_ (.Y(_01279_),
    .A(_01275_),
    .B(_01278_));
 sg13g2_inv_2 _07473_ (.Y(_01280_),
    .A(_01279_));
 sg13g2_nand2_1 _07474_ (.Y(_01281_),
    .A(_01274_),
    .B(_01280_));
 sg13g2_inv_1 _07475_ (.Y(_01282_),
    .A(_01194_));
 sg13g2_inv_2 _07476_ (.Y(_01283_),
    .A(_00046_));
 sg13g2_inv_1 _07477_ (.Y(_01284_),
    .A(_00045_));
 sg13g2_nor2_1 _07478_ (.A(\r1[13] ),
    .B(_01179_),
    .Y(_01285_));
 sg13g2_nand2_1 _07479_ (.Y(_01286_),
    .A(_01071_),
    .B(_01285_));
 sg13g2_nor2_1 _07480_ (.A(_01286_),
    .B(_00873_),
    .Y(_01287_));
 sg13g2_nand2_1 _07481_ (.Y(_01288_),
    .A(_00871_),
    .B(_01287_));
 sg13g2_xnor2_1 _07482_ (.Y(_01289_),
    .A(_01284_),
    .B(_01288_));
 sg13g2_xnor2_1 _07483_ (.Y(_01290_),
    .A(_01283_),
    .B(_01289_));
 sg13g2_xnor2_1 _07484_ (.Y(_01291_),
    .A(_01282_),
    .B(_01290_));
 sg13g2_nand2_1 _07485_ (.Y(_01292_),
    .A(_01281_),
    .B(_01291_));
 sg13g2_nand2_1 _07486_ (.Y(_01293_),
    .A(_01290_),
    .B(_01194_));
 sg13g2_xnor2_1 _07487_ (.Y(_01294_),
    .A(_00046_),
    .B(_01289_));
 sg13g2_nand2_1 _07488_ (.Y(_01295_),
    .A(_01294_),
    .B(_01282_));
 sg13g2_nand2_1 _07489_ (.Y(_01296_),
    .A(_01293_),
    .B(_01295_));
 sg13g2_nand3_1 _07490_ (.B(_01296_),
    .C(_01280_),
    .A(_01274_),
    .Y(_01297_));
 sg13g2_nand2_1 _07491_ (.Y(_01298_),
    .A(_01292_),
    .B(_01297_));
 sg13g2_buf_2 _07492_ (.A(_01298_),
    .X(_01299_));
 sg13g2_nor2_1 _07493_ (.A(_05490_),
    .B(_01299_),
    .Y(_01300_));
 sg13g2_nand2_1 _07494_ (.Y(_01301_),
    .A(_01300_),
    .B(_01205_));
 sg13g2_nand3_1 _07495_ (.B(_01297_),
    .C(_03300_),
    .A(_01292_),
    .Y(_01302_));
 sg13g2_nand2_1 _07496_ (.Y(_01303_),
    .A(_01302_),
    .B(_01269_));
 sg13g2_nand2_1 _07497_ (.Y(_01304_),
    .A(_01301_),
    .B(_01303_));
 sg13g2_nand2b_1 _07498_ (.Y(_01305_),
    .B(_01304_),
    .A_N(_01272_));
 sg13g2_nand3_1 _07499_ (.B(_01303_),
    .C(_01272_),
    .A(_01301_),
    .Y(_01306_));
 sg13g2_nand2_1 _07500_ (.Y(_01307_),
    .A(_01305_),
    .B(_01306_));
 sg13g2_nand2b_1 _07501_ (.Y(_01308_),
    .B(_01307_),
    .A_N(_01271_));
 sg13g2_nand3_1 _07502_ (.B(_01306_),
    .C(_01271_),
    .A(_01305_),
    .Y(_01309_));
 sg13g2_nand2_1 _07503_ (.Y(_01310_),
    .A(_01308_),
    .B(_01309_));
 sg13g2_nor2_1 _07504_ (.A(net44),
    .B(_00805_),
    .Y(_01311_));
 sg13g2_nand2_1 _07505_ (.Y(_01312_),
    .A(_01008_),
    .B(net65));
 sg13g2_nand2_1 _07506_ (.Y(_01313_),
    .A(_01008_),
    .B(_05565_));
 sg13g2_nand2_1 _07507_ (.Y(_01314_),
    .A(_01313_),
    .B(_01223_));
 sg13g2_o21ai_1 _07508_ (.B1(_01314_),
    .Y(_01315_),
    .A1(_01312_),
    .A2(_01227_));
 sg13g2_xnor2_1 _07509_ (.Y(_01316_),
    .A(_01311_),
    .B(_01315_));
 sg13g2_nand2_1 _07510_ (.Y(_01317_),
    .A(_01310_),
    .B(_01316_));
 sg13g2_inv_2 _07511_ (.Y(_01318_),
    .A(_01316_));
 sg13g2_nand3_1 _07512_ (.B(_01309_),
    .C(_01318_),
    .A(_01308_),
    .Y(_01319_));
 sg13g2_nand2_1 _07513_ (.Y(_01320_),
    .A(_01317_),
    .B(_01319_));
 sg13g2_nand2b_1 _07514_ (.Y(_01321_),
    .B(_01320_),
    .A_N(_01268_));
 sg13g2_nand3_1 _07515_ (.B(_01319_),
    .C(_01268_),
    .A(_01317_),
    .Y(_01322_));
 sg13g2_nand2_1 _07516_ (.Y(_01323_),
    .A(_01321_),
    .B(_01322_));
 sg13g2_nor3_1 _07517_ (.A(net45),
    .B(_00462_),
    .C(_01129_),
    .Y(_01324_));
 sg13g2_nor2_1 _07518_ (.A(net45),
    .B(_00702_),
    .Y(_01325_));
 sg13g2_nand2_1 _07519_ (.Y(_01326_),
    .A(_01325_),
    .B(_01241_));
 sg13g2_inv_1 _07520_ (.Y(_01327_),
    .A(_01326_));
 sg13g2_nor2_1 _07521_ (.A(net49),
    .B(_00702_),
    .Y(_01328_));
 sg13g2_a21oi_1 _07522_ (.A1(net50),
    .A2(_00706_),
    .Y(_01329_),
    .B1(_01328_));
 sg13g2_nor2_1 _07523_ (.A(_01327_),
    .B(_01329_),
    .Y(_01330_));
 sg13g2_a21oi_1 _07524_ (.A1(_01228_),
    .A2(_01221_),
    .Y(_01331_),
    .B1(_01225_));
 sg13g2_xnor2_1 _07525_ (.Y(_01332_),
    .A(_01330_),
    .B(_01331_));
 sg13g2_xor2_1 _07526_ (.B(_01332_),
    .A(_01324_),
    .X(_01333_));
 sg13g2_nand2_1 _07527_ (.Y(_01334_),
    .A(_01323_),
    .B(_01333_));
 sg13g2_inv_1 _07528_ (.Y(_01335_),
    .A(_01333_));
 sg13g2_nand3_1 _07529_ (.B(_01322_),
    .C(_01335_),
    .A(_01321_),
    .Y(_01336_));
 sg13g2_nand2_1 _07530_ (.Y(_01337_),
    .A(_01334_),
    .B(_01336_));
 sg13g2_nand2b_1 _07531_ (.Y(_01338_),
    .B(_01337_),
    .A_N(_01266_));
 sg13g2_nand3_1 _07532_ (.B(_01336_),
    .C(_01266_),
    .A(_01334_),
    .Y(_01339_));
 sg13g2_nand2_1 _07533_ (.Y(_01340_),
    .A(_01338_),
    .B(_01339_));
 sg13g2_nor2b_1 _07534_ (.A(_01244_),
    .B_N(_01242_),
    .Y(_01341_));
 sg13g2_a21oi_1 _07535_ (.A1(_01245_),
    .A2(_01239_),
    .Y(_01342_),
    .B1(_01341_));
 sg13g2_inv_1 _07536_ (.Y(_01343_),
    .A(_01342_));
 sg13g2_nand2_1 _07537_ (.Y(_01344_),
    .A(_01340_),
    .B(_01343_));
 sg13g2_nand3_1 _07538_ (.B(_01339_),
    .C(_01342_),
    .A(_01338_),
    .Y(_01345_));
 sg13g2_nand2_1 _07539_ (.Y(_01346_),
    .A(_01344_),
    .B(_01345_));
 sg13g2_xnor2_1 _07540_ (.Y(_01347_),
    .A(_01264_),
    .B(_01346_));
 sg13g2_inv_2 _07541_ (.Y(_01348_),
    .A(_01347_));
 sg13g2_nor2_1 _07542_ (.A(_01261_),
    .B(_01348_),
    .Y(_01349_));
 sg13g2_nand2_1 _07543_ (.Y(_01350_),
    .A(_01155_),
    .B(_01349_));
 sg13g2_nand3_1 _07544_ (.B(_01344_),
    .C(_01345_),
    .A(_01264_),
    .Y(_01351_));
 sg13g2_nand3_1 _07545_ (.B(_01256_),
    .C(_01258_),
    .A(_01158_),
    .Y(_01352_));
 sg13g2_nand2_1 _07546_ (.Y(_01353_),
    .A(_01351_),
    .B(_01352_));
 sg13g2_nand2_1 _07547_ (.Y(_01354_),
    .A(_01346_),
    .B(_01263_));
 sg13g2_nand2_1 _07548_ (.Y(_01355_),
    .A(_01353_),
    .B(_01354_));
 sg13g2_nand2_1 _07549_ (.Y(_01356_),
    .A(_01350_),
    .B(_01355_));
 sg13g2_nand2_1 _07550_ (.Y(_01357_),
    .A(_01320_),
    .B(_01268_));
 sg13g2_nor2_1 _07551_ (.A(_01268_),
    .B(_01320_),
    .Y(_01358_));
 sg13g2_a21oi_2 _07552_ (.B1(_01358_),
    .Y(_01359_),
    .A2(_01333_),
    .A1(_01357_));
 sg13g2_nand2_1 _07553_ (.Y(_01360_),
    .A(_01307_),
    .B(_01271_));
 sg13g2_nor2_1 _07554_ (.A(_01271_),
    .B(_01307_),
    .Y(_01361_));
 sg13g2_a21oi_2 _07555_ (.B1(_01361_),
    .Y(_01362_),
    .A2(_01316_),
    .A1(_01360_));
 sg13g2_inv_1 _07556_ (.Y(_01363_),
    .A(_01301_));
 sg13g2_a21oi_2 _07557_ (.B1(_01363_),
    .Y(_01364_),
    .A2(_01272_),
    .A1(_01303_));
 sg13g2_inv_1 _07558_ (.Y(_01365_),
    .A(_01295_));
 sg13g2_a21oi_1 _07559_ (.A1(_01199_),
    .A2(_01293_),
    .Y(_01366_),
    .B1(_01365_));
 sg13g2_nor2_1 _07560_ (.A(_01296_),
    .B(_01201_),
    .Y(_01367_));
 sg13g2_nand2_1 _07561_ (.Y(_01368_),
    .A(_01367_),
    .B(_01166_));
 sg13g2_nand2b_1 _07562_ (.Y(_01369_),
    .B(_01368_),
    .A_N(_01366_));
 sg13g2_nand2_1 _07563_ (.Y(_01370_),
    .A(_01367_),
    .B(_01167_));
 sg13g2_nor2_1 _07564_ (.A(_01370_),
    .B(_01002_),
    .Y(_01371_));
 sg13g2_nor2_1 _07565_ (.A(_01369_),
    .B(_01371_),
    .Y(_01372_));
 sg13g2_nand2_1 _07566_ (.Y(_01373_),
    .A(_00997_),
    .B(_00757_));
 sg13g2_nor2_1 _07567_ (.A(_01373_),
    .B(_01370_),
    .Y(_01374_));
 sg13g2_nand2_1 _07568_ (.Y(_01375_),
    .A(_01374_),
    .B(_00424_));
 sg13g2_nand2_1 _07569_ (.Y(_01376_),
    .A(_01372_),
    .B(_01375_));
 sg13g2_inv_1 _07570_ (.Y(_01377_),
    .A(\r2[15] ));
 sg13g2_nand2b_1 _07571_ (.Y(_01378_),
    .B(_01377_),
    .A_N(_01289_));
 sg13g2_buf_1 _07572_ (.A(_00038_),
    .X(_01379_));
 sg13g2_buf_1 _07573_ (.A(\r1[14] ),
    .X(_01380_));
 sg13g2_inv_1 _07574_ (.Y(_01381_),
    .A(_01380_));
 sg13g2_inv_2 _07575_ (.Y(_01382_),
    .A(\r1[13] ));
 sg13g2_nand3_1 _07576_ (.B(_01381_),
    .C(_01382_),
    .A(_01180_),
    .Y(_01383_));
 sg13g2_nor3_1 _07577_ (.A(_00979_),
    .B(_01383_),
    .C(_00980_),
    .Y(_01384_));
 sg13g2_nor4_1 _07578_ (.A(_00674_),
    .B(_01383_),
    .C(_00975_),
    .D(_00435_),
    .Y(_01385_));
 sg13g2_nand2_1 _07579_ (.Y(_01386_),
    .A(_01385_),
    .B(_00443_));
 sg13g2_nand2_1 _07580_ (.Y(_01387_),
    .A(_01384_),
    .B(_01386_));
 sg13g2_nand2_1 _07581_ (.Y(_01388_),
    .A(_01387_),
    .B(_00039_));
 sg13g2_inv_1 _07582_ (.Y(_01389_),
    .A(_00039_));
 sg13g2_nand3_1 _07583_ (.B(_01386_),
    .C(_01389_),
    .A(_01384_),
    .Y(_01390_));
 sg13g2_nand2_1 _07584_ (.Y(_01391_),
    .A(_01388_),
    .B(_01390_));
 sg13g2_xnor2_1 _07585_ (.Y(_01392_),
    .A(_01379_),
    .B(_01391_));
 sg13g2_xnor2_1 _07586_ (.Y(_01393_),
    .A(_01378_),
    .B(_01392_));
 sg13g2_inv_1 _07587_ (.Y(_01394_),
    .A(_01393_));
 sg13g2_nand2_1 _07588_ (.Y(_01395_),
    .A(_01376_),
    .B(_01394_));
 sg13g2_nand3_1 _07589_ (.B(_01375_),
    .C(_01393_),
    .A(_01372_),
    .Y(_01396_));
 sg13g2_nand2_1 _07590_ (.Y(_01397_),
    .A(_01395_),
    .B(_01396_));
 sg13g2_buf_8 _07591_ (.A(_01397_),
    .X(_01398_));
 sg13g2_nor2_1 _07592_ (.A(net101),
    .B(_01398_),
    .Y(_01399_));
 sg13g2_xnor2_1 _07593_ (.Y(_01400_),
    .A(_01296_),
    .B(_01281_));
 sg13g2_nand2_1 _07594_ (.Y(_01401_),
    .A(_01400_),
    .B(net68));
 sg13g2_nand2_1 _07595_ (.Y(_01402_),
    .A(_01399_),
    .B(_01401_));
 sg13g2_nand3_1 _07596_ (.B(_01396_),
    .C(net90),
    .A(_01395_),
    .Y(_01403_));
 sg13g2_nor2_1 _07597_ (.A(net62),
    .B(_01299_),
    .Y(_01404_));
 sg13g2_nand2_1 _07598_ (.Y(_01405_),
    .A(_01403_),
    .B(_01404_));
 sg13g2_nand2_1 _07599_ (.Y(_01406_),
    .A(_01402_),
    .B(_01405_));
 sg13g2_nor2_1 _07600_ (.A(net69),
    .B(_01204_),
    .Y(_01407_));
 sg13g2_nand2_1 _07601_ (.Y(_01408_),
    .A(_01406_),
    .B(_01407_));
 sg13g2_inv_1 _07602_ (.Y(_01409_),
    .A(_01407_));
 sg13g2_nand3_1 _07603_ (.B(_01405_),
    .C(_01409_),
    .A(_01402_),
    .Y(_01410_));
 sg13g2_nand2_1 _07604_ (.Y(_01411_),
    .A(_01408_),
    .B(_01410_));
 sg13g2_nand2b_1 _07605_ (.Y(_01412_),
    .B(_01411_),
    .A_N(_01364_));
 sg13g2_nand3_1 _07606_ (.B(_01410_),
    .C(_01364_),
    .A(_01408_),
    .Y(_01413_));
 sg13g2_nand2_1 _07607_ (.Y(_01414_),
    .A(_01412_),
    .B(_01413_));
 sg13g2_nor2_1 _07608_ (.A(net51),
    .B(_00903_),
    .Y(_01415_));
 sg13g2_nand2_1 _07609_ (.Y(_01416_),
    .A(_01208_),
    .B(net71));
 sg13g2_nor2_1 _07610_ (.A(_01312_),
    .B(_01416_),
    .Y(_01417_));
 sg13g2_nand2_1 _07611_ (.Y(_01418_),
    .A(_01416_),
    .B(_01312_));
 sg13g2_nor2b_1 _07612_ (.A(_01417_),
    .B_N(_01418_),
    .Y(_01419_));
 sg13g2_xor2_1 _07613_ (.B(_01419_),
    .A(_01415_),
    .X(_01420_));
 sg13g2_nand2_1 _07614_ (.Y(_01421_),
    .A(_01414_),
    .B(_01420_));
 sg13g2_inv_1 _07615_ (.Y(_01422_),
    .A(_01420_));
 sg13g2_nand3_1 _07616_ (.B(_01413_),
    .C(_01422_),
    .A(_01412_),
    .Y(_01423_));
 sg13g2_nand2_1 _07617_ (.Y(_01424_),
    .A(_01421_),
    .B(_01423_));
 sg13g2_nand2b_1 _07618_ (.Y(_01425_),
    .B(_01424_),
    .A_N(_01362_));
 sg13g2_nand3_1 _07619_ (.B(_01423_),
    .C(_01362_),
    .A(_01421_),
    .Y(_01426_));
 sg13g2_nand2_1 _07620_ (.Y(_01427_),
    .A(_01425_),
    .B(_01426_));
 sg13g2_inv_1 _07621_ (.Y(_01428_),
    .A(_00805_));
 sg13g2_nand2_1 _07622_ (.Y(_01429_),
    .A(_01428_),
    .B(_00223_));
 sg13g2_xnor2_1 _07623_ (.Y(_01430_),
    .A(_01325_),
    .B(_01429_));
 sg13g2_nor2_1 _07624_ (.A(_01223_),
    .B(_01313_),
    .Y(_01431_));
 sg13g2_a21oi_1 _07625_ (.A1(_01314_),
    .A2(_01311_),
    .Y(_01432_),
    .B1(_01431_));
 sg13g2_xnor2_1 _07626_ (.Y(_01433_),
    .A(_01430_),
    .B(_01432_));
 sg13g2_xnor2_1 _07627_ (.Y(_01434_),
    .A(_01326_),
    .B(_01433_));
 sg13g2_nand2_1 _07628_ (.Y(_01435_),
    .A(_01427_),
    .B(_01434_));
 sg13g2_inv_1 _07629_ (.Y(_01436_),
    .A(_01434_));
 sg13g2_nand3_1 _07630_ (.B(_01426_),
    .C(_01436_),
    .A(_01425_),
    .Y(_01437_));
 sg13g2_nand2_1 _07631_ (.Y(_01438_),
    .A(_01435_),
    .B(_01437_));
 sg13g2_nand2b_1 _07632_ (.Y(_01439_),
    .B(_01438_),
    .A_N(_01359_));
 sg13g2_nand3_1 _07633_ (.B(_01437_),
    .C(_01359_),
    .A(_01435_),
    .Y(_01440_));
 sg13g2_nand2_1 _07634_ (.Y(_01441_),
    .A(_01439_),
    .B(_01440_));
 sg13g2_nor2b_1 _07635_ (.A(_01331_),
    .B_N(_01330_),
    .Y(_01442_));
 sg13g2_a21oi_1 _07636_ (.A1(_01332_),
    .A2(_01324_),
    .Y(_01443_),
    .B1(_01442_));
 sg13g2_inv_1 _07637_ (.Y(_01444_),
    .A(_01443_));
 sg13g2_nand2_1 _07638_ (.Y(_01445_),
    .A(_01441_),
    .B(_01444_));
 sg13g2_nand3_1 _07639_ (.B(_01440_),
    .C(_01443_),
    .A(_01439_),
    .Y(_01446_));
 sg13g2_nand2_1 _07640_ (.Y(_01447_),
    .A(_01445_),
    .B(_01446_));
 sg13g2_nand2_1 _07641_ (.Y(_01448_),
    .A(_01337_),
    .B(_01266_));
 sg13g2_nor2_1 _07642_ (.A(_01266_),
    .B(_01337_),
    .Y(_01449_));
 sg13g2_a21oi_1 _07643_ (.A1(_01448_),
    .A2(_01343_),
    .Y(_01450_),
    .B1(_01449_));
 sg13g2_inv_1 _07644_ (.Y(_01451_),
    .A(_01450_));
 sg13g2_nand2_1 _07645_ (.Y(_01452_),
    .A(_01447_),
    .B(_01451_));
 sg13g2_nand3_1 _07646_ (.B(_01446_),
    .C(_01450_),
    .A(_01445_),
    .Y(_01453_));
 sg13g2_nand2_1 _07647_ (.Y(_01454_),
    .A(_01452_),
    .B(_01453_));
 sg13g2_nand2_1 _07648_ (.Y(_01455_),
    .A(_01356_),
    .B(_01454_));
 sg13g2_inv_1 _07649_ (.Y(_01456_),
    .A(_01454_));
 sg13g2_nand3_1 _07650_ (.B(_01456_),
    .C(_01355_),
    .A(_01350_),
    .Y(_01457_));
 sg13g2_nand2_1 _07651_ (.Y(_01458_),
    .A(_01455_),
    .B(_01457_));
 sg13g2_nand2_1 _07652_ (.Y(_01459_),
    .A(_01458_),
    .B(net64));
 sg13g2_xnor2_1 _07653_ (.Y(_01460_),
    .A(_00648_),
    .B(_00742_));
 sg13g2_xnor2_1 _07654_ (.Y(_01461_),
    .A(_00241_),
    .B(_00539_));
 sg13g2_nand2_1 _07655_ (.Y(_01462_),
    .A(_00645_),
    .B(_01461_));
 sg13g2_nand2_1 _07656_ (.Y(_01463_),
    .A(_01462_),
    .B(_00580_));
 sg13g2_o21ai_1 _07657_ (.B1(_00542_),
    .Y(_01464_),
    .A1(_00586_),
    .A2(_00644_));
 sg13g2_nand2_1 _07658_ (.Y(_01465_),
    .A(_01463_),
    .B(_01464_));
 sg13g2_nor2_1 _07659_ (.A(_01460_),
    .B(_01465_),
    .Y(_01466_));
 sg13g2_inv_1 _07660_ (.Y(_01467_),
    .A(_00859_));
 sg13g2_nand2_1 _07661_ (.Y(_01468_),
    .A(_01466_),
    .B(_01467_));
 sg13g2_o21ai_1 _07662_ (.B1(_00856_),
    .Y(_01469_),
    .A1(_00743_),
    .A2(_00963_));
 sg13g2_nand2_1 _07663_ (.Y(_01470_),
    .A(_01468_),
    .B(_01469_));
 sg13g2_nor2_1 _07664_ (.A(_00960_),
    .B(_01060_),
    .Y(_01471_));
 sg13g2_nand2_1 _07665_ (.Y(_01472_),
    .A(_01470_),
    .B(_01471_));
 sg13g2_nand2_1 _07666_ (.Y(_01473_),
    .A(_01057_),
    .B(_00957_));
 sg13g2_nand2_1 _07667_ (.Y(_01474_),
    .A(_01473_),
    .B(_01059_));
 sg13g2_nand2_1 _07668_ (.Y(_01475_),
    .A(_01472_),
    .B(_01474_));
 sg13g2_inv_1 _07669_ (.Y(_01476_),
    .A(_01150_));
 sg13g2_nand2_1 _07670_ (.Y(_01477_),
    .A(_01260_),
    .B(_01476_));
 sg13g2_inv_1 _07671_ (.Y(_01478_),
    .A(_01477_));
 sg13g2_nand2_1 _07672_ (.Y(_01479_),
    .A(_01475_),
    .B(_01478_));
 sg13g2_a21oi_1 _07673_ (.A1(_01259_),
    .A2(_01157_),
    .Y(_01480_),
    .B1(_01147_));
 sg13g2_nor2b_1 _07674_ (.A(_01480_),
    .B_N(_01352_),
    .Y(_01481_));
 sg13g2_nand2_1 _07675_ (.Y(_01482_),
    .A(_01479_),
    .B(_01481_));
 sg13g2_xnor2_1 _07676_ (.Y(_01483_),
    .A(_01347_),
    .B(_01482_));
 sg13g2_nand2_1 _07677_ (.Y(_01484_),
    .A(_01483_),
    .B(net70));
 sg13g2_nand2_1 _07678_ (.Y(_01485_),
    .A(_01459_),
    .B(_01484_));
 sg13g2_inv_2 _07679_ (.Y(_01486_),
    .A(_03673_));
 sg13g2_buf_1 _07680_ (.A(_01486_),
    .X(_01487_));
 sg13g2_nand2_1 _07681_ (.Y(_01488_),
    .A(_01485_),
    .B(net67));
 sg13g2_xnor2_1 _07682_ (.Y(_01489_),
    .A(_01261_),
    .B(_01155_));
 sg13g2_xnor2_1 _07683_ (.Y(_01490_),
    .A(_01150_),
    .B(_01475_));
 sg13g2_inv_1 _07684_ (.Y(_01491_),
    .A(_01490_));
 sg13g2_nor2_1 _07685_ (.A(net64),
    .B(_01491_),
    .Y(_01492_));
 sg13g2_a21oi_1 _07686_ (.A1(net64),
    .A2(_01489_),
    .Y(_01493_),
    .B1(_01492_));
 sg13g2_nand2_1 _07687_ (.Y(_01494_),
    .A(_01493_),
    .B(net78));
 sg13g2_nand3_1 _07688_ (.B(_03965_),
    .C(_01494_),
    .A(_01488_),
    .Y(_01495_));
 sg13g2_xnor2_1 _07689_ (.Y(_01496_),
    .A(_01060_),
    .B(_00966_));
 sg13g2_xnor2_1 _07690_ (.Y(_01497_),
    .A(_00960_),
    .B(_01470_));
 sg13g2_nor2b_1 _07691_ (.A(net64),
    .B_N(_01497_),
    .Y(_01498_));
 sg13g2_a21oi_1 _07692_ (.A1(net64),
    .A2(_01496_),
    .Y(_01499_),
    .B1(_01498_));
 sg13g2_nand2_1 _07693_ (.Y(_01500_),
    .A(_01499_),
    .B(net67));
 sg13g2_inv_2 _07694_ (.Y(_01501_),
    .A(_03965_));
 sg13g2_buf_1 _07695_ (.A(net64),
    .X(_01502_));
 sg13g2_xnor2_1 _07696_ (.Y(_01503_),
    .A(_01460_),
    .B(_01465_));
 sg13g2_xnor2_1 _07697_ (.Y(_01504_),
    .A(_00859_),
    .B(_00747_));
 sg13g2_a21oi_1 _07698_ (.A1(_01504_),
    .A2(net56),
    .Y(_01505_),
    .B1(_01486_));
 sg13g2_o21ai_1 _07699_ (.B1(_01505_),
    .Y(_01506_),
    .A1(net56),
    .A2(_01503_));
 sg13g2_nand3_1 _07700_ (.B(_01501_),
    .C(_01506_),
    .A(_01500_),
    .Y(_01507_));
 sg13g2_nand2_1 _07701_ (.Y(_01508_),
    .A(_01495_),
    .B(_01507_));
 sg13g2_buf_8 _07702_ (.A(_01508_),
    .X(_01509_));
 sg13g2_inv_4 _07703_ (.A(_01509_),
    .Y(_01510_));
 sg13g2_nand2_1 _07704_ (.Y(_01511_),
    .A(_01454_),
    .B(_01347_));
 sg13g2_inv_1 _07705_ (.Y(_01512_),
    .A(_01328_));
 sg13g2_nand2_1 _07706_ (.Y(_01513_),
    .A(_01428_),
    .B(net50));
 sg13g2_nor2_1 _07707_ (.A(_01512_),
    .B(_01513_),
    .Y(_01514_));
 sg13g2_nor2_1 _07708_ (.A(net49),
    .B(_00903_),
    .Y(_01515_));
 sg13g2_xnor2_1 _07709_ (.Y(_01516_),
    .A(_01515_),
    .B(_01513_));
 sg13g2_a21oi_1 _07710_ (.A1(_01418_),
    .A2(_01415_),
    .Y(_01517_),
    .B1(_01417_));
 sg13g2_xnor2_1 _07711_ (.Y(_01518_),
    .A(_01516_),
    .B(_01517_));
 sg13g2_xor2_1 _07712_ (.B(_01518_),
    .A(_01514_),
    .X(_01519_));
 sg13g2_nand2_1 _07713_ (.Y(_01520_),
    .A(_01401_),
    .B(_01403_));
 sg13g2_nor2_1 _07714_ (.A(_01403_),
    .B(_01401_),
    .Y(_01521_));
 sg13g2_a21oi_2 _07715_ (.B1(_01521_),
    .Y(_01522_),
    .A2(_01407_),
    .A1(_01520_));
 sg13g2_inv_1 _07716_ (.Y(_01523_),
    .A(\r2[16] ));
 sg13g2_nand2_1 _07717_ (.Y(_01524_),
    .A(_01391_),
    .B(_01523_));
 sg13g2_buf_1 _07718_ (.A(\r1[15] ),
    .X(_01525_));
 sg13g2_nor4_1 _07719_ (.A(_01380_),
    .B(_01525_),
    .C(_01286_),
    .D(_00873_),
    .Y(_01526_));
 sg13g2_nand2_1 _07720_ (.Y(_01527_),
    .A(_01074_),
    .B(_01526_));
 sg13g2_nand2_1 _07721_ (.Y(_01528_),
    .A(_01527_),
    .B(_00014_));
 sg13g2_inv_1 _07722_ (.Y(_01529_),
    .A(_00014_));
 sg13g2_nand3_1 _07723_ (.B(_01526_),
    .C(_01529_),
    .A(_01074_),
    .Y(_01530_));
 sg13g2_nand2_1 _07724_ (.Y(_01531_),
    .A(_01528_),
    .B(_01530_));
 sg13g2_nand2b_1 _07725_ (.Y(_01532_),
    .B(_01531_),
    .A_N(_00013_));
 sg13g2_nand3_1 _07726_ (.B(_01530_),
    .C(_00013_),
    .A(_01528_),
    .Y(_01533_));
 sg13g2_nand2_1 _07727_ (.Y(_01534_),
    .A(_01532_),
    .B(_01533_));
 sg13g2_nand2b_1 _07728_ (.Y(_01535_),
    .B(_01534_),
    .A_N(_01524_));
 sg13g2_nand3_1 _07729_ (.B(_01524_),
    .C(_01533_),
    .A(_01532_),
    .Y(_01536_));
 sg13g2_buf_2 _07730_ (.A(_01536_),
    .X(_01537_));
 sg13g2_nand2_2 _07731_ (.Y(_01538_),
    .A(_01535_),
    .B(_01537_));
 sg13g2_nand2_1 _07732_ (.Y(_01539_),
    .A(_01394_),
    .B(_01291_));
 sg13g2_nor2b_1 _07733_ (.A(_01539_),
    .B_N(_01273_),
    .Y(_01540_));
 sg13g2_nand2_1 _07734_ (.Y(_01541_),
    .A(_01095_),
    .B(_01540_));
 sg13g2_inv_1 _07735_ (.Y(_01542_),
    .A(_01539_));
 sg13g2_inv_1 _07736_ (.Y(_01543_),
    .A(_01278_));
 sg13g2_nand2_1 _07737_ (.Y(_01544_),
    .A(_01392_),
    .B(_01378_));
 sg13g2_nor2_1 _07738_ (.A(_01378_),
    .B(_01392_),
    .Y(_01545_));
 sg13g2_a21oi_1 _07739_ (.A1(_01293_),
    .A2(_01544_),
    .Y(_01546_),
    .B1(_01545_));
 sg13g2_a21oi_1 _07740_ (.A1(_01542_),
    .A2(_01543_),
    .Y(_01547_),
    .B1(_01546_));
 sg13g2_nand2_1 _07741_ (.Y(_01548_),
    .A(_01541_),
    .B(_01547_));
 sg13g2_xnor2_1 _07742_ (.Y(_01549_),
    .A(_01538_),
    .B(_01548_));
 sg13g2_nand3_1 _07743_ (.B(_01396_),
    .C(net68),
    .A(_01395_),
    .Y(_01550_));
 sg13g2_buf_1 _07744_ (.A(_01550_),
    .X(_01551_));
 sg13g2_nand3_1 _07745_ (.B(_01551_),
    .C(net90),
    .A(_01549_),
    .Y(_01552_));
 sg13g2_inv_1 _07746_ (.Y(_01553_),
    .A(_01538_));
 sg13g2_nand2_1 _07747_ (.Y(_01554_),
    .A(_01548_),
    .B(_01553_));
 sg13g2_nand3_1 _07748_ (.B(_01547_),
    .C(_01538_),
    .A(_01541_),
    .Y(_01555_));
 sg13g2_nand3_1 _07749_ (.B(_01555_),
    .C(net90),
    .A(_01554_),
    .Y(_01556_));
 sg13g2_buf_1 _07750_ (.A(_01556_),
    .X(_01557_));
 sg13g2_nand2b_1 _07751_ (.Y(_01558_),
    .B(_01557_),
    .A_N(_01551_));
 sg13g2_nand2_1 _07752_ (.Y(_01559_),
    .A(_01552_),
    .B(_01558_));
 sg13g2_nor2_1 _07753_ (.A(net69),
    .B(_01299_),
    .Y(_01560_));
 sg13g2_nand2_1 _07754_ (.Y(_01561_),
    .A(_01559_),
    .B(_01560_));
 sg13g2_inv_1 _07755_ (.Y(_01562_),
    .A(_01560_));
 sg13g2_nand3_1 _07756_ (.B(_01558_),
    .C(_01562_),
    .A(_01552_),
    .Y(_01563_));
 sg13g2_nand2_1 _07757_ (.Y(_01564_),
    .A(_01561_),
    .B(_01563_));
 sg13g2_nand2b_1 _07758_ (.Y(_01565_),
    .B(_01564_),
    .A_N(_01522_));
 sg13g2_nand3_1 _07759_ (.B(_01563_),
    .C(_01522_),
    .A(_01561_),
    .Y(_01566_));
 sg13g2_nand2_1 _07760_ (.Y(_01567_),
    .A(_01565_),
    .B(_01566_));
 sg13g2_nor2_1 _07761_ (.A(net44),
    .B(_01005_),
    .Y(_01568_));
 sg13g2_inv_1 _07762_ (.Y(_01569_),
    .A(_01204_));
 sg13g2_nand2_1 _07763_ (.Y(_01570_),
    .A(_01569_),
    .B(net65));
 sg13g2_nor2_1 _07764_ (.A(_01416_),
    .B(_01570_),
    .Y(_01571_));
 sg13g2_nor2_1 _07765_ (.A(net57),
    .B(_01204_),
    .Y(_01572_));
 sg13g2_inv_1 _07766_ (.Y(_01573_),
    .A(_01572_));
 sg13g2_o21ai_1 _07767_ (.B1(_01573_),
    .Y(_01574_),
    .A1(_01099_),
    .A2(net63));
 sg13g2_nand2b_1 _07768_ (.Y(_01575_),
    .B(_01574_),
    .A_N(_01571_));
 sg13g2_xor2_1 _07769_ (.B(_01575_),
    .A(_01568_),
    .X(_01576_));
 sg13g2_inv_1 _07770_ (.Y(_01577_),
    .A(_01576_));
 sg13g2_nand2_1 _07771_ (.Y(_01578_),
    .A(_01567_),
    .B(_01577_));
 sg13g2_nand3_1 _07772_ (.B(_01566_),
    .C(_01576_),
    .A(_01565_),
    .Y(_01579_));
 sg13g2_nand2_1 _07773_ (.Y(_01580_),
    .A(_01578_),
    .B(_01579_));
 sg13g2_nand2_1 _07774_ (.Y(_01581_),
    .A(_01411_),
    .B(_01364_));
 sg13g2_nor2_1 _07775_ (.A(_01364_),
    .B(_01411_),
    .Y(_01582_));
 sg13g2_a21oi_2 _07776_ (.B1(_01582_),
    .Y(_01583_),
    .A2(_01420_),
    .A1(_01581_));
 sg13g2_inv_1 _07777_ (.Y(_01584_),
    .A(_01583_));
 sg13g2_nand2_1 _07778_ (.Y(_01585_),
    .A(_01580_),
    .B(_01584_));
 sg13g2_nand3_1 _07779_ (.B(_01579_),
    .C(_01583_),
    .A(_01578_),
    .Y(_01586_));
 sg13g2_nand3b_1 _07780_ (.B(_01585_),
    .C(_01586_),
    .Y(_01587_),
    .A_N(_01519_));
 sg13g2_nand2_1 _07781_ (.Y(_01588_),
    .A(_01585_),
    .B(_01586_));
 sg13g2_nand2_1 _07782_ (.Y(_01589_),
    .A(_01588_),
    .B(_01519_));
 sg13g2_nand2_1 _07783_ (.Y(_01590_),
    .A(_01587_),
    .B(_01589_));
 sg13g2_nand2_1 _07784_ (.Y(_01591_),
    .A(_01424_),
    .B(_01362_));
 sg13g2_nor2_1 _07785_ (.A(_01362_),
    .B(_01424_),
    .Y(_01592_));
 sg13g2_a21oi_2 _07786_ (.B1(_01592_),
    .Y(_01593_),
    .A2(_01434_),
    .A1(_01591_));
 sg13g2_nand2_1 _07787_ (.Y(_01594_),
    .A(_01590_),
    .B(_01593_));
 sg13g2_nor2b_1 _07788_ (.A(_01432_),
    .B_N(_01430_),
    .Y(_01595_));
 sg13g2_a21oi_1 _07789_ (.A1(_01433_),
    .A2(_01327_),
    .Y(_01596_),
    .B1(_01595_));
 sg13g2_inv_1 _07790_ (.Y(_01597_),
    .A(_01596_));
 sg13g2_nor2_1 _07791_ (.A(_01593_),
    .B(_01590_),
    .Y(_01598_));
 sg13g2_a21oi_1 _07792_ (.A1(_01594_),
    .A2(_01597_),
    .Y(_01599_),
    .B1(_01598_));
 sg13g2_nand2_1 _07793_ (.Y(_01600_),
    .A(_01580_),
    .B(_01583_));
 sg13g2_nor2_1 _07794_ (.A(_01583_),
    .B(_01580_),
    .Y(_01601_));
 sg13g2_a21oi_2 _07795_ (.B1(_01601_),
    .Y(_01602_),
    .A2(_01519_),
    .A1(_01600_));
 sg13g2_nor2_1 _07796_ (.A(net45),
    .B(_00903_),
    .Y(_01603_));
 sg13g2_inv_1 _07797_ (.Y(_01604_),
    .A(_01603_));
 sg13g2_nor2_1 _07798_ (.A(_01604_),
    .B(_01429_),
    .Y(_01605_));
 sg13g2_nand2_1 _07799_ (.Y(_01606_),
    .A(_01008_),
    .B(net50));
 sg13g2_nor2b_1 _07800_ (.A(_01606_),
    .B_N(_01515_),
    .Y(_01607_));
 sg13g2_nor2_1 _07801_ (.A(net49),
    .B(_01005_),
    .Y(_01608_));
 sg13g2_nor2_1 _07802_ (.A(_01603_),
    .B(_01608_),
    .Y(_01609_));
 sg13g2_nor2_1 _07803_ (.A(_01607_),
    .B(_01609_),
    .Y(_01610_));
 sg13g2_a21oi_1 _07804_ (.A1(_01574_),
    .A2(_01568_),
    .Y(_01611_),
    .B1(_01571_));
 sg13g2_xnor2_1 _07805_ (.Y(_01612_),
    .A(_01610_),
    .B(_01611_));
 sg13g2_xor2_1 _07806_ (.B(_01612_),
    .A(_01605_),
    .X(_01613_));
 sg13g2_nand2_1 _07807_ (.Y(_01614_),
    .A(_01564_),
    .B(_01522_));
 sg13g2_nor2_1 _07808_ (.A(_01522_),
    .B(_01564_),
    .Y(_01615_));
 sg13g2_a21oi_2 _07809_ (.B1(_01615_),
    .Y(_01616_),
    .A2(_01577_),
    .A1(_01614_));
 sg13g2_nand2_1 _07810_ (.Y(_01617_),
    .A(_01557_),
    .B(_01551_));
 sg13g2_nor2_1 _07811_ (.A(_01551_),
    .B(_01557_),
    .Y(_01618_));
 sg13g2_a21oi_2 _07812_ (.B1(_01618_),
    .Y(_01619_),
    .A2(_01560_),
    .A1(_01617_));
 sg13g2_nor2_1 _07813_ (.A(net69),
    .B(_01398_),
    .Y(_01620_));
 sg13g2_nand2_1 _07814_ (.Y(_01621_),
    .A(_01549_),
    .B(net68));
 sg13g2_nand2_1 _07815_ (.Y(_01622_),
    .A(_01197_),
    .B(_01291_));
 sg13g2_nor2_1 _07816_ (.A(_01538_),
    .B(_01393_),
    .Y(_01623_));
 sg13g2_nor2b_1 _07817_ (.A(_01622_),
    .B_N(_01623_),
    .Y(_01624_));
 sg13g2_nand4_1 _07818_ (.B(_01624_),
    .C(_01167_),
    .A(_00773_),
    .Y(_01625_),
    .D(_00997_));
 sg13g2_o21ai_1 _07819_ (.B1(_01537_),
    .Y(_01626_),
    .A1(_01544_),
    .A2(_01538_));
 sg13g2_nand2_1 _07820_ (.Y(_01627_),
    .A(_01366_),
    .B(_01623_));
 sg13g2_nand2b_1 _07821_ (.Y(_01628_),
    .B(_01627_),
    .A_N(_01626_));
 sg13g2_a21oi_1 _07822_ (.A1(_01169_),
    .A2(_01624_),
    .Y(_01629_),
    .B1(_01628_));
 sg13g2_nand2_1 _07823_ (.Y(_01630_),
    .A(_01625_),
    .B(_01629_));
 sg13g2_inv_1 _07824_ (.Y(_01631_),
    .A(\r2[17] ));
 sg13g2_nand2_1 _07825_ (.Y(_01632_),
    .A(_01531_),
    .B(_01631_));
 sg13g2_buf_1 _07826_ (.A(_00016_),
    .X(_01633_));
 sg13g2_xor2_1 _07827_ (.B(_00015_),
    .A(_01633_),
    .X(_01634_));
 sg13g2_nor2_1 _07828_ (.A(_01380_),
    .B(_01525_),
    .Y(_01635_));
 sg13g2_buf_1 _07829_ (.A(\r1[16] ),
    .X(_01636_));
 sg13g2_inv_1 _07830_ (.Y(_01637_),
    .A(_01636_));
 sg13g2_nand3_1 _07831_ (.B(_01382_),
    .C(_01637_),
    .A(_01635_),
    .Y(_01638_));
 sg13g2_nor3_1 _07832_ (.A(_01181_),
    .B(_01638_),
    .C(_00975_),
    .Y(_01639_));
 sg13g2_nand2_1 _07833_ (.Y(_01640_),
    .A(_00782_),
    .B(_01639_));
 sg13g2_nor3_1 _07834_ (.A(_01181_),
    .B(_01638_),
    .C(_00979_),
    .Y(_01641_));
 sg13g2_nand2_1 _07835_ (.Y(_01642_),
    .A(_01640_),
    .B(_01641_));
 sg13g2_xnor2_1 _07836_ (.Y(_01643_),
    .A(_01634_),
    .B(_01642_));
 sg13g2_xnor2_1 _07837_ (.Y(_01644_),
    .A(_01632_),
    .B(_01643_));
 sg13g2_nand2_1 _07838_ (.Y(_01645_),
    .A(_01630_),
    .B(_01644_));
 sg13g2_inv_1 _07839_ (.Y(_01646_),
    .A(_01644_));
 sg13g2_nand3_1 _07840_ (.B(_01629_),
    .C(_01646_),
    .A(_01625_),
    .Y(_01647_));
 sg13g2_nand2_1 _07841_ (.Y(_01648_),
    .A(_01645_),
    .B(_01647_));
 sg13g2_buf_8 _07842_ (.A(_01648_),
    .X(_01649_));
 sg13g2_nor2_1 _07843_ (.A(_00412_),
    .B(_01649_),
    .Y(_01650_));
 sg13g2_nand2_1 _07844_ (.Y(_01651_),
    .A(_01621_),
    .B(_01650_));
 sg13g2_nand2_2 _07845_ (.Y(_01652_),
    .A(_01554_),
    .B(_01555_));
 sg13g2_nor2_1 _07846_ (.A(net62),
    .B(_01652_),
    .Y(_01653_));
 sg13g2_nand3_1 _07847_ (.B(_01647_),
    .C(_01009_),
    .A(_01645_),
    .Y(_01654_));
 sg13g2_nand2_1 _07848_ (.Y(_01655_),
    .A(_01653_),
    .B(_01654_));
 sg13g2_nand3b_1 _07849_ (.B(_01651_),
    .C(_01655_),
    .Y(_01656_),
    .A_N(_01620_));
 sg13g2_nand2_1 _07850_ (.Y(_01657_),
    .A(_01651_),
    .B(_01655_));
 sg13g2_nand2_1 _07851_ (.Y(_01658_),
    .A(_01657_),
    .B(_01620_));
 sg13g2_nand2_1 _07852_ (.Y(_01659_),
    .A(_01656_),
    .B(_01658_));
 sg13g2_nand2b_1 _07853_ (.Y(_01660_),
    .B(_01659_),
    .A_N(_01619_));
 sg13g2_nand3_1 _07854_ (.B(_01658_),
    .C(_01619_),
    .A(_01656_),
    .Y(_01661_));
 sg13g2_nand2_1 _07855_ (.Y(_01662_),
    .A(_01660_),
    .B(_01661_));
 sg13g2_nor2_1 _07856_ (.A(net44),
    .B(_01099_),
    .Y(_01663_));
 sg13g2_nor2_1 _07857_ (.A(net63),
    .B(_01299_),
    .Y(_01664_));
 sg13g2_inv_1 _07858_ (.Y(_01665_),
    .A(_01664_));
 sg13g2_nand2_1 _07859_ (.Y(_01666_),
    .A(_01400_),
    .B(net71));
 sg13g2_nand2_1 _07860_ (.Y(_01667_),
    .A(_01666_),
    .B(_01570_));
 sg13g2_o21ai_1 _07861_ (.B1(_01667_),
    .Y(_01668_),
    .A1(_01665_),
    .A2(_01573_));
 sg13g2_xnor2_1 _07862_ (.Y(_01669_),
    .A(_01663_),
    .B(_01668_));
 sg13g2_nand2_1 _07863_ (.Y(_01670_),
    .A(_01662_),
    .B(_01669_));
 sg13g2_inv_1 _07864_ (.Y(_01671_),
    .A(_01669_));
 sg13g2_nand3_1 _07865_ (.B(_01661_),
    .C(_01671_),
    .A(_01660_),
    .Y(_01672_));
 sg13g2_nand2_1 _07866_ (.Y(_01673_),
    .A(_01670_),
    .B(_01672_));
 sg13g2_nand2b_1 _07867_ (.Y(_01674_),
    .B(_01673_),
    .A_N(_01616_));
 sg13g2_nand3_1 _07868_ (.B(_01672_),
    .C(_01616_),
    .A(_01670_),
    .Y(_01675_));
 sg13g2_nand3b_1 _07869_ (.B(_01674_),
    .C(_01675_),
    .Y(_01676_),
    .A_N(_01613_));
 sg13g2_nand2_1 _07870_ (.Y(_01677_),
    .A(_01674_),
    .B(_01675_));
 sg13g2_nand2_1 _07871_ (.Y(_01678_),
    .A(_01677_),
    .B(_01613_));
 sg13g2_nand2_1 _07872_ (.Y(_01679_),
    .A(_01676_),
    .B(_01678_));
 sg13g2_nand2b_1 _07873_ (.Y(_01680_),
    .B(_01679_),
    .A_N(_01602_));
 sg13g2_nand3_1 _07874_ (.B(_01678_),
    .C(_01602_),
    .A(_01676_),
    .Y(_01681_));
 sg13g2_nand2_1 _07875_ (.Y(_01682_),
    .A(_01680_),
    .B(_01681_));
 sg13g2_nor2b_1 _07876_ (.A(_01517_),
    .B_N(_01516_),
    .Y(_01683_));
 sg13g2_a21oi_1 _07877_ (.A1(_01518_),
    .A2(_01514_),
    .Y(_01684_),
    .B1(_01683_));
 sg13g2_inv_1 _07878_ (.Y(_01685_),
    .A(_01684_));
 sg13g2_nand2_1 _07879_ (.Y(_01686_),
    .A(_01682_),
    .B(_01685_));
 sg13g2_nand3_1 _07880_ (.B(_01681_),
    .C(_01684_),
    .A(_01680_),
    .Y(_01687_));
 sg13g2_nand2_1 _07881_ (.Y(_01688_),
    .A(_01686_),
    .B(_01687_));
 sg13g2_nor2_1 _07882_ (.A(_01599_),
    .B(_01688_),
    .Y(_01689_));
 sg13g2_inv_1 _07883_ (.Y(_01690_),
    .A(_01599_));
 sg13g2_a21oi_1 _07884_ (.A1(_01686_),
    .A2(_01687_),
    .Y(_01691_),
    .B1(_01690_));
 sg13g2_nor2_1 _07885_ (.A(_01689_),
    .B(_01691_),
    .Y(_01692_));
 sg13g2_nand2_1 _07886_ (.Y(_01693_),
    .A(_01438_),
    .B(_01359_));
 sg13g2_nor2_1 _07887_ (.A(_01359_),
    .B(_01438_),
    .Y(_01694_));
 sg13g2_a21oi_1 _07888_ (.A1(_01693_),
    .A2(_01444_),
    .Y(_01695_),
    .B1(_01694_));
 sg13g2_inv_1 _07889_ (.Y(_01696_),
    .A(_01695_));
 sg13g2_nand2b_1 _07890_ (.Y(_01697_),
    .B(_01590_),
    .A_N(_01593_));
 sg13g2_nand3_1 _07891_ (.B(_01589_),
    .C(_01593_),
    .A(_01587_),
    .Y(_01698_));
 sg13g2_nand2_1 _07892_ (.Y(_01699_),
    .A(_01697_),
    .B(_01698_));
 sg13g2_nand2_1 _07893_ (.Y(_01700_),
    .A(_01699_),
    .B(_01597_));
 sg13g2_nand3_1 _07894_ (.B(_01698_),
    .C(_01596_),
    .A(_01697_),
    .Y(_01701_));
 sg13g2_nand2_1 _07895_ (.Y(_01702_),
    .A(_01700_),
    .B(_01701_));
 sg13g2_xnor2_1 _07896_ (.Y(_01703_),
    .A(_01696_),
    .B(_01702_));
 sg13g2_nand2_1 _07897_ (.Y(_01704_),
    .A(_01692_),
    .B(_01703_));
 sg13g2_nor2_1 _07898_ (.A(_01511_),
    .B(_01704_),
    .Y(_01705_));
 sg13g2_nand2_1 _07899_ (.Y(_01706_),
    .A(_01482_),
    .B(_01705_));
 sg13g2_nand2_1 _07900_ (.Y(_01707_),
    .A(_01702_),
    .B(_01695_));
 sg13g2_nand3_1 _07901_ (.B(_01701_),
    .C(_01696_),
    .A(_01700_),
    .Y(_01708_));
 sg13g2_buf_1 _07902_ (.A(_01708_),
    .X(_01709_));
 sg13g2_nand2_1 _07903_ (.Y(_01710_),
    .A(_01707_),
    .B(_01709_));
 sg13g2_nand3_1 _07904_ (.B(_01686_),
    .C(_01687_),
    .A(_01690_),
    .Y(_01711_));
 sg13g2_nand2_1 _07905_ (.Y(_01712_),
    .A(_01688_),
    .B(_01599_));
 sg13g2_nand2_1 _07906_ (.Y(_01713_),
    .A(_01711_),
    .B(_01712_));
 sg13g2_nor2_1 _07907_ (.A(_01710_),
    .B(_01713_),
    .Y(_01714_));
 sg13g2_nand3_1 _07908_ (.B(_01445_),
    .C(_01446_),
    .A(_01451_),
    .Y(_01715_));
 sg13g2_nand2_1 _07909_ (.Y(_01716_),
    .A(_01447_),
    .B(_01450_));
 sg13g2_inv_1 _07910_ (.Y(_01717_),
    .A(_01716_));
 sg13g2_a21oi_1 _07911_ (.A1(_01715_),
    .A2(_01351_),
    .Y(_01718_),
    .B1(_01717_));
 sg13g2_nand2_1 _07912_ (.Y(_01719_),
    .A(_01711_),
    .B(_01709_));
 sg13g2_nand2_1 _07913_ (.Y(_01720_),
    .A(_01719_),
    .B(_01712_));
 sg13g2_inv_1 _07914_ (.Y(_01721_),
    .A(_01720_));
 sg13g2_a21oi_1 _07915_ (.A1(_01714_),
    .A2(_01718_),
    .Y(_01722_),
    .B1(_01721_));
 sg13g2_nand2_1 _07916_ (.Y(_01723_),
    .A(_01706_),
    .B(_01722_));
 sg13g2_nand2_1 _07917_ (.Y(_01724_),
    .A(_01679_),
    .B(_01602_));
 sg13g2_nor2_1 _07918_ (.A(_01602_),
    .B(_01679_),
    .Y(_01725_));
 sg13g2_a21oi_1 _07919_ (.A1(_01724_),
    .A2(_01685_),
    .Y(_01726_),
    .B1(_01725_));
 sg13g2_nand2_1 _07920_ (.Y(_01727_),
    .A(_01673_),
    .B(_01616_));
 sg13g2_nor2_1 _07921_ (.A(_01616_),
    .B(_01673_),
    .Y(_01728_));
 sg13g2_a21oi_1 _07922_ (.A1(_01727_),
    .A2(_01613_),
    .Y(_01729_),
    .B1(_01728_));
 sg13g2_nand2_1 _07923_ (.Y(_01730_),
    .A(_01659_),
    .B(_01619_));
 sg13g2_nor2_1 _07924_ (.A(_01619_),
    .B(_01659_),
    .Y(_01731_));
 sg13g2_a21oi_1 _07925_ (.A1(_01730_),
    .A2(_01669_),
    .Y(_01732_),
    .B1(_01731_));
 sg13g2_nand2_1 _07926_ (.Y(_01733_),
    .A(_01621_),
    .B(_01654_));
 sg13g2_nand3_1 _07927_ (.B(_01647_),
    .C(_00610_),
    .A(_01645_),
    .Y(_01734_));
 sg13g2_nor2_1 _07928_ (.A(_01557_),
    .B(_01734_),
    .Y(_01735_));
 sg13g2_a21oi_2 _07929_ (.B1(_01735_),
    .Y(_01736_),
    .A2(_01620_),
    .A1(_01733_));
 sg13g2_nor2_1 _07930_ (.A(_00555_),
    .B(_01652_),
    .Y(_01737_));
 sg13g2_nand3_1 _07931_ (.B(_01535_),
    .C(_01537_),
    .A(_01644_),
    .Y(_01738_));
 sg13g2_nor2_1 _07932_ (.A(_01738_),
    .B(_01539_),
    .Y(_01739_));
 sg13g2_nand4_1 _07933_ (.B(_01739_),
    .C(_01089_),
    .A(_00899_),
    .Y(_01740_),
    .D(_01273_));
 sg13g2_nand2b_1 _07934_ (.Y(_01741_),
    .B(_01632_),
    .A_N(_01643_));
 sg13g2_o21ai_1 _07935_ (.B1(_01741_),
    .Y(_01742_),
    .A1(_01537_),
    .A2(_01646_));
 sg13g2_nand2b_1 _07936_ (.Y(_01743_),
    .B(_01546_),
    .A_N(_01738_));
 sg13g2_nand2b_1 _07937_ (.Y(_01744_),
    .B(_01743_),
    .A_N(_01742_));
 sg13g2_a21oi_1 _07938_ (.A1(_01279_),
    .A2(_01739_),
    .Y(_01745_),
    .B1(_01744_));
 sg13g2_nand2_1 _07939_ (.Y(_01746_),
    .A(_01740_),
    .B(_01745_));
 sg13g2_buf_1 _07940_ (.A(\r1[17] ),
    .X(_01747_));
 sg13g2_nor3_1 _07941_ (.A(_01636_),
    .B(_01747_),
    .C(_01527_),
    .Y(_01748_));
 sg13g2_xnor2_1 _07942_ (.Y(_01749_),
    .A(_01634_),
    .B(_01748_));
 sg13g2_inv_1 _07943_ (.Y(_01750_),
    .A(_01633_));
 sg13g2_a21oi_1 _07944_ (.A1(_01642_),
    .A2(_01750_),
    .Y(_01751_),
    .B1(\r2[18] ));
 sg13g2_o21ai_1 _07945_ (.B1(_01751_),
    .Y(_01752_),
    .A1(_01750_),
    .A2(_01642_));
 sg13g2_xor2_1 _07946_ (.B(_01752_),
    .A(_01749_),
    .X(_01753_));
 sg13g2_nand2_1 _07947_ (.Y(_01754_),
    .A(_01746_),
    .B(_01753_));
 sg13g2_inv_1 _07948_ (.Y(_01755_),
    .A(_01753_));
 sg13g2_nand3_1 _07949_ (.B(_01745_),
    .C(_01755_),
    .A(_01740_),
    .Y(_01756_));
 sg13g2_nand2_1 _07950_ (.Y(_01757_),
    .A(_01754_),
    .B(_01756_));
 sg13g2_nor2_1 _07951_ (.A(net62),
    .B(_01757_),
    .Y(_01758_));
 sg13g2_nand2_1 _07952_ (.Y(_01759_),
    .A(_01650_),
    .B(_01758_));
 sg13g2_nand3_1 _07953_ (.B(_01756_),
    .C(_01009_),
    .A(_01754_),
    .Y(_01760_));
 sg13g2_nand2_1 _07954_ (.Y(_01761_),
    .A(_01734_),
    .B(_01760_));
 sg13g2_nand2_1 _07955_ (.Y(_01762_),
    .A(_01759_),
    .B(_01761_));
 sg13g2_nand2b_1 _07956_ (.Y(_01763_),
    .B(_01762_),
    .A_N(_01737_));
 sg13g2_nand3_1 _07957_ (.B(_01761_),
    .C(_01737_),
    .A(_01759_),
    .Y(_01764_));
 sg13g2_nand2_1 _07958_ (.Y(_01765_),
    .A(_01763_),
    .B(_01764_));
 sg13g2_nand2b_1 _07959_ (.Y(_01766_),
    .B(_01765_),
    .A_N(_01736_));
 sg13g2_nand3_1 _07960_ (.B(_01763_),
    .C(_01764_),
    .A(_01736_),
    .Y(_01767_));
 sg13g2_nand2_1 _07961_ (.Y(_01768_),
    .A(_01766_),
    .B(_01767_));
 sg13g2_nor2_1 _07962_ (.A(net44),
    .B(_01204_),
    .Y(_01769_));
 sg13g2_inv_2 _07963_ (.Y(_01770_),
    .A(_01398_));
 sg13g2_nand2_1 _07964_ (.Y(_01771_),
    .A(_01770_),
    .B(_00193_));
 sg13g2_nor2_1 _07965_ (.A(_01666_),
    .B(_01771_),
    .Y(_01772_));
 sg13g2_nor2_1 _07966_ (.A(_05567_),
    .B(_01398_),
    .Y(_01773_));
 sg13g2_inv_1 _07967_ (.Y(_01774_),
    .A(_01773_));
 sg13g2_nand2_1 _07968_ (.Y(_01775_),
    .A(_01774_),
    .B(_01665_));
 sg13g2_nand2b_1 _07969_ (.Y(_01776_),
    .B(_01775_),
    .A_N(_01772_));
 sg13g2_xnor2_1 _07970_ (.Y(_01777_),
    .A(_01769_),
    .B(_01776_));
 sg13g2_nand2_1 _07971_ (.Y(_01778_),
    .A(_01768_),
    .B(_01777_));
 sg13g2_inv_1 _07972_ (.Y(_01779_),
    .A(_01777_));
 sg13g2_nand3_1 _07973_ (.B(_01767_),
    .C(_01779_),
    .A(_01766_),
    .Y(_01780_));
 sg13g2_nand2_1 _07974_ (.Y(_01781_),
    .A(_01778_),
    .B(_01780_));
 sg13g2_nand2b_1 _07975_ (.Y(_01782_),
    .B(_01781_),
    .A_N(_01732_));
 sg13g2_nand3_1 _07976_ (.B(_01778_),
    .C(_01780_),
    .A(_01732_),
    .Y(_01783_));
 sg13g2_nand2_1 _07977_ (.Y(_01784_),
    .A(_01782_),
    .B(_01783_));
 sg13g2_nor2_1 _07978_ (.A(_00649_),
    .B(_01099_),
    .Y(_01785_));
 sg13g2_xnor2_1 _07979_ (.Y(_01786_),
    .A(_01606_),
    .B(_01785_));
 sg13g2_a22oi_1 _07980_ (.Y(_01787_),
    .B1(_01663_),
    .B2(_01667_),
    .A2(_01572_),
    .A1(_01664_));
 sg13g2_xnor2_1 _07981_ (.Y(_01788_),
    .A(_01786_),
    .B(_01787_));
 sg13g2_xor2_1 _07982_ (.B(_01788_),
    .A(_01607_),
    .X(_01789_));
 sg13g2_nand2_1 _07983_ (.Y(_01790_),
    .A(_01784_),
    .B(_01789_));
 sg13g2_inv_1 _07984_ (.Y(_01791_),
    .A(_01789_));
 sg13g2_nand3_1 _07985_ (.B(_01783_),
    .C(_01791_),
    .A(_01782_),
    .Y(_01792_));
 sg13g2_nand2_1 _07986_ (.Y(_01793_),
    .A(_01790_),
    .B(_01792_));
 sg13g2_nand2b_1 _07987_ (.Y(_01794_),
    .B(_01793_),
    .A_N(_01729_));
 sg13g2_nand3_1 _07988_ (.B(_01790_),
    .C(_01792_),
    .A(_01729_),
    .Y(_01795_));
 sg13g2_nand2_1 _07989_ (.Y(_01796_),
    .A(_01794_),
    .B(_01795_));
 sg13g2_nor2b_1 _07990_ (.A(_01611_),
    .B_N(_01610_),
    .Y(_01797_));
 sg13g2_a21oi_1 _07991_ (.A1(_01612_),
    .A2(_01605_),
    .Y(_01798_),
    .B1(_01797_));
 sg13g2_inv_1 _07992_ (.Y(_01799_),
    .A(_01798_));
 sg13g2_nand2_1 _07993_ (.Y(_01800_),
    .A(_01796_),
    .B(_01799_));
 sg13g2_nand3_1 _07994_ (.B(_01795_),
    .C(_01798_),
    .A(_01794_),
    .Y(_01801_));
 sg13g2_nand2_1 _07995_ (.Y(_01802_),
    .A(_01800_),
    .B(_01801_));
 sg13g2_xor2_1 _07996_ (.B(_01802_),
    .A(_01726_),
    .X(_01803_));
 sg13g2_buf_2 _07997_ (.A(_01803_),
    .X(_01804_));
 sg13g2_nand2_1 _07998_ (.Y(_01805_),
    .A(_01723_),
    .B(_01804_));
 sg13g2_inv_1 _07999_ (.Y(_01806_),
    .A(_01804_));
 sg13g2_nand3_1 _08000_ (.B(_01722_),
    .C(_01806_),
    .A(_01706_),
    .Y(_01807_));
 sg13g2_nand3_1 _08001_ (.B(_01807_),
    .C(net56),
    .A(_01805_),
    .Y(_01808_));
 sg13g2_nor2_1 _08002_ (.A(_01456_),
    .B(_01710_),
    .Y(_01809_));
 sg13g2_nand3_1 _08003_ (.B(_01809_),
    .C(_01349_),
    .A(_01155_),
    .Y(_01810_));
 sg13g2_inv_1 _08004_ (.Y(_01811_),
    .A(_01355_));
 sg13g2_inv_1 _08005_ (.Y(_01812_),
    .A(_01707_));
 sg13g2_a21oi_1 _08006_ (.A1(_01709_),
    .A2(_01715_),
    .Y(_01813_),
    .B1(_01812_));
 sg13g2_a21oi_1 _08007_ (.A1(_01809_),
    .A2(_01811_),
    .Y(_01814_),
    .B1(_01813_));
 sg13g2_nand2_1 _08008_ (.Y(_01815_),
    .A(_01810_),
    .B(_01814_));
 sg13g2_xnor2_1 _08009_ (.Y(_01816_),
    .A(_01713_),
    .B(_01815_));
 sg13g2_buf_8 _08010_ (.A(net70),
    .X(_01817_));
 sg13g2_nand2_1 _08011_ (.Y(_01818_),
    .A(_01816_),
    .B(net61));
 sg13g2_nand2_1 _08012_ (.Y(_01819_),
    .A(_01808_),
    .B(_01818_));
 sg13g2_a21oi_1 _08013_ (.A1(_01819_),
    .A2(_03640_),
    .Y(_01820_),
    .B1(_01501_));
 sg13g2_nand2_1 _08014_ (.Y(_01821_),
    .A(_01804_),
    .B(_01692_));
 sg13g2_nor2b_1 _08015_ (.A(_01821_),
    .B_N(_01809_),
    .Y(_01822_));
 sg13g2_nand2_1 _08016_ (.Y(_01823_),
    .A(_01356_),
    .B(_01822_));
 sg13g2_nor2_1 _08017_ (.A(_01726_),
    .B(_01802_),
    .Y(_01824_));
 sg13g2_nand2_1 _08018_ (.Y(_01825_),
    .A(_01804_),
    .B(_01689_));
 sg13g2_nand2b_1 _08019_ (.Y(_01826_),
    .B(_01825_),
    .A_N(_01824_));
 sg13g2_nor2b_1 _08020_ (.A(_01821_),
    .B_N(_01813_),
    .Y(_01827_));
 sg13g2_nor2_1 _08021_ (.A(_01826_),
    .B(_01827_),
    .Y(_01828_));
 sg13g2_nand2_1 _08022_ (.Y(_01829_),
    .A(_01823_),
    .B(_01828_));
 sg13g2_nand2_1 _08023_ (.Y(_01830_),
    .A(_01793_),
    .B(_01729_));
 sg13g2_nor2_1 _08024_ (.A(_01729_),
    .B(_01793_),
    .Y(_01831_));
 sg13g2_a21oi_1 _08025_ (.A1(_01830_),
    .A2(_01799_),
    .Y(_01832_),
    .B1(_01831_));
 sg13g2_nand2_1 _08026_ (.Y(_01833_),
    .A(_01781_),
    .B(_01732_));
 sg13g2_nor2_1 _08027_ (.A(_01732_),
    .B(_01781_),
    .Y(_01834_));
 sg13g2_a21oi_2 _08028_ (.B1(_01834_),
    .Y(_01835_),
    .A2(_01789_),
    .A1(_01833_));
 sg13g2_nor2_1 _08029_ (.A(_00555_),
    .B(_01649_),
    .Y(_01836_));
 sg13g2_nand2_1 _08030_ (.Y(_01837_),
    .A(_01758_),
    .B(net90));
 sg13g2_a21oi_2 _08031_ (.B1(_01757_),
    .Y(_01838_),
    .A2(_00551_),
    .A1(_00412_));
 sg13g2_nand2_1 _08032_ (.Y(_01839_),
    .A(_01837_),
    .B(_01838_));
 sg13g2_xnor2_1 _08033_ (.Y(_01840_),
    .A(_01836_),
    .B(_01839_));
 sg13g2_a22oi_1 _08034_ (.Y(_01841_),
    .B1(_01737_),
    .B2(_01761_),
    .A2(_01758_),
    .A1(_01650_));
 sg13g2_buf_1 _08035_ (.A(_01841_),
    .X(_01842_));
 sg13g2_nand2_1 _08036_ (.Y(_01843_),
    .A(_01840_),
    .B(_01842_));
 sg13g2_inv_1 _08037_ (.Y(_01844_),
    .A(_01836_));
 sg13g2_xnor2_1 _08038_ (.Y(_01845_),
    .A(_01844_),
    .B(_01839_));
 sg13g2_inv_1 _08039_ (.Y(_01846_),
    .A(_01842_));
 sg13g2_nand2_1 _08040_ (.Y(_01847_),
    .A(_01845_),
    .B(_01846_));
 sg13g2_nand2_1 _08041_ (.Y(_01848_),
    .A(_01843_),
    .B(_01847_));
 sg13g2_nor2_1 _08042_ (.A(net44),
    .B(_01299_),
    .Y(_01849_));
 sg13g2_nand2_1 _08043_ (.Y(_01850_),
    .A(_01549_),
    .B(net71));
 sg13g2_xor2_1 _08044_ (.B(_01850_),
    .A(_01771_),
    .X(_01851_));
 sg13g2_xnor2_1 _08045_ (.Y(_01852_),
    .A(_01849_),
    .B(_01851_));
 sg13g2_inv_2 _08046_ (.Y(_01853_),
    .A(_01852_));
 sg13g2_nand2_1 _08047_ (.Y(_01854_),
    .A(_01848_),
    .B(_01853_));
 sg13g2_nand3_1 _08048_ (.B(_01847_),
    .C(_01852_),
    .A(_01843_),
    .Y(_01855_));
 sg13g2_nand2_1 _08049_ (.Y(_01856_),
    .A(_01854_),
    .B(_01855_));
 sg13g2_nand2_1 _08050_ (.Y(_01857_),
    .A(_01765_),
    .B(_01736_));
 sg13g2_nor2_1 _08051_ (.A(_01736_),
    .B(_01765_),
    .Y(_01858_));
 sg13g2_a21oi_2 _08052_ (.B1(_01858_),
    .Y(_01859_),
    .A2(_01777_),
    .A1(_01857_));
 sg13g2_inv_1 _08053_ (.Y(_01860_),
    .A(_01859_));
 sg13g2_nand2_1 _08054_ (.Y(_01861_),
    .A(_01856_),
    .B(_01860_));
 sg13g2_nand3_1 _08055_ (.B(_01859_),
    .C(_01855_),
    .A(_01854_),
    .Y(_01862_));
 sg13g2_nand2_1 _08056_ (.Y(_01863_),
    .A(_01861_),
    .B(_01862_));
 sg13g2_nor2_1 _08057_ (.A(_00232_),
    .B(_01099_),
    .Y(_01864_));
 sg13g2_nand2_1 _08058_ (.Y(_01865_),
    .A(_01864_),
    .B(_01608_));
 sg13g2_a21oi_1 _08059_ (.A1(_01569_),
    .A2(_00223_),
    .Y(_01866_),
    .B1(_01864_));
 sg13g2_nor2_1 _08060_ (.A(_00232_),
    .B(_01204_),
    .Y(_01867_));
 sg13g2_inv_1 _08061_ (.Y(_01868_),
    .A(_01867_));
 sg13g2_nor2b_1 _08062_ (.A(_01868_),
    .B_N(_01785_),
    .Y(_01869_));
 sg13g2_nor2_1 _08063_ (.A(_01866_),
    .B(_01869_),
    .Y(_01870_));
 sg13g2_a21oi_1 _08064_ (.A1(_01775_),
    .A2(_01769_),
    .Y(_01871_),
    .B1(_01772_));
 sg13g2_xnor2_1 _08065_ (.Y(_01872_),
    .A(_01870_),
    .B(_01871_));
 sg13g2_xnor2_1 _08066_ (.Y(_01873_),
    .A(_01865_),
    .B(_01872_));
 sg13g2_nand2_1 _08067_ (.Y(_01874_),
    .A(_01863_),
    .B(_01873_));
 sg13g2_inv_1 _08068_ (.Y(_01875_),
    .A(_01873_));
 sg13g2_nand3_1 _08069_ (.B(_01862_),
    .C(_01875_),
    .A(_01861_),
    .Y(_01876_));
 sg13g2_nand3_1 _08070_ (.B(_01874_),
    .C(_01876_),
    .A(_01835_),
    .Y(_01877_));
 sg13g2_nand2_1 _08071_ (.Y(_01878_),
    .A(_01874_),
    .B(_01876_));
 sg13g2_inv_1 _08072_ (.Y(_01879_),
    .A(_01835_));
 sg13g2_nand2_1 _08073_ (.Y(_01880_),
    .A(_01878_),
    .B(_01879_));
 sg13g2_nand2_1 _08074_ (.Y(_01881_),
    .A(_01877_),
    .B(_01880_));
 sg13g2_nor2b_1 _08075_ (.A(_01787_),
    .B_N(_01786_),
    .Y(_01882_));
 sg13g2_a21oi_1 _08076_ (.A1(_01788_),
    .A2(_01607_),
    .Y(_01883_),
    .B1(_01882_));
 sg13g2_inv_1 _08077_ (.Y(_01884_),
    .A(_01883_));
 sg13g2_nand2_1 _08078_ (.Y(_01885_),
    .A(_01881_),
    .B(_01884_));
 sg13g2_nand3_1 _08079_ (.B(_01880_),
    .C(_01883_),
    .A(_01877_),
    .Y(_01886_));
 sg13g2_nand2_1 _08080_ (.Y(_01887_),
    .A(_01885_),
    .B(_01886_));
 sg13g2_nor2_1 _08081_ (.A(_01832_),
    .B(_01887_),
    .Y(_01888_));
 sg13g2_nand2_1 _08082_ (.Y(_01889_),
    .A(_01887_),
    .B(_01832_));
 sg13g2_inv_4 _08083_ (.A(_01889_),
    .Y(_01890_));
 sg13g2_nor2_2 _08084_ (.A(_01888_),
    .B(_01890_),
    .Y(_01891_));
 sg13g2_inv_2 _08085_ (.Y(_01892_),
    .A(_01891_));
 sg13g2_nand2_1 _08086_ (.Y(_01893_),
    .A(_01829_),
    .B(_01892_));
 sg13g2_nand3_1 _08087_ (.B(_01891_),
    .C(_01828_),
    .A(_01823_),
    .Y(_01894_));
 sg13g2_nand3_1 _08088_ (.B(_01894_),
    .C(net61),
    .A(_01893_),
    .Y(_01895_));
 sg13g2_nor2_1 _08089_ (.A(_01481_),
    .B(_01511_),
    .Y(_01896_));
 sg13g2_nor2_1 _08090_ (.A(_01718_),
    .B(_01896_),
    .Y(_01897_));
 sg13g2_nor2_1 _08091_ (.A(_01477_),
    .B(_01511_),
    .Y(_01898_));
 sg13g2_nand2_1 _08092_ (.Y(_01899_),
    .A(_01898_),
    .B(_01475_));
 sg13g2_nand2_1 _08093_ (.Y(_01900_),
    .A(_01897_),
    .B(_01899_));
 sg13g2_nand2_1 _08094_ (.Y(_01901_),
    .A(_01891_),
    .B(_01804_));
 sg13g2_nor2_1 _08095_ (.A(_01704_),
    .B(_01901_),
    .Y(_01902_));
 sg13g2_nand2_1 _08096_ (.Y(_01903_),
    .A(_01900_),
    .B(_01902_));
 sg13g2_nor2_1 _08097_ (.A(_01888_),
    .B(_01824_),
    .Y(_01904_));
 sg13g2_nor2_1 _08098_ (.A(_01890_),
    .B(_01904_),
    .Y(_01905_));
 sg13g2_nor2_1 _08099_ (.A(_01720_),
    .B(_01901_),
    .Y(_01906_));
 sg13g2_nor2_1 _08100_ (.A(_01905_),
    .B(_01906_),
    .Y(_01907_));
 sg13g2_nand2_1 _08101_ (.Y(_01908_),
    .A(_01903_),
    .B(_01907_));
 sg13g2_nand2_1 _08102_ (.Y(_01909_),
    .A(_01878_),
    .B(_01835_));
 sg13g2_nor2_1 _08103_ (.A(_01835_),
    .B(_01878_),
    .Y(_01910_));
 sg13g2_a21oi_1 _08104_ (.A1(_01909_),
    .A2(_01884_),
    .Y(_01911_),
    .B1(_01910_));
 sg13g2_inv_1 _08105_ (.Y(_01912_),
    .A(_01865_));
 sg13g2_nor2b_1 _08106_ (.A(_01871_),
    .B_N(_01870_),
    .Y(_01913_));
 sg13g2_a21oi_1 _08107_ (.A1(_01872_),
    .A2(_01912_),
    .Y(_01914_),
    .B1(_01913_));
 sg13g2_nand2_1 _08108_ (.Y(_01915_),
    .A(_01856_),
    .B(_01859_));
 sg13g2_nor2_1 _08109_ (.A(_01859_),
    .B(_01856_),
    .Y(_01916_));
 sg13g2_a21oi_1 _08110_ (.A1(_01915_),
    .A2(_01873_),
    .Y(_01917_),
    .B1(_01916_));
 sg13g2_inv_1 _08111_ (.Y(_01918_),
    .A(_01917_));
 sg13g2_nand2_1 _08112_ (.Y(_01919_),
    .A(_01845_),
    .B(_01842_));
 sg13g2_nor2_1 _08113_ (.A(_01842_),
    .B(_01845_),
    .Y(_01920_));
 sg13g2_a21oi_1 _08114_ (.A1(_01853_),
    .A2(_01919_),
    .Y(_01921_),
    .B1(_01920_));
 sg13g2_nor2_1 _08115_ (.A(net44),
    .B(_01398_),
    .Y(_01922_));
 sg13g2_nor2_2 _08116_ (.A(_05567_),
    .B(_01649_),
    .Y(_01923_));
 sg13g2_nand2_1 _08117_ (.Y(_01924_),
    .A(_01549_),
    .B(_00193_));
 sg13g2_xnor2_1 _08118_ (.Y(_01925_),
    .A(_01923_),
    .B(_01924_));
 sg13g2_xor2_1 _08119_ (.B(_01925_),
    .A(_01922_),
    .X(_01926_));
 sg13g2_xnor2_1 _08120_ (.Y(_01927_),
    .A(_01755_),
    .B(_01746_));
 sg13g2_nand2_1 _08121_ (.Y(_01928_),
    .A(_01927_),
    .B(_00332_));
 sg13g2_inv_1 _08122_ (.Y(_01929_),
    .A(_01928_));
 sg13g2_nand2_1 _08123_ (.Y(_01930_),
    .A(_01839_),
    .B(_01929_));
 sg13g2_nand3_1 _08124_ (.B(_01838_),
    .C(_01928_),
    .A(_01837_),
    .Y(_01931_));
 sg13g2_nor2_1 _08125_ (.A(_00551_),
    .B(_01760_),
    .Y(_01932_));
 sg13g2_a21oi_1 _08126_ (.A1(_01838_),
    .A2(_01836_),
    .Y(_01933_),
    .B1(_01932_));
 sg13g2_nand3_1 _08127_ (.B(_01931_),
    .C(_01933_),
    .A(_01930_),
    .Y(_01934_));
 sg13g2_nor2_1 _08128_ (.A(_03267_),
    .B(_01837_),
    .Y(_01935_));
 sg13g2_inv_2 _08129_ (.Y(_01936_),
    .A(_01935_));
 sg13g2_nand2_1 _08130_ (.Y(_01937_),
    .A(_01934_),
    .B(_01936_));
 sg13g2_xor2_1 _08131_ (.B(_01937_),
    .A(_01926_),
    .X(_01938_));
 sg13g2_nand2b_1 _08132_ (.Y(_01939_),
    .B(_01938_),
    .A_N(_01921_));
 sg13g2_xnor2_1 _08133_ (.Y(_01940_),
    .A(_01926_),
    .B(_01937_));
 sg13g2_nand2_1 _08134_ (.Y(_01941_),
    .A(_01940_),
    .B(_01921_));
 sg13g2_nand2_1 _08135_ (.Y(_01942_),
    .A(_01939_),
    .B(_01941_));
 sg13g2_nand2_1 _08136_ (.Y(_01943_),
    .A(_01400_),
    .B(_00223_));
 sg13g2_xnor2_1 _08137_ (.Y(_01944_),
    .A(_01867_),
    .B(_01943_));
 sg13g2_nand2_1 _08138_ (.Y(_01945_),
    .A(_01850_),
    .B(_01771_));
 sg13g2_nor2_1 _08139_ (.A(_01774_),
    .B(_01924_),
    .Y(_01946_));
 sg13g2_a21oi_1 _08140_ (.A1(_01945_),
    .A2(_01849_),
    .Y(_01947_),
    .B1(_01946_));
 sg13g2_xnor2_1 _08141_ (.Y(_01948_),
    .A(_01944_),
    .B(_01947_));
 sg13g2_xor2_1 _08142_ (.B(_01948_),
    .A(_01869_),
    .X(_01949_));
 sg13g2_nand2_1 _08143_ (.Y(_01950_),
    .A(_01942_),
    .B(_01949_));
 sg13g2_inv_1 _08144_ (.Y(_01951_),
    .A(_01949_));
 sg13g2_nand3_1 _08145_ (.B(_01941_),
    .C(_01951_),
    .A(_01939_),
    .Y(_01952_));
 sg13g2_nand2_1 _08146_ (.Y(_01953_),
    .A(_01950_),
    .B(_01952_));
 sg13g2_xnor2_1 _08147_ (.Y(_01954_),
    .A(_01918_),
    .B(_01953_));
 sg13g2_xnor2_1 _08148_ (.Y(_01955_),
    .A(_01914_),
    .B(_01954_));
 sg13g2_nand2b_1 _08149_ (.Y(_01956_),
    .B(_01955_),
    .A_N(_01911_));
 sg13g2_inv_1 _08150_ (.Y(_01957_),
    .A(_01914_));
 sg13g2_xnor2_1 _08151_ (.Y(_01958_),
    .A(_01957_),
    .B(_01954_));
 sg13g2_nand2_1 _08152_ (.Y(_01959_),
    .A(_01958_),
    .B(_01911_));
 sg13g2_nand2_2 _08153_ (.Y(_01960_),
    .A(_01956_),
    .B(_01959_));
 sg13g2_nand2_1 _08154_ (.Y(_01961_),
    .A(_01908_),
    .B(_01960_));
 sg13g2_inv_1 _08155_ (.Y(_01962_),
    .A(_01960_));
 sg13g2_nand3_1 _08156_ (.B(_01907_),
    .C(_01962_),
    .A(_01903_),
    .Y(_01963_));
 sg13g2_nand3_1 _08157_ (.B(_01963_),
    .C(net56),
    .A(_01961_),
    .Y(_01964_));
 sg13g2_nand3_1 _08158_ (.B(_01964_),
    .C(net67),
    .A(_01895_),
    .Y(_01965_));
 sg13g2_xnor2_1 _08159_ (.Y(_01966_),
    .A(_01710_),
    .B(_01900_));
 sg13g2_nand2_1 _08160_ (.Y(_01967_),
    .A(_01966_),
    .B(net64));
 sg13g2_nand3_1 _08161_ (.B(_01457_),
    .C(net70),
    .A(_01455_),
    .Y(_01968_));
 sg13g2_nand3_1 _08162_ (.B(_01968_),
    .C(_01486_),
    .A(_01967_),
    .Y(_01969_));
 sg13g2_xnor2_1 _08163_ (.Y(_01970_),
    .A(_01348_),
    .B(_01482_));
 sg13g2_nand2_1 _08164_ (.Y(_01971_),
    .A(_01970_),
    .B(net64));
 sg13g2_nand2_1 _08165_ (.Y(_01972_),
    .A(_01489_),
    .B(net70));
 sg13g2_nand3_1 _08166_ (.B(net78),
    .C(_01972_),
    .A(_01971_),
    .Y(_01973_));
 sg13g2_a21oi_1 _08167_ (.A1(_01969_),
    .A2(_01973_),
    .Y(_01974_),
    .B1(net72));
 sg13g2_a21oi_1 _08168_ (.A1(_01820_),
    .A2(_01965_),
    .Y(_01975_),
    .B1(_01974_));
 sg13g2_buf_8 _08169_ (.A(_01975_),
    .X(_01976_));
 sg13g2_inv_4 _08170_ (.A(net20),
    .Y(_01977_));
 sg13g2_nor2_1 _08171_ (.A(_01510_),
    .B(_01977_),
    .Y(_01978_));
 sg13g2_nand2_1 _08172_ (.Y(_01979_),
    .A(_01816_),
    .B(_00202_));
 sg13g2_nand2_1 _08173_ (.Y(_01980_),
    .A(_01966_),
    .B(net70));
 sg13g2_nand2_1 _08174_ (.Y(_01981_),
    .A(_01979_),
    .B(_01980_));
 sg13g2_a21oi_1 _08175_ (.A1(_01981_),
    .A2(net78),
    .Y(_01982_),
    .B1(_01501_));
 sg13g2_nand3_1 _08176_ (.B(_01894_),
    .C(net56),
    .A(_01893_),
    .Y(_01983_));
 sg13g2_nand2_1 _08177_ (.Y(_01984_),
    .A(_01805_),
    .B(_01807_));
 sg13g2_nand2_1 _08178_ (.Y(_01985_),
    .A(_01984_),
    .B(net61));
 sg13g2_nand3_1 _08179_ (.B(_01487_),
    .C(_01985_),
    .A(_01983_),
    .Y(_01986_));
 sg13g2_nand2_1 _08180_ (.Y(_01987_),
    .A(_01982_),
    .B(_01986_));
 sg13g2_a21o_1 _08181_ (.A2(_01494_),
    .A1(_01488_),
    .B1(net72),
    .X(_01988_));
 sg13g2_nand3_1 _08182_ (.B(_03965_),
    .C(_01973_),
    .A(_01969_),
    .Y(_01989_));
 sg13g2_nor2_1 _08183_ (.A(_00201_),
    .B(_01491_),
    .Y(_01990_));
 sg13g2_a21oi_1 _08184_ (.A1(_00201_),
    .A2(_01496_),
    .Y(_01991_),
    .B1(_01990_));
 sg13g2_nand2_1 _08185_ (.Y(_01992_),
    .A(_01991_),
    .B(net67));
 sg13g2_nand2_1 _08186_ (.Y(_01993_),
    .A(_01497_),
    .B(net56));
 sg13g2_a21oi_1 _08187_ (.A1(_01504_),
    .A2(net61),
    .Y(_01994_),
    .B1(_01486_));
 sg13g2_nand2_1 _08188_ (.Y(_01995_),
    .A(_01993_),
    .B(_01994_));
 sg13g2_nand3_1 _08189_ (.B(_01501_),
    .C(_01995_),
    .A(_01992_),
    .Y(_01996_));
 sg13g2_nand2_1 _08190_ (.Y(_01997_),
    .A(_01989_),
    .B(_01996_));
 sg13g2_buf_8 _08191_ (.A(_01997_),
    .X(_01998_));
 sg13g2_nand3_1 _08192_ (.B(_01988_),
    .C(_01998_),
    .A(_01987_),
    .Y(_01999_));
 sg13g2_nand2_1 _08193_ (.Y(_02000_),
    .A(_01819_),
    .B(net67));
 sg13g2_a21o_1 _08194_ (.A2(_01968_),
    .A1(_01967_),
    .B1(net67),
    .X(_02001_));
 sg13g2_nand2_1 _08195_ (.Y(_02002_),
    .A(_02000_),
    .B(_02001_));
 sg13g2_nand2_1 _08196_ (.Y(_02003_),
    .A(_02002_),
    .B(net72));
 sg13g2_a21oi_1 _08197_ (.A1(_01991_),
    .A2(net78),
    .Y(_02004_),
    .B1(net72));
 sg13g2_nand3_1 _08198_ (.B(net67),
    .C(_01972_),
    .A(_01971_),
    .Y(_02005_));
 sg13g2_nand2_1 _08199_ (.Y(_02006_),
    .A(_02004_),
    .B(_02005_));
 sg13g2_nand2_1 _08200_ (.Y(_02007_),
    .A(_02003_),
    .B(_02006_));
 sg13g2_buf_8 _08201_ (.A(_02007_),
    .X(_02008_));
 sg13g2_nand2_1 _08202_ (.Y(_02009_),
    .A(_01981_),
    .B(net67));
 sg13g2_inv_1 _08203_ (.Y(_02010_),
    .A(_01485_));
 sg13g2_nand2_1 _08204_ (.Y(_02011_),
    .A(_02010_),
    .B(net78));
 sg13g2_nand2_1 _08205_ (.Y(_02012_),
    .A(_02009_),
    .B(_02011_));
 sg13g2_nand2_1 _08206_ (.Y(_02013_),
    .A(_02012_),
    .B(_03976_));
 sg13g2_inv_1 _08207_ (.Y(_02014_),
    .A(_01493_));
 sg13g2_a21oi_1 _08208_ (.A1(_01499_),
    .A2(net78),
    .Y(_02015_),
    .B1(_03965_));
 sg13g2_o21ai_1 _08209_ (.B1(_02015_),
    .Y(_02016_),
    .A1(net78),
    .A2(_02014_));
 sg13g2_nand2_1 _08210_ (.Y(_02017_),
    .A(_02013_),
    .B(_02016_));
 sg13g2_buf_8 _08211_ (.A(_02017_),
    .X(_02018_));
 sg13g2_nand2_2 _08212_ (.Y(_02019_),
    .A(_02008_),
    .B(net19));
 sg13g2_nor2_1 _08213_ (.A(_01999_),
    .B(_02019_),
    .Y(_02020_));
 sg13g2_inv_1 _08214_ (.Y(_02021_),
    .A(_02020_));
 sg13g2_nand2_1 _08215_ (.Y(_02022_),
    .A(_02019_),
    .B(_01999_));
 sg13g2_nand2_1 _08216_ (.Y(_02023_),
    .A(_02021_),
    .B(_02022_));
 sg13g2_xnor2_1 _08217_ (.Y(_02024_),
    .A(_01978_),
    .B(_02023_));
 sg13g2_inv_1 _08218_ (.Y(_02025_),
    .A(_02024_));
 sg13g2_nand2_1 _08219_ (.Y(_02026_),
    .A(net20),
    .B(_01998_));
 sg13g2_inv_1 _08220_ (.Y(_02027_),
    .A(_02026_));
 sg13g2_nand2_2 _08221_ (.Y(_02028_),
    .A(_01987_),
    .B(_01988_));
 sg13g2_nor2_1 _08222_ (.A(_02028_),
    .B(_02019_),
    .Y(_02029_));
 sg13g2_inv_8 _08223_ (.Y(_02030_),
    .A(_02028_));
 sg13g2_nand2_1 _08224_ (.Y(_02031_),
    .A(_02030_),
    .B(net19));
 sg13g2_inv_4 _08225_ (.A(_02008_),
    .Y(_02032_));
 sg13g2_nand2_1 _08226_ (.Y(_02033_),
    .A(_02031_),
    .B(_02032_));
 sg13g2_nand2b_1 _08227_ (.Y(_02034_),
    .B(_02033_),
    .A_N(_02029_));
 sg13g2_xnor2_1 _08228_ (.Y(_02035_),
    .A(_02027_),
    .B(_02034_));
 sg13g2_a21oi_2 _08229_ (.B1(_02020_),
    .Y(_02036_),
    .A2(_01978_),
    .A1(_02022_));
 sg13g2_inv_2 _08230_ (.Y(_02037_),
    .A(_02036_));
 sg13g2_nand2_1 _08231_ (.Y(_02038_),
    .A(_01908_),
    .B(_01962_));
 sg13g2_nand3_1 _08232_ (.B(_01907_),
    .C(_01960_),
    .A(_01903_),
    .Y(_02039_));
 sg13g2_nand2_1 _08233_ (.Y(_02040_),
    .A(_02038_),
    .B(_02039_));
 sg13g2_a21oi_1 _08234_ (.A1(_02040_),
    .A2(_01817_),
    .Y(_02041_),
    .B1(_03684_));
 sg13g2_nor3_1 _08235_ (.A(_01892_),
    .B(_01960_),
    .C(_01821_),
    .Y(_02042_));
 sg13g2_nand2_1 _08236_ (.Y(_02043_),
    .A(_01815_),
    .B(_02042_));
 sg13g2_nor2_1 _08237_ (.A(_01960_),
    .B(_01892_),
    .Y(_02044_));
 sg13g2_inv_1 _08238_ (.Y(_02045_),
    .A(_01956_));
 sg13g2_a21o_1 _08239_ (.A2(_01959_),
    .A1(_01888_),
    .B1(_02045_),
    .X(_02046_));
 sg13g2_a21oi_1 _08240_ (.A1(_01826_),
    .A2(_02044_),
    .Y(_02047_),
    .B1(_02046_));
 sg13g2_nand2_1 _08241_ (.Y(_02048_),
    .A(_02043_),
    .B(_02047_));
 sg13g2_nand2_1 _08242_ (.Y(_02049_),
    .A(_01953_),
    .B(_01917_));
 sg13g2_nor2_1 _08243_ (.A(_01917_),
    .B(_01953_),
    .Y(_02050_));
 sg13g2_a21oi_1 _08244_ (.A1(_02049_),
    .A2(_01957_),
    .Y(_02051_),
    .B1(_02050_));
 sg13g2_nor2_1 _08245_ (.A(_01943_),
    .B(_01868_),
    .Y(_02052_));
 sg13g2_nand2_1 _08246_ (.Y(_02053_),
    .A(_01400_),
    .B(net50));
 sg13g2_nor2_1 _08247_ (.A(_00649_),
    .B(_01398_),
    .Y(_02054_));
 sg13g2_xnor2_1 _08248_ (.Y(_02055_),
    .A(_02053_),
    .B(_02054_));
 sg13g2_inv_1 _08249_ (.Y(_02056_),
    .A(_01923_));
 sg13g2_nor2_1 _08250_ (.A(_01924_),
    .B(_02056_),
    .Y(_02057_));
 sg13g2_a21oi_1 _08251_ (.A1(_01925_),
    .A2(_01922_),
    .Y(_02058_),
    .B1(_02057_));
 sg13g2_xnor2_1 _08252_ (.Y(_02059_),
    .A(_02055_),
    .B(_02058_));
 sg13g2_xor2_1 _08253_ (.B(_02059_),
    .A(_02052_),
    .X(_02060_));
 sg13g2_o21ai_1 _08254_ (.B1(_01936_),
    .Y(_02061_),
    .A1(_01838_),
    .A2(_01929_));
 sg13g2_buf_8 _08255_ (.A(_02061_),
    .X(_02062_));
 sg13g2_nor2_1 _08256_ (.A(_01112_),
    .B(_01652_),
    .Y(_02063_));
 sg13g2_nand2_1 _08257_ (.Y(_02064_),
    .A(_01927_),
    .B(net71));
 sg13g2_o21ai_1 _08258_ (.B1(_02064_),
    .Y(_02065_),
    .A1(_01649_),
    .A2(net63));
 sg13g2_nor2_1 _08259_ (.A(_00325_),
    .B(_01757_),
    .Y(_02066_));
 sg13g2_nand2_1 _08260_ (.Y(_02067_),
    .A(_01923_),
    .B(_02066_));
 sg13g2_nand2_1 _08261_ (.Y(_02068_),
    .A(_02065_),
    .B(_02067_));
 sg13g2_xor2_1 _08262_ (.B(_02068_),
    .A(_02063_),
    .X(_02069_));
 sg13g2_xor2_1 _08263_ (.B(_02069_),
    .A(_02062_),
    .X(_02070_));
 sg13g2_a21oi_1 _08264_ (.A1(_01926_),
    .A2(_01934_),
    .Y(_02071_),
    .B1(_01935_));
 sg13g2_inv_1 _08265_ (.Y(_02072_),
    .A(_02071_));
 sg13g2_nand2_1 _08266_ (.Y(_02073_),
    .A(_02070_),
    .B(_02072_));
 sg13g2_xnor2_1 _08267_ (.Y(_02074_),
    .A(_02062_),
    .B(_02069_));
 sg13g2_nand2_1 _08268_ (.Y(_02075_),
    .A(_02074_),
    .B(_02071_));
 sg13g2_nand2_1 _08269_ (.Y(_02076_),
    .A(_02073_),
    .B(_02075_));
 sg13g2_xnor2_1 _08270_ (.Y(_02077_),
    .A(_02060_),
    .B(_02076_));
 sg13g2_inv_1 _08271_ (.Y(_02078_),
    .A(_02077_));
 sg13g2_nand2_1 _08272_ (.Y(_02079_),
    .A(_01938_),
    .B(_01921_));
 sg13g2_nor2_1 _08273_ (.A(_01921_),
    .B(_01938_),
    .Y(_02080_));
 sg13g2_a21oi_1 _08274_ (.A1(_02079_),
    .A2(_01949_),
    .Y(_02081_),
    .B1(_02080_));
 sg13g2_nand2_1 _08275_ (.Y(_02082_),
    .A(_02078_),
    .B(_02081_));
 sg13g2_nand2b_1 _08276_ (.Y(_02083_),
    .B(_02077_),
    .A_N(_02081_));
 sg13g2_nand2_1 _08277_ (.Y(_02084_),
    .A(_02082_),
    .B(_02083_));
 sg13g2_nor2b_1 _08278_ (.A(_01947_),
    .B_N(_01944_),
    .Y(_02085_));
 sg13g2_a21oi_1 _08279_ (.A1(_01948_),
    .A2(_01869_),
    .Y(_02086_),
    .B1(_02085_));
 sg13g2_nand2_1 _08280_ (.Y(_02087_),
    .A(_02084_),
    .B(_02086_));
 sg13g2_inv_1 _08281_ (.Y(_02088_),
    .A(_02086_));
 sg13g2_nand3_1 _08282_ (.B(_02083_),
    .C(_02088_),
    .A(_02082_),
    .Y(_02089_));
 sg13g2_nand2_1 _08283_ (.Y(_02090_),
    .A(_02087_),
    .B(_02089_));
 sg13g2_xnor2_1 _08284_ (.Y(_02091_),
    .A(_02051_),
    .B(_02090_));
 sg13g2_nand2_1 _08285_ (.Y(_02092_),
    .A(_02048_),
    .B(_02091_));
 sg13g2_inv_1 _08286_ (.Y(_02093_),
    .A(_02091_));
 sg13g2_nand3_1 _08287_ (.B(_02093_),
    .C(_02047_),
    .A(_02043_),
    .Y(_02094_));
 sg13g2_nand3_1 _08288_ (.B(_02094_),
    .C(_01502_),
    .A(_02092_),
    .Y(_02095_));
 sg13g2_nand2_1 _08289_ (.Y(_02096_),
    .A(_02041_),
    .B(_02095_));
 sg13g2_nand3_1 _08290_ (.B(_03684_),
    .C(_01985_),
    .A(_01983_),
    .Y(_02097_));
 sg13g2_nand2_1 _08291_ (.Y(_02098_),
    .A(_02096_),
    .B(_02097_));
 sg13g2_nand2_1 _08292_ (.Y(_02099_),
    .A(_02098_),
    .B(net72));
 sg13g2_nand2_1 _08293_ (.Y(_02100_),
    .A(_02012_),
    .B(_01501_));
 sg13g2_nand2_1 _08294_ (.Y(_02101_),
    .A(_02099_),
    .B(_02100_));
 sg13g2_buf_8 _08295_ (.A(_02101_),
    .X(_02102_));
 sg13g2_inv_8 _08296_ (.Y(_02103_),
    .A(_01998_));
 sg13g2_nor2_1 _08297_ (.A(_02103_),
    .B(_01510_),
    .Y(_02104_));
 sg13g2_nand3_1 _08298_ (.B(_02104_),
    .C(net20),
    .A(net18),
    .Y(_02105_));
 sg13g2_nand3_1 _08299_ (.B(_02097_),
    .C(net72),
    .A(_02096_),
    .Y(_02106_));
 sg13g2_nand3_1 _08300_ (.B(_01501_),
    .C(_02011_),
    .A(_02009_),
    .Y(_02107_));
 sg13g2_nand3_1 _08301_ (.B(_02107_),
    .C(_01509_),
    .A(_02106_),
    .Y(_02108_));
 sg13g2_buf_1 _08302_ (.A(_02108_),
    .X(_02109_));
 sg13g2_nand2_1 _08303_ (.Y(_02110_),
    .A(_02109_),
    .B(_02026_));
 sg13g2_nand2_1 _08304_ (.Y(_02111_),
    .A(_02105_),
    .B(_02110_));
 sg13g2_nand2_1 _08305_ (.Y(_02112_),
    .A(_02111_),
    .B(_02031_));
 sg13g2_inv_1 _08306_ (.Y(_02113_),
    .A(_02031_));
 sg13g2_nand3_1 _08307_ (.B(_02110_),
    .C(_02113_),
    .A(_02105_),
    .Y(_02114_));
 sg13g2_nand3_1 _08308_ (.B(_02112_),
    .C(_02114_),
    .A(_02037_),
    .Y(_02115_));
 sg13g2_nand2_1 _08309_ (.Y(_02116_),
    .A(_02111_),
    .B(_02113_));
 sg13g2_nand3_1 _08310_ (.B(_02110_),
    .C(_02031_),
    .A(_02105_),
    .Y(_02117_));
 sg13g2_nand3_1 _08311_ (.B(_02117_),
    .C(_02036_),
    .A(_02116_),
    .Y(_02118_));
 sg13g2_buf_1 _08312_ (.A(_02118_),
    .X(_02119_));
 sg13g2_nand2_1 _08313_ (.Y(_02120_),
    .A(_02115_),
    .B(_02119_));
 sg13g2_nand2b_1 _08314_ (.Y(_02121_),
    .B(_02120_),
    .A_N(_02035_));
 sg13g2_nand3_1 _08315_ (.B(_02119_),
    .C(_02035_),
    .A(_02115_),
    .Y(_02122_));
 sg13g2_nand2_1 _08316_ (.Y(_02123_),
    .A(_02121_),
    .B(_02122_));
 sg13g2_nor2_1 _08317_ (.A(_02025_),
    .B(_02123_),
    .Y(_02124_));
 sg13g2_inv_1 _08318_ (.Y(_02125_),
    .A(_02124_));
 sg13g2_nand2_1 _08319_ (.Y(_02126_),
    .A(_02123_),
    .B(_02025_));
 sg13g2_nand2_1 _08320_ (.Y(_02127_),
    .A(_02125_),
    .B(_02126_));
 sg13g2_xor2_1 _08321_ (.B(_02036_),
    .A(_02109_),
    .X(_02128_));
 sg13g2_nand2_1 _08322_ (.Y(_02129_),
    .A(_02127_),
    .B(_02128_));
 sg13g2_inv_1 _08323_ (.Y(_02130_),
    .A(_02128_));
 sg13g2_nand3_1 _08324_ (.B(_02126_),
    .C(_02130_),
    .A(_02125_),
    .Y(_02131_));
 sg13g2_nand2_1 _08325_ (.Y(_02132_),
    .A(_02030_),
    .B(_01509_));
 sg13g2_nor4_1 _08326_ (.A(_02103_),
    .B(_02018_),
    .C(_02032_),
    .D(_02132_),
    .Y(_02133_));
 sg13g2_a221oi_1 _08327_ (.B2(_02032_),
    .C1(_02103_),
    .B1(_02132_),
    .A1(_02016_),
    .Y(_02134_),
    .A2(_02013_));
 sg13g2_nor2_1 _08328_ (.A(_02133_),
    .B(_02134_),
    .Y(_02135_));
 sg13g2_nand3_1 _08329_ (.B(_02131_),
    .C(_02135_),
    .A(_02129_),
    .Y(_02136_));
 sg13g2_nor2_1 _08330_ (.A(_01510_),
    .B(_02032_),
    .Y(_02137_));
 sg13g2_nand2_1 _08331_ (.Y(_02138_),
    .A(_02137_),
    .B(net19));
 sg13g2_nand2b_1 _08332_ (.Y(_02139_),
    .B(_02032_),
    .A_N(_02018_));
 sg13g2_nand3_1 _08333_ (.B(_01998_),
    .C(_02019_),
    .A(_02139_),
    .Y(_02140_));
 sg13g2_xnor2_1 _08334_ (.Y(_02141_),
    .A(_02132_),
    .B(_02140_));
 sg13g2_nor2_1 _08335_ (.A(_02138_),
    .B(_02141_),
    .Y(_02142_));
 sg13g2_xnor2_1 _08336_ (.Y(_02143_),
    .A(_02130_),
    .B(_02127_));
 sg13g2_nor2_1 _08337_ (.A(_02135_),
    .B(_02143_),
    .Y(_02144_));
 sg13g2_a21oi_2 _08338_ (.B1(_02144_),
    .Y(_02145_),
    .A2(_02142_),
    .A1(_02136_));
 sg13g2_nor2_1 _08339_ (.A(_02109_),
    .B(_02036_),
    .Y(_02146_));
 sg13g2_a21oi_1 _08340_ (.A1(_02126_),
    .A2(_02128_),
    .Y(_02147_),
    .B1(_02124_));
 sg13g2_inv_1 _08341_ (.Y(_02148_),
    .A(_02147_));
 sg13g2_nor2_1 _08342_ (.A(net72),
    .B(_02002_),
    .Y(_02149_));
 sg13g2_nand3_1 _08343_ (.B(_01964_),
    .C(_03640_),
    .A(_01895_),
    .Y(_02150_));
 sg13g2_nand2_1 _08344_ (.Y(_02151_),
    .A(_02150_),
    .B(net72));
 sg13g2_nand3_1 _08345_ (.B(_02094_),
    .C(_01817_),
    .A(_02092_),
    .Y(_02152_));
 sg13g2_nand2_1 _08346_ (.Y(_02153_),
    .A(_02152_),
    .B(_01487_));
 sg13g2_nand3_1 _08347_ (.B(_01718_),
    .C(_01703_),
    .A(_01692_),
    .Y(_02154_));
 sg13g2_nand2_1 _08348_ (.Y(_02155_),
    .A(_02154_),
    .B(_01720_));
 sg13g2_nor2_1 _08349_ (.A(_02091_),
    .B(_01960_),
    .Y(_02156_));
 sg13g2_nand2_1 _08350_ (.Y(_02157_),
    .A(_01905_),
    .B(_02156_));
 sg13g2_nor2_1 _08351_ (.A(_02051_),
    .B(_02090_),
    .Y(_02158_));
 sg13g2_a21oi_1 _08352_ (.A1(_02093_),
    .A2(_02045_),
    .Y(_02159_),
    .B1(_02158_));
 sg13g2_nand2_1 _08353_ (.Y(_02160_),
    .A(_02157_),
    .B(_02159_));
 sg13g2_nor2_1 _08354_ (.A(_02155_),
    .B(_02160_),
    .Y(_02161_));
 sg13g2_nand2_1 _08355_ (.Y(_02162_),
    .A(_02161_),
    .B(_01706_));
 sg13g2_nand3_1 _08356_ (.B(_01891_),
    .C(_01804_),
    .A(_02156_),
    .Y(_02163_));
 sg13g2_nand3_1 _08357_ (.B(_02157_),
    .C(_02159_),
    .A(_02163_),
    .Y(_02164_));
 sg13g2_nand2_1 _08358_ (.Y(_02165_),
    .A(_02162_),
    .B(_02164_));
 sg13g2_inv_1 _08359_ (.Y(_02166_),
    .A(_02073_));
 sg13g2_a21oi_1 _08360_ (.A1(_02060_),
    .A2(_02075_),
    .Y(_02167_),
    .B1(_02166_));
 sg13g2_nor2_1 _08361_ (.A(_01112_),
    .B(_01649_),
    .Y(_02168_));
 sg13g2_xnor2_1 _08362_ (.Y(_02169_),
    .A(_02066_),
    .B(_02064_));
 sg13g2_xnor2_1 _08363_ (.Y(_02170_),
    .A(_02168_),
    .B(_02169_));
 sg13g2_nor2b_1 _08364_ (.A(_02058_),
    .B_N(_02055_),
    .Y(_02171_));
 sg13g2_a21oi_1 _08365_ (.A1(_02059_),
    .A2(_02052_),
    .Y(_02172_),
    .B1(_02171_));
 sg13g2_xnor2_1 _08366_ (.Y(_02173_),
    .A(_02170_),
    .B(_02172_));
 sg13g2_nand2_1 _08367_ (.Y(_02174_),
    .A(_01549_),
    .B(_00223_));
 sg13g2_nand3_1 _08368_ (.B(_01770_),
    .C(_00231_),
    .A(_01943_),
    .Y(_02175_));
 sg13g2_xnor2_1 _08369_ (.Y(_02176_),
    .A(_02174_),
    .B(_02175_));
 sg13g2_a22oi_1 _08370_ (.Y(_02177_),
    .B1(_02063_),
    .B2(_02065_),
    .A2(_02066_),
    .A1(_01923_));
 sg13g2_xnor2_1 _08371_ (.Y(_02178_),
    .A(_02062_),
    .B(_02177_));
 sg13g2_o21ai_1 _08372_ (.B1(_01936_),
    .Y(_02179_),
    .A1(_02062_),
    .A2(_02069_));
 sg13g2_xnor2_1 _08373_ (.Y(_02180_),
    .A(_02178_),
    .B(_02179_));
 sg13g2_xnor2_1 _08374_ (.Y(_02181_),
    .A(_02176_),
    .B(_02180_));
 sg13g2_xnor2_1 _08375_ (.Y(_02182_),
    .A(_02173_),
    .B(_02181_));
 sg13g2_xor2_1 _08376_ (.B(_02182_),
    .A(_02167_),
    .X(_02183_));
 sg13g2_and2_1 _08377_ (.A(_02089_),
    .B(_02083_),
    .X(_02184_));
 sg13g2_xor2_1 _08378_ (.B(_02184_),
    .A(_02183_),
    .X(_02185_));
 sg13g2_nand2_1 _08379_ (.Y(_02186_),
    .A(_02165_),
    .B(_02185_));
 sg13g2_inv_1 _08380_ (.Y(_02187_),
    .A(_02185_));
 sg13g2_nand3_1 _08381_ (.B(_02164_),
    .C(_02187_),
    .A(_02162_),
    .Y(_02188_));
 sg13g2_nand3_1 _08382_ (.B(_02188_),
    .C(_01502_),
    .A(_02186_),
    .Y(_02189_));
 sg13g2_nor2b_1 _08383_ (.A(_02153_),
    .B_N(_02189_),
    .Y(_02190_));
 sg13g2_nor2_1 _08384_ (.A(_02151_),
    .B(_02190_),
    .Y(_02191_));
 sg13g2_nor2_1 _08385_ (.A(_02149_),
    .B(_02191_),
    .Y(_02192_));
 sg13g2_buf_8 _08386_ (.A(_02192_),
    .X(_02193_));
 sg13g2_nand2_1 _08387_ (.Y(_02194_),
    .A(_02193_),
    .B(_01509_));
 sg13g2_inv_1 _08388_ (.Y(_02195_),
    .A(_02194_));
 sg13g2_nand2_2 _08389_ (.Y(_02196_),
    .A(net18),
    .B(_01998_));
 sg13g2_a21oi_1 _08390_ (.A1(_02033_),
    .A2(_02027_),
    .Y(_02197_),
    .B1(_02029_));
 sg13g2_xnor2_1 _08391_ (.Y(_02198_),
    .A(_02196_),
    .B(_02197_));
 sg13g2_xnor2_1 _08392_ (.Y(_02199_),
    .A(_02195_),
    .B(_02198_));
 sg13g2_nand2_1 _08393_ (.Y(_02200_),
    .A(_02194_),
    .B(_02196_));
 sg13g2_nand3_1 _08394_ (.B(net18),
    .C(_02104_),
    .A(_02193_),
    .Y(_02201_));
 sg13g2_and2_1 _08395_ (.A(_02200_),
    .B(_02201_),
    .X(_02202_));
 sg13g2_buf_8 _08396_ (.A(_02202_),
    .X(_02203_));
 sg13g2_inv_8 _08397_ (.Y(_02204_),
    .A(net18));
 sg13g2_nor2_1 _08398_ (.A(_01977_),
    .B(_02204_),
    .Y(_02205_));
 sg13g2_a22oi_1 _08399_ (.Y(_02206_),
    .B1(_02113_),
    .B2(_02110_),
    .A2(_02104_),
    .A1(_02205_));
 sg13g2_xor2_1 _08400_ (.B(_02206_),
    .A(_02203_),
    .X(_02207_));
 sg13g2_a21oi_1 _08401_ (.A1(_02116_),
    .A2(_02117_),
    .Y(_02208_),
    .B1(_02036_));
 sg13g2_a21oi_2 _08402_ (.B1(_02208_),
    .Y(_02209_),
    .A2(_02035_),
    .A1(_02119_));
 sg13g2_xnor2_1 _08403_ (.Y(_02210_),
    .A(_02207_),
    .B(_02209_));
 sg13g2_xnor2_1 _08404_ (.Y(_02211_),
    .A(_02199_),
    .B(_02210_));
 sg13g2_nand2_1 _08405_ (.Y(_02212_),
    .A(_02148_),
    .B(_02211_));
 sg13g2_xor2_1 _08406_ (.B(_02209_),
    .A(_02207_),
    .X(_02213_));
 sg13g2_nand2_1 _08407_ (.Y(_02214_),
    .A(_02213_),
    .B(_02199_));
 sg13g2_inv_1 _08408_ (.Y(_02215_),
    .A(_02199_));
 sg13g2_nand2_1 _08409_ (.Y(_02216_),
    .A(_02210_),
    .B(_02215_));
 sg13g2_nand2_1 _08410_ (.Y(_02217_),
    .A(_02214_),
    .B(_02216_));
 sg13g2_nand2_1 _08411_ (.Y(_02218_),
    .A(_02217_),
    .B(_02147_));
 sg13g2_nand2_1 _08412_ (.Y(_02219_),
    .A(_02212_),
    .B(_02218_));
 sg13g2_nand2b_1 _08413_ (.Y(_02220_),
    .B(_02219_),
    .A_N(_02146_));
 sg13g2_nand3_1 _08414_ (.B(_02218_),
    .C(_02146_),
    .A(_02212_),
    .Y(_02221_));
 sg13g2_nand2_1 _08415_ (.Y(_02222_),
    .A(_02220_),
    .B(_02221_));
 sg13g2_nor2_2 _08416_ (.A(_02145_),
    .B(_02222_),
    .Y(_02223_));
 sg13g2_nand2_1 _08417_ (.Y(_02224_),
    .A(_02209_),
    .B(_02207_));
 sg13g2_nor2_1 _08418_ (.A(_02207_),
    .B(_02209_),
    .Y(_02225_));
 sg13g2_a21oi_1 _08419_ (.A1(_02224_),
    .A2(_02199_),
    .Y(_02226_),
    .B1(_02225_));
 sg13g2_nand2_1 _08420_ (.Y(_02227_),
    .A(net18),
    .B(net19));
 sg13g2_nor3_2 _08421_ (.A(_02103_),
    .B(_02149_),
    .C(_02191_),
    .Y(_02228_));
 sg13g2_xnor2_1 _08422_ (.Y(_02229_),
    .A(_02227_),
    .B(_02228_));
 sg13g2_nand2_1 _08423_ (.Y(_02230_),
    .A(net20),
    .B(net19));
 sg13g2_nand2_1 _08424_ (.Y(_02231_),
    .A(_02201_),
    .B(_02230_));
 sg13g2_nand3_1 _08425_ (.B(_02200_),
    .C(_02231_),
    .A(_02229_),
    .Y(_02232_));
 sg13g2_nand2_1 _08426_ (.Y(_02233_),
    .A(_02231_),
    .B(_02200_));
 sg13g2_inv_2 _08427_ (.Y(_02234_),
    .A(_02229_));
 sg13g2_nand2_1 _08428_ (.Y(_02235_),
    .A(_02233_),
    .B(_02234_));
 sg13g2_nand2_1 _08429_ (.Y(_02236_),
    .A(_02232_),
    .B(_02235_));
 sg13g2_nand2_1 _08430_ (.Y(_02237_),
    .A(_02236_),
    .B(_02030_));
 sg13g2_nand3_1 _08431_ (.B(_02235_),
    .C(_02028_),
    .A(_02232_),
    .Y(_02238_));
 sg13g2_nand2_1 _08432_ (.Y(_02239_),
    .A(_02237_),
    .B(_02238_));
 sg13g2_nor2b_1 _08433_ (.A(_02203_),
    .B_N(_02230_),
    .Y(_02240_));
 sg13g2_nand2_1 _08434_ (.Y(_02241_),
    .A(_02206_),
    .B(_02203_));
 sg13g2_nand2b_1 _08435_ (.Y(_02242_),
    .B(_02241_),
    .A_N(_02240_));
 sg13g2_inv_1 _08436_ (.Y(_02243_),
    .A(_02242_));
 sg13g2_nand2_1 _08437_ (.Y(_02244_),
    .A(_02239_),
    .B(_02243_));
 sg13g2_nand3_1 _08438_ (.B(_02238_),
    .C(_02242_),
    .A(_02237_),
    .Y(_02245_));
 sg13g2_buf_8 _08439_ (.A(_02245_),
    .X(_02246_));
 sg13g2_nand2_1 _08440_ (.Y(_02247_),
    .A(_02244_),
    .B(_02246_));
 sg13g2_nor2_1 _08441_ (.A(_02028_),
    .B(_02032_),
    .Y(_02248_));
 sg13g2_xor2_1 _08442_ (.B(_02227_),
    .A(_02248_),
    .X(_02249_));
 sg13g2_xnor2_1 _08443_ (.Y(_02250_),
    .A(_02228_),
    .B(_02249_));
 sg13g2_nand2_1 _08444_ (.Y(_02251_),
    .A(_02247_),
    .B(_02250_));
 sg13g2_inv_1 _08445_ (.Y(_02252_),
    .A(_02250_));
 sg13g2_nand3_1 _08446_ (.B(_02246_),
    .C(_02252_),
    .A(_02244_),
    .Y(_02253_));
 sg13g2_nand2_1 _08447_ (.Y(_02254_),
    .A(_02251_),
    .B(_02253_));
 sg13g2_nand2b_1 _08448_ (.Y(_02255_),
    .B(_02254_),
    .A_N(_02226_));
 sg13g2_nand3_1 _08449_ (.B(_02253_),
    .C(_02226_),
    .A(_02251_),
    .Y(_02256_));
 sg13g2_nand2_1 _08450_ (.Y(_02257_),
    .A(_02255_),
    .B(_02256_));
 sg13g2_nor2_1 _08451_ (.A(_02196_),
    .B(_02197_),
    .Y(_02258_));
 sg13g2_nand2b_1 _08452_ (.Y(_02259_),
    .B(_02195_),
    .A_N(_02198_));
 sg13g2_nor2b_1 _08453_ (.A(_02258_),
    .B_N(_02259_),
    .Y(_02260_));
 sg13g2_nand2_1 _08454_ (.Y(_02261_),
    .A(_02257_),
    .B(_02260_));
 sg13g2_inv_1 _08455_ (.Y(_02262_),
    .A(_02260_));
 sg13g2_nand3_1 _08456_ (.B(_02256_),
    .C(_02262_),
    .A(_02255_),
    .Y(_02263_));
 sg13g2_nand2_1 _08457_ (.Y(_02264_),
    .A(_02261_),
    .B(_02263_));
 sg13g2_nor2_1 _08458_ (.A(_02147_),
    .B(_02217_),
    .Y(_02265_));
 sg13g2_a21oi_2 _08459_ (.B1(_02265_),
    .Y(_02266_),
    .A2(_02146_),
    .A1(_02218_));
 sg13g2_nand2_1 _08460_ (.Y(_02267_),
    .A(_02264_),
    .B(_02266_));
 sg13g2_nand2_1 _08461_ (.Y(_02268_),
    .A(_02223_),
    .B(_02267_));
 sg13g2_inv_1 _08462_ (.Y(_02269_),
    .A(_02266_));
 sg13g2_nand3_1 _08463_ (.B(_02263_),
    .C(_02261_),
    .A(_02269_),
    .Y(_02270_));
 sg13g2_buf_1 _08464_ (.A(_02270_),
    .X(_02271_));
 sg13g2_nand2_1 _08465_ (.Y(_02272_),
    .A(_02268_),
    .B(_02271_));
 sg13g2_a21oi_1 _08466_ (.A1(_02251_),
    .A2(_02253_),
    .Y(_02273_),
    .B1(_02226_));
 sg13g2_a21oi_2 _08467_ (.B1(_02273_),
    .Y(_02274_),
    .A2(_02262_),
    .A1(_02256_));
 sg13g2_inv_2 _08468_ (.Y(_02275_),
    .A(_02274_));
 sg13g2_nand2_1 _08469_ (.Y(_02276_),
    .A(_02193_),
    .B(net19));
 sg13g2_inv_2 _08470_ (.Y(_02277_),
    .A(_02276_));
 sg13g2_xnor2_1 _08471_ (.Y(_02278_),
    .A(_01977_),
    .B(net18));
 sg13g2_nand2_1 _08472_ (.Y(_02279_),
    .A(_02278_),
    .B(_02008_));
 sg13g2_xnor2_1 _08473_ (.Y(_02280_),
    .A(_02277_),
    .B(_02279_));
 sg13g2_nor2_1 _08474_ (.A(_02032_),
    .B(_02204_),
    .Y(_02281_));
 sg13g2_nand2_1 _08475_ (.Y(_02282_),
    .A(_02277_),
    .B(_02196_));
 sg13g2_xnor2_1 _08476_ (.Y(_02283_),
    .A(_02281_),
    .B(_02282_));
 sg13g2_inv_2 _08477_ (.Y(_02284_),
    .A(_02283_));
 sg13g2_nor2_1 _08478_ (.A(_02234_),
    .B(_02233_),
    .Y(_02285_));
 sg13g2_a21oi_2 _08479_ (.B1(_02285_),
    .Y(_02286_),
    .A2(_02030_),
    .A1(_02235_));
 sg13g2_xnor2_1 _08480_ (.Y(_02287_),
    .A(_02284_),
    .B(_02286_));
 sg13g2_xnor2_1 _08481_ (.Y(_02288_),
    .A(_02280_),
    .B(_02287_));
 sg13g2_a21oi_1 _08482_ (.A1(_02237_),
    .A2(_02238_),
    .Y(_02289_),
    .B1(_02242_));
 sg13g2_a21oi_1 _08483_ (.A1(_02246_),
    .A2(_02250_),
    .Y(_02290_),
    .B1(_02289_));
 sg13g2_inv_1 _08484_ (.Y(_02291_),
    .A(_02290_));
 sg13g2_nand2_1 _08485_ (.Y(_02292_),
    .A(_02288_),
    .B(_02291_));
 sg13g2_xnor2_1 _08486_ (.Y(_02293_),
    .A(_02283_),
    .B(_02286_));
 sg13g2_nand2_1 _08487_ (.Y(_02294_),
    .A(_02293_),
    .B(_02280_));
 sg13g2_inv_1 _08488_ (.Y(_02295_),
    .A(_02280_));
 sg13g2_nand2_1 _08489_ (.Y(_02296_),
    .A(_02287_),
    .B(_02295_));
 sg13g2_nand2_1 _08490_ (.Y(_02297_),
    .A(_02294_),
    .B(_02296_));
 sg13g2_nand2_1 _08491_ (.Y(_02298_),
    .A(_02297_),
    .B(_02290_));
 sg13g2_nand2_1 _08492_ (.Y(_02299_),
    .A(_02292_),
    .B(_02298_));
 sg13g2_nand2_2 _08493_ (.Y(_02300_),
    .A(net18),
    .B(_02030_));
 sg13g2_nor2_1 _08494_ (.A(_02019_),
    .B(_02300_),
    .Y(_02301_));
 sg13g2_nor2b_1 _08495_ (.A(_02249_),
    .B_N(_02228_),
    .Y(_02302_));
 sg13g2_nor2_1 _08496_ (.A(_02301_),
    .B(_02302_),
    .Y(_02303_));
 sg13g2_nand2_1 _08497_ (.Y(_02304_),
    .A(_02299_),
    .B(_02303_));
 sg13g2_inv_1 _08498_ (.Y(_02305_),
    .A(_02303_));
 sg13g2_nand3_1 _08499_ (.B(_02298_),
    .C(_02305_),
    .A(_02292_),
    .Y(_02306_));
 sg13g2_nand2_1 _08500_ (.Y(_02307_),
    .A(_02304_),
    .B(_02306_));
 sg13g2_xnor2_1 _08501_ (.Y(_02308_),
    .A(_02275_),
    .B(_02307_));
 sg13g2_nand2_1 _08502_ (.Y(_02309_),
    .A(_02272_),
    .B(_02308_));
 sg13g2_inv_1 _08503_ (.Y(_02310_),
    .A(_02307_));
 sg13g2_nand2_1 _08504_ (.Y(_02311_),
    .A(_02310_),
    .B(_02275_));
 sg13g2_nand2_1 _08505_ (.Y(_02312_),
    .A(_02307_),
    .B(_02274_));
 sg13g2_nand2_1 _08506_ (.Y(_02313_),
    .A(_02311_),
    .B(_02312_));
 sg13g2_nand3_1 _08507_ (.B(_02313_),
    .C(_02271_),
    .A(_02268_),
    .Y(_02314_));
 sg13g2_nand2_1 _08508_ (.Y(_02315_),
    .A(_02309_),
    .B(_02314_));
 sg13g2_buf_8 _08509_ (.A(_02315_),
    .X(_02316_));
 sg13g2_nor2_1 _08510_ (.A(net92),
    .B(_02316_),
    .Y(_02317_));
 sg13g2_nor2_1 _08511_ (.A(_02290_),
    .B(_02297_),
    .Y(_02318_));
 sg13g2_a21oi_2 _08512_ (.B1(_02318_),
    .Y(_02319_),
    .A2(_02305_),
    .A1(_02298_));
 sg13g2_nand2_1 _08513_ (.Y(_02320_),
    .A(_02286_),
    .B(_02284_));
 sg13g2_nor2_1 _08514_ (.A(_02284_),
    .B(_02286_),
    .Y(_02321_));
 sg13g2_a21oi_1 _08515_ (.A1(_02320_),
    .A2(_02280_),
    .Y(_02322_),
    .B1(_02321_));
 sg13g2_inv_1 _08516_ (.Y(_02323_),
    .A(_02322_));
 sg13g2_inv_1 _08517_ (.Y(_02324_),
    .A(_02281_));
 sg13g2_a21oi_1 _08518_ (.A1(_02324_),
    .A2(_02196_),
    .Y(_02325_),
    .B1(_02276_));
 sg13g2_inv_8 _08519_ (.Y(_02326_),
    .A(_02193_));
 sg13g2_nor2_1 _08520_ (.A(_02028_),
    .B(_02326_),
    .Y(_02327_));
 sg13g2_nand2_1 _08521_ (.Y(_02328_),
    .A(_02327_),
    .B(_02281_));
 sg13g2_nand2_1 _08522_ (.Y(_02329_),
    .A(_02193_),
    .B(_02008_));
 sg13g2_nand2_1 _08523_ (.Y(_02330_),
    .A(_02329_),
    .B(_02300_));
 sg13g2_nand2_1 _08524_ (.Y(_02331_),
    .A(_02328_),
    .B(_02330_));
 sg13g2_nand2_1 _08525_ (.Y(_02332_),
    .A(_02331_),
    .B(_01977_));
 sg13g2_nand3_1 _08526_ (.B(net20),
    .C(_02330_),
    .A(_02328_),
    .Y(_02333_));
 sg13g2_nand2_1 _08527_ (.Y(_02334_),
    .A(_02332_),
    .B(_02333_));
 sg13g2_nand2b_1 _08528_ (.Y(_02335_),
    .B(_02334_),
    .A_N(_02325_));
 sg13g2_nand3_1 _08529_ (.B(_02333_),
    .C(_02325_),
    .A(_02332_),
    .Y(_02336_));
 sg13g2_nand2_1 _08530_ (.Y(_02337_),
    .A(_02335_),
    .B(_02336_));
 sg13g2_nand2_1 _08531_ (.Y(_02338_),
    .A(_02278_),
    .B(_02030_));
 sg13g2_xor2_1 _08532_ (.B(_02338_),
    .A(_02329_),
    .X(_02339_));
 sg13g2_nand2_1 _08533_ (.Y(_02340_),
    .A(_02337_),
    .B(_02339_));
 sg13g2_inv_1 _08534_ (.Y(_02341_),
    .A(_02339_));
 sg13g2_nand3_1 _08535_ (.B(_02336_),
    .C(_02341_),
    .A(_02335_),
    .Y(_02342_));
 sg13g2_nand2_1 _08536_ (.Y(_02343_),
    .A(_02340_),
    .B(_02342_));
 sg13g2_nand2_1 _08537_ (.Y(_02344_),
    .A(_02323_),
    .B(_02343_));
 sg13g2_inv_2 _08538_ (.Y(_02345_),
    .A(_02343_));
 sg13g2_nand2_1 _08539_ (.Y(_02346_),
    .A(_02322_),
    .B(_02345_));
 sg13g2_nand2_1 _08540_ (.Y(_02347_),
    .A(_02344_),
    .B(_02346_));
 sg13g2_nor2_1 _08541_ (.A(_02276_),
    .B(_02279_),
    .Y(_02348_));
 sg13g2_nand2_1 _08542_ (.Y(_02349_),
    .A(_02205_),
    .B(_02008_));
 sg13g2_nor2b_1 _08543_ (.A(_02348_),
    .B_N(_02349_),
    .Y(_02350_));
 sg13g2_nand2_1 _08544_ (.Y(_02351_),
    .A(_02347_),
    .B(_02350_));
 sg13g2_inv_1 _08545_ (.Y(_02352_),
    .A(_02350_));
 sg13g2_nand3_1 _08546_ (.B(_02346_),
    .C(_02352_),
    .A(_02344_),
    .Y(_02353_));
 sg13g2_nand2_1 _08547_ (.Y(_02354_),
    .A(_02351_),
    .B(_02353_));
 sg13g2_xnor2_1 _08548_ (.Y(_02355_),
    .A(_02319_),
    .B(_02354_));
 sg13g2_buf_1 _08549_ (.A(_02355_),
    .X(_02356_));
 sg13g2_nand2_1 _08550_ (.Y(_02357_),
    .A(_02264_),
    .B(_02269_));
 sg13g2_nand3_1 _08551_ (.B(_02266_),
    .C(_02263_),
    .A(_02261_),
    .Y(_02358_));
 sg13g2_nand2_1 _08552_ (.Y(_02359_),
    .A(_02357_),
    .B(_02358_));
 sg13g2_nand3_1 _08553_ (.B(_02308_),
    .C(_02223_),
    .A(_02359_),
    .Y(_02360_));
 sg13g2_nor2_1 _08554_ (.A(_02266_),
    .B(_02264_),
    .Y(_02361_));
 sg13g2_nand2_1 _08555_ (.Y(_02362_),
    .A(_02361_),
    .B(_02312_));
 sg13g2_nand2_1 _08556_ (.Y(_02363_),
    .A(_02362_),
    .B(_02311_));
 sg13g2_inv_1 _08557_ (.Y(_02364_),
    .A(_02363_));
 sg13g2_nand2_1 _08558_ (.Y(_02365_),
    .A(_02360_),
    .B(_02364_));
 sg13g2_nand2b_1 _08559_ (.Y(_02366_),
    .B(_02365_),
    .A_N(_02356_));
 sg13g2_nand3_1 _08560_ (.B(_02364_),
    .C(_02356_),
    .A(_02360_),
    .Y(_02367_));
 sg13g2_buf_1 _08561_ (.A(_02367_),
    .X(_02368_));
 sg13g2_buf_8 _08562_ (.A(net90),
    .X(_02369_));
 sg13g2_nand3_1 _08563_ (.B(_02368_),
    .C(net73),
    .A(_02366_),
    .Y(_02370_));
 sg13g2_nand2b_1 _08564_ (.Y(_02371_),
    .B(_02370_),
    .A_N(_02317_));
 sg13g2_nand2_1 _08565_ (.Y(_02372_),
    .A(_02271_),
    .B(_02267_));
 sg13g2_nand2b_1 _08566_ (.Y(_02373_),
    .B(_02372_),
    .A_N(_02223_));
 sg13g2_nand2_1 _08567_ (.Y(_02374_),
    .A(_02359_),
    .B(_02223_));
 sg13g2_nand2_1 _08568_ (.Y(_02375_),
    .A(_02373_),
    .B(_02374_));
 sg13g2_buf_8 _08569_ (.A(_02375_),
    .X(_02376_));
 sg13g2_nor2_1 _08570_ (.A(net91),
    .B(_02376_),
    .Y(_02377_));
 sg13g2_nand3_1 _08571_ (.B(_02314_),
    .C(net73),
    .A(_02309_),
    .Y(_02378_));
 sg13g2_nand3_1 _08572_ (.B(_02368_),
    .C(net110),
    .A(_02366_),
    .Y(_02379_));
 sg13g2_nor2_1 _08573_ (.A(_02378_),
    .B(_02379_),
    .Y(_02380_));
 sg13g2_a21oi_1 _08574_ (.A1(_02371_),
    .A2(_02377_),
    .Y(_02381_),
    .B1(_02380_));
 sg13g2_nand3_1 _08575_ (.B(_02221_),
    .C(_02144_),
    .A(_02220_),
    .Y(_02382_));
 sg13g2_inv_1 _08576_ (.Y(_02383_),
    .A(_02267_));
 sg13g2_a21oi_1 _08577_ (.A1(_02271_),
    .A2(_02382_),
    .Y(_02384_),
    .B1(_02383_));
 sg13g2_nor2_1 _08578_ (.A(_02356_),
    .B(_02313_),
    .Y(_02385_));
 sg13g2_nand2_1 _08579_ (.Y(_02386_),
    .A(_02384_),
    .B(_02385_));
 sg13g2_nor2_1 _08580_ (.A(_02274_),
    .B(_02307_),
    .Y(_02387_));
 sg13g2_nand2_1 _08581_ (.Y(_02388_),
    .A(_02354_),
    .B(_02319_));
 sg13g2_nand2_1 _08582_ (.Y(_02390_),
    .A(_02387_),
    .B(_02388_));
 sg13g2_nor2_1 _08583_ (.A(_02319_),
    .B(_02354_),
    .Y(_02391_));
 sg13g2_inv_1 _08584_ (.Y(_02392_),
    .A(_02391_));
 sg13g2_nand2_1 _08585_ (.Y(_02393_),
    .A(_02390_),
    .B(_02392_));
 sg13g2_inv_1 _08586_ (.Y(_02394_),
    .A(_02393_));
 sg13g2_nand2_1 _08587_ (.Y(_02395_),
    .A(_02386_),
    .B(_02394_));
 sg13g2_inv_1 _08588_ (.Y(_02396_),
    .A(_02344_));
 sg13g2_a21oi_1 _08589_ (.A1(_02346_),
    .A2(_02352_),
    .Y(_02397_),
    .B1(_02396_));
 sg13g2_inv_1 _08590_ (.Y(_02398_),
    .A(_02300_));
 sg13g2_inv_1 _08591_ (.Y(_02399_),
    .A(_02327_));
 sg13g2_nor2_1 _08592_ (.A(_02399_),
    .B(_02279_),
    .Y(_02401_));
 sg13g2_a21oi_1 _08593_ (.A1(net20),
    .A2(_02398_),
    .Y(_02402_),
    .B1(_02401_));
 sg13g2_inv_1 _08594_ (.Y(_02403_),
    .A(_02402_));
 sg13g2_nor2_1 _08595_ (.A(_02204_),
    .B(_02326_),
    .Y(_02404_));
 sg13g2_a22oi_1 _08596_ (.Y(_02405_),
    .B1(net20),
    .B2(_02330_),
    .A2(_02248_),
    .A1(_02404_));
 sg13g2_inv_2 _08597_ (.Y(_02406_),
    .A(_02336_));
 sg13g2_a21oi_1 _08598_ (.A1(_02335_),
    .A2(_02339_),
    .Y(_02407_),
    .B1(_02406_));
 sg13g2_nor2_1 _08599_ (.A(_02405_),
    .B(_02407_),
    .Y(_02408_));
 sg13g2_nand2_1 _08600_ (.Y(_02409_),
    .A(_02407_),
    .B(_02405_));
 sg13g2_nor2b_1 _08601_ (.A(_02408_),
    .B_N(_02409_),
    .Y(_02410_));
 sg13g2_xnor2_1 _08602_ (.Y(_02412_),
    .A(_02403_),
    .B(_02410_));
 sg13g2_xor2_1 _08603_ (.B(_02412_),
    .A(_02397_),
    .X(_02413_));
 sg13g2_nand2_1 _08604_ (.Y(_02414_),
    .A(_02395_),
    .B(_02413_));
 sg13g2_inv_1 _08605_ (.Y(_02415_),
    .A(_02413_));
 sg13g2_nand3_1 _08606_ (.B(_02394_),
    .C(_02415_),
    .A(_02386_),
    .Y(_02416_));
 sg13g2_buf_8 _08607_ (.A(_02416_),
    .X(_02417_));
 sg13g2_nand2_2 _08608_ (.Y(_02418_),
    .A(_02414_),
    .B(_02417_));
 sg13g2_nor2_2 _08609_ (.A(net92),
    .B(_02418_),
    .Y(_02419_));
 sg13g2_inv_4 _08610_ (.A(_02370_),
    .Y(_02420_));
 sg13g2_nand2_1 _08611_ (.Y(_02421_),
    .A(_02419_),
    .B(_02420_));
 sg13g2_nand3_1 _08612_ (.B(_02417_),
    .C(net73),
    .A(_02414_),
    .Y(_02423_));
 sg13g2_nand2_1 _08613_ (.Y(_02424_),
    .A(_02423_),
    .B(_02379_));
 sg13g2_nand2_1 _08614_ (.Y(_02425_),
    .A(_02421_),
    .B(_02424_));
 sg13g2_nor2_1 _08615_ (.A(net91),
    .B(_02316_),
    .Y(_02426_));
 sg13g2_nand2_1 _08616_ (.Y(_02427_),
    .A(_02425_),
    .B(_02426_));
 sg13g2_inv_1 _08617_ (.Y(_02428_),
    .A(_02426_));
 sg13g2_nand3_1 _08618_ (.B(_02424_),
    .C(_02428_),
    .A(_02421_),
    .Y(_02429_));
 sg13g2_nand2_1 _08619_ (.Y(_02430_),
    .A(_02427_),
    .B(_02429_));
 sg13g2_nand2b_1 _08620_ (.Y(_02431_),
    .B(_02430_),
    .A_N(_02381_));
 sg13g2_nand3_1 _08621_ (.B(_02429_),
    .C(_02381_),
    .A(_02427_),
    .Y(_02432_));
 sg13g2_nand2_1 _08622_ (.Y(_02434_),
    .A(_02431_),
    .B(_02432_));
 sg13g2_nand3b_1 _08623_ (.B(_02136_),
    .C(_02142_),
    .Y(_02435_),
    .A_N(_02144_));
 sg13g2_inv_1 _08624_ (.Y(_02436_),
    .A(_02143_));
 sg13g2_nand2_1 _08625_ (.Y(_02437_),
    .A(_02436_),
    .B(_02135_));
 sg13g2_nand2b_1 _08626_ (.Y(_02438_),
    .B(_02143_),
    .A_N(_02135_));
 sg13g2_nand3b_1 _08627_ (.B(_02437_),
    .C(_02438_),
    .Y(_02439_),
    .A_N(_02142_));
 sg13g2_nand2_2 _08628_ (.Y(_02440_),
    .A(_02435_),
    .B(_02439_));
 sg13g2_nor2_1 _08629_ (.A(_00198_),
    .B(_02440_),
    .Y(_02441_));
 sg13g2_xnor2_1 _08630_ (.Y(_02442_),
    .A(_02145_),
    .B(_02222_));
 sg13g2_buf_8 _08631_ (.A(_02442_),
    .X(_02443_));
 sg13g2_nor2_1 _08632_ (.A(net104),
    .B(_02443_),
    .Y(_02445_));
 sg13g2_nor2_1 _08633_ (.A(net111),
    .B(_02376_),
    .Y(_02446_));
 sg13g2_xnor2_1 _08634_ (.Y(_02447_),
    .A(_02445_),
    .B(_02446_));
 sg13g2_xnor2_1 _08635_ (.Y(_02448_),
    .A(_02441_),
    .B(_02447_));
 sg13g2_nand2_1 _08636_ (.Y(_02449_),
    .A(_02434_),
    .B(_02448_));
 sg13g2_inv_1 _08637_ (.Y(_02450_),
    .A(_02448_));
 sg13g2_nand3_1 _08638_ (.B(_02432_),
    .C(_02450_),
    .A(_02431_),
    .Y(_02451_));
 sg13g2_nand2_1 _08639_ (.Y(_02452_),
    .A(_02420_),
    .B(_02317_));
 sg13g2_nand2_1 _08640_ (.Y(_02453_),
    .A(_02452_),
    .B(_02371_));
 sg13g2_nand2_1 _08641_ (.Y(_02454_),
    .A(_02453_),
    .B(_02377_));
 sg13g2_inv_1 _08642_ (.Y(_02456_),
    .A(_02377_));
 sg13g2_nand3_1 _08643_ (.B(_02371_),
    .C(_02456_),
    .A(_02452_),
    .Y(_02457_));
 sg13g2_buf_8 _08644_ (.A(net101),
    .X(_02458_));
 sg13g2_nor2_1 _08645_ (.A(net89),
    .B(_02376_),
    .Y(_02459_));
 sg13g2_nor2_1 _08646_ (.A(net91),
    .B(_02443_),
    .Y(_02460_));
 sg13g2_inv_1 _08647_ (.Y(_02461_),
    .A(_02376_));
 sg13g2_nand2_1 _08648_ (.Y(_02462_),
    .A(_02461_),
    .B(net110));
 sg13g2_nand2_1 _08649_ (.Y(_02463_),
    .A(_02378_),
    .B(_02462_));
 sg13g2_a22oi_1 _08650_ (.Y(_02464_),
    .B1(_02460_),
    .B2(_02463_),
    .A2(_02459_),
    .A1(_02317_));
 sg13g2_nand3_1 _08651_ (.B(_02457_),
    .C(_02464_),
    .A(_02454_),
    .Y(_02465_));
 sg13g2_buf_8 _08652_ (.A(_00198_),
    .X(_02467_));
 sg13g2_xnor2_1 _08653_ (.Y(_02468_),
    .A(_02138_),
    .B(_02141_));
 sg13g2_buf_8 _08654_ (.A(_02468_),
    .X(_02469_));
 sg13g2_nor2_1 _08655_ (.A(net88),
    .B(_02469_),
    .Y(_02470_));
 sg13g2_inv_1 _08656_ (.Y(_02471_),
    .A(_02440_));
 sg13g2_nand2_1 _08657_ (.Y(_02472_),
    .A(_02471_),
    .B(net119));
 sg13g2_nor2_1 _08658_ (.A(net111),
    .B(_02443_),
    .Y(_02473_));
 sg13g2_inv_1 _08659_ (.Y(_02474_),
    .A(_02473_));
 sg13g2_nor2_1 _08660_ (.A(_02472_),
    .B(_02474_),
    .Y(_02475_));
 sg13g2_nand2_1 _08661_ (.Y(_02476_),
    .A(_02474_),
    .B(_02472_));
 sg13g2_nand2b_1 _08662_ (.Y(_02478_),
    .B(_02476_),
    .A_N(_02475_));
 sg13g2_xnor2_1 _08663_ (.Y(_02479_),
    .A(_02470_),
    .B(_02478_));
 sg13g2_a21oi_1 _08664_ (.A1(_02454_),
    .A2(_02457_),
    .Y(_02480_),
    .B1(_02464_));
 sg13g2_a21oi_1 _08665_ (.A1(_02465_),
    .A2(_02479_),
    .Y(_02481_),
    .B1(_02480_));
 sg13g2_nand3_1 _08666_ (.B(_02451_),
    .C(_02481_),
    .A(_02449_),
    .Y(_02482_));
 sg13g2_a21oi_1 _08667_ (.A1(_02476_),
    .A2(_02470_),
    .Y(_02483_),
    .B1(_02475_));
 sg13g2_inv_1 _08668_ (.Y(_02484_),
    .A(_02483_));
 sg13g2_nand2_1 _08669_ (.Y(_02485_),
    .A(_02449_),
    .B(_02451_));
 sg13g2_nand2b_1 _08670_ (.Y(_02486_),
    .B(_02485_),
    .A_N(_02481_));
 sg13g2_inv_1 _08671_ (.Y(_02487_),
    .A(_02486_));
 sg13g2_a21oi_1 _08672_ (.A1(_02482_),
    .A2(_02484_),
    .Y(_02489_),
    .B1(_02487_));
 sg13g2_inv_1 _08673_ (.Y(_02490_),
    .A(_02431_));
 sg13g2_a21oi_1 _08674_ (.A1(_02432_),
    .A2(_02448_),
    .Y(_02491_),
    .B1(_02490_));
 sg13g2_a22oi_1 _08675_ (.Y(_02492_),
    .B1(_02426_),
    .B2(_02424_),
    .A2(_02420_),
    .A1(_02419_));
 sg13g2_nor2_1 _08676_ (.A(_02415_),
    .B(_02356_),
    .Y(_02493_));
 sg13g2_nand2_1 _08677_ (.Y(_02494_),
    .A(_02413_),
    .B(_02391_));
 sg13g2_or2_1 _08678_ (.X(_02495_),
    .B(_02412_),
    .A(_02397_));
 sg13g2_buf_1 _08679_ (.A(_02495_),
    .X(_02496_));
 sg13g2_nand2_1 _08680_ (.Y(_02497_),
    .A(_02494_),
    .B(_02496_));
 sg13g2_a21oi_1 _08681_ (.A1(_02363_),
    .A2(_02493_),
    .Y(_02498_),
    .B1(_02497_));
 sg13g2_nand4_1 _08682_ (.B(_02308_),
    .C(_02493_),
    .A(_02359_),
    .Y(_02500_),
    .D(_02223_));
 sg13g2_nand2_1 _08683_ (.Y(_02501_),
    .A(_02498_),
    .B(_02500_));
 sg13g2_nor2_1 _08684_ (.A(_02205_),
    .B(_02327_),
    .Y(_02502_));
 sg13g2_nor3_1 _08685_ (.A(_02326_),
    .B(_01977_),
    .C(_02300_),
    .Y(_02503_));
 sg13g2_nor3_2 _08686_ (.A(_02204_),
    .B(_02502_),
    .C(_02503_),
    .Y(_02504_));
 sg13g2_a21oi_1 _08687_ (.A1(_02204_),
    .A2(_02399_),
    .Y(_02505_),
    .B1(_02504_));
 sg13g2_inv_1 _08688_ (.Y(_02506_),
    .A(_02505_));
 sg13g2_a21oi_1 _08689_ (.A1(_02409_),
    .A2(_02403_),
    .Y(_02507_),
    .B1(_02408_));
 sg13g2_nor2_1 _08690_ (.A(_02506_),
    .B(_02507_),
    .Y(_02508_));
 sg13g2_inv_2 _08691_ (.Y(_02509_),
    .A(_02508_));
 sg13g2_nand2_1 _08692_ (.Y(_02511_),
    .A(_02507_),
    .B(_02506_));
 sg13g2_nand2_1 _08693_ (.Y(_02512_),
    .A(_02509_),
    .B(_02511_));
 sg13g2_inv_2 _08694_ (.Y(_02513_),
    .A(_02512_));
 sg13g2_nand2_2 _08695_ (.Y(_02514_),
    .A(_02501_),
    .B(_02513_));
 sg13g2_nand3_1 _08696_ (.B(_02512_),
    .C(_02500_),
    .A(_02498_),
    .Y(_02515_));
 sg13g2_buf_8 _08697_ (.A(_02515_),
    .X(_02516_));
 sg13g2_nand2_2 _08698_ (.Y(_02517_),
    .A(_02514_),
    .B(_02516_));
 sg13g2_nor2_1 _08699_ (.A(net89),
    .B(_02517_),
    .Y(_02518_));
 sg13g2_nand2_1 _08700_ (.Y(_02519_),
    .A(_02518_),
    .B(_02419_));
 sg13g2_nand3_1 _08701_ (.B(_02516_),
    .C(_02369_),
    .A(_02514_),
    .Y(_02520_));
 sg13g2_inv_2 _08702_ (.Y(_02522_),
    .A(_02419_));
 sg13g2_nand2_1 _08703_ (.Y(_02523_),
    .A(_02520_),
    .B(_02522_));
 sg13g2_nand2_1 _08704_ (.Y(_02524_),
    .A(_02519_),
    .B(_02523_));
 sg13g2_nand2_2 _08705_ (.Y(_02525_),
    .A(_02366_),
    .B(_02368_));
 sg13g2_nor2_1 _08706_ (.A(net76),
    .B(_02525_),
    .Y(_02526_));
 sg13g2_nand2_1 _08707_ (.Y(_02527_),
    .A(_02524_),
    .B(_02526_));
 sg13g2_inv_1 _08708_ (.Y(_02528_),
    .A(_02526_));
 sg13g2_nand3_1 _08709_ (.B(_02523_),
    .C(_02528_),
    .A(_02519_),
    .Y(_02529_));
 sg13g2_nand2_1 _08710_ (.Y(_02530_),
    .A(_02527_),
    .B(_02529_));
 sg13g2_nand2b_1 _08711_ (.Y(_02531_),
    .B(_02530_),
    .A_N(_02492_));
 sg13g2_nand3_1 _08712_ (.B(_02529_),
    .C(_02492_),
    .A(_02527_),
    .Y(_02533_));
 sg13g2_nand2_1 _08713_ (.Y(_02534_),
    .A(_02531_),
    .B(_02533_));
 sg13g2_nor2_1 _08714_ (.A(net88),
    .B(_02443_),
    .Y(_02535_));
 sg13g2_nand2_1 _08715_ (.Y(_02536_),
    .A(_02461_),
    .B(net119));
 sg13g2_o21ai_1 _08716_ (.B1(_02536_),
    .Y(_02537_),
    .A1(net111),
    .A2(_02316_));
 sg13g2_nor2_1 _08717_ (.A(net104),
    .B(_02316_),
    .Y(_02538_));
 sg13g2_nand2_1 _08718_ (.Y(_02539_),
    .A(_02538_),
    .B(_02446_));
 sg13g2_nand2_1 _08719_ (.Y(_02540_),
    .A(_02537_),
    .B(_02539_));
 sg13g2_xnor2_1 _08720_ (.Y(_02541_),
    .A(_02535_),
    .B(_02540_));
 sg13g2_nand2_1 _08721_ (.Y(_02542_),
    .A(_02534_),
    .B(_02541_));
 sg13g2_inv_1 _08722_ (.Y(_02544_),
    .A(_02541_));
 sg13g2_nand3_1 _08723_ (.B(_02533_),
    .C(_02544_),
    .A(_02531_),
    .Y(_02545_));
 sg13g2_nand2_1 _08724_ (.Y(_02546_),
    .A(_02542_),
    .B(_02545_));
 sg13g2_nand2b_1 _08725_ (.Y(_02547_),
    .B(_02546_),
    .A_N(_02491_));
 sg13g2_nand3_1 _08726_ (.B(_02545_),
    .C(_02491_),
    .A(_02542_),
    .Y(_02548_));
 sg13g2_nand2_1 _08727_ (.Y(_02549_),
    .A(_02547_),
    .B(_02548_));
 sg13g2_nor2_1 _08728_ (.A(_02474_),
    .B(_02536_),
    .Y(_02550_));
 sg13g2_nand2b_1 _08729_ (.Y(_02551_),
    .B(_02441_),
    .A_N(_02447_));
 sg13g2_nor2b_1 _08730_ (.A(_02550_),
    .B_N(_02551_),
    .Y(_02552_));
 sg13g2_inv_1 _08731_ (.Y(_02553_),
    .A(_02552_));
 sg13g2_nand2_1 _08732_ (.Y(_02555_),
    .A(_02549_),
    .B(_02553_));
 sg13g2_nand3_1 _08733_ (.B(_02548_),
    .C(_02552_),
    .A(_02547_),
    .Y(_02556_));
 sg13g2_nand2_1 _08734_ (.Y(_02557_),
    .A(_02555_),
    .B(_02556_));
 sg13g2_nand2b_1 _08735_ (.Y(_02558_),
    .B(_02557_),
    .A_N(_02489_));
 sg13g2_nand3_1 _08736_ (.B(_02556_),
    .C(_02489_),
    .A(_02555_),
    .Y(_02559_));
 sg13g2_nand2_1 _08737_ (.Y(_02560_),
    .A(_02558_),
    .B(_02559_));
 sg13g2_inv_4 _08738_ (.A(net118),
    .Y(_02561_));
 sg13g2_buf_8 _08739_ (.A(_02561_),
    .X(_02562_));
 sg13g2_nor2_1 _08740_ (.A(net87),
    .B(_02440_),
    .Y(_02563_));
 sg13g2_inv_1 _08741_ (.Y(_02564_),
    .A(_02563_));
 sg13g2_nand2_1 _08742_ (.Y(_02566_),
    .A(_02560_),
    .B(_02564_));
 sg13g2_nand3_1 _08743_ (.B(_02559_),
    .C(_02563_),
    .A(_02558_),
    .Y(_02567_));
 sg13g2_nand2_1 _08744_ (.Y(_02568_),
    .A(_02566_),
    .B(_02567_));
 sg13g2_nand2_1 _08745_ (.Y(_02569_),
    .A(_02486_),
    .B(_02482_));
 sg13g2_nand2_1 _08746_ (.Y(_02570_),
    .A(_02569_),
    .B(_02484_));
 sg13g2_nand3_1 _08747_ (.B(_02482_),
    .C(_02483_),
    .A(_02486_),
    .Y(_02571_));
 sg13g2_nand2_1 _08748_ (.Y(_02572_),
    .A(_02454_),
    .B(_02457_));
 sg13g2_nand2b_1 _08749_ (.Y(_02573_),
    .B(_02572_),
    .A_N(_02464_));
 sg13g2_nand2_1 _08750_ (.Y(_02574_),
    .A(_02573_),
    .B(_02465_));
 sg13g2_nand2_1 _08751_ (.Y(_02575_),
    .A(_02574_),
    .B(_02479_));
 sg13g2_inv_1 _08752_ (.Y(_02576_),
    .A(_02479_));
 sg13g2_nand3_1 _08753_ (.B(_02465_),
    .C(_02576_),
    .A(_02573_),
    .Y(_02577_));
 sg13g2_nand2_1 _08754_ (.Y(_02578_),
    .A(_02317_),
    .B(_02459_));
 sg13g2_nand2_1 _08755_ (.Y(_02579_),
    .A(_02578_),
    .B(_02463_));
 sg13g2_nand2b_1 _08756_ (.Y(_02580_),
    .B(_02579_),
    .A_N(_02460_));
 sg13g2_nand3_1 _08757_ (.B(_02463_),
    .C(_02460_),
    .A(_02578_),
    .Y(_02581_));
 sg13g2_nand2_1 _08758_ (.Y(_02582_),
    .A(_02580_),
    .B(_02581_));
 sg13g2_nor2_1 _08759_ (.A(net92),
    .B(_02443_),
    .Y(_02583_));
 sg13g2_inv_1 _08760_ (.Y(_02584_),
    .A(_02583_));
 sg13g2_o21ai_1 _08761_ (.B1(_02584_),
    .Y(_02585_),
    .A1(net89),
    .A2(_02376_));
 sg13g2_nor2_1 _08762_ (.A(_05494_),
    .B(_02440_),
    .Y(_02587_));
 sg13g2_nand2_1 _08763_ (.Y(_02588_),
    .A(_02459_),
    .B(_02583_));
 sg13g2_inv_1 _08764_ (.Y(_02589_),
    .A(_02588_));
 sg13g2_a21oi_1 _08765_ (.A1(_02585_),
    .A2(_02587_),
    .Y(_02590_),
    .B1(_02589_));
 sg13g2_nand2_1 _08766_ (.Y(_02591_),
    .A(_02582_),
    .B(_02590_));
 sg13g2_nor2_2 _08767_ (.A(_01509_),
    .B(_02103_),
    .Y(_02592_));
 sg13g2_nor2b_1 _08768_ (.A(_02592_),
    .B_N(net19),
    .Y(_02593_));
 sg13g2_o21ai_1 _08769_ (.B1(_02138_),
    .Y(_02594_),
    .A1(_02137_),
    .A2(_02593_));
 sg13g2_buf_2 _08770_ (.A(_02594_),
    .X(_02595_));
 sg13g2_nor2_1 _08771_ (.A(net88),
    .B(_02595_),
    .Y(_02596_));
 sg13g2_nand2b_1 _08772_ (.Y(_02598_),
    .B(net102),
    .A_N(_02469_));
 sg13g2_nand2_1 _08773_ (.Y(_02599_),
    .A(_02471_),
    .B(net102));
 sg13g2_nor2_1 _08774_ (.A(net104),
    .B(_02469_),
    .Y(_02600_));
 sg13g2_inv_1 _08775_ (.Y(_02601_),
    .A(_02600_));
 sg13g2_nand2_1 _08776_ (.Y(_02602_),
    .A(_02599_),
    .B(_02601_));
 sg13g2_o21ai_1 _08777_ (.B1(_02602_),
    .Y(_02603_),
    .A1(_02472_),
    .A2(_02598_));
 sg13g2_xnor2_1 _08778_ (.Y(_02604_),
    .A(_02596_),
    .B(_02603_));
 sg13g2_inv_1 _08779_ (.Y(_02605_),
    .A(_02590_));
 sg13g2_nand3_1 _08780_ (.B(_02581_),
    .C(_02605_),
    .A(_02580_),
    .Y(_02606_));
 sg13g2_inv_1 _08781_ (.Y(_02607_),
    .A(_02606_));
 sg13g2_a21oi_1 _08782_ (.A1(_02591_),
    .A2(_02604_),
    .Y(_02609_),
    .B1(_02607_));
 sg13g2_nand3_1 _08783_ (.B(_02577_),
    .C(_02609_),
    .A(_02575_),
    .Y(_02610_));
 sg13g2_nor2_1 _08784_ (.A(_02601_),
    .B(_02599_),
    .Y(_02611_));
 sg13g2_a21oi_1 _08785_ (.A1(_02602_),
    .A2(_02596_),
    .Y(_02612_),
    .B1(_02611_));
 sg13g2_inv_1 _08786_ (.Y(_02613_),
    .A(_02612_));
 sg13g2_a21oi_1 _08787_ (.A1(_02575_),
    .A2(_02577_),
    .Y(_02614_),
    .B1(_02609_));
 sg13g2_a21oi_1 _08788_ (.A1(_02610_),
    .A2(_02613_),
    .Y(_02615_),
    .B1(_02614_));
 sg13g2_nand3_1 _08789_ (.B(_02571_),
    .C(_02615_),
    .A(_02570_),
    .Y(_02616_));
 sg13g2_nor2_1 _08790_ (.A(_02561_),
    .B(_02469_),
    .Y(_02617_));
 sg13g2_nand2_1 _08791_ (.Y(_02618_),
    .A(_02570_),
    .B(_02571_));
 sg13g2_nand2b_1 _08792_ (.Y(_02620_),
    .B(_02618_),
    .A_N(_02615_));
 sg13g2_inv_1 _08793_ (.Y(_02621_),
    .A(_02620_));
 sg13g2_a21oi_1 _08794_ (.A1(_02616_),
    .A2(_02617_),
    .Y(_02622_),
    .B1(_02621_));
 sg13g2_nand2_1 _08795_ (.Y(_02623_),
    .A(_02568_),
    .B(_02622_));
 sg13g2_inv_1 _08796_ (.Y(_02624_),
    .A(_02622_));
 sg13g2_nand3_1 _08797_ (.B(_02567_),
    .C(_02624_),
    .A(_02566_),
    .Y(_02625_));
 sg13g2_buf_1 _08798_ (.A(_02625_),
    .X(_02626_));
 sg13g2_nand2_1 _08799_ (.Y(_02627_),
    .A(_02623_),
    .B(_02626_));
 sg13g2_inv_1 _08800_ (.Y(_02628_),
    .A(_02558_));
 sg13g2_a21oi_1 _08801_ (.A1(_02559_),
    .A2(_02563_),
    .Y(_02629_),
    .B1(_02628_));
 sg13g2_inv_1 _08802_ (.Y(_02631_),
    .A(_02629_));
 sg13g2_nor2_1 _08803_ (.A(net87),
    .B(_02443_),
    .Y(_02632_));
 sg13g2_a21oi_1 _08804_ (.A1(_02542_),
    .A2(_02545_),
    .Y(_02633_),
    .B1(_02491_));
 sg13g2_a21oi_1 _08805_ (.A1(_02548_),
    .A2(_02553_),
    .Y(_02634_),
    .B1(_02633_));
 sg13g2_a21oi_1 _08806_ (.A1(_02527_),
    .A2(_02529_),
    .Y(_02635_),
    .B1(_02492_));
 sg13g2_a21oi_1 _08807_ (.A1(_02533_),
    .A2(_02541_),
    .Y(_02636_),
    .B1(_02635_));
 sg13g2_nand3_1 _08808_ (.B(_02516_),
    .C(net110),
    .A(_02514_),
    .Y(_02637_));
 sg13g2_nor2_1 _08809_ (.A(_02423_),
    .B(_02637_),
    .Y(_02638_));
 sg13g2_a21oi_1 _08810_ (.A1(_02523_),
    .A2(_02526_),
    .Y(_02639_),
    .B1(_02638_));
 sg13g2_nand2_1 _08811_ (.Y(_02640_),
    .A(_02413_),
    .B(_02513_));
 sg13g2_nor3_1 _08812_ (.A(_02356_),
    .B(_02640_),
    .C(_02313_),
    .Y(_02642_));
 sg13g2_nand2_1 _08813_ (.Y(_02643_),
    .A(_02642_),
    .B(_02272_));
 sg13g2_inv_1 _08814_ (.Y(_02644_),
    .A(_02640_));
 sg13g2_o21ai_1 _08815_ (.B1(_02509_),
    .Y(_02645_),
    .A1(_02512_),
    .A2(_02496_));
 sg13g2_a21oi_1 _08816_ (.A1(_02393_),
    .A2(_02644_),
    .Y(_02646_),
    .B1(_02645_));
 sg13g2_nand2_1 _08817_ (.Y(_02647_),
    .A(_02643_),
    .B(_02646_));
 sg13g2_nand3_1 _08818_ (.B(_02193_),
    .C(net20),
    .A(_02300_),
    .Y(_02648_));
 sg13g2_xnor2_1 _08819_ (.Y(_02649_),
    .A(_02648_),
    .B(_02504_));
 sg13g2_nand2_1 _08820_ (.Y(_02650_),
    .A(_02647_),
    .B(_02649_));
 sg13g2_inv_1 _08821_ (.Y(_02651_),
    .A(_02649_));
 sg13g2_nand3_1 _08822_ (.B(_02646_),
    .C(_02651_),
    .A(_02643_),
    .Y(_02653_));
 sg13g2_buf_1 _08823_ (.A(_02653_),
    .X(_02654_));
 sg13g2_nand2_2 _08824_ (.Y(_02655_),
    .A(_02650_),
    .B(_02654_));
 sg13g2_nor2_1 _08825_ (.A(net92),
    .B(_02655_),
    .Y(_02656_));
 sg13g2_nand2_1 _08826_ (.Y(_02657_),
    .A(_02518_),
    .B(_02656_));
 sg13g2_nand3_1 _08827_ (.B(_02654_),
    .C(net73),
    .A(_02650_),
    .Y(_02658_));
 sg13g2_nand2_1 _08828_ (.Y(_02659_),
    .A(_02637_),
    .B(_02658_));
 sg13g2_nand2_1 _08829_ (.Y(_02660_),
    .A(_02657_),
    .B(_02659_));
 sg13g2_nor2_1 _08830_ (.A(net91),
    .B(_02418_),
    .Y(_02661_));
 sg13g2_nand2_1 _08831_ (.Y(_02662_),
    .A(_02660_),
    .B(_02661_));
 sg13g2_inv_1 _08832_ (.Y(_02664_),
    .A(_02661_));
 sg13g2_nand3_1 _08833_ (.B(_02659_),
    .C(_02664_),
    .A(_02657_),
    .Y(_02665_));
 sg13g2_nand2_1 _08834_ (.Y(_02666_),
    .A(_02662_),
    .B(_02665_));
 sg13g2_nand2b_1 _08835_ (.Y(_02667_),
    .B(_02666_),
    .A_N(_02639_));
 sg13g2_nand3_1 _08836_ (.B(_02639_),
    .C(_02665_),
    .A(_02662_),
    .Y(_02668_));
 sg13g2_nand2_1 _08837_ (.Y(_02669_),
    .A(_02667_),
    .B(_02668_));
 sg13g2_nor2_1 _08838_ (.A(_00198_),
    .B(_02376_),
    .Y(_02670_));
 sg13g2_inv_4 _08839_ (.A(_02525_),
    .Y(_02671_));
 sg13g2_nand2_1 _08840_ (.Y(_02672_),
    .A(_02671_),
    .B(net102));
 sg13g2_xnor2_1 _08841_ (.Y(_02673_),
    .A(_02538_),
    .B(_02672_));
 sg13g2_xor2_1 _08842_ (.B(_02673_),
    .A(_02670_),
    .X(_02675_));
 sg13g2_nand2_1 _08843_ (.Y(_02676_),
    .A(_02669_),
    .B(_02675_));
 sg13g2_inv_1 _08844_ (.Y(_02677_),
    .A(_02675_));
 sg13g2_nand3_1 _08845_ (.B(_02668_),
    .C(_02677_),
    .A(_02667_),
    .Y(_02678_));
 sg13g2_nand2_1 _08846_ (.Y(_02679_),
    .A(_02676_),
    .B(_02678_));
 sg13g2_nand2b_1 _08847_ (.Y(_02680_),
    .B(_02679_),
    .A_N(_02636_));
 sg13g2_nand3_1 _08848_ (.B(_02678_),
    .C(_02636_),
    .A(_02676_),
    .Y(_02681_));
 sg13g2_nand2_1 _08849_ (.Y(_02682_),
    .A(_02680_),
    .B(_02681_));
 sg13g2_inv_1 _08850_ (.Y(_02683_),
    .A(_02539_));
 sg13g2_a21oi_1 _08851_ (.A1(_02537_),
    .A2(_02535_),
    .Y(_02684_),
    .B1(_02683_));
 sg13g2_inv_1 _08852_ (.Y(_02686_),
    .A(_02684_));
 sg13g2_nand2_1 _08853_ (.Y(_02687_),
    .A(_02682_),
    .B(_02686_));
 sg13g2_nand3_1 _08854_ (.B(_02681_),
    .C(_02684_),
    .A(_02680_),
    .Y(_02688_));
 sg13g2_nand2_1 _08855_ (.Y(_02689_),
    .A(_02687_),
    .B(_02688_));
 sg13g2_nand2b_1 _08856_ (.Y(_02690_),
    .B(_02689_),
    .A_N(_02634_));
 sg13g2_nand3_1 _08857_ (.B(_02688_),
    .C(_02634_),
    .A(_02687_),
    .Y(_02691_));
 sg13g2_nand2_1 _08858_ (.Y(_02692_),
    .A(_02690_),
    .B(_02691_));
 sg13g2_nand2b_1 _08859_ (.Y(_02693_),
    .B(_02692_),
    .A_N(_02632_));
 sg13g2_nand3_1 _08860_ (.B(_02691_),
    .C(_02632_),
    .A(_02690_),
    .Y(_02694_));
 sg13g2_nand3_1 _08861_ (.B(_02693_),
    .C(_02694_),
    .A(_02631_),
    .Y(_02695_));
 sg13g2_buf_8 _08862_ (.A(_02695_),
    .X(_02697_));
 sg13g2_nand2_1 _08863_ (.Y(_02698_),
    .A(_02693_),
    .B(_02694_));
 sg13g2_nand2_1 _08864_ (.Y(_02699_),
    .A(_02698_),
    .B(_02629_));
 sg13g2_nand2_1 _08865_ (.Y(_02700_),
    .A(_02697_),
    .B(_02699_));
 sg13g2_nor2_1 _08866_ (.A(_02627_),
    .B(_02700_),
    .Y(_02701_));
 sg13g2_nand2_1 _08867_ (.Y(_02702_),
    .A(_02620_),
    .B(_02616_));
 sg13g2_nand2b_1 _08868_ (.Y(_02703_),
    .B(_02702_),
    .A_N(_02617_));
 sg13g2_nand3_1 _08869_ (.B(_02616_),
    .C(_02617_),
    .A(_02620_),
    .Y(_02704_));
 sg13g2_buf_1 _08870_ (.A(_02704_),
    .X(_02705_));
 sg13g2_nand2_1 _08871_ (.Y(_02706_),
    .A(_02703_),
    .B(_02705_));
 sg13g2_nand2_1 _08872_ (.Y(_02708_),
    .A(_02575_),
    .B(_02577_));
 sg13g2_nand2b_1 _08873_ (.Y(_02709_),
    .B(_02708_),
    .A_N(_02609_));
 sg13g2_nand2_1 _08874_ (.Y(_02710_),
    .A(_02709_),
    .B(_02610_));
 sg13g2_nand2_1 _08875_ (.Y(_02711_),
    .A(_02710_),
    .B(_02612_));
 sg13g2_nand3_1 _08876_ (.B(_02610_),
    .C(_02613_),
    .A(_02709_),
    .Y(_02712_));
 sg13g2_nand2_1 _08877_ (.Y(_02713_),
    .A(_02711_),
    .B(_02712_));
 sg13g2_nand2_1 _08878_ (.Y(_02714_),
    .A(_02591_),
    .B(_02606_));
 sg13g2_nand2b_1 _08879_ (.Y(_02715_),
    .B(_02714_),
    .A_N(_02604_));
 sg13g2_nand3_1 _08880_ (.B(_02606_),
    .C(_02604_),
    .A(_02591_),
    .Y(_02716_));
 sg13g2_nand2_1 _08881_ (.Y(_02717_),
    .A(_02715_),
    .B(_02716_));
 sg13g2_nand2_1 _08882_ (.Y(_02719_),
    .A(_02585_),
    .B(_02588_));
 sg13g2_nand2_1 _08883_ (.Y(_02720_),
    .A(_02719_),
    .B(_02587_));
 sg13g2_inv_1 _08884_ (.Y(_02721_),
    .A(_02587_));
 sg13g2_nand3_1 _08885_ (.B(_02588_),
    .C(_02721_),
    .A(_02585_),
    .Y(_02722_));
 sg13g2_nand2_1 _08886_ (.Y(_02723_),
    .A(_02471_),
    .B(net110));
 sg13g2_o21ai_1 _08887_ (.B1(_02723_),
    .Y(_02724_),
    .A1(net89),
    .A2(_02443_));
 sg13g2_nor2_1 _08888_ (.A(net76),
    .B(_02469_),
    .Y(_02725_));
 sg13g2_nor2_1 _08889_ (.A(net101),
    .B(_02440_),
    .Y(_02726_));
 sg13g2_inv_1 _08890_ (.Y(_02727_),
    .A(_02726_));
 sg13g2_nor2_1 _08891_ (.A(_02727_),
    .B(_02584_),
    .Y(_02728_));
 sg13g2_a21oi_1 _08892_ (.A1(_02724_),
    .A2(_02725_),
    .Y(_02730_),
    .B1(_02728_));
 sg13g2_nand3_1 _08893_ (.B(_02722_),
    .C(_02730_),
    .A(_02720_),
    .Y(_02731_));
 sg13g2_xnor2_1 _08894_ (.Y(_02732_),
    .A(_02103_),
    .B(net19));
 sg13g2_nand2_2 _08895_ (.Y(_02733_),
    .A(_02732_),
    .B(_01509_));
 sg13g2_nor2_1 _08896_ (.A(net88),
    .B(_02733_),
    .Y(_02734_));
 sg13g2_nor2_1 _08897_ (.A(net111),
    .B(_02595_),
    .Y(_02735_));
 sg13g2_nor2b_1 _08898_ (.A(_02601_),
    .B_N(_02735_),
    .Y(_02736_));
 sg13g2_buf_8 _08899_ (.A(net104),
    .X(_02737_));
 sg13g2_o21ai_1 _08900_ (.B1(_02598_),
    .Y(_02738_),
    .A1(net86),
    .A2(_02595_));
 sg13g2_nand2b_1 _08901_ (.Y(_02739_),
    .B(_02738_),
    .A_N(_02736_));
 sg13g2_xnor2_1 _08902_ (.Y(_02741_),
    .A(_02734_),
    .B(_02739_));
 sg13g2_a21oi_1 _08903_ (.A1(_02720_),
    .A2(_02722_),
    .Y(_02742_),
    .B1(_02730_));
 sg13g2_a21oi_1 _08904_ (.A1(_02731_),
    .A2(_02741_),
    .Y(_02743_),
    .B1(_02742_));
 sg13g2_nand2_1 _08905_ (.Y(_02744_),
    .A(_02717_),
    .B(_02743_));
 sg13g2_a21oi_1 _08906_ (.A1(_02738_),
    .A2(_02734_),
    .Y(_02745_),
    .B1(_02736_));
 sg13g2_inv_1 _08907_ (.Y(_02746_),
    .A(_02745_));
 sg13g2_nand3b_1 _08908_ (.B(_02715_),
    .C(_02716_),
    .Y(_02747_),
    .A_N(_02743_));
 sg13g2_inv_1 _08909_ (.Y(_02748_),
    .A(_02747_));
 sg13g2_a21oi_1 _08910_ (.A1(_02744_),
    .A2(_02746_),
    .Y(_02749_),
    .B1(_02748_));
 sg13g2_nand2_1 _08911_ (.Y(_02750_),
    .A(_02713_),
    .B(_02749_));
 sg13g2_nor2_1 _08912_ (.A(net87),
    .B(_02595_),
    .Y(_02752_));
 sg13g2_nor2_1 _08913_ (.A(_02749_),
    .B(_02713_),
    .Y(_02753_));
 sg13g2_a21oi_2 _08914_ (.B1(_02753_),
    .Y(_02754_),
    .A2(_02752_),
    .A1(_02750_));
 sg13g2_inv_4 _08915_ (.A(_02754_),
    .Y(_02755_));
 sg13g2_nand2_1 _08916_ (.Y(_02756_),
    .A(_02706_),
    .B(_02755_));
 sg13g2_nand3_1 _08917_ (.B(_02705_),
    .C(_02754_),
    .A(_02703_),
    .Y(_02757_));
 sg13g2_nand2_1 _08918_ (.Y(_02758_),
    .A(_02756_),
    .B(_02757_));
 sg13g2_nand2_1 _08919_ (.Y(_02759_),
    .A(_02747_),
    .B(_02744_));
 sg13g2_nand2_1 _08920_ (.Y(_02760_),
    .A(_02759_),
    .B(_02745_));
 sg13g2_nand3_1 _08921_ (.B(_02744_),
    .C(_02746_),
    .A(_02747_),
    .Y(_02761_));
 sg13g2_nand2_1 _08922_ (.Y(_02763_),
    .A(_02760_),
    .B(_02761_));
 sg13g2_inv_1 _08923_ (.Y(_02764_),
    .A(_02742_));
 sg13g2_nand2_1 _08924_ (.Y(_02765_),
    .A(_02764_),
    .B(_02731_));
 sg13g2_nand2b_1 _08925_ (.Y(_02766_),
    .B(_02765_),
    .A_N(_02741_));
 sg13g2_nand3_1 _08926_ (.B(_02731_),
    .C(_02741_),
    .A(_02764_),
    .Y(_02767_));
 sg13g2_nand2_1 _08927_ (.Y(_02768_),
    .A(_02766_),
    .B(_02767_));
 sg13g2_nand2b_1 _08928_ (.Y(_02769_),
    .B(_02724_),
    .A_N(_02728_));
 sg13g2_xor2_1 _08929_ (.B(_02769_),
    .A(_02725_),
    .X(_02770_));
 sg13g2_nor2_1 _08930_ (.A(_05485_),
    .B(_02469_),
    .Y(_02771_));
 sg13g2_nand2b_1 _08931_ (.Y(_02772_),
    .B(_02727_),
    .A_N(_02771_));
 sg13g2_nand2_1 _08932_ (.Y(_02774_),
    .A(_02726_),
    .B(_02771_));
 sg13g2_nor2_1 _08933_ (.A(_05493_),
    .B(_02595_),
    .Y(_02775_));
 sg13g2_nand3_1 _08934_ (.B(_02774_),
    .C(_02775_),
    .A(_02772_),
    .Y(_02776_));
 sg13g2_and2_1 _08935_ (.A(_02776_),
    .B(_02774_),
    .X(_02777_));
 sg13g2_nand2_1 _08936_ (.Y(_02778_),
    .A(_02770_),
    .B(_02777_));
 sg13g2_nor2_1 _08937_ (.A(net86),
    .B(_02733_),
    .Y(_02779_));
 sg13g2_nor2_1 _08938_ (.A(_02779_),
    .B(_02735_),
    .Y(_02780_));
 sg13g2_nand2_1 _08939_ (.Y(_02781_),
    .A(_02735_),
    .B(_02779_));
 sg13g2_inv_1 _08940_ (.Y(_02782_),
    .A(_02781_));
 sg13g2_buf_8 _08941_ (.A(_03651_),
    .X(_02783_));
 sg13g2_nand2_1 _08942_ (.Y(_02785_),
    .A(_02592_),
    .B(net100));
 sg13g2_o21ai_1 _08943_ (.B1(_02785_),
    .Y(_02786_),
    .A1(_02780_),
    .A2(_02782_));
 sg13g2_nor2_1 _08944_ (.A(_02777_),
    .B(_02770_),
    .Y(_02787_));
 sg13g2_a21oi_1 _08945_ (.A1(_02778_),
    .A2(_02786_),
    .Y(_02788_),
    .B1(_02787_));
 sg13g2_nand2_1 _08946_ (.Y(_02789_),
    .A(_02768_),
    .B(_02788_));
 sg13g2_nand3b_1 _08947_ (.B(_02766_),
    .C(_02767_),
    .Y(_02790_),
    .A_N(_02788_));
 sg13g2_inv_1 _08948_ (.Y(_02791_),
    .A(_02790_));
 sg13g2_a21oi_1 _08949_ (.A1(_02789_),
    .A2(_02782_),
    .Y(_02792_),
    .B1(_02791_));
 sg13g2_nand2_1 _08950_ (.Y(_02793_),
    .A(_02763_),
    .B(_02792_));
 sg13g2_nor2_1 _08951_ (.A(_02561_),
    .B(_02733_),
    .Y(_02794_));
 sg13g2_nand3b_1 _08952_ (.B(_02760_),
    .C(_02761_),
    .Y(_02796_),
    .A_N(_02792_));
 sg13g2_inv_1 _08953_ (.Y(_02797_),
    .A(_02796_));
 sg13g2_a21oi_1 _08954_ (.A1(_02793_),
    .A2(_02794_),
    .Y(_02798_),
    .B1(_02797_));
 sg13g2_nand3b_1 _08955_ (.B(_02711_),
    .C(_02712_),
    .Y(_02799_),
    .A_N(_02749_));
 sg13g2_nand2_1 _08956_ (.Y(_02800_),
    .A(_02799_),
    .B(_02750_));
 sg13g2_xor2_1 _08957_ (.B(_02800_),
    .A(_02752_),
    .X(_02801_));
 sg13g2_nor2_2 _08958_ (.A(_02798_),
    .B(_02801_),
    .Y(_02802_));
 sg13g2_nand2_1 _08959_ (.Y(_02803_),
    .A(_02758_),
    .B(_02802_));
 sg13g2_nand3_1 _08960_ (.B(_02703_),
    .C(_02705_),
    .A(_02755_),
    .Y(_02804_));
 sg13g2_buf_1 _08961_ (.A(_02804_),
    .X(_02805_));
 sg13g2_nand2_1 _08962_ (.Y(_02807_),
    .A(_02803_),
    .B(_02805_));
 sg13g2_nand2_1 _08963_ (.Y(_02808_),
    .A(_02701_),
    .B(_02807_));
 sg13g2_inv_1 _08964_ (.Y(_02809_),
    .A(_02699_));
 sg13g2_a21oi_1 _08965_ (.A1(_02697_),
    .A2(_02626_),
    .Y(_02810_),
    .B1(_02809_));
 sg13g2_inv_1 _08966_ (.Y(_02811_),
    .A(_02810_));
 sg13g2_nand2_1 _08967_ (.Y(_02812_),
    .A(_02808_),
    .B(_02811_));
 sg13g2_nand2_1 _08968_ (.Y(_02813_),
    .A(_02513_),
    .B(_02649_));
 sg13g2_nor3_1 _08969_ (.A(_02813_),
    .B(_02415_),
    .C(_02356_),
    .Y(_02814_));
 sg13g2_nand2_1 _08970_ (.Y(_02815_),
    .A(_02365_),
    .B(_02814_));
 sg13g2_inv_1 _08971_ (.Y(_02816_),
    .A(_02504_));
 sg13g2_a21oi_1 _08972_ (.A1(_02509_),
    .A2(_02816_),
    .Y(_02818_),
    .B1(_02648_));
 sg13g2_a21oi_2 _08973_ (.B1(_02813_),
    .Y(_02819_),
    .A2(_02496_),
    .A1(_02494_));
 sg13g2_nor2_1 _08974_ (.A(_02818_),
    .B(_02819_),
    .Y(_02820_));
 sg13g2_nand2_1 _08975_ (.Y(_02821_),
    .A(_02815_),
    .B(_02820_));
 sg13g2_nor2_1 _08976_ (.A(net18),
    .B(_02326_),
    .Y(_02822_));
 sg13g2_nor2_1 _08977_ (.A(_02822_),
    .B(_02503_),
    .Y(_02823_));
 sg13g2_nand2_1 _08978_ (.Y(_02824_),
    .A(_02821_),
    .B(_02823_));
 sg13g2_inv_1 _08979_ (.Y(_02825_),
    .A(_02823_));
 sg13g2_nand3_1 _08980_ (.B(_02825_),
    .C(_02820_),
    .A(_02815_),
    .Y(_02826_));
 sg13g2_nand2_2 _08981_ (.Y(_02827_),
    .A(_02824_),
    .B(_02826_));
 sg13g2_nand3_1 _08982_ (.B(_02656_),
    .C(net73),
    .A(_02827_),
    .Y(_02829_));
 sg13g2_nand3_1 _08983_ (.B(_02823_),
    .C(_02820_),
    .A(_02815_),
    .Y(_02830_));
 sg13g2_buf_1 _08984_ (.A(_02830_),
    .X(_02831_));
 sg13g2_nor2_1 _08985_ (.A(_02651_),
    .B(_02509_),
    .Y(_02832_));
 sg13g2_nor2_1 _08986_ (.A(_02832_),
    .B(_02819_),
    .Y(_02833_));
 sg13g2_nand3_1 _08987_ (.B(net73),
    .C(_02833_),
    .A(_02831_),
    .Y(_02834_));
 sg13g2_inv_2 _08988_ (.Y(_02835_),
    .A(_02656_));
 sg13g2_nand2_1 _08989_ (.Y(_02836_),
    .A(_02834_),
    .B(_02835_));
 sg13g2_nand2_1 _08990_ (.Y(_02837_),
    .A(_02829_),
    .B(_02836_));
 sg13g2_nor2_1 _08991_ (.A(net91),
    .B(_02517_),
    .Y(_02838_));
 sg13g2_nand2_1 _08992_ (.Y(_02840_),
    .A(_02837_),
    .B(_02838_));
 sg13g2_inv_1 _08993_ (.Y(_02841_),
    .A(_02838_));
 sg13g2_nand3_1 _08994_ (.B(_02836_),
    .C(_02841_),
    .A(_02829_),
    .Y(_02842_));
 sg13g2_inv_1 _08995_ (.Y(_02843_),
    .A(_02657_));
 sg13g2_a21oi_1 _08996_ (.A1(_02659_),
    .A2(_02661_),
    .Y(_02844_),
    .B1(_02843_));
 sg13g2_nand3_1 _08997_ (.B(_02842_),
    .C(_02844_),
    .A(_02840_),
    .Y(_02845_));
 sg13g2_buf_1 _08998_ (.A(_02845_),
    .X(_02846_));
 sg13g2_nor2_1 _08999_ (.A(net88),
    .B(_02316_),
    .Y(_02847_));
 sg13g2_nand3_1 _09000_ (.B(_02417_),
    .C(net102),
    .A(_02414_),
    .Y(_02848_));
 sg13g2_buf_1 _09001_ (.A(_02848_),
    .X(_02849_));
 sg13g2_nand2_1 _09002_ (.Y(_02851_),
    .A(_02671_),
    .B(_03432_));
 sg13g2_xnor2_1 _09003_ (.Y(_02852_),
    .A(_02849_),
    .B(_02851_));
 sg13g2_xnor2_1 _09004_ (.Y(_02853_),
    .A(_02847_),
    .B(_02852_));
 sg13g2_a21oi_1 _09005_ (.A1(_02840_),
    .A2(_02842_),
    .Y(_02854_),
    .B1(_02844_));
 sg13g2_a21oi_1 _09006_ (.A1(_02846_),
    .A2(_02853_),
    .Y(_02855_),
    .B1(_02854_));
 sg13g2_nor2_1 _09007_ (.A(net91),
    .B(_02655_),
    .Y(_02856_));
 sg13g2_inv_1 _09008_ (.Y(_02857_),
    .A(_02856_));
 sg13g2_nand3_1 _09009_ (.B(net110),
    .C(_02833_),
    .A(_02831_),
    .Y(_02858_));
 sg13g2_nor3_2 _09010_ (.A(_02404_),
    .B(_02832_),
    .C(_02819_),
    .Y(_02859_));
 sg13g2_inv_1 _09011_ (.Y(_02860_),
    .A(_02859_));
 sg13g2_nand2_1 _09012_ (.Y(_02862_),
    .A(_02860_),
    .B(net73));
 sg13g2_nand2_1 _09013_ (.Y(_02863_),
    .A(_02858_),
    .B(_02862_));
 sg13g2_nor2_2 _09014_ (.A(net92),
    .B(_02859_),
    .Y(_02864_));
 sg13g2_nand4_1 _09015_ (.B(net73),
    .C(_02833_),
    .A(_02831_),
    .Y(_02865_),
    .D(_02864_));
 sg13g2_nand2_1 _09016_ (.Y(_02866_),
    .A(_02863_),
    .B(_02865_));
 sg13g2_xnor2_1 _09017_ (.Y(_02867_),
    .A(_02857_),
    .B(_02866_));
 sg13g2_inv_2 _09018_ (.Y(_02868_),
    .A(_02829_));
 sg13g2_a21oi_1 _09019_ (.A1(_02836_),
    .A2(_02838_),
    .Y(_02869_),
    .B1(_02868_));
 sg13g2_nand2_1 _09020_ (.Y(_02870_),
    .A(_02867_),
    .B(_02869_));
 sg13g2_nand2_1 _09021_ (.Y(_02871_),
    .A(_02866_),
    .B(_02856_));
 sg13g2_nand3_1 _09022_ (.B(_02865_),
    .C(_02857_),
    .A(_02863_),
    .Y(_02872_));
 sg13g2_nand2_1 _09023_ (.Y(_02873_),
    .A(_02871_),
    .B(_02872_));
 sg13g2_nand2b_1 _09024_ (.Y(_02874_),
    .B(_02873_),
    .A_N(_02869_));
 sg13g2_nand2_1 _09025_ (.Y(_02875_),
    .A(_02870_),
    .B(_02874_));
 sg13g2_nor2_1 _09026_ (.A(_00198_),
    .B(_02525_),
    .Y(_02876_));
 sg13g2_nand3_1 _09027_ (.B(_02516_),
    .C(_03432_),
    .A(_02514_),
    .Y(_02877_));
 sg13g2_nor2_1 _09028_ (.A(_02849_),
    .B(_02877_),
    .Y(_02878_));
 sg13g2_inv_1 _09029_ (.Y(_02879_),
    .A(_02418_));
 sg13g2_nor2_1 _09030_ (.A(net111),
    .B(_02517_),
    .Y(_02880_));
 sg13g2_a21oi_1 _09031_ (.A1(net106),
    .A2(_02879_),
    .Y(_02881_),
    .B1(_02880_));
 sg13g2_nor2_1 _09032_ (.A(_02878_),
    .B(_02881_),
    .Y(_02883_));
 sg13g2_xnor2_1 _09033_ (.Y(_02884_),
    .A(_02876_),
    .B(_02883_));
 sg13g2_inv_1 _09034_ (.Y(_02885_),
    .A(_02884_));
 sg13g2_nand2_1 _09035_ (.Y(_02886_),
    .A(_02875_),
    .B(_02885_));
 sg13g2_nand3_1 _09036_ (.B(_02874_),
    .C(_02884_),
    .A(_02870_),
    .Y(_02887_));
 sg13g2_nand2_1 _09037_ (.Y(_02888_),
    .A(_02886_),
    .B(_02887_));
 sg13g2_nand2b_1 _09038_ (.Y(_02889_),
    .B(_02888_),
    .A_N(_02855_));
 sg13g2_nand3_1 _09039_ (.B(_02887_),
    .C(_02855_),
    .A(_02886_),
    .Y(_02890_));
 sg13g2_nand2_1 _09040_ (.Y(_02891_),
    .A(_02889_),
    .B(_02890_));
 sg13g2_nor2_1 _09041_ (.A(_02849_),
    .B(_02851_),
    .Y(_02892_));
 sg13g2_nand2b_1 _09042_ (.Y(_02894_),
    .B(_02847_),
    .A_N(_02852_));
 sg13g2_nor2b_1 _09043_ (.A(_02892_),
    .B_N(_02894_),
    .Y(_02895_));
 sg13g2_inv_1 _09044_ (.Y(_02896_),
    .A(_02895_));
 sg13g2_nand2_1 _09045_ (.Y(_02897_),
    .A(_02891_),
    .B(_02896_));
 sg13g2_nand3_1 _09046_ (.B(_02890_),
    .C(_02895_),
    .A(_02889_),
    .Y(_02898_));
 sg13g2_nand2_1 _09047_ (.Y(_02899_),
    .A(_02840_),
    .B(_02842_));
 sg13g2_nand2b_1 _09048_ (.Y(_02900_),
    .B(_02899_),
    .A_N(_02844_));
 sg13g2_nand2_1 _09049_ (.Y(_02901_),
    .A(_02900_),
    .B(_02846_));
 sg13g2_nand2_1 _09050_ (.Y(_02902_),
    .A(_02901_),
    .B(_02853_));
 sg13g2_inv_1 _09051_ (.Y(_02903_),
    .A(_02853_));
 sg13g2_nand3_1 _09052_ (.B(_02846_),
    .C(_02903_),
    .A(_02900_),
    .Y(_02905_));
 sg13g2_a21oi_1 _09053_ (.A1(_02662_),
    .A2(_02665_),
    .Y(_02906_),
    .B1(_02639_));
 sg13g2_a21oi_1 _09054_ (.A1(_02668_),
    .A2(_02675_),
    .Y(_02907_),
    .B1(_02906_));
 sg13g2_nand3_1 _09055_ (.B(_02905_),
    .C(_02907_),
    .A(_02902_),
    .Y(_02908_));
 sg13g2_nor2b_1 _09056_ (.A(_02672_),
    .B_N(_02538_),
    .Y(_02909_));
 sg13g2_a21oi_1 _09057_ (.A1(_02673_),
    .A2(_02670_),
    .Y(_02910_),
    .B1(_02909_));
 sg13g2_inv_1 _09058_ (.Y(_02911_),
    .A(_02910_));
 sg13g2_nand2_1 _09059_ (.Y(_02912_),
    .A(_02901_),
    .B(_02903_));
 sg13g2_nand3_1 _09060_ (.B(_02846_),
    .C(_02853_),
    .A(_02900_),
    .Y(_02913_));
 sg13g2_inv_1 _09061_ (.Y(_02914_),
    .A(_02907_));
 sg13g2_nand3_1 _09062_ (.B(_02913_),
    .C(_02914_),
    .A(_02912_),
    .Y(_02916_));
 sg13g2_inv_1 _09063_ (.Y(_02917_),
    .A(_02916_));
 sg13g2_a21oi_1 _09064_ (.A1(_02908_),
    .A2(_02911_),
    .Y(_02918_),
    .B1(_02917_));
 sg13g2_nand3_1 _09065_ (.B(_02898_),
    .C(_02918_),
    .A(_02897_),
    .Y(_02919_));
 sg13g2_nor2_1 _09066_ (.A(_02561_),
    .B(_02316_),
    .Y(_02920_));
 sg13g2_nand2_1 _09067_ (.Y(_02921_),
    .A(_02897_),
    .B(_02898_));
 sg13g2_nand2b_1 _09068_ (.Y(_02922_),
    .B(_02921_),
    .A_N(_02918_));
 sg13g2_inv_1 _09069_ (.Y(_02923_),
    .A(_02922_));
 sg13g2_a21oi_2 _09070_ (.B1(_02923_),
    .Y(_02924_),
    .A2(_02920_),
    .A1(_02919_));
 sg13g2_inv_4 _09071_ (.A(_02924_),
    .Y(_02925_));
 sg13g2_nor2_2 _09072_ (.A(net87),
    .B(_02525_),
    .Y(_02927_));
 sg13g2_inv_1 _09073_ (.Y(_02928_),
    .A(_02889_));
 sg13g2_a21oi_1 _09074_ (.A1(_02890_),
    .A2(_02896_),
    .Y(_02929_),
    .B1(_02928_));
 sg13g2_inv_1 _09075_ (.Y(_02930_),
    .A(_02874_));
 sg13g2_a21oi_1 _09076_ (.A1(_02870_),
    .A2(_02885_),
    .Y(_02931_),
    .B1(_02930_));
 sg13g2_nor2_1 _09077_ (.A(_00198_),
    .B(_02418_),
    .Y(_02932_));
 sg13g2_nor2_1 _09078_ (.A(net104),
    .B(_02655_),
    .Y(_02933_));
 sg13g2_nand2_1 _09079_ (.Y(_02934_),
    .A(_02880_),
    .B(_02933_));
 sg13g2_nand3_1 _09080_ (.B(_02654_),
    .C(net102),
    .A(_02650_),
    .Y(_02935_));
 sg13g2_nand2_1 _09081_ (.Y(_02936_),
    .A(_02877_),
    .B(_02935_));
 sg13g2_nand2_1 _09082_ (.Y(_02938_),
    .A(_02934_),
    .B(_02936_));
 sg13g2_xnor2_1 _09083_ (.Y(_02939_),
    .A(_02932_),
    .B(_02938_));
 sg13g2_nand2_1 _09084_ (.Y(_02940_),
    .A(_02831_),
    .B(_02833_));
 sg13g2_nor2_1 _09085_ (.A(net91),
    .B(_02940_),
    .Y(_02941_));
 sg13g2_xnor2_1 _09086_ (.Y(_02942_),
    .A(_02864_),
    .B(_02941_));
 sg13g2_inv_1 _09087_ (.Y(_02943_),
    .A(_02865_));
 sg13g2_a21oi_1 _09088_ (.A1(_02863_),
    .A2(_02856_),
    .Y(_02944_),
    .B1(_02943_));
 sg13g2_nor2_1 _09089_ (.A(_02942_),
    .B(_02944_),
    .Y(_02945_));
 sg13g2_inv_2 _09090_ (.Y(_02946_),
    .A(_02945_));
 sg13g2_nand2_1 _09091_ (.Y(_02947_),
    .A(_02944_),
    .B(_02942_));
 sg13g2_nand2_1 _09092_ (.Y(_02949_),
    .A(_02946_),
    .B(_02947_));
 sg13g2_xnor2_1 _09093_ (.Y(_02950_),
    .A(_02939_),
    .B(_02949_));
 sg13g2_nand2b_1 _09094_ (.Y(_02951_),
    .B(_02950_),
    .A_N(_02931_));
 sg13g2_nand2b_1 _09095_ (.Y(_02952_),
    .B(_02949_),
    .A_N(_02939_));
 sg13g2_nand3_1 _09096_ (.B(_02947_),
    .C(_02939_),
    .A(_02946_),
    .Y(_02953_));
 sg13g2_nand2_1 _09097_ (.Y(_02954_),
    .A(_02952_),
    .B(_02953_));
 sg13g2_nand2_2 _09098_ (.Y(_02955_),
    .A(_02954_),
    .B(_02931_));
 sg13g2_nand2_1 _09099_ (.Y(_02956_),
    .A(_02951_),
    .B(_02955_));
 sg13g2_a21oi_2 _09100_ (.B1(_02878_),
    .Y(_02957_),
    .A2(_02876_),
    .A1(_02883_));
 sg13g2_inv_2 _09101_ (.Y(_02958_),
    .A(_02957_));
 sg13g2_nand2_1 _09102_ (.Y(_02960_),
    .A(_02956_),
    .B(_02958_));
 sg13g2_nand3_1 _09103_ (.B(_02955_),
    .C(_02957_),
    .A(_02951_),
    .Y(_02961_));
 sg13g2_nand2_1 _09104_ (.Y(_02962_),
    .A(_02960_),
    .B(_02961_));
 sg13g2_nand2b_1 _09105_ (.Y(_02963_),
    .B(_02962_),
    .A_N(_02929_));
 sg13g2_nand2_1 _09106_ (.Y(_02964_),
    .A(_02956_),
    .B(_02957_));
 sg13g2_nand3_1 _09107_ (.B(_02955_),
    .C(_02958_),
    .A(_02951_),
    .Y(_02965_));
 sg13g2_nand2_1 _09108_ (.Y(_02966_),
    .A(_02964_),
    .B(_02965_));
 sg13g2_nand2_1 _09109_ (.Y(_02967_),
    .A(_02966_),
    .B(_02929_));
 sg13g2_nand2_1 _09110_ (.Y(_02968_),
    .A(_02963_),
    .B(_02967_));
 sg13g2_nand2b_1 _09111_ (.Y(_02969_),
    .B(_02968_),
    .A_N(_02927_));
 sg13g2_nand3_1 _09112_ (.B(_02967_),
    .C(_02927_),
    .A(_02963_),
    .Y(_02971_));
 sg13g2_nand2_1 _09113_ (.Y(_02972_),
    .A(_02969_),
    .B(_02971_));
 sg13g2_xnor2_1 _09114_ (.Y(_02973_),
    .A(_02925_),
    .B(_02972_));
 sg13g2_inv_2 _09115_ (.Y(_02974_),
    .A(_02963_));
 sg13g2_a21oi_1 _09116_ (.A1(_02967_),
    .A2(_02927_),
    .Y(_02975_),
    .B1(_02974_));
 sg13g2_nor2_1 _09117_ (.A(_02562_),
    .B(_02418_),
    .Y(_02976_));
 sg13g2_nor2_1 _09118_ (.A(_02931_),
    .B(_02954_),
    .Y(_02977_));
 sg13g2_a21oi_2 _09119_ (.B1(_02977_),
    .Y(_02978_),
    .A2(_02958_),
    .A1(_02955_));
 sg13g2_a21oi_1 _09120_ (.A1(_02947_),
    .A2(_02939_),
    .Y(_02979_),
    .B1(_02945_));
 sg13g2_nand2_1 _09121_ (.Y(_02980_),
    .A(_02941_),
    .B(_02864_));
 sg13g2_inv_2 _09122_ (.Y(_02982_),
    .A(_05568_));
 sg13g2_nand2_1 _09123_ (.Y(_02983_),
    .A(_02860_),
    .B(_02982_));
 sg13g2_nand2_1 _09124_ (.Y(_02984_),
    .A(_02980_),
    .B(_02983_));
 sg13g2_nand3_1 _09125_ (.B(_02982_),
    .C(_02864_),
    .A(_02941_),
    .Y(_02985_));
 sg13g2_buf_1 _09126_ (.A(_02985_),
    .X(_02986_));
 sg13g2_nand2_1 _09127_ (.Y(_02987_),
    .A(_02984_),
    .B(_02986_));
 sg13g2_nand2_1 _09128_ (.Y(_02988_),
    .A(_02827_),
    .B(_03542_));
 sg13g2_nand2b_1 _09129_ (.Y(_02989_),
    .B(_02988_),
    .A_N(_02933_));
 sg13g2_nand3_1 _09130_ (.B(_02933_),
    .C(_03542_),
    .A(_02827_),
    .Y(_02990_));
 sg13g2_buf_1 _09131_ (.A(_02990_),
    .X(_02991_));
 sg13g2_nand2_1 _09132_ (.Y(_02993_),
    .A(_02989_),
    .B(_02991_));
 sg13g2_nor2_1 _09133_ (.A(_00198_),
    .B(_02517_),
    .Y(_02994_));
 sg13g2_nand2_1 _09134_ (.Y(_02995_),
    .A(_02993_),
    .B(_02994_));
 sg13g2_inv_1 _09135_ (.Y(_02996_),
    .A(_02994_));
 sg13g2_nand3_1 _09136_ (.B(_02991_),
    .C(_02996_),
    .A(_02989_),
    .Y(_02997_));
 sg13g2_nand2_1 _09137_ (.Y(_02998_),
    .A(_02995_),
    .B(_02997_));
 sg13g2_xnor2_1 _09138_ (.Y(_02999_),
    .A(_02987_),
    .B(_02998_));
 sg13g2_nand2b_1 _09139_ (.Y(_03000_),
    .B(_02999_),
    .A_N(_02979_));
 sg13g2_xor2_1 _09140_ (.B(_02998_),
    .A(_02987_),
    .X(_03001_));
 sg13g2_nand2_1 _09141_ (.Y(_03002_),
    .A(_03001_),
    .B(_02979_));
 sg13g2_nand2_1 _09142_ (.Y(_03004_),
    .A(_03000_),
    .B(_03002_));
 sg13g2_inv_1 _09143_ (.Y(_03005_),
    .A(_02934_));
 sg13g2_nor2b_1 _09144_ (.A(_02938_),
    .B_N(_02932_),
    .Y(_03006_));
 sg13g2_nor2_1 _09145_ (.A(_03005_),
    .B(_03006_),
    .Y(_03007_));
 sg13g2_nand2_1 _09146_ (.Y(_03008_),
    .A(_03004_),
    .B(_03007_));
 sg13g2_inv_1 _09147_ (.Y(_03009_),
    .A(_03007_));
 sg13g2_nand3_1 _09148_ (.B(_03002_),
    .C(_03009_),
    .A(_03000_),
    .Y(_03010_));
 sg13g2_nand2_1 _09149_ (.Y(_03011_),
    .A(_03008_),
    .B(_03010_));
 sg13g2_xnor2_1 _09150_ (.Y(_03012_),
    .A(_02978_),
    .B(_03011_));
 sg13g2_xnor2_1 _09151_ (.Y(_03013_),
    .A(_02976_),
    .B(_03012_));
 sg13g2_xnor2_1 _09152_ (.Y(_03015_),
    .A(_02975_),
    .B(_03013_));
 sg13g2_nand2_1 _09153_ (.Y(_03016_),
    .A(_02973_),
    .B(_03015_));
 sg13g2_nand2_1 _09154_ (.Y(_03017_),
    .A(_02908_),
    .B(_02916_));
 sg13g2_nand2_1 _09155_ (.Y(_03018_),
    .A(_03017_),
    .B(_02911_));
 sg13g2_nand3_1 _09156_ (.B(_02916_),
    .C(_02910_),
    .A(_02908_),
    .Y(_03019_));
 sg13g2_inv_1 _09157_ (.Y(_03020_),
    .A(_02680_));
 sg13g2_a21oi_1 _09158_ (.A1(_02681_),
    .A2(_02686_),
    .Y(_03021_),
    .B1(_03020_));
 sg13g2_nand3_1 _09159_ (.B(_03019_),
    .C(_03021_),
    .A(_03018_),
    .Y(_03022_));
 sg13g2_buf_2 _09160_ (.A(_03022_),
    .X(_03023_));
 sg13g2_nor2_2 _09161_ (.A(net87),
    .B(_02376_),
    .Y(_03024_));
 sg13g2_nand2_1 _09162_ (.Y(_03026_),
    .A(_03018_),
    .B(_03019_));
 sg13g2_nand2b_1 _09163_ (.Y(_03027_),
    .B(_03026_),
    .A_N(_03021_));
 sg13g2_inv_2 _09164_ (.Y(_03028_),
    .A(_03027_));
 sg13g2_a21oi_2 _09165_ (.B1(_03028_),
    .Y(_03029_),
    .A2(_03024_),
    .A1(_03023_));
 sg13g2_inv_2 _09166_ (.Y(_03030_),
    .A(_03029_));
 sg13g2_nand2_1 _09167_ (.Y(_03031_),
    .A(_02922_),
    .B(_02919_));
 sg13g2_nand2b_1 _09168_ (.Y(_03032_),
    .B(_03031_),
    .A_N(_02920_));
 sg13g2_nand3_1 _09169_ (.B(_02919_),
    .C(_02920_),
    .A(_02922_),
    .Y(_03033_));
 sg13g2_nand2_1 _09170_ (.Y(_03034_),
    .A(_03032_),
    .B(_03033_));
 sg13g2_xnor2_1 _09171_ (.Y(_03035_),
    .A(_03030_),
    .B(_03034_));
 sg13g2_a21oi_1 _09172_ (.A1(_02687_),
    .A2(_02688_),
    .Y(_03037_),
    .B1(_02634_));
 sg13g2_a21oi_1 _09173_ (.A1(_02691_),
    .A2(_02632_),
    .Y(_03038_),
    .B1(_03037_));
 sg13g2_nand2_1 _09174_ (.Y(_03039_),
    .A(_03027_),
    .B(_03023_));
 sg13g2_inv_1 _09175_ (.Y(_03040_),
    .A(_03024_));
 sg13g2_nand2_1 _09176_ (.Y(_03041_),
    .A(_03039_),
    .B(_03040_));
 sg13g2_nand3_1 _09177_ (.B(_03023_),
    .C(_03024_),
    .A(_03027_),
    .Y(_03042_));
 sg13g2_nand2_1 _09178_ (.Y(_03043_),
    .A(_03041_),
    .B(_03042_));
 sg13g2_nor2_1 _09179_ (.A(_03038_),
    .B(_03043_),
    .Y(_03044_));
 sg13g2_nand2_1 _09180_ (.Y(_03045_),
    .A(_03039_),
    .B(_03024_));
 sg13g2_nand3_1 _09181_ (.B(_03023_),
    .C(_03040_),
    .A(_03027_),
    .Y(_03046_));
 sg13g2_nand3_1 _09182_ (.B(_03046_),
    .C(_03038_),
    .A(_03045_),
    .Y(_03048_));
 sg13g2_inv_2 _09183_ (.Y(_03049_),
    .A(_03048_));
 sg13g2_nor2_1 _09184_ (.A(_03044_),
    .B(_03049_),
    .Y(_03050_));
 sg13g2_nand2_1 _09185_ (.Y(_03051_),
    .A(_03035_),
    .B(_03050_));
 sg13g2_nor2_1 _09186_ (.A(_03016_),
    .B(_03051_),
    .Y(_03052_));
 sg13g2_nand2_1 _09187_ (.Y(_03053_),
    .A(_03034_),
    .B(_03029_));
 sg13g2_nand2_1 _09188_ (.Y(_03054_),
    .A(_03053_),
    .B(_03044_));
 sg13g2_nand3_1 _09189_ (.B(_03032_),
    .C(_03033_),
    .A(_03030_),
    .Y(_03055_));
 sg13g2_nand2_1 _09190_ (.Y(_03056_),
    .A(_03054_),
    .B(_03055_));
 sg13g2_xnor2_1 _09191_ (.Y(_03057_),
    .A(_02927_),
    .B(_02968_));
 sg13g2_nand2_1 _09192_ (.Y(_03059_),
    .A(_03057_),
    .B(_02925_));
 sg13g2_nand2_1 _09193_ (.Y(_03060_),
    .A(_02972_),
    .B(_02924_));
 sg13g2_nand2_1 _09194_ (.Y(_03061_),
    .A(_03059_),
    .B(_03060_));
 sg13g2_nor2b_1 _09195_ (.A(_03061_),
    .B_N(_03015_),
    .Y(_03062_));
 sg13g2_nand2_1 _09196_ (.Y(_03063_),
    .A(_03056_),
    .B(_03062_));
 sg13g2_nor2_1 _09197_ (.A(_02924_),
    .B(_02972_),
    .Y(_03064_));
 sg13g2_nand2b_1 _09198_ (.Y(_03065_),
    .B(_03013_),
    .A_N(_02975_));
 sg13g2_inv_1 _09199_ (.Y(_03066_),
    .A(_03065_));
 sg13g2_a21oi_1 _09200_ (.A1(_03015_),
    .A2(_03064_),
    .Y(_03067_),
    .B1(_03066_));
 sg13g2_nand2_1 _09201_ (.Y(_03068_),
    .A(_03063_),
    .B(_03067_));
 sg13g2_a21oi_1 _09202_ (.A1(_02812_),
    .A2(_03052_),
    .Y(_03070_),
    .B1(_03068_));
 sg13g2_nand2_1 _09203_ (.Y(_03071_),
    .A(_02801_),
    .B(_02798_));
 sg13g2_nor2b_1 _09204_ (.A(_02802_),
    .B_N(_03071_),
    .Y(_03072_));
 sg13g2_nand2_1 _09205_ (.Y(_03073_),
    .A(_03072_),
    .B(_02758_));
 sg13g2_nor2b_1 _09206_ (.A(_03073_),
    .B_N(_02701_),
    .Y(_03074_));
 sg13g2_nand2_1 _09207_ (.Y(_03075_),
    .A(_02796_),
    .B(_02793_));
 sg13g2_nand2b_1 _09208_ (.Y(_03076_),
    .B(_03075_),
    .A_N(_02794_));
 sg13g2_nor2_1 _09209_ (.A(net89),
    .B(_02469_),
    .Y(_03077_));
 sg13g2_nor2_2 _09210_ (.A(_05485_),
    .B(_02595_),
    .Y(_03078_));
 sg13g2_xnor2_1 _09211_ (.Y(_03079_),
    .A(_03078_),
    .B(_03077_));
 sg13g2_nor2_1 _09212_ (.A(_05494_),
    .B(_02733_),
    .Y(_03081_));
 sg13g2_nor2b_1 _09213_ (.A(_03079_),
    .B_N(_03081_),
    .Y(_03082_));
 sg13g2_a21oi_1 _09214_ (.A1(_03077_),
    .A2(_03078_),
    .Y(_03083_),
    .B1(_03082_));
 sg13g2_nand2_1 _09215_ (.Y(_03084_),
    .A(_02772_),
    .B(_02774_));
 sg13g2_nand2b_1 _09216_ (.Y(_03085_),
    .B(_03084_),
    .A_N(_02775_));
 sg13g2_nand2_1 _09217_ (.Y(_03086_),
    .A(_03085_),
    .B(_02776_));
 sg13g2_inv_1 _09218_ (.Y(_03087_),
    .A(_03086_));
 sg13g2_nand2b_1 _09219_ (.Y(_03088_),
    .B(_03087_),
    .A_N(_03083_));
 sg13g2_nand2_1 _09220_ (.Y(_03089_),
    .A(_03086_),
    .B(_03083_));
 sg13g2_nand2_1 _09221_ (.Y(_03090_),
    .A(_03088_),
    .B(_03089_));
 sg13g2_inv_1 _09222_ (.Y(_03092_),
    .A(_03090_));
 sg13g2_inv_1 _09223_ (.Y(_03093_),
    .A(_02733_));
 sg13g2_a22oi_1 _09224_ (.Y(_03094_),
    .B1(net102),
    .B2(_03093_),
    .A2(_02592_),
    .A1(net106));
 sg13g2_inv_1 _09225_ (.Y(_03095_),
    .A(_03094_));
 sg13g2_nand2_1 _09226_ (.Y(_03096_),
    .A(_03092_),
    .B(_03095_));
 sg13g2_and2_1 _09227_ (.A(_03096_),
    .B(_03088_),
    .X(_03097_));
 sg13g2_nor2b_1 _09228_ (.A(_02787_),
    .B_N(_02778_),
    .Y(_03098_));
 sg13g2_xnor2_1 _09229_ (.Y(_03099_),
    .A(_02786_),
    .B(_03098_));
 sg13g2_nor2_1 _09230_ (.A(_03097_),
    .B(_03099_),
    .Y(_03100_));
 sg13g2_nand2_1 _09231_ (.Y(_03101_),
    .A(_02790_),
    .B(_02789_));
 sg13g2_nand2_1 _09232_ (.Y(_03103_),
    .A(_03101_),
    .B(_02781_));
 sg13g2_nand3_1 _09233_ (.B(_02789_),
    .C(_02782_),
    .A(_02790_),
    .Y(_03104_));
 sg13g2_nand2_1 _09234_ (.Y(_03105_),
    .A(_03103_),
    .B(_03104_));
 sg13g2_nand2b_1 _09235_ (.Y(_03106_),
    .B(_03105_),
    .A_N(_03100_));
 sg13g2_inv_1 _09236_ (.Y(_03107_),
    .A(_02592_));
 sg13g2_nor2_1 _09237_ (.A(_02561_),
    .B(_03107_),
    .Y(_03108_));
 sg13g2_nand3_1 _09238_ (.B(_03104_),
    .C(_03100_),
    .A(_03103_),
    .Y(_03109_));
 sg13g2_inv_1 _09239_ (.Y(_03110_),
    .A(_03109_));
 sg13g2_a21oi_1 _09240_ (.A1(_03106_),
    .A2(_03108_),
    .Y(_03111_),
    .B1(_03110_));
 sg13g2_inv_1 _09241_ (.Y(_03112_),
    .A(_03111_));
 sg13g2_nand3_1 _09242_ (.B(_02793_),
    .C(_02794_),
    .A(_02796_),
    .Y(_03114_));
 sg13g2_nand3_1 _09243_ (.B(_03112_),
    .C(_03114_),
    .A(_03076_),
    .Y(_03115_));
 sg13g2_nor2_1 _09244_ (.A(_02561_),
    .B(_01510_),
    .Y(_03116_));
 sg13g2_nor2_1 _09245_ (.A(net89),
    .B(_02595_),
    .Y(_03117_));
 sg13g2_a21o_1 _09246_ (.A2(_03093_),
    .A1(net110),
    .B1(_03117_),
    .X(_03118_));
 sg13g2_nor2_1 _09247_ (.A(net89),
    .B(_02733_),
    .Y(_03119_));
 sg13g2_nand2_2 _09248_ (.Y(_03120_),
    .A(_03078_),
    .B(_03119_));
 sg13g2_nand2_1 _09249_ (.Y(_03121_),
    .A(_03118_),
    .B(_03120_));
 sg13g2_o21ai_1 _09250_ (.B1(_03121_),
    .Y(_03122_),
    .A1(net76),
    .A2(_03107_));
 sg13g2_nor2_1 _09251_ (.A(net86),
    .B(_01510_),
    .Y(_03123_));
 sg13g2_nand2_1 _09252_ (.Y(_03125_),
    .A(_03122_),
    .B(_03123_));
 sg13g2_nand2_1 _09253_ (.Y(_03126_),
    .A(_02592_),
    .B(net102));
 sg13g2_o21ai_1 _09254_ (.B1(_03126_),
    .Y(_03127_),
    .A1(net88),
    .A2(_01510_));
 sg13g2_xor2_1 _09255_ (.B(_03079_),
    .A(_03081_),
    .X(_03128_));
 sg13g2_xnor2_1 _09256_ (.Y(_03129_),
    .A(_03120_),
    .B(_03128_));
 sg13g2_xor2_1 _09257_ (.B(_03129_),
    .A(_03127_),
    .X(_03130_));
 sg13g2_nor2_1 _09258_ (.A(_03125_),
    .B(_03130_),
    .Y(_03131_));
 sg13g2_nand2_1 _09259_ (.Y(_03132_),
    .A(_03128_),
    .B(_03120_));
 sg13g2_nor2_1 _09260_ (.A(_03120_),
    .B(_03128_),
    .Y(_03133_));
 sg13g2_a21oi_1 _09261_ (.A1(_03132_),
    .A2(_03127_),
    .Y(_03134_),
    .B1(_03133_));
 sg13g2_nand2_1 _09262_ (.Y(_03136_),
    .A(_03090_),
    .B(_03094_));
 sg13g2_nand3b_1 _09263_ (.B(_03096_),
    .C(_03136_),
    .Y(_03137_),
    .A_N(_03134_));
 sg13g2_buf_1 _09264_ (.A(_03137_),
    .X(_03138_));
 sg13g2_nand2_1 _09265_ (.Y(_03139_),
    .A(_03096_),
    .B(_03136_));
 sg13g2_nand2_1 _09266_ (.Y(_03140_),
    .A(_03139_),
    .B(_03134_));
 sg13g2_nand2_1 _09267_ (.Y(_03141_),
    .A(_03138_),
    .B(_03140_));
 sg13g2_nand2b_1 _09268_ (.Y(_03142_),
    .B(_03141_),
    .A_N(_03131_));
 sg13g2_nand3_1 _09269_ (.B(_03140_),
    .C(_03131_),
    .A(_03138_),
    .Y(_03143_));
 sg13g2_nand2_1 _09270_ (.Y(_03144_),
    .A(_03142_),
    .B(_03143_));
 sg13g2_nand2b_1 _09271_ (.Y(_03145_),
    .B(_03144_),
    .A_N(_03116_));
 sg13g2_inv_1 _09272_ (.Y(_03147_),
    .A(_03125_));
 sg13g2_nor2_1 _09273_ (.A(_03123_),
    .B(_03122_),
    .Y(_03148_));
 sg13g2_nand3_1 _09274_ (.B(net93),
    .C(_01509_),
    .A(_03119_),
    .Y(_03149_));
 sg13g2_nor4_1 _09275_ (.A(_03147_),
    .B(_03148_),
    .C(_03149_),
    .D(_03130_),
    .Y(_03150_));
 sg13g2_nand2_1 _09276_ (.Y(_03151_),
    .A(_03145_),
    .B(_03150_));
 sg13g2_inv_1 _09277_ (.Y(_03152_),
    .A(_03143_));
 sg13g2_a21oi_1 _09278_ (.A1(_03142_),
    .A2(_03116_),
    .Y(_03153_),
    .B1(_03152_));
 sg13g2_nand2_1 _09279_ (.Y(_03154_),
    .A(_03151_),
    .B(_03153_));
 sg13g2_xnor2_1 _09280_ (.Y(_03155_),
    .A(_03097_),
    .B(_03099_));
 sg13g2_nand2_1 _09281_ (.Y(_03156_),
    .A(_03155_),
    .B(_03138_));
 sg13g2_nand2_1 _09282_ (.Y(_03158_),
    .A(_03154_),
    .B(_03156_));
 sg13g2_nor2_1 _09283_ (.A(_03138_),
    .B(_03155_),
    .Y(_03159_));
 sg13g2_inv_1 _09284_ (.Y(_03160_),
    .A(_03159_));
 sg13g2_nand2_1 _09285_ (.Y(_03161_),
    .A(_03158_),
    .B(_03160_));
 sg13g2_nand2_1 _09286_ (.Y(_03162_),
    .A(_03106_),
    .B(_03109_));
 sg13g2_nand2b_1 _09287_ (.Y(_03163_),
    .B(_03162_),
    .A_N(_03108_));
 sg13g2_nand3_1 _09288_ (.B(_03109_),
    .C(_03108_),
    .A(_03106_),
    .Y(_03164_));
 sg13g2_nand3_1 _09289_ (.B(_03163_),
    .C(_03164_),
    .A(_03161_),
    .Y(_03165_));
 sg13g2_a21oi_2 _09290_ (.B1(_03112_),
    .Y(_03166_),
    .A2(_03114_),
    .A1(_03076_));
 sg13g2_a21oi_1 _09291_ (.A1(_03115_),
    .A2(_03165_),
    .Y(_03167_),
    .B1(_03166_));
 sg13g2_nand3_1 _09292_ (.B(_03074_),
    .C(_03167_),
    .A(_03052_),
    .Y(_03169_));
 sg13g2_nand2_1 _09293_ (.Y(_03170_),
    .A(_03070_),
    .B(_03169_));
 sg13g2_nor2_1 _09294_ (.A(net87),
    .B(_02517_),
    .Y(_03171_));
 sg13g2_inv_1 _09295_ (.Y(_03172_),
    .A(_03000_));
 sg13g2_a21oi_1 _09296_ (.A1(_03002_),
    .A2(_03009_),
    .Y(_03173_),
    .B1(_03172_));
 sg13g2_inv_1 _09297_ (.Y(_03174_),
    .A(_03173_));
 sg13g2_nand3_1 _09298_ (.B(_02991_),
    .C(_02994_),
    .A(_02989_),
    .Y(_03175_));
 sg13g2_inv_1 _09299_ (.Y(_03176_),
    .A(_03175_));
 sg13g2_nor2b_1 _09300_ (.A(_03176_),
    .B_N(_02991_),
    .Y(_03177_));
 sg13g2_nor2_1 _09301_ (.A(net88),
    .B(_02655_),
    .Y(_03178_));
 sg13g2_nor2_1 _09302_ (.A(_03531_),
    .B(_02859_),
    .Y(_03180_));
 sg13g2_nor2_2 _09303_ (.A(net86),
    .B(_02940_),
    .Y(_03181_));
 sg13g2_xnor2_1 _09304_ (.Y(_03182_),
    .A(_03180_),
    .B(_03181_));
 sg13g2_xnor2_1 _09305_ (.Y(_03183_),
    .A(_03178_),
    .B(_03182_));
 sg13g2_nand2b_1 _09306_ (.Y(_03184_),
    .B(_02998_),
    .A_N(_02987_));
 sg13g2_nand3b_1 _09307_ (.B(_03184_),
    .C(_02986_),
    .Y(_03185_),
    .A_N(_03183_));
 sg13g2_nand2_1 _09308_ (.Y(_03186_),
    .A(_03184_),
    .B(_02986_));
 sg13g2_nand2_1 _09309_ (.Y(_03187_),
    .A(_03186_),
    .B(_03183_));
 sg13g2_nand3b_1 _09310_ (.B(_03185_),
    .C(_03187_),
    .Y(_03188_),
    .A_N(_03177_));
 sg13g2_nand2_1 _09311_ (.Y(_03189_),
    .A(_03185_),
    .B(_03187_));
 sg13g2_nand2_1 _09312_ (.Y(_03191_),
    .A(_03189_),
    .B(_03177_));
 sg13g2_nand2_1 _09313_ (.Y(_03192_),
    .A(_03188_),
    .B(_03191_));
 sg13g2_xnor2_1 _09314_ (.Y(_03193_),
    .A(_03174_),
    .B(_03192_));
 sg13g2_xnor2_1 _09315_ (.Y(_03194_),
    .A(_03171_),
    .B(_03193_));
 sg13g2_inv_2 _09316_ (.Y(_03195_),
    .A(_03194_));
 sg13g2_nand2_1 _09317_ (.Y(_03196_),
    .A(_03011_),
    .B(_02978_));
 sg13g2_nor2_1 _09318_ (.A(_02978_),
    .B(_03011_),
    .Y(_03197_));
 sg13g2_a21oi_1 _09319_ (.A1(_03196_),
    .A2(_02976_),
    .Y(_03198_),
    .B1(_03197_));
 sg13g2_inv_1 _09320_ (.Y(_03199_),
    .A(_03198_));
 sg13g2_nand2_1 _09321_ (.Y(_03200_),
    .A(_03195_),
    .B(_03199_));
 sg13g2_nand2_1 _09322_ (.Y(_03202_),
    .A(_03194_),
    .B(_03198_));
 sg13g2_nand2_1 _09323_ (.Y(_03203_),
    .A(_03200_),
    .B(_03202_));
 sg13g2_inv_1 _09324_ (.Y(_03204_),
    .A(_03203_));
 sg13g2_nand2_1 _09325_ (.Y(_03205_),
    .A(_03170_),
    .B(_03204_));
 sg13g2_nand3_1 _09326_ (.B(_03169_),
    .C(_03203_),
    .A(_03070_),
    .Y(_03206_));
 sg13g2_inv_4 _09327_ (.A(_05529_),
    .Y(_03207_));
 sg13g2_nor2_1 _09328_ (.A(_05528_),
    .B(_03207_),
    .Y(_03208_));
 sg13g2_nor2_1 _09329_ (.A(_05529_),
    .B(_05543_),
    .Y(_03209_));
 sg13g2_inv_1 _09330_ (.Y(_03210_),
    .A(_03209_));
 sg13g2_nor2_1 _09331_ (.A(_05542_),
    .B(_03210_),
    .Y(_03211_));
 sg13g2_buf_2 _09332_ (.A(_03211_),
    .X(_03213_));
 sg13g2_a21oi_2 _09333_ (.B1(_03213_),
    .Y(_03214_),
    .A2(_03208_),
    .A1(\frame_counter[9] ));
 sg13g2_buf_8 _09334_ (.A(_03214_),
    .X(_03215_));
 sg13g2_buf_1 _09335_ (.A(_03215_),
    .X(_03216_));
 sg13g2_nand3_1 _09336_ (.B(_03206_),
    .C(net48),
    .A(_03205_),
    .Y(_03217_));
 sg13g2_buf_1 _09337_ (.A(_03217_),
    .X(_03218_));
 sg13g2_a21oi_1 _09338_ (.A1(_05529_),
    .A2(_00018_),
    .Y(_03219_),
    .B1(_05531_));
 sg13g2_buf_8 _09339_ (.A(_03219_),
    .X(_03220_));
 sg13g2_inv_1 _09340_ (.Y(_03221_),
    .A(_03213_));
 sg13g2_nor2_1 _09341_ (.A(_05526_),
    .B(_03221_),
    .Y(_03222_));
 sg13g2_nand2_1 _09342_ (.Y(_03224_),
    .A(_03222_),
    .B(_00216_));
 sg13g2_inv_1 _09343_ (.Y(_03225_),
    .A(_03208_));
 sg13g2_nor3_1 _09344_ (.A(_05530_),
    .B(_05526_),
    .C(_03225_),
    .Y(_03226_));
 sg13g2_buf_1 _09345_ (.A(_03226_),
    .X(_03227_));
 sg13g2_a21oi_1 _09346_ (.A1(_03227_),
    .A2(net110),
    .Y(_03228_),
    .B1(net127));
 sg13g2_nand3_1 _09347_ (.B(net127),
    .C(_03245_),
    .A(_03227_),
    .Y(_03229_));
 sg13g2_nor2b_1 _09348_ (.A(_03228_),
    .B_N(_03229_),
    .Y(_03230_));
 sg13g2_xor2_1 _09349_ (.B(_03230_),
    .A(_03224_),
    .X(_03231_));
 sg13g2_nand2_1 _09350_ (.Y(_03232_),
    .A(_03222_),
    .B(net89));
 sg13g2_a21oi_1 _09351_ (.A1(_03227_),
    .A2(net108),
    .Y(_03233_),
    .B1(net128));
 sg13g2_nand3_1 _09352_ (.B(\hvsync_gen.vpos[1] ),
    .C(net108),
    .A(_03227_),
    .Y(_03235_));
 sg13g2_o21ai_1 _09353_ (.B1(_03235_),
    .Y(_03236_),
    .A1(_03232_),
    .A2(_03233_));
 sg13g2_nor2b_1 _09354_ (.A(_03231_),
    .B_N(_03236_),
    .Y(_03237_));
 sg13g2_xor2_1 _09355_ (.B(_03231_),
    .A(_03236_),
    .X(_03238_));
 sg13g2_nor2_1 _09356_ (.A(_02982_),
    .B(_03238_),
    .Y(_03239_));
 sg13g2_nor2_1 _09357_ (.A(_03237_),
    .B(_03239_),
    .Y(_03240_));
 sg13g2_nand2b_1 _09358_ (.Y(_03241_),
    .B(_03230_),
    .A_N(_03224_));
 sg13g2_nand2_1 _09359_ (.Y(_03242_),
    .A(_03222_),
    .B(_05568_));
 sg13g2_nand2_2 _09360_ (.Y(_03243_),
    .A(_03227_),
    .B(_05568_));
 sg13g2_xnor2_1 _09361_ (.Y(_03244_),
    .A(_04374_),
    .B(_03243_));
 sg13g2_xnor2_1 _09362_ (.Y(_03246_),
    .A(_03242_),
    .B(_03244_));
 sg13g2_a21oi_1 _09363_ (.A1(_03229_),
    .A2(_03241_),
    .Y(_03247_),
    .B1(_03246_));
 sg13g2_nand3_1 _09364_ (.B(_03229_),
    .C(_03241_),
    .A(_03246_),
    .Y(_03248_));
 sg13g2_nand2b_1 _09365_ (.Y(_03249_),
    .B(_03248_),
    .A_N(_03247_));
 sg13g2_xnor2_1 _09366_ (.Y(_03250_),
    .A(_03542_),
    .B(_03249_));
 sg13g2_xor2_1 _09367_ (.B(_03250_),
    .A(_03240_),
    .X(_03251_));
 sg13g2_nor2b_1 _09368_ (.A(_03233_),
    .B_N(_03235_),
    .Y(_03252_));
 sg13g2_xor2_1 _09369_ (.B(_03252_),
    .A(_03232_),
    .X(_03253_));
 sg13g2_nand2_1 _09370_ (.Y(_03254_),
    .A(_03222_),
    .B(\envelopeA[0] ));
 sg13g2_nand2_1 _09371_ (.Y(_03255_),
    .A(_03254_),
    .B(_00061_));
 sg13g2_nor2b_1 _09372_ (.A(_03253_),
    .B_N(_03255_),
    .Y(_03257_));
 sg13g2_xor2_1 _09373_ (.B(_03253_),
    .A(_03255_),
    .X(_03258_));
 sg13g2_nor2b_1 _09374_ (.A(_03258_),
    .B_N(_00216_),
    .Y(_03259_));
 sg13g2_nor2_1 _09375_ (.A(_03257_),
    .B(_03259_),
    .Y(_03260_));
 sg13g2_xnor2_1 _09376_ (.Y(_03261_),
    .A(_02982_),
    .B(_03238_));
 sg13g2_nor2_1 _09377_ (.A(_03260_),
    .B(_03261_),
    .Y(_03262_));
 sg13g2_xnor2_1 _09378_ (.Y(_03263_),
    .A(_03260_),
    .B(_03261_));
 sg13g2_nand2_1 _09379_ (.Y(_03264_),
    .A(_03227_),
    .B(_03311_));
 sg13g2_xnor2_1 _09380_ (.Y(_03265_),
    .A(_02499_),
    .B(_03254_));
 sg13g2_xor2_1 _09381_ (.B(_03265_),
    .A(_03264_),
    .X(_03266_));
 sg13g2_nor2_1 _09382_ (.A(_03264_),
    .B(_03265_),
    .Y(_03268_));
 sg13g2_a21oi_1 _09383_ (.A1(_03266_),
    .A2(_02458_),
    .Y(_03269_),
    .B1(_03268_));
 sg13g2_xor2_1 _09384_ (.B(_03258_),
    .A(_00216_),
    .X(_03270_));
 sg13g2_nor2_1 _09385_ (.A(_03269_),
    .B(_03270_),
    .Y(_03271_));
 sg13g2_nand2b_1 _09386_ (.Y(_03272_),
    .B(_03271_),
    .A_N(_03263_));
 sg13g2_nor2b_1 _09387_ (.A(_03262_),
    .B_N(_03272_),
    .Y(_03273_));
 sg13g2_xnor2_1 _09388_ (.Y(_03274_),
    .A(_03251_),
    .B(_03273_));
 sg13g2_inv_2 _09389_ (.Y(_03275_),
    .A(_03274_));
 sg13g2_nor2_1 _09390_ (.A(_03220_),
    .B(_03275_),
    .Y(_03276_));
 sg13g2_inv_1 _09391_ (.Y(_03277_),
    .A(_03276_));
 sg13g2_a21oi_1 _09392_ (.A1(_02703_),
    .A2(_02705_),
    .Y(_03279_),
    .B1(_02755_));
 sg13g2_nor2_1 _09393_ (.A(_03279_),
    .B(_02627_),
    .Y(_03280_));
 sg13g2_inv_2 _09394_ (.Y(_03281_),
    .A(_02700_));
 sg13g2_inv_1 _09395_ (.Y(_03282_),
    .A(_02805_));
 sg13g2_nor2_1 _09396_ (.A(_02802_),
    .B(_03282_),
    .Y(_03283_));
 sg13g2_nand2_1 _09397_ (.Y(_03284_),
    .A(_03167_),
    .B(_03071_));
 sg13g2_nand2_1 _09398_ (.Y(_03285_),
    .A(_03283_),
    .B(_03284_));
 sg13g2_nand3_1 _09399_ (.B(_03281_),
    .C(_03285_),
    .A(_03280_),
    .Y(_03286_));
 sg13g2_nand2_1 _09400_ (.Y(_03287_),
    .A(_03286_),
    .B(_02811_));
 sg13g2_inv_1 _09401_ (.Y(_03288_),
    .A(_03038_));
 sg13g2_nand3_1 _09402_ (.B(_03042_),
    .C(_03288_),
    .A(_03041_),
    .Y(_03290_));
 sg13g2_nand2_1 _09403_ (.Y(_03291_),
    .A(_03290_),
    .B(_03048_));
 sg13g2_nand2_1 _09404_ (.Y(_03292_),
    .A(_03055_),
    .B(_03053_));
 sg13g2_nor2_1 _09405_ (.A(_03291_),
    .B(_03292_),
    .Y(_03293_));
 sg13g2_nand2_1 _09406_ (.Y(_03294_),
    .A(_03287_),
    .B(_03293_));
 sg13g2_inv_4 _09407_ (.A(_03056_),
    .Y(_03295_));
 sg13g2_nand2_1 _09408_ (.Y(_03296_),
    .A(_03294_),
    .B(_03295_));
 sg13g2_nand2_1 _09409_ (.Y(_03297_),
    .A(_03296_),
    .B(_02973_));
 sg13g2_nand3_1 _09410_ (.B(_03061_),
    .C(_03295_),
    .A(_03294_),
    .Y(_03298_));
 sg13g2_inv_4 _09411_ (.A(_03215_),
    .Y(_03299_));
 sg13g2_nand3_1 _09412_ (.B(_03298_),
    .C(_03299_),
    .A(_03297_),
    .Y(_03301_));
 sg13g2_buf_1 _09413_ (.A(_03301_),
    .X(_03302_));
 sg13g2_nand3_1 _09414_ (.B(_03277_),
    .C(_03302_),
    .A(_03218_),
    .Y(_03303_));
 sg13g2_buf_1 _09415_ (.A(_03943_),
    .X(_03304_));
 sg13g2_nor2_1 _09416_ (.A(net124),
    .B(_05486_),
    .Y(_03305_));
 sg13g2_nor2_1 _09417_ (.A(_03245_),
    .B(_04715_),
    .Y(_03306_));
 sg13g2_nor2_1 _09418_ (.A(_03305_),
    .B(_03306_),
    .Y(_03307_));
 sg13g2_buf_8 _09419_ (.A(_03307_),
    .X(_03308_));
 sg13g2_inv_1 _09420_ (.Y(_03309_),
    .A(_03943_));
 sg13g2_nor2_1 _09421_ (.A(_00226_),
    .B(_03309_),
    .Y(_03310_));
 sg13g2_buf_2 _09422_ (.A(_03310_),
    .X(_03312_));
 sg13g2_inv_1 _09423_ (.Y(_03313_),
    .A(_03312_));
 sg13g2_inv_1 _09424_ (.Y(_03314_),
    .A(net123));
 sg13g2_nor2_1 _09425_ (.A(net109),
    .B(_03314_),
    .Y(_03315_));
 sg13g2_nor2_1 _09426_ (.A(net123),
    .B(net76),
    .Y(_03316_));
 sg13g2_nor2_1 _09427_ (.A(_03315_),
    .B(_03316_),
    .Y(_03317_));
 sg13g2_inv_1 _09428_ (.Y(_03318_),
    .A(_03317_));
 sg13g2_nor2_1 _09429_ (.A(_03305_),
    .B(_03318_),
    .Y(_03319_));
 sg13g2_inv_1 _09430_ (.Y(_03320_),
    .A(_03319_));
 sg13g2_nand2_1 _09431_ (.Y(_03321_),
    .A(_03318_),
    .B(_03305_));
 sg13g2_nand2_2 _09432_ (.Y(_03323_),
    .A(_03320_),
    .B(_03321_));
 sg13g2_nor2_1 _09433_ (.A(net60),
    .B(_03323_),
    .Y(_03324_));
 sg13g2_inv_1 _09434_ (.Y(_03325_),
    .A(_03324_));
 sg13g2_nor2_1 _09435_ (.A(net122),
    .B(net111),
    .Y(_03326_));
 sg13g2_nor2_1 _09436_ (.A(net93),
    .B(_02970_),
    .Y(_03327_));
 sg13g2_nor2_1 _09437_ (.A(_03326_),
    .B(_03327_),
    .Y(_03328_));
 sg13g2_o21ai_1 _09438_ (.B1(_03328_),
    .Y(_03329_),
    .A1(_03315_),
    .A2(_03319_));
 sg13g2_nor2_1 _09439_ (.A(_03315_),
    .B(_03319_),
    .Y(_03330_));
 sg13g2_nand2b_1 _09440_ (.Y(_03331_),
    .B(_03330_),
    .A_N(_03328_));
 sg13g2_nand2_2 _09441_ (.Y(_03332_),
    .A(_03329_),
    .B(_03331_));
 sg13g2_inv_1 _09442_ (.Y(_03334_),
    .A(_03332_));
 sg13g2_nand2_1 _09443_ (.Y(_03335_),
    .A(_03334_),
    .B(_02467_));
 sg13g2_xnor2_1 _09444_ (.Y(_03336_),
    .A(_03325_),
    .B(_03335_));
 sg13g2_o21ai_1 _09445_ (.B1(_03336_),
    .Y(_03337_),
    .A1(net85),
    .A2(_03308_));
 sg13g2_nor3_2 _09446_ (.A(net107),
    .B(_03308_),
    .C(_03325_),
    .Y(_03338_));
 sg13g2_nand2_1 _09447_ (.Y(_03339_),
    .A(_03337_),
    .B(_03338_));
 sg13g2_nor2_1 _09448_ (.A(_03325_),
    .B(_03335_),
    .Y(_03340_));
 sg13g2_nor2_1 _09449_ (.A(_03943_),
    .B(_03323_),
    .Y(_03341_));
 sg13g2_nand2_1 _09450_ (.Y(_03342_),
    .A(_03334_),
    .B(_03312_));
 sg13g2_nor2_1 _09451_ (.A(_02981_),
    .B(net86),
    .Y(_03343_));
 sg13g2_nor2_1 _09452_ (.A(_03443_),
    .B(net112),
    .Y(_03345_));
 sg13g2_nor2_1 _09453_ (.A(_03343_),
    .B(_03345_),
    .Y(_03346_));
 sg13g2_nor2_1 _09454_ (.A(_03315_),
    .B(_03327_),
    .Y(_03347_));
 sg13g2_a21oi_1 _09455_ (.A1(_03320_),
    .A2(_03347_),
    .Y(_03348_),
    .B1(_03326_));
 sg13g2_xnor2_1 _09456_ (.Y(_03349_),
    .A(_03346_),
    .B(_03348_));
 sg13g2_buf_2 _09457_ (.A(_03349_),
    .X(_03350_));
 sg13g2_nor2_1 _09458_ (.A(net107),
    .B(_03350_),
    .Y(_03351_));
 sg13g2_inv_1 _09459_ (.Y(_03352_),
    .A(_03351_));
 sg13g2_nor2_1 _09460_ (.A(_03342_),
    .B(_03352_),
    .Y(_03353_));
 sg13g2_nand2_1 _09461_ (.Y(_03354_),
    .A(_03352_),
    .B(_03342_));
 sg13g2_nor2b_1 _09462_ (.A(_03353_),
    .B_N(_03354_),
    .Y(_03356_));
 sg13g2_xnor2_1 _09463_ (.Y(_03357_),
    .A(_03341_),
    .B(_03356_));
 sg13g2_xnor2_1 _09464_ (.Y(_03358_),
    .A(_03340_),
    .B(_03357_));
 sg13g2_inv_1 _09465_ (.Y(_03359_),
    .A(_03358_));
 sg13g2_nor2_1 _09466_ (.A(_03339_),
    .B(_03359_),
    .Y(_03360_));
 sg13g2_inv_1 _09467_ (.Y(_03361_),
    .A(_03360_));
 sg13g2_nand2_1 _09468_ (.Y(_03362_),
    .A(_03359_),
    .B(_03339_));
 sg13g2_nor2_1 _09469_ (.A(_05528_),
    .B(_03210_),
    .Y(_03363_));
 sg13g2_nor2_1 _09470_ (.A(_05533_),
    .B(_03363_),
    .Y(_03364_));
 sg13g2_buf_1 _09471_ (.A(_03364_),
    .X(_03365_));
 sg13g2_inv_4 _09472_ (.A(net59),
    .Y(_03367_));
 sg13g2_nand3_1 _09473_ (.B(_03362_),
    .C(_03367_),
    .A(_03361_),
    .Y(_03368_));
 sg13g2_buf_1 _09474_ (.A(_03368_),
    .X(_03369_));
 sg13g2_a21oi_1 _09475_ (.A1(_03218_),
    .A2(_03302_),
    .Y(_03370_),
    .B1(_03277_));
 sg13g2_a21oi_2 _09476_ (.B1(_03370_),
    .Y(_03371_),
    .A2(_03369_),
    .A1(_03303_));
 sg13g2_inv_1 _09477_ (.Y(_03372_),
    .A(_03340_));
 sg13g2_nor2_1 _09478_ (.A(_03372_),
    .B(_03357_),
    .Y(_03373_));
 sg13g2_nor2_1 _09479_ (.A(_03373_),
    .B(_03360_),
    .Y(_03374_));
 sg13g2_a21oi_1 _09480_ (.A1(_03354_),
    .A2(_03341_),
    .Y(_03375_),
    .B1(_03353_));
 sg13g2_nor2_1 _09481_ (.A(net85),
    .B(_03332_),
    .Y(_03376_));
 sg13g2_inv_1 _09482_ (.Y(_03378_),
    .A(_03343_));
 sg13g2_a21oi_1 _09483_ (.A1(_03348_),
    .A2(_03378_),
    .Y(_03379_),
    .B1(_03345_));
 sg13g2_nor2_1 _09484_ (.A(net100),
    .B(net115),
    .Y(_03380_));
 sg13g2_nor2_1 _09485_ (.A(_02718_),
    .B(_02467_),
    .Y(_03381_));
 sg13g2_nor2_1 _09486_ (.A(_03380_),
    .B(_03381_),
    .Y(_03382_));
 sg13g2_nor2b_1 _09487_ (.A(_03379_),
    .B_N(_03382_),
    .Y(_03383_));
 sg13g2_nor2b_1 _09488_ (.A(_03382_),
    .B_N(_03379_),
    .Y(_03384_));
 sg13g2_nor2_2 _09489_ (.A(_03383_),
    .B(_03384_),
    .Y(_03385_));
 sg13g2_inv_1 _09490_ (.Y(_03386_),
    .A(_03385_));
 sg13g2_nor2_1 _09491_ (.A(net60),
    .B(_03386_),
    .Y(_03387_));
 sg13g2_inv_1 _09492_ (.Y(_03389_),
    .A(_03387_));
 sg13g2_nor2_1 _09493_ (.A(_03352_),
    .B(_03389_),
    .Y(_03390_));
 sg13g2_nand2_1 _09494_ (.Y(_03391_),
    .A(_03385_),
    .B(_03410_));
 sg13g2_o21ai_1 _09495_ (.B1(_03391_),
    .Y(_03392_),
    .A1(_03350_),
    .A2(net60));
 sg13g2_nor2b_1 _09496_ (.A(_03390_),
    .B_N(_03392_),
    .Y(_03393_));
 sg13g2_xnor2_1 _09497_ (.Y(_03394_),
    .A(_03376_),
    .B(_03393_));
 sg13g2_xnor2_1 _09498_ (.Y(_03395_),
    .A(_03375_),
    .B(_03394_));
 sg13g2_nor2_1 _09499_ (.A(_03374_),
    .B(_03395_),
    .Y(_03396_));
 sg13g2_nand2_1 _09500_ (.Y(_03397_),
    .A(_03395_),
    .B(_03374_));
 sg13g2_nand3b_1 _09501_ (.B(_03367_),
    .C(_03397_),
    .Y(_03398_),
    .A_N(_03396_));
 sg13g2_buf_1 _09502_ (.A(_03398_),
    .X(_03400_));
 sg13g2_nor2_1 _09503_ (.A(_02700_),
    .B(_03291_),
    .Y(_03401_));
 sg13g2_inv_1 _09504_ (.Y(_03402_),
    .A(_02623_));
 sg13g2_a21oi_1 _09505_ (.A1(_02626_),
    .A2(_02805_),
    .Y(_03403_),
    .B1(_03402_));
 sg13g2_nand2_1 _09506_ (.Y(_03404_),
    .A(_03401_),
    .B(_03403_));
 sg13g2_a21oi_1 _09507_ (.A1(_03290_),
    .A2(_02697_),
    .Y(_03405_),
    .B1(_03049_));
 sg13g2_inv_2 _09508_ (.Y(_03406_),
    .A(_03405_));
 sg13g2_nand2_1 _09509_ (.Y(_03407_),
    .A(_03404_),
    .B(_03406_));
 sg13g2_nor2_1 _09510_ (.A(_03061_),
    .B(_03292_),
    .Y(_03408_));
 sg13g2_inv_2 _09511_ (.Y(_03409_),
    .A(_03408_));
 sg13g2_inv_2 _09512_ (.Y(_03411_),
    .A(_03015_));
 sg13g2_nor2_1 _09513_ (.A(_03203_),
    .B(_03411_),
    .Y(_03412_));
 sg13g2_nor2b_1 _09514_ (.A(_03409_),
    .B_N(_03412_),
    .Y(_03413_));
 sg13g2_o21ai_1 _09515_ (.B1(_03200_),
    .Y(_03414_),
    .A1(_03065_),
    .A2(_03203_));
 sg13g2_nor2_1 _09516_ (.A(_03029_),
    .B(_03034_),
    .Y(_03415_));
 sg13g2_nand2_1 _09517_ (.Y(_03416_),
    .A(_03415_),
    .B(_03060_));
 sg13g2_nand2_1 _09518_ (.Y(_03417_),
    .A(_03416_),
    .B(_03059_));
 sg13g2_nand2_1 _09519_ (.Y(_03418_),
    .A(_03417_),
    .B(_03412_));
 sg13g2_nand2b_1 _09520_ (.Y(_03419_),
    .B(_03418_),
    .A_N(_03414_));
 sg13g2_a21oi_1 _09521_ (.A1(_03407_),
    .A2(_03413_),
    .Y(_03420_),
    .B1(_03419_));
 sg13g2_nor2b_1 _09522_ (.A(_02627_),
    .B_N(_02758_),
    .Y(_03422_));
 sg13g2_and2_1 _09523_ (.A(_03401_),
    .B(_03422_),
    .X(_03423_));
 sg13g2_nor2_1 _09524_ (.A(_03165_),
    .B(_03166_),
    .Y(_03424_));
 sg13g2_nand3_1 _09525_ (.B(_03115_),
    .C(_03424_),
    .A(_03072_),
    .Y(_03425_));
 sg13g2_inv_1 _09526_ (.Y(_03426_),
    .A(_03115_));
 sg13g2_o21ai_1 _09527_ (.B1(_03071_),
    .Y(_03427_),
    .A1(_03426_),
    .A2(_02802_));
 sg13g2_nand2_1 _09528_ (.Y(_03428_),
    .A(_03425_),
    .B(_03427_));
 sg13g2_nand3_1 _09529_ (.B(_03423_),
    .C(_03428_),
    .A(_03413_),
    .Y(_03429_));
 sg13g2_nand2_1 _09530_ (.Y(_03430_),
    .A(_03420_),
    .B(_03429_));
 sg13g2_nor2_1 _09531_ (.A(_03173_),
    .B(_03192_),
    .Y(_03431_));
 sg13g2_a21oi_1 _09532_ (.A1(_03193_),
    .A2(_03171_),
    .Y(_03433_),
    .B1(_03431_));
 sg13g2_nor2_1 _09533_ (.A(net87),
    .B(_02655_),
    .Y(_03434_));
 sg13g2_a22oi_1 _09534_ (.Y(_03435_),
    .B1(net100),
    .B2(_02827_),
    .A2(_02860_),
    .A1(net106));
 sg13g2_nor2_2 _09535_ (.A(net88),
    .B(_02859_),
    .Y(_03436_));
 sg13g2_nand2_1 _09536_ (.Y(_03437_),
    .A(_03181_),
    .B(_03436_));
 sg13g2_nand2b_1 _09537_ (.Y(_03438_),
    .B(_03437_),
    .A_N(_03435_));
 sg13g2_nor2b_1 _09538_ (.A(_03182_),
    .B_N(_03178_),
    .Y(_03439_));
 sg13g2_a21oi_1 _09539_ (.A1(_03181_),
    .A2(_03180_),
    .Y(_03440_),
    .B1(_03439_));
 sg13g2_xnor2_1 _09540_ (.Y(_03441_),
    .A(_03438_),
    .B(_03440_));
 sg13g2_and2_1 _09541_ (.A(_03188_),
    .B(_03187_),
    .X(_03442_));
 sg13g2_buf_1 _09542_ (.A(_03442_),
    .X(_03444_));
 sg13g2_xnor2_1 _09543_ (.Y(_03445_),
    .A(_03441_),
    .B(_03444_));
 sg13g2_xor2_1 _09544_ (.B(_03445_),
    .A(_03434_),
    .X(_03446_));
 sg13g2_xor2_1 _09545_ (.B(_03446_),
    .A(_03433_),
    .X(_03447_));
 sg13g2_nand2_1 _09546_ (.Y(_03448_),
    .A(_03430_),
    .B(_03447_));
 sg13g2_inv_1 _09547_ (.Y(_03449_),
    .A(_03447_));
 sg13g2_nand3_1 _09548_ (.B(_03429_),
    .C(_03449_),
    .A(_03420_),
    .Y(_03450_));
 sg13g2_nand3_1 _09549_ (.B(_03450_),
    .C(_03215_),
    .A(_03448_),
    .Y(_03451_));
 sg13g2_nand2_1 _09550_ (.Y(_03452_),
    .A(_03408_),
    .B(_03401_));
 sg13g2_nand2_1 _09551_ (.Y(_03453_),
    .A(_03071_),
    .B(_02805_));
 sg13g2_nor2_1 _09552_ (.A(_02802_),
    .B(_03167_),
    .Y(_03455_));
 sg13g2_nor2_1 _09553_ (.A(_03453_),
    .B(_03455_),
    .Y(_03456_));
 sg13g2_nor2b_1 _09554_ (.A(_03279_),
    .B_N(_02626_),
    .Y(_03457_));
 sg13g2_nand2_1 _09555_ (.Y(_03458_),
    .A(_03456_),
    .B(_03457_));
 sg13g2_nor2b_1 _09556_ (.A(_03282_),
    .B_N(_02626_),
    .Y(_03459_));
 sg13g2_a21oi_2 _09557_ (.B1(_03402_),
    .Y(_03460_),
    .A2(_03459_),
    .A1(_03458_));
 sg13g2_nand2b_1 _09558_ (.Y(_03461_),
    .B(_03460_),
    .A_N(_03452_));
 sg13g2_nand2_1 _09559_ (.Y(_03462_),
    .A(_03408_),
    .B(_03405_));
 sg13g2_inv_1 _09560_ (.Y(_03463_),
    .A(_03417_));
 sg13g2_nand2_1 _09561_ (.Y(_03464_),
    .A(_03462_),
    .B(_03463_));
 sg13g2_inv_1 _09562_ (.Y(_03466_),
    .A(_03464_));
 sg13g2_nand2_1 _09563_ (.Y(_03467_),
    .A(_03461_),
    .B(_03466_));
 sg13g2_nand2_1 _09564_ (.Y(_03468_),
    .A(_03467_),
    .B(_03015_));
 sg13g2_nand3_1 _09565_ (.B(_03411_),
    .C(_03466_),
    .A(_03461_),
    .Y(_03469_));
 sg13g2_nand3_1 _09566_ (.B(_03469_),
    .C(_03299_),
    .A(_03468_),
    .Y(_03470_));
 sg13g2_nand2_1 _09567_ (.Y(_03471_),
    .A(_03451_),
    .B(_03470_));
 sg13g2_a21oi_1 _09568_ (.A1(_03248_),
    .A2(_03531_),
    .Y(_03472_),
    .B1(_03247_));
 sg13g2_xnor2_1 _09569_ (.Y(_03473_),
    .A(_00019_),
    .B(_03243_));
 sg13g2_inv_1 _09570_ (.Y(_03474_),
    .A(_03243_));
 sg13g2_nor2_1 _09571_ (.A(_03242_),
    .B(_03244_),
    .Y(_03475_));
 sg13g2_a21oi_1 _09572_ (.A1(net129),
    .A2(_03474_),
    .Y(_03477_),
    .B1(_03475_));
 sg13g2_xnor2_1 _09573_ (.Y(_03478_),
    .A(_03473_),
    .B(_03477_));
 sg13g2_xnor2_1 _09574_ (.Y(_03479_),
    .A(net86),
    .B(_03478_));
 sg13g2_xor2_1 _09575_ (.B(_03479_),
    .A(_03472_),
    .X(_03480_));
 sg13g2_nand2b_1 _09576_ (.Y(_03481_),
    .B(_03251_),
    .A_N(_03273_));
 sg13g2_o21ai_1 _09577_ (.B1(_03481_),
    .Y(_03482_),
    .A1(_03240_),
    .A2(_03250_));
 sg13g2_or2_1 _09578_ (.X(_03483_),
    .B(_03482_),
    .A(_03480_));
 sg13g2_nand2_1 _09579_ (.Y(_03484_),
    .A(_03482_),
    .B(_03480_));
 sg13g2_nand2_2 _09580_ (.Y(_03485_),
    .A(_03483_),
    .B(_03484_));
 sg13g2_nor2_1 _09581_ (.A(_03220_),
    .B(_03485_),
    .Y(_03486_));
 sg13g2_nand2_1 _09582_ (.Y(_03488_),
    .A(_03471_),
    .B(_03486_));
 sg13g2_inv_1 _09583_ (.Y(_03489_),
    .A(_03486_));
 sg13g2_nand3_1 _09584_ (.B(_03489_),
    .C(_03470_),
    .A(_03451_),
    .Y(_03490_));
 sg13g2_buf_1 _09585_ (.A(_03490_),
    .X(_03491_));
 sg13g2_nand2_1 _09586_ (.Y(_03492_),
    .A(_03488_),
    .B(_03491_));
 sg13g2_nand2b_1 _09587_ (.Y(_03493_),
    .B(_03492_),
    .A_N(_03400_));
 sg13g2_nand3_1 _09588_ (.B(_03491_),
    .C(_03400_),
    .A(_03488_),
    .Y(_03494_));
 sg13g2_nand2_1 _09589_ (.Y(_03495_),
    .A(_03493_),
    .B(_03494_));
 sg13g2_nand2b_1 _09590_ (.Y(_03496_),
    .B(_03495_),
    .A_N(_03371_));
 sg13g2_nand3_1 _09591_ (.B(_03494_),
    .C(_03371_),
    .A(_03493_),
    .Y(_03497_));
 sg13g2_nand2_1 _09592_ (.Y(_03499_),
    .A(_03496_),
    .B(_03497_));
 sg13g2_xnor2_1 _09593_ (.Y(_03500_),
    .A(_03269_),
    .B(_03270_));
 sg13g2_buf_1 _09594_ (.A(_03500_),
    .X(_03501_));
 sg13g2_nor2_1 _09595_ (.A(net85),
    .B(_03501_),
    .Y(_03502_));
 sg13g2_xor2_1 _09596_ (.B(_03263_),
    .A(_03271_),
    .X(_03503_));
 sg13g2_buf_8 _09597_ (.A(_03503_),
    .X(_03504_));
 sg13g2_nor2_1 _09598_ (.A(net60),
    .B(_03504_),
    .Y(_03505_));
 sg13g2_nor2_1 _09599_ (.A(net107),
    .B(_03275_),
    .Y(_03506_));
 sg13g2_xnor2_1 _09600_ (.Y(_03507_),
    .A(_03505_),
    .B(_03506_));
 sg13g2_xor2_1 _09601_ (.B(_03507_),
    .A(_03502_),
    .X(_03508_));
 sg13g2_nor2_1 _09602_ (.A(_03313_),
    .B(_03501_),
    .Y(_03510_));
 sg13g2_inv_1 _09603_ (.Y(_03511_),
    .A(_03510_));
 sg13g2_nor2_1 _09604_ (.A(net100),
    .B(_03504_),
    .Y(_03512_));
 sg13g2_inv_1 _09605_ (.Y(_03513_),
    .A(_03512_));
 sg13g2_nor2_1 _09606_ (.A(_03511_),
    .B(_03513_),
    .Y(_03514_));
 sg13g2_nor2b_1 _09607_ (.A(_03508_),
    .B_N(_03514_),
    .Y(_03515_));
 sg13g2_xnor2_1 _09608_ (.Y(_03516_),
    .A(_03514_),
    .B(_03508_));
 sg13g2_nand2b_1 _09609_ (.Y(_03517_),
    .B(_02369_),
    .A_N(_03266_));
 sg13g2_nand2_1 _09610_ (.Y(_03518_),
    .A(_03266_),
    .B(_02458_));
 sg13g2_nand2_2 _09611_ (.Y(_03519_),
    .A(_03517_),
    .B(_03518_));
 sg13g2_xnor2_1 _09612_ (.Y(_03521_),
    .A(_03510_),
    .B(_03512_));
 sg13g2_o21ai_1 _09613_ (.B1(_03521_),
    .Y(_03522_),
    .A1(_03304_),
    .A2(_03519_));
 sg13g2_nor2_1 _09614_ (.A(net107),
    .B(_03501_),
    .Y(_03523_));
 sg13g2_nor2_1 _09615_ (.A(_03313_),
    .B(_03519_),
    .Y(_03524_));
 sg13g2_nand2_1 _09616_ (.Y(_03525_),
    .A(_03523_),
    .B(_03524_));
 sg13g2_inv_1 _09617_ (.Y(_03526_),
    .A(_03525_));
 sg13g2_nand2_1 _09618_ (.Y(_03527_),
    .A(_03522_),
    .B(_03526_));
 sg13g2_inv_2 _09619_ (.Y(_03528_),
    .A(_03527_));
 sg13g2_nand2_1 _09620_ (.Y(_03529_),
    .A(_03516_),
    .B(_03528_));
 sg13g2_inv_1 _09621_ (.Y(_03530_),
    .A(_03529_));
 sg13g2_nor2_1 _09622_ (.A(_03515_),
    .B(_03530_),
    .Y(_03532_));
 sg13g2_nor2b_1 _09623_ (.A(_03507_),
    .B_N(_03502_),
    .Y(_03533_));
 sg13g2_a21oi_1 _09624_ (.A1(_03505_),
    .A2(_03506_),
    .Y(_03534_),
    .B1(_03533_));
 sg13g2_nor2_1 _09625_ (.A(net85),
    .B(_03504_),
    .Y(_03535_));
 sg13g2_nand3_1 _09626_ (.B(_03410_),
    .C(_03484_),
    .A(_03483_),
    .Y(_03536_));
 sg13g2_nor3_1 _09627_ (.A(net60),
    .B(_03275_),
    .C(_03536_),
    .Y(_03537_));
 sg13g2_o21ai_1 _09628_ (.B1(_03536_),
    .Y(_03538_),
    .A1(net60),
    .A2(_03275_));
 sg13g2_nor2b_1 _09629_ (.A(_03537_),
    .B_N(_03538_),
    .Y(_03539_));
 sg13g2_xnor2_1 _09630_ (.Y(_03540_),
    .A(_03535_),
    .B(_03539_));
 sg13g2_nor2_1 _09631_ (.A(_03534_),
    .B(_03540_),
    .Y(_03541_));
 sg13g2_inv_1 _09632_ (.Y(_03543_),
    .A(_03541_));
 sg13g2_nand2_1 _09633_ (.Y(_03544_),
    .A(_03540_),
    .B(_03534_));
 sg13g2_nand2_1 _09634_ (.Y(_03545_),
    .A(_03543_),
    .B(_03544_));
 sg13g2_nor2_1 _09635_ (.A(_03532_),
    .B(_03545_),
    .Y(_03546_));
 sg13g2_and2_1 _09636_ (.A(_03545_),
    .B(_03532_),
    .X(_03547_));
 sg13g2_nor3_1 _09637_ (.A(_03365_),
    .B(_03546_),
    .C(_03547_),
    .Y(_03548_));
 sg13g2_nand2_1 _09638_ (.Y(_03549_),
    .A(_03499_),
    .B(_03548_));
 sg13g2_inv_1 _09639_ (.Y(_03550_),
    .A(_03548_));
 sg13g2_nand3_1 _09640_ (.B(_03497_),
    .C(_03550_),
    .A(_03496_),
    .Y(_03551_));
 sg13g2_nand2_1 _09641_ (.Y(_03552_),
    .A(_03549_),
    .B(_03551_));
 sg13g2_nand2_1 _09642_ (.Y(_03554_),
    .A(_03218_),
    .B(_03302_));
 sg13g2_nand2_1 _09643_ (.Y(_03555_),
    .A(_03554_),
    .B(_03277_));
 sg13g2_nand3_1 _09644_ (.B(_03276_),
    .C(_03302_),
    .A(_03218_),
    .Y(_03556_));
 sg13g2_nand2_1 _09645_ (.Y(_03557_),
    .A(_03555_),
    .B(_03556_));
 sg13g2_nand2_1 _09646_ (.Y(_03558_),
    .A(_03557_),
    .B(_03369_));
 sg13g2_inv_1 _09647_ (.Y(_03559_),
    .A(_03369_));
 sg13g2_nand3_1 _09648_ (.B(_03556_),
    .C(_03559_),
    .A(_03555_),
    .Y(_03560_));
 sg13g2_nand2_1 _09649_ (.Y(_03561_),
    .A(_03558_),
    .B(_03560_));
 sg13g2_nand3_1 _09650_ (.B(_03469_),
    .C(net48),
    .A(_03468_),
    .Y(_03562_));
 sg13g2_nand2_1 _09651_ (.Y(_03563_),
    .A(_03458_),
    .B(_03459_));
 sg13g2_nand3_1 _09652_ (.B(_03401_),
    .C(_02623_),
    .A(_03563_),
    .Y(_03565_));
 sg13g2_nand2_1 _09653_ (.Y(_03566_),
    .A(_03565_),
    .B(_03406_));
 sg13g2_nand2_1 _09654_ (.Y(_03567_),
    .A(_03566_),
    .B(_03035_));
 sg13g2_nand3_1 _09655_ (.B(_03292_),
    .C(_03406_),
    .A(_03565_),
    .Y(_03568_));
 sg13g2_nand3_1 _09656_ (.B(_03568_),
    .C(_03299_),
    .A(_03567_),
    .Y(_03569_));
 sg13g2_nor2_1 _09657_ (.A(_03220_),
    .B(_03504_),
    .Y(_03570_));
 sg13g2_inv_1 _09658_ (.Y(_03571_),
    .A(_03570_));
 sg13g2_nand3_1 _09659_ (.B(_03569_),
    .C(_03571_),
    .A(_03562_),
    .Y(_03572_));
 sg13g2_buf_1 _09660_ (.A(_03572_),
    .X(_03573_));
 sg13g2_nor2_1 _09661_ (.A(_03338_),
    .B(_03337_),
    .Y(_03574_));
 sg13g2_inv_1 _09662_ (.Y(_03576_),
    .A(_03339_));
 sg13g2_nor3_1 _09663_ (.A(net59),
    .B(_03574_),
    .C(_03576_),
    .Y(_03577_));
 sg13g2_inv_1 _09664_ (.Y(_03578_),
    .A(_03577_));
 sg13g2_nand2_1 _09665_ (.Y(_03579_),
    .A(_03468_),
    .B(_03469_));
 sg13g2_nand2_1 _09666_ (.Y(_03580_),
    .A(_03579_),
    .B(net48));
 sg13g2_nand2_1 _09667_ (.Y(_03581_),
    .A(_03567_),
    .B(_03568_));
 sg13g2_nand2_1 _09668_ (.Y(_03582_),
    .A(_03581_),
    .B(_03299_));
 sg13g2_nand3_1 _09669_ (.B(_03582_),
    .C(_03570_),
    .A(_03580_),
    .Y(_03583_));
 sg13g2_inv_1 _09670_ (.Y(_03584_),
    .A(_03583_));
 sg13g2_a21oi_1 _09671_ (.A1(_03573_),
    .A2(_03578_),
    .Y(_03585_),
    .B1(_03584_));
 sg13g2_nand2_1 _09672_ (.Y(_03587_),
    .A(_03561_),
    .B(_03585_));
 sg13g2_nor2_1 _09673_ (.A(_03528_),
    .B(_03516_),
    .Y(_03588_));
 sg13g2_nor3_2 _09674_ (.A(net59),
    .B(_03588_),
    .C(_03530_),
    .Y(_03589_));
 sg13g2_nor2_1 _09675_ (.A(_03585_),
    .B(_03561_),
    .Y(_03590_));
 sg13g2_a21oi_2 _09676_ (.B1(_03590_),
    .Y(_03591_),
    .A2(_03589_),
    .A1(_03587_));
 sg13g2_nand2_1 _09677_ (.Y(_03592_),
    .A(_03552_),
    .B(_03591_));
 sg13g2_buf_8 _09678_ (.A(_03220_),
    .X(_03593_));
 sg13g2_nor2_1 _09679_ (.A(_02740_),
    .B(_02562_),
    .Y(_03594_));
 sg13g2_nor2_1 _09680_ (.A(_03932_),
    .B(_02751_),
    .Y(_03595_));
 sg13g2_nor2_1 _09681_ (.A(_03594_),
    .B(_03595_),
    .Y(_03596_));
 sg13g2_inv_1 _09682_ (.Y(_03598_),
    .A(_03380_));
 sg13g2_o21ai_1 _09683_ (.B1(_03598_),
    .Y(_03599_),
    .A1(_03381_),
    .A2(_03379_));
 sg13g2_or2_1 _09684_ (.X(_03600_),
    .B(_03599_),
    .A(_03596_));
 sg13g2_nand2_1 _09685_ (.Y(_03601_),
    .A(_03599_),
    .B(_03596_));
 sg13g2_nand2_1 _09686_ (.Y(_03602_),
    .A(_03600_),
    .B(_03601_));
 sg13g2_buf_8 _09687_ (.A(_03602_),
    .X(_03603_));
 sg13g2_nor2_1 _09688_ (.A(net66),
    .B(_03603_),
    .Y(_03604_));
 sg13g2_inv_1 _09689_ (.Y(_03605_),
    .A(_03604_));
 sg13g2_nor2_1 _09690_ (.A(_03591_),
    .B(_03552_),
    .Y(_03606_));
 sg13g2_a21oi_1 _09691_ (.A1(_03592_),
    .A2(_03605_),
    .Y(_03607_),
    .B1(_03606_));
 sg13g2_inv_1 _09692_ (.Y(_03609_),
    .A(_03607_));
 sg13g2_nand2_1 _09693_ (.Y(_03610_),
    .A(_03495_),
    .B(_03371_));
 sg13g2_nor2_1 _09694_ (.A(_03371_),
    .B(_03495_),
    .Y(_03611_));
 sg13g2_a21oi_1 _09695_ (.A1(_03610_),
    .A2(_03548_),
    .Y(_03612_),
    .B1(_03611_));
 sg13g2_a21oi_1 _09696_ (.A1(_03451_),
    .A2(_03470_),
    .Y(_03613_),
    .B1(_03489_));
 sg13g2_a21oi_2 _09697_ (.B1(_03613_),
    .Y(_03614_),
    .A2(_03400_),
    .A1(_03491_));
 sg13g2_nor2_1 _09698_ (.A(_03375_),
    .B(_03394_),
    .Y(_03615_));
 sg13g2_a21oi_1 _09699_ (.A1(_03392_),
    .A2(_03376_),
    .Y(_03616_),
    .B1(_03390_));
 sg13g2_nor2_1 _09700_ (.A(net85),
    .B(_03350_),
    .Y(_03617_));
 sg13g2_nand3_1 _09701_ (.B(_03312_),
    .C(_03601_),
    .A(_03600_),
    .Y(_03618_));
 sg13g2_nor2_1 _09702_ (.A(_03391_),
    .B(_03618_),
    .Y(_03619_));
 sg13g2_nor2_1 _09703_ (.A(net107),
    .B(_03603_),
    .Y(_03620_));
 sg13g2_inv_1 _09704_ (.Y(_03621_),
    .A(_03620_));
 sg13g2_nand2_1 _09705_ (.Y(_03622_),
    .A(_03621_),
    .B(_03389_));
 sg13g2_nand2b_1 _09706_ (.Y(_03623_),
    .B(_03622_),
    .A_N(_03619_));
 sg13g2_xor2_1 _09707_ (.B(_03623_),
    .A(_03617_),
    .X(_03624_));
 sg13g2_xor2_1 _09708_ (.B(_03624_),
    .A(_03616_),
    .X(_03625_));
 sg13g2_nor3_1 _09709_ (.A(_03615_),
    .B(_03396_),
    .C(_03625_),
    .Y(_03626_));
 sg13g2_o21ai_1 _09710_ (.B1(_03625_),
    .Y(_03627_),
    .A1(_03615_),
    .A2(_03396_));
 sg13g2_nand3b_1 _09711_ (.B(_03367_),
    .C(_03627_),
    .Y(_03628_),
    .A_N(_03626_));
 sg13g2_nand2_1 _09712_ (.Y(_03630_),
    .A(_03293_),
    .B(_02810_));
 sg13g2_nand2_1 _09713_ (.Y(_03631_),
    .A(_03630_),
    .B(_03295_));
 sg13g2_nand2_1 _09714_ (.Y(_03632_),
    .A(_03447_),
    .B(_03204_));
 sg13g2_nor2_1 _09715_ (.A(_03632_),
    .B(_03016_),
    .Y(_03633_));
 sg13g2_inv_1 _09716_ (.Y(_03634_),
    .A(_03200_));
 sg13g2_nor2_1 _09717_ (.A(_03433_),
    .B(_03446_),
    .Y(_03635_));
 sg13g2_a21oi_1 _09718_ (.A1(_03447_),
    .A2(_03634_),
    .Y(_03636_),
    .B1(_03635_));
 sg13g2_o21ai_1 _09719_ (.B1(_03636_),
    .Y(_03637_),
    .A1(_03632_),
    .A2(_03067_));
 sg13g2_a21oi_1 _09720_ (.A1(_03631_),
    .A2(_03633_),
    .Y(_03638_),
    .B1(_03637_));
 sg13g2_nand2_1 _09721_ (.Y(_03639_),
    .A(_03293_),
    .B(_02701_));
 sg13g2_nor2b_1 _09722_ (.A(_03639_),
    .B_N(_03633_),
    .Y(_03641_));
 sg13g2_inv_1 _09723_ (.Y(_03642_),
    .A(_03166_));
 sg13g2_and3_1 _09724_ (.X(_03643_),
    .A(_03163_),
    .B(_03164_),
    .C(_03159_));
 sg13g2_a21oi_1 _09725_ (.A1(_03642_),
    .A2(_03643_),
    .Y(_03644_),
    .B1(_03426_));
 sg13g2_nor2_1 _09726_ (.A(_03644_),
    .B(_03073_),
    .Y(_03645_));
 sg13g2_nor2_1 _09727_ (.A(_02807_),
    .B(_03645_),
    .Y(_03646_));
 sg13g2_a21oi_1 _09728_ (.A1(_03163_),
    .A2(_03164_),
    .Y(_03647_),
    .B1(_03159_));
 sg13g2_nor4_1 _09729_ (.A(_03647_),
    .B(_03166_),
    .C(_03426_),
    .D(_03643_),
    .Y(_03648_));
 sg13g2_nand3_1 _09730_ (.B(_03143_),
    .C(_03116_),
    .A(_03142_),
    .Y(_03649_));
 sg13g2_nand3_1 _09731_ (.B(_03649_),
    .C(_03150_),
    .A(_03145_),
    .Y(_03650_));
 sg13g2_inv_1 _09732_ (.Y(_03652_),
    .A(_03153_));
 sg13g2_nor2b_1 _09733_ (.A(_03159_),
    .B_N(_03156_),
    .Y(_03653_));
 sg13g2_nor2_1 _09734_ (.A(_03652_),
    .B(_03653_),
    .Y(_03654_));
 sg13g2_nand2_1 _09735_ (.Y(_03655_),
    .A(_03653_),
    .B(_03652_));
 sg13g2_o21ai_1 _09736_ (.B1(_03655_),
    .Y(_03656_),
    .A1(_03650_),
    .A2(_03654_));
 sg13g2_nand4_1 _09737_ (.B(_03072_),
    .C(_03656_),
    .A(_03648_),
    .Y(_03657_),
    .D(_02758_));
 sg13g2_nand2_1 _09738_ (.Y(_03658_),
    .A(_03646_),
    .B(_03657_));
 sg13g2_nand2_1 _09739_ (.Y(_03659_),
    .A(_03641_),
    .B(_03658_));
 sg13g2_nand2_1 _09740_ (.Y(_03660_),
    .A(_03638_),
    .B(_03659_));
 sg13g2_nor2_1 _09741_ (.A(net87),
    .B(_02940_),
    .Y(_03661_));
 sg13g2_nand2_1 _09742_ (.Y(_03663_),
    .A(_03437_),
    .B(_03436_));
 sg13g2_nor2_1 _09743_ (.A(_03438_),
    .B(_03440_),
    .Y(_03664_));
 sg13g2_xnor2_1 _09744_ (.Y(_03665_),
    .A(_03663_),
    .B(_03664_));
 sg13g2_xor2_1 _09745_ (.B(_03665_),
    .A(_03661_),
    .X(_03666_));
 sg13g2_inv_1 _09746_ (.Y(_03667_),
    .A(_03666_));
 sg13g2_nand2_1 _09747_ (.Y(_03668_),
    .A(_03444_),
    .B(_03441_));
 sg13g2_nor2_1 _09748_ (.A(_03441_),
    .B(_03444_),
    .Y(_03669_));
 sg13g2_a21oi_1 _09749_ (.A1(_03668_),
    .A2(_03434_),
    .Y(_03670_),
    .B1(_03669_));
 sg13g2_nor2_1 _09750_ (.A(_03667_),
    .B(_03670_),
    .Y(_03671_));
 sg13g2_inv_1 _09751_ (.Y(_03672_),
    .A(_03671_));
 sg13g2_nand2_1 _09752_ (.Y(_03674_),
    .A(_03670_),
    .B(_03667_));
 sg13g2_nand2_1 _09753_ (.Y(_03675_),
    .A(_03672_),
    .B(_03674_));
 sg13g2_inv_1 _09754_ (.Y(_03676_),
    .A(_03675_));
 sg13g2_nand2_1 _09755_ (.Y(_03677_),
    .A(_03660_),
    .B(_03676_));
 sg13g2_nand3_1 _09756_ (.B(_03675_),
    .C(_03659_),
    .A(_03638_),
    .Y(_03678_));
 sg13g2_nand3_1 _09757_ (.B(_03678_),
    .C(_03215_),
    .A(_03677_),
    .Y(_03679_));
 sg13g2_nand3_1 _09758_ (.B(_03206_),
    .C(_03299_),
    .A(_03205_),
    .Y(_03680_));
 sg13g2_nand2_1 _09759_ (.Y(_03681_),
    .A(_03679_),
    .B(_03680_));
 sg13g2_inv_1 _09760_ (.Y(_03682_),
    .A(_00020_));
 sg13g2_nand2_1 _09761_ (.Y(_03683_),
    .A(_03474_),
    .B(_00019_));
 sg13g2_xnor2_1 _09762_ (.Y(_03685_),
    .A(_03682_),
    .B(_03683_));
 sg13g2_xnor2_1 _09763_ (.Y(_03686_),
    .A(net61),
    .B(_03685_));
 sg13g2_nor2_1 _09764_ (.A(_03473_),
    .B(_03477_),
    .Y(_03687_));
 sg13g2_nor2_1 _09765_ (.A(_02737_),
    .B(_03478_),
    .Y(_03688_));
 sg13g2_nor2_1 _09766_ (.A(_03687_),
    .B(_03688_),
    .Y(_03689_));
 sg13g2_xnor2_1 _09767_ (.Y(_03690_),
    .A(_03686_),
    .B(_03689_));
 sg13g2_o21ai_1 _09768_ (.B1(_03484_),
    .Y(_03691_),
    .A1(_03472_),
    .A2(_03479_));
 sg13g2_or2_1 _09769_ (.X(_03692_),
    .B(_03691_),
    .A(_03690_));
 sg13g2_nand2_1 _09770_ (.Y(_03693_),
    .A(_03691_),
    .B(_03690_));
 sg13g2_nand2_2 _09771_ (.Y(_03694_),
    .A(_03692_),
    .B(_03693_));
 sg13g2_nor2_1 _09772_ (.A(_03220_),
    .B(_03694_),
    .Y(_03696_));
 sg13g2_nand2_1 _09773_ (.Y(_03697_),
    .A(_03681_),
    .B(_03696_));
 sg13g2_inv_1 _09774_ (.Y(_03698_),
    .A(_03696_));
 sg13g2_nand3_1 _09775_ (.B(_03698_),
    .C(_03680_),
    .A(_03679_),
    .Y(_03699_));
 sg13g2_nand2_1 _09776_ (.Y(_03700_),
    .A(_03697_),
    .B(_03699_));
 sg13g2_nand2b_1 _09777_ (.Y(_03701_),
    .B(_03700_),
    .A_N(_03628_));
 sg13g2_nand3_1 _09778_ (.B(_03699_),
    .C(_03628_),
    .A(_03697_),
    .Y(_03702_));
 sg13g2_nand2_1 _09779_ (.Y(_03703_),
    .A(_03701_),
    .B(_03702_));
 sg13g2_nand2b_1 _09780_ (.Y(_03704_),
    .B(_03703_),
    .A_N(_03614_));
 sg13g2_nand3_1 _09781_ (.B(_03702_),
    .C(_03614_),
    .A(_03701_),
    .Y(_03705_));
 sg13g2_nand2_1 _09782_ (.Y(_03707_),
    .A(_03704_),
    .B(_03705_));
 sg13g2_a21oi_1 _09783_ (.A1(_03538_),
    .A2(_03535_),
    .Y(_03708_),
    .B1(_03537_));
 sg13g2_nor2_1 _09784_ (.A(_03304_),
    .B(_03275_),
    .Y(_03709_));
 sg13g2_nor2_1 _09785_ (.A(net60),
    .B(_03485_),
    .Y(_03710_));
 sg13g2_nor2_1 _09786_ (.A(net107),
    .B(_03694_),
    .Y(_03711_));
 sg13g2_xnor2_1 _09787_ (.Y(_03712_),
    .A(_03710_),
    .B(_03711_));
 sg13g2_xor2_1 _09788_ (.B(_03712_),
    .A(_03709_),
    .X(_03713_));
 sg13g2_xor2_1 _09789_ (.B(_03713_),
    .A(_03708_),
    .X(_03714_));
 sg13g2_or3_1 _09790_ (.A(_03541_),
    .B(_03546_),
    .C(_03714_),
    .X(_03715_));
 sg13g2_o21ai_1 _09791_ (.B1(_03714_),
    .Y(_03716_),
    .A1(_03541_),
    .A2(_03546_));
 sg13g2_nand3_1 _09792_ (.B(_03367_),
    .C(_03716_),
    .A(_03715_),
    .Y(_03718_));
 sg13g2_inv_1 _09793_ (.Y(_03719_),
    .A(_03718_));
 sg13g2_nand2_1 _09794_ (.Y(_03720_),
    .A(_03707_),
    .B(_03719_));
 sg13g2_nand3_1 _09795_ (.B(_03705_),
    .C(_03718_),
    .A(_03704_),
    .Y(_03721_));
 sg13g2_nand2_1 _09796_ (.Y(_03722_),
    .A(_03720_),
    .B(_03721_));
 sg13g2_nand2b_1 _09797_ (.Y(_03723_),
    .B(_03722_),
    .A_N(_03612_));
 sg13g2_nand3_1 _09798_ (.B(_03721_),
    .C(_03612_),
    .A(_03720_),
    .Y(_03724_));
 sg13g2_nand2_1 _09799_ (.Y(_03725_),
    .A(_03723_),
    .B(_03724_));
 sg13g2_a21oi_1 _09800_ (.A1(_03599_),
    .A2(_03596_),
    .Y(_03726_),
    .B1(_03595_));
 sg13g2_xnor2_1 _09801_ (.Y(_03727_),
    .A(_02597_),
    .B(_03726_));
 sg13g2_inv_2 _09802_ (.Y(_03729_),
    .A(_03727_));
 sg13g2_nor2_1 _09803_ (.A(net66),
    .B(_03729_),
    .Y(_03730_));
 sg13g2_inv_1 _09804_ (.Y(_03731_),
    .A(_03730_));
 sg13g2_nand2_1 _09805_ (.Y(_03732_),
    .A(_03725_),
    .B(_03731_));
 sg13g2_nand3_1 _09806_ (.B(_03724_),
    .C(_03730_),
    .A(_03723_),
    .Y(_03733_));
 sg13g2_nand3_1 _09807_ (.B(_03732_),
    .C(_03733_),
    .A(_03609_),
    .Y(_03734_));
 sg13g2_nand2_1 _09808_ (.Y(_03735_),
    .A(_03732_),
    .B(_03733_));
 sg13g2_nand2_1 _09809_ (.Y(_03736_),
    .A(_03735_),
    .B(_03607_));
 sg13g2_nand2_1 _09810_ (.Y(_03737_),
    .A(_03734_),
    .B(_03736_));
 sg13g2_nand2_1 _09811_ (.Y(_03738_),
    .A(_03722_),
    .B(_03612_));
 sg13g2_nor2_1 _09812_ (.A(_03612_),
    .B(_03722_),
    .Y(_03740_));
 sg13g2_a21oi_1 _09813_ (.A1(_03738_),
    .A2(_03731_),
    .Y(_03741_),
    .B1(_03740_));
 sg13g2_inv_1 _09814_ (.Y(_03742_),
    .A(_03741_));
 sg13g2_a21oi_1 _09815_ (.A1(_03679_),
    .A2(_03680_),
    .Y(_03743_),
    .B1(_03698_));
 sg13g2_a21oi_2 _09816_ (.B1(_03743_),
    .Y(_03744_),
    .A2(_03628_),
    .A1(_03699_));
 sg13g2_inv_2 _09817_ (.Y(_03745_),
    .A(_03744_));
 sg13g2_a21oi_1 _09818_ (.A1(_03622_),
    .A2(_03617_),
    .Y(_03746_),
    .B1(_03619_));
 sg13g2_nor2_1 _09819_ (.A(net85),
    .B(_03386_),
    .Y(_03747_));
 sg13g2_nor2_1 _09820_ (.A(net60),
    .B(_03729_),
    .Y(_03748_));
 sg13g2_inv_1 _09821_ (.Y(_03749_),
    .A(_03748_));
 sg13g2_o21ai_1 _09822_ (.B1(_03618_),
    .Y(_03751_),
    .A1(_03421_),
    .A2(_03729_));
 sg13g2_o21ai_1 _09823_ (.B1(_03751_),
    .Y(_03752_),
    .A1(_03621_),
    .A2(_03749_));
 sg13g2_xor2_1 _09824_ (.B(_03752_),
    .A(_03747_),
    .X(_03753_));
 sg13g2_xor2_1 _09825_ (.B(_03753_),
    .A(_03746_),
    .X(_03754_));
 sg13g2_o21ai_1 _09826_ (.B1(_03627_),
    .Y(_03755_),
    .A1(_03616_),
    .A2(_03624_));
 sg13g2_or2_1 _09827_ (.X(_03756_),
    .B(_03755_),
    .A(_03754_));
 sg13g2_nand2_1 _09828_ (.Y(_03757_),
    .A(_03755_),
    .B(_03754_));
 sg13g2_nand3_1 _09829_ (.B(_03367_),
    .C(_03757_),
    .A(_03756_),
    .Y(_03758_));
 sg13g2_nor2_1 _09830_ (.A(_03675_),
    .B(_03449_),
    .Y(_03759_));
 sg13g2_nand2_1 _09831_ (.Y(_03760_),
    .A(_03759_),
    .B(_03412_));
 sg13g2_inv_2 _09832_ (.Y(_03762_),
    .A(_03760_));
 sg13g2_nand2_1 _09833_ (.Y(_03763_),
    .A(_03414_),
    .B(_03759_));
 sg13g2_a21oi_1 _09834_ (.A1(_03676_),
    .A2(_03635_),
    .Y(_03764_),
    .B1(_03671_));
 sg13g2_nand2_1 _09835_ (.Y(_03765_),
    .A(_03763_),
    .B(_03764_));
 sg13g2_a21oi_1 _09836_ (.A1(_03464_),
    .A2(_03762_),
    .Y(_03766_),
    .B1(_03765_));
 sg13g2_inv_1 _09837_ (.Y(_03767_),
    .A(_03452_));
 sg13g2_nand3_1 _09838_ (.B(_03767_),
    .C(_03762_),
    .A(_03460_),
    .Y(_03768_));
 sg13g2_nand2_1 _09839_ (.Y(_03769_),
    .A(_03766_),
    .B(_03768_));
 sg13g2_a22oi_1 _09840_ (.Y(_03770_),
    .B1(_03436_),
    .B2(_03181_),
    .A2(_02860_),
    .A1(net118));
 sg13g2_nand3_1 _09841_ (.B(net118),
    .C(_03436_),
    .A(_03181_),
    .Y(_03771_));
 sg13g2_nor2b_1 _09842_ (.A(_03770_),
    .B_N(_03771_),
    .Y(_03773_));
 sg13g2_nor3_1 _09843_ (.A(_03438_),
    .B(_03663_),
    .C(_03440_),
    .Y(_03774_));
 sg13g2_a21oi_1 _09844_ (.A1(_03665_),
    .A2(_03661_),
    .Y(_03775_),
    .B1(_03774_));
 sg13g2_nor2b_1 _09845_ (.A(_03773_),
    .B_N(_03775_),
    .Y(_03776_));
 sg13g2_nand2b_1 _09846_ (.Y(_03777_),
    .B(_03773_),
    .A_N(_03775_));
 sg13g2_nor2b_1 _09847_ (.A(_03776_),
    .B_N(_03777_),
    .Y(_03778_));
 sg13g2_nand2_1 _09848_ (.Y(_03779_),
    .A(_03769_),
    .B(_03778_));
 sg13g2_inv_1 _09849_ (.Y(_03780_),
    .A(_03778_));
 sg13g2_nand3_1 _09850_ (.B(_03768_),
    .C(_03780_),
    .A(_03766_),
    .Y(_03781_));
 sg13g2_nand2_1 _09851_ (.Y(_03782_),
    .A(_03779_),
    .B(_03781_));
 sg13g2_nand2_1 _09852_ (.Y(_03783_),
    .A(_03782_),
    .B(net48));
 sg13g2_nand2_1 _09853_ (.Y(_03784_),
    .A(_03448_),
    .B(_03450_));
 sg13g2_nand2_1 _09854_ (.Y(_03785_),
    .A(_03784_),
    .B(_03299_));
 sg13g2_nand2_1 _09855_ (.Y(_03786_),
    .A(_03474_),
    .B(_00020_));
 sg13g2_nor2_1 _09856_ (.A(_00019_),
    .B(_03786_),
    .Y(_03787_));
 sg13g2_a21oi_1 _09857_ (.A1(_03685_),
    .A2(net56),
    .Y(_03788_),
    .B1(_03787_));
 sg13g2_nand2_1 _09858_ (.Y(_03789_),
    .A(_00429_),
    .B(net74));
 sg13g2_inv_1 _09859_ (.Y(_03790_),
    .A(_03789_));
 sg13g2_inv_1 _09860_ (.Y(_03791_),
    .A(_00023_));
 sg13g2_xnor2_1 _09861_ (.Y(_03792_),
    .A(_03791_),
    .B(_03786_));
 sg13g2_xnor2_1 _09862_ (.Y(_03794_),
    .A(_03790_),
    .B(_03792_));
 sg13g2_xor2_1 _09863_ (.B(_03794_),
    .A(_03788_),
    .X(_03795_));
 sg13g2_o21ai_1 _09864_ (.B1(_03686_),
    .Y(_03796_),
    .A1(_03687_),
    .A2(_03688_));
 sg13g2_nand2_1 _09865_ (.Y(_03797_),
    .A(_03693_),
    .B(_03796_));
 sg13g2_or2_1 _09866_ (.X(_03798_),
    .B(_03797_),
    .A(_03795_));
 sg13g2_nand2_1 _09867_ (.Y(_03799_),
    .A(_03797_),
    .B(_03795_));
 sg13g2_nand2_2 _09868_ (.Y(_03800_),
    .A(_03798_),
    .B(_03799_));
 sg13g2_nor2_1 _09869_ (.A(_03593_),
    .B(_03800_),
    .Y(_03801_));
 sg13g2_nand3_1 _09870_ (.B(_03785_),
    .C(_03801_),
    .A(_03783_),
    .Y(_03802_));
 sg13g2_nand3_1 _09871_ (.B(_03781_),
    .C(net48),
    .A(_03779_),
    .Y(_03803_));
 sg13g2_nand3_1 _09872_ (.B(_03450_),
    .C(_03299_),
    .A(_03448_),
    .Y(_03804_));
 sg13g2_inv_1 _09873_ (.Y(_03805_),
    .A(_03801_));
 sg13g2_nand3_1 _09874_ (.B(_03804_),
    .C(_03805_),
    .A(_03803_),
    .Y(_03806_));
 sg13g2_nand2_1 _09875_ (.Y(_03807_),
    .A(_03802_),
    .B(_03806_));
 sg13g2_nand2b_1 _09876_ (.Y(_03808_),
    .B(_03807_),
    .A_N(_03758_));
 sg13g2_nand3_1 _09877_ (.B(_03806_),
    .C(_03758_),
    .A(_03802_),
    .Y(_03809_));
 sg13g2_buf_1 _09878_ (.A(_03809_),
    .X(_03810_));
 sg13g2_nand3_1 _09879_ (.B(_03808_),
    .C(_03810_),
    .A(_03745_),
    .Y(_03811_));
 sg13g2_nand2_1 _09880_ (.Y(_03812_),
    .A(_03808_),
    .B(_03810_));
 sg13g2_nand2_1 _09881_ (.Y(_03813_),
    .A(_03812_),
    .B(_03744_));
 sg13g2_inv_1 _09882_ (.Y(_03815_),
    .A(_03694_));
 sg13g2_nand2_1 _09883_ (.Y(_03816_),
    .A(_03815_),
    .B(_03312_));
 sg13g2_nor2_1 _09884_ (.A(_03536_),
    .B(_03816_),
    .Y(_03817_));
 sg13g2_nand2b_1 _09885_ (.Y(_03818_),
    .B(_03709_),
    .A_N(_03712_));
 sg13g2_nor2b_1 _09886_ (.A(_03817_),
    .B_N(_03818_),
    .Y(_03819_));
 sg13g2_nor2_1 _09887_ (.A(net85),
    .B(_03485_),
    .Y(_03820_));
 sg13g2_inv_1 _09888_ (.Y(_03821_),
    .A(_03800_));
 sg13g2_nand2_1 _09889_ (.Y(_03822_),
    .A(_03821_),
    .B(_03410_));
 sg13g2_nor2_1 _09890_ (.A(_03816_),
    .B(_03822_),
    .Y(_03823_));
 sg13g2_nand2_1 _09891_ (.Y(_03824_),
    .A(_03822_),
    .B(_03816_));
 sg13g2_nor2b_1 _09892_ (.A(_03823_),
    .B_N(_03824_),
    .Y(_03826_));
 sg13g2_xnor2_1 _09893_ (.Y(_03827_),
    .A(_03820_),
    .B(_03826_));
 sg13g2_xor2_1 _09894_ (.B(_03827_),
    .A(_03819_),
    .X(_03828_));
 sg13g2_o21ai_1 _09895_ (.B1(_03716_),
    .Y(_03829_),
    .A1(_03708_),
    .A2(_03713_));
 sg13g2_or2_1 _09896_ (.X(_03830_),
    .B(_03829_),
    .A(_03828_));
 sg13g2_nand2_1 _09897_ (.Y(_03831_),
    .A(_03829_),
    .B(_03828_));
 sg13g2_nand3_1 _09898_ (.B(_03367_),
    .C(_03831_),
    .A(_03830_),
    .Y(_03832_));
 sg13g2_inv_1 _09899_ (.Y(_03833_),
    .A(_03832_));
 sg13g2_nand3_1 _09900_ (.B(_03813_),
    .C(_03833_),
    .A(_03811_),
    .Y(_03834_));
 sg13g2_nand2_1 _09901_ (.Y(_03835_),
    .A(_03812_),
    .B(_03745_));
 sg13g2_nand3_1 _09902_ (.B(_03744_),
    .C(_03810_),
    .A(_03808_),
    .Y(_03836_));
 sg13g2_nand3_1 _09903_ (.B(_03836_),
    .C(_03832_),
    .A(_03835_),
    .Y(_03837_));
 sg13g2_nand2_1 _09904_ (.Y(_03838_),
    .A(_03834_),
    .B(_03837_));
 sg13g2_nand2_1 _09905_ (.Y(_03839_),
    .A(_03703_),
    .B(_03614_));
 sg13g2_nor2_1 _09906_ (.A(_03614_),
    .B(_03703_),
    .Y(_03840_));
 sg13g2_a21oi_2 _09907_ (.B1(_03840_),
    .Y(_03841_),
    .A2(_03719_),
    .A1(_03839_));
 sg13g2_inv_2 _09908_ (.Y(_03842_),
    .A(_03841_));
 sg13g2_nand2_1 _09909_ (.Y(_03843_),
    .A(_03838_),
    .B(_03842_));
 sg13g2_nand3_1 _09910_ (.B(_03834_),
    .C(_03837_),
    .A(_03841_),
    .Y(_03844_));
 sg13g2_nor2_1 _09911_ (.A(_00021_),
    .B(_03726_),
    .Y(_03845_));
 sg13g2_inv_1 _09912_ (.Y(_03847_),
    .A(_03845_));
 sg13g2_nand2_1 _09913_ (.Y(_03848_),
    .A(_03847_),
    .B(_05513_));
 sg13g2_nand2_1 _09914_ (.Y(_03849_),
    .A(_03845_),
    .B(_05512_));
 sg13g2_nand2_2 _09915_ (.Y(_03850_),
    .A(_03848_),
    .B(_03849_));
 sg13g2_nor2_1 _09916_ (.A(net66),
    .B(_03850_),
    .Y(_03851_));
 sg13g2_nand3_1 _09917_ (.B(_03844_),
    .C(_03851_),
    .A(_03843_),
    .Y(_03852_));
 sg13g2_nand3_1 _09918_ (.B(_03837_),
    .C(_03834_),
    .A(_03842_),
    .Y(_03853_));
 sg13g2_nand2_1 _09919_ (.Y(_03854_),
    .A(_03838_),
    .B(_03841_));
 sg13g2_inv_1 _09920_ (.Y(_03855_),
    .A(_03851_));
 sg13g2_nand3_1 _09921_ (.B(_03854_),
    .C(_03855_),
    .A(_03853_),
    .Y(_03856_));
 sg13g2_nand3_1 _09922_ (.B(_03852_),
    .C(_03856_),
    .A(_03742_),
    .Y(_03858_));
 sg13g2_nand2_1 _09923_ (.Y(_03859_),
    .A(_03856_),
    .B(_03852_));
 sg13g2_nand2_1 _09924_ (.Y(_03860_),
    .A(_03859_),
    .B(_03741_));
 sg13g2_nand2_1 _09925_ (.Y(_03861_),
    .A(_03858_),
    .B(_03860_));
 sg13g2_nor2_1 _09926_ (.A(_03737_),
    .B(_03861_),
    .Y(_03862_));
 sg13g2_inv_1 _09927_ (.Y(_03863_),
    .A(_03591_));
 sg13g2_nand2_1 _09928_ (.Y(_03864_),
    .A(_03552_),
    .B(_03863_));
 sg13g2_nand3_1 _09929_ (.B(_03551_),
    .C(_03591_),
    .A(_03549_),
    .Y(_03865_));
 sg13g2_nand2_1 _09930_ (.Y(_03866_),
    .A(_03864_),
    .B(_03865_));
 sg13g2_nand2_1 _09931_ (.Y(_03867_),
    .A(_03866_),
    .B(_03605_));
 sg13g2_nand3_1 _09932_ (.B(_03865_),
    .C(_03604_),
    .A(_03864_),
    .Y(_03869_));
 sg13g2_nand2_1 _09933_ (.Y(_03870_),
    .A(_03867_),
    .B(_03869_));
 sg13g2_nand2b_1 _09934_ (.Y(_03871_),
    .B(_03561_),
    .A_N(_03585_));
 sg13g2_nand3_1 _09935_ (.B(_03560_),
    .C(_03585_),
    .A(_03558_),
    .Y(_03872_));
 sg13g2_nand2_1 _09936_ (.Y(_03873_),
    .A(_03871_),
    .B(_03872_));
 sg13g2_nand2_1 _09937_ (.Y(_03874_),
    .A(_03873_),
    .B(_03589_));
 sg13g2_inv_1 _09938_ (.Y(_03875_),
    .A(_03589_));
 sg13g2_nand3_1 _09939_ (.B(_03872_),
    .C(_03875_),
    .A(_03871_),
    .Y(_03876_));
 sg13g2_nand2_1 _09940_ (.Y(_03877_),
    .A(_03874_),
    .B(_03876_));
 sg13g2_nand2_1 _09941_ (.Y(_03878_),
    .A(_03583_),
    .B(_03573_));
 sg13g2_nand2_1 _09942_ (.Y(_03879_),
    .A(_03878_),
    .B(_03577_));
 sg13g2_nand3_1 _09943_ (.B(_03573_),
    .C(_03578_),
    .A(_03583_),
    .Y(_03880_));
 sg13g2_nand2_1 _09944_ (.Y(_03881_),
    .A(_03879_),
    .B(_03880_));
 sg13g2_nor2_1 _09945_ (.A(net66),
    .B(_03501_),
    .Y(_03882_));
 sg13g2_nand2_1 _09946_ (.Y(_03883_),
    .A(_03297_),
    .B(_03298_));
 sg13g2_nand2_1 _09947_ (.Y(_03884_),
    .A(_03287_),
    .B(_03050_));
 sg13g2_nand3_1 _09948_ (.B(_03291_),
    .C(_02811_),
    .A(_03286_),
    .Y(_03885_));
 sg13g2_a21oi_1 _09949_ (.A1(_03884_),
    .A2(_03885_),
    .Y(_03886_),
    .B1(net48));
 sg13g2_a21oi_1 _09950_ (.A1(_03883_),
    .A2(_03216_),
    .Y(_03887_),
    .B1(_03886_));
 sg13g2_nor2_1 _09951_ (.A(_03882_),
    .B(_03887_),
    .Y(_03888_));
 sg13g2_nand2_1 _09952_ (.Y(_03889_),
    .A(_03881_),
    .B(_03888_));
 sg13g2_nor2_1 _09953_ (.A(_03526_),
    .B(_03522_),
    .Y(_03890_));
 sg13g2_nor3_1 _09954_ (.A(net59),
    .B(_03890_),
    .C(_03528_),
    .Y(_03891_));
 sg13g2_nand3b_1 _09955_ (.B(_03879_),
    .C(_03880_),
    .Y(_03892_),
    .A_N(_03888_));
 sg13g2_inv_1 _09956_ (.Y(_03893_),
    .A(_03892_));
 sg13g2_a21oi_1 _09957_ (.A1(_03889_),
    .A2(_03891_),
    .Y(_03894_),
    .B1(_03893_));
 sg13g2_nand2_1 _09958_ (.Y(_03895_),
    .A(_03877_),
    .B(_03894_));
 sg13g2_nor2_1 _09959_ (.A(net66),
    .B(_03386_),
    .Y(_03896_));
 sg13g2_inv_1 _09960_ (.Y(_03897_),
    .A(_03896_));
 sg13g2_nor2_1 _09961_ (.A(_03894_),
    .B(_03877_),
    .Y(_03898_));
 sg13g2_a21oi_2 _09962_ (.B1(_03898_),
    .Y(_03900_),
    .A2(_03897_),
    .A1(_03895_));
 sg13g2_nand2_1 _09963_ (.Y(_03901_),
    .A(_03870_),
    .B(_03900_));
 sg13g2_nand2_1 _09964_ (.Y(_03902_),
    .A(_03892_),
    .B(_03889_));
 sg13g2_nand2_1 _09965_ (.Y(_03903_),
    .A(_03902_),
    .B(_03891_));
 sg13g2_inv_1 _09966_ (.Y(_03904_),
    .A(_03891_));
 sg13g2_nand3_1 _09967_ (.B(_03889_),
    .C(_03904_),
    .A(_03892_),
    .Y(_03905_));
 sg13g2_nand3_1 _09968_ (.B(_03568_),
    .C(_03216_),
    .A(_03567_),
    .Y(_03906_));
 sg13g2_inv_1 _09969_ (.Y(_03907_),
    .A(_03220_));
 sg13g2_nand3_1 _09970_ (.B(_03907_),
    .C(_03518_),
    .A(_03517_),
    .Y(_03908_));
 sg13g2_a21oi_1 _09971_ (.A1(_03460_),
    .A2(_03281_),
    .Y(_03909_),
    .B1(net48));
 sg13g2_o21ai_1 _09972_ (.B1(_03909_),
    .Y(_03911_),
    .A1(_03281_),
    .A2(_03460_));
 sg13g2_nand3_1 _09973_ (.B(_03908_),
    .C(_03911_),
    .A(_03906_),
    .Y(_03912_));
 sg13g2_nor3_1 _09974_ (.A(_03421_),
    .B(_03308_),
    .C(net59),
    .Y(_03913_));
 sg13g2_inv_1 _09975_ (.Y(_03914_),
    .A(_03913_));
 sg13g2_a21oi_1 _09976_ (.A1(_03906_),
    .A2(_03911_),
    .Y(_03915_),
    .B1(_03908_));
 sg13g2_a21oi_1 _09977_ (.A1(_03912_),
    .A2(_03914_),
    .Y(_03916_),
    .B1(_03915_));
 sg13g2_xor2_1 _09978_ (.B(_03887_),
    .A(_03882_),
    .X(_03917_));
 sg13g2_nand2_1 _09979_ (.Y(_03918_),
    .A(_03916_),
    .B(_03917_));
 sg13g2_or2_1 _09980_ (.X(_03919_),
    .B(_03523_),
    .A(_03524_));
 sg13g2_nand3_1 _09981_ (.B(_03367_),
    .C(_03525_),
    .A(_03919_),
    .Y(_03920_));
 sg13g2_inv_1 _09982_ (.Y(_03922_),
    .A(_03920_));
 sg13g2_nor2_1 _09983_ (.A(_03917_),
    .B(_03916_),
    .Y(_03923_));
 sg13g2_a21oi_1 _09984_ (.A1(_03918_),
    .A2(_03922_),
    .Y(_03924_),
    .B1(_03923_));
 sg13g2_nand3_1 _09985_ (.B(_03905_),
    .C(_03924_),
    .A(_03903_),
    .Y(_03925_));
 sg13g2_buf_1 _09986_ (.A(_03925_),
    .X(_03926_));
 sg13g2_nor2_1 _09987_ (.A(net66),
    .B(_03350_),
    .Y(_03927_));
 sg13g2_inv_1 _09988_ (.Y(_03928_),
    .A(_03927_));
 sg13g2_nand2_1 _09989_ (.Y(_03929_),
    .A(_03903_),
    .B(_03905_));
 sg13g2_nand2b_1 _09990_ (.Y(_03930_),
    .B(_03929_),
    .A_N(_03924_));
 sg13g2_inv_1 _09991_ (.Y(_03931_),
    .A(_03930_));
 sg13g2_a21oi_2 _09992_ (.B1(_03931_),
    .Y(_03933_),
    .A2(_03928_),
    .A1(_03926_));
 sg13g2_nand2b_1 _09993_ (.Y(_03934_),
    .B(_03877_),
    .A_N(_03894_));
 sg13g2_nand3_1 _09994_ (.B(_03876_),
    .C(_03894_),
    .A(_03874_),
    .Y(_03935_));
 sg13g2_nand2_1 _09995_ (.Y(_03936_),
    .A(_03934_),
    .B(_03935_));
 sg13g2_nand2_1 _09996_ (.Y(_03937_),
    .A(_03936_),
    .B(_03897_));
 sg13g2_nand3_1 _09997_ (.B(_03935_),
    .C(_03896_),
    .A(_03934_),
    .Y(_03938_));
 sg13g2_nand2_1 _09998_ (.Y(_03939_),
    .A(_03937_),
    .B(_03938_));
 sg13g2_nor2_1 _09999_ (.A(_03933_),
    .B(_03939_),
    .Y(_03940_));
 sg13g2_nor2_1 _10000_ (.A(_03900_),
    .B(_03870_),
    .Y(_03941_));
 sg13g2_a21oi_1 _10001_ (.A1(_03901_),
    .A2(_03940_),
    .Y(_03942_),
    .B1(_03941_));
 sg13g2_inv_1 _10002_ (.Y(_03944_),
    .A(_03942_));
 sg13g2_inv_2 _10003_ (.Y(_03945_),
    .A(_03734_));
 sg13g2_nand2_1 _10004_ (.Y(_03946_),
    .A(_03945_),
    .B(_03860_));
 sg13g2_nand2_1 _10005_ (.Y(_03947_),
    .A(_03946_),
    .B(_03858_));
 sg13g2_a21oi_1 _10006_ (.A1(_03862_),
    .A2(_03944_),
    .Y(_03948_),
    .B1(_03947_));
 sg13g2_nor2_1 _10007_ (.A(_03593_),
    .B(_03332_),
    .Y(_03949_));
 sg13g2_nand2b_1 _10008_ (.Y(_03950_),
    .B(_03912_),
    .A_N(_03915_));
 sg13g2_nand2_1 _10009_ (.Y(_03951_),
    .A(_03950_),
    .B(_03914_));
 sg13g2_nand3b_1 _10010_ (.B(_03913_),
    .C(_03912_),
    .Y(_03952_),
    .A_N(_03915_));
 sg13g2_inv_1 _10011_ (.Y(_03953_),
    .A(_03308_));
 sg13g2_inv_2 _10012_ (.Y(_03955_),
    .A(_03323_));
 sg13g2_a22oi_1 _10013_ (.Y(_03956_),
    .B1(_03410_),
    .B2(_03955_),
    .A2(_03312_),
    .A1(_03953_));
 sg13g2_nor3_2 _10014_ (.A(_03956_),
    .B(net59),
    .C(_03338_),
    .Y(_03957_));
 sg13g2_nand3_1 _10015_ (.B(_03952_),
    .C(_03957_),
    .A(_03951_),
    .Y(_03958_));
 sg13g2_nor3_1 _10016_ (.A(net100),
    .B(net59),
    .C(_03519_),
    .Y(_03959_));
 sg13g2_a21oi_1 _10017_ (.A1(_03951_),
    .A2(_03952_),
    .Y(_03960_),
    .B1(_03957_));
 sg13g2_a21oi_1 _10018_ (.A1(_03958_),
    .A2(_03959_),
    .Y(_03961_),
    .B1(_03960_));
 sg13g2_nor2b_1 _10019_ (.A(_03923_),
    .B_N(_03918_),
    .Y(_03962_));
 sg13g2_xnor2_1 _10020_ (.Y(_03963_),
    .A(_03922_),
    .B(_03962_));
 sg13g2_nor2_1 _10021_ (.A(_03961_),
    .B(_03963_),
    .Y(_03964_));
 sg13g2_inv_1 _10022_ (.Y(_03966_),
    .A(_03964_));
 sg13g2_nand2_1 _10023_ (.Y(_03967_),
    .A(_03963_),
    .B(_03961_));
 sg13g2_nand2_1 _10024_ (.Y(_03968_),
    .A(_03966_),
    .B(_03967_));
 sg13g2_xnor2_1 _10025_ (.Y(_03969_),
    .A(_03949_),
    .B(_03968_));
 sg13g2_nand2b_1 _10026_ (.Y(_03970_),
    .B(_03958_),
    .A_N(_03960_));
 sg13g2_xor2_1 _10027_ (.B(_03970_),
    .A(_03959_),
    .X(_03971_));
 sg13g2_nand2_1 _10028_ (.Y(_03972_),
    .A(_03971_),
    .B(_03957_));
 sg13g2_nand2_1 _10029_ (.Y(_03973_),
    .A(_03955_),
    .B(_03907_));
 sg13g2_nor2_1 _10030_ (.A(_03957_),
    .B(_03971_),
    .Y(_03974_));
 sg13g2_a21oi_1 _10031_ (.A1(_03972_),
    .A2(_03973_),
    .Y(_03975_),
    .B1(_03974_));
 sg13g2_nor2_2 _10032_ (.A(_03969_),
    .B(_03975_),
    .Y(_03977_));
 sg13g2_nand2_1 _10033_ (.Y(_03978_),
    .A(_03930_),
    .B(_03926_));
 sg13g2_nand2_1 _10034_ (.Y(_03979_),
    .A(_03978_),
    .B(_03927_));
 sg13g2_nand3_1 _10035_ (.B(_03926_),
    .C(_03928_),
    .A(_03930_),
    .Y(_03980_));
 sg13g2_nand2_1 _10036_ (.Y(_03981_),
    .A(_03979_),
    .B(_03980_));
 sg13g2_inv_1 _10037_ (.Y(_03982_),
    .A(_03949_));
 sg13g2_a21oi_1 _10038_ (.A1(_03967_),
    .A2(_03982_),
    .Y(_03983_),
    .B1(_03964_));
 sg13g2_nand2_1 _10039_ (.Y(_03984_),
    .A(_03981_),
    .B(_03983_));
 sg13g2_nor2_1 _10040_ (.A(_03983_),
    .B(_03981_),
    .Y(_03985_));
 sg13g2_a21oi_1 _10041_ (.A1(_03977_),
    .A2(_03984_),
    .Y(_03986_),
    .B1(_03985_));
 sg13g2_inv_1 _10042_ (.Y(_03988_),
    .A(_03986_));
 sg13g2_xnor2_1 _10043_ (.Y(_03989_),
    .A(_03933_),
    .B(_03939_));
 sg13g2_xnor2_1 _10044_ (.Y(_03990_),
    .A(_03900_),
    .B(_03870_));
 sg13g2_nor2_1 _10045_ (.A(_03989_),
    .B(_03990_),
    .Y(_03991_));
 sg13g2_nand3_1 _10046_ (.B(_03988_),
    .C(_03991_),
    .A(_03862_),
    .Y(_03992_));
 sg13g2_nand2_1 _10047_ (.Y(_03993_),
    .A(_03948_),
    .B(_03992_));
 sg13g2_inv_1 _10048_ (.Y(_03994_),
    .A(_03853_));
 sg13g2_a21oi_1 _10049_ (.A1(_03854_),
    .A2(_03855_),
    .Y(_03995_),
    .B1(_03994_));
 sg13g2_o21ai_1 _10050_ (.B1(_03757_),
    .Y(_03996_),
    .A1(_03746_),
    .A2(_03753_));
 sg13g2_a22oi_1 _10051_ (.Y(_03997_),
    .B1(_03747_),
    .B2(_03751_),
    .A2(_03748_),
    .A1(_03620_));
 sg13g2_nor2_1 _10052_ (.A(_02783_),
    .B(_03850_),
    .Y(_03999_));
 sg13g2_o21ai_1 _10053_ (.B1(_03749_),
    .Y(_04000_),
    .A1(net85),
    .A2(_03603_));
 sg13g2_xor2_1 _10054_ (.B(_04000_),
    .A(_03999_),
    .X(_04001_));
 sg13g2_xnor2_1 _10055_ (.Y(_04002_),
    .A(_03997_),
    .B(_04001_));
 sg13g2_a21oi_1 _10056_ (.A1(_03996_),
    .A2(_04002_),
    .Y(_04003_),
    .B1(net59));
 sg13g2_o21ai_1 _10057_ (.B1(_04003_),
    .Y(_04004_),
    .A1(_03996_),
    .A2(_04002_));
 sg13g2_inv_1 _10058_ (.Y(_04005_),
    .A(_00228_));
 sg13g2_nor2_1 _10059_ (.A(_03791_),
    .B(_03243_),
    .Y(_04006_));
 sg13g2_xnor2_1 _10060_ (.Y(_04007_),
    .A(_00025_),
    .B(_04006_));
 sg13g2_xnor2_1 _10061_ (.Y(_04008_),
    .A(_04005_),
    .B(_04007_));
 sg13g2_inv_1 _10062_ (.Y(_04010_),
    .A(_04008_));
 sg13g2_a22oi_1 _10063_ (.Y(_04011_),
    .B1(_03790_),
    .B2(_03792_),
    .A2(_04006_),
    .A1(_03682_));
 sg13g2_nor2_1 _10064_ (.A(_04010_),
    .B(_04011_),
    .Y(_04012_));
 sg13g2_nand2_1 _10065_ (.Y(_04013_),
    .A(_04011_),
    .B(_04010_));
 sg13g2_inv_1 _10066_ (.Y(_04014_),
    .A(_04013_));
 sg13g2_nor2_1 _10067_ (.A(_04012_),
    .B(_04014_),
    .Y(_04015_));
 sg13g2_inv_1 _10068_ (.Y(_04016_),
    .A(_04015_));
 sg13g2_nor2_1 _10069_ (.A(_03788_),
    .B(_03794_),
    .Y(_04017_));
 sg13g2_a21oi_1 _10070_ (.A1(_03797_),
    .A2(_03795_),
    .Y(_04018_),
    .B1(_04017_));
 sg13g2_xnor2_1 _10071_ (.Y(_04019_),
    .A(_04016_),
    .B(_04018_));
 sg13g2_nor2_1 _10072_ (.A(net66),
    .B(_04019_),
    .Y(_04021_));
 sg13g2_xor2_1 _10073_ (.B(_04021_),
    .A(_04004_),
    .X(_04022_));
 sg13g2_nand3_1 _10074_ (.B(_03676_),
    .C(_03778_),
    .A(_03660_),
    .Y(_04023_));
 sg13g2_nand2_1 _10075_ (.Y(_04024_),
    .A(_03671_),
    .B(_03778_));
 sg13g2_nand4_1 _10076_ (.B(_03771_),
    .C(_03777_),
    .A(_04023_),
    .Y(_04025_),
    .D(_04024_));
 sg13g2_nand2_1 _10077_ (.Y(_04026_),
    .A(_04025_),
    .B(net48));
 sg13g2_nand3_1 _10078_ (.B(_03678_),
    .C(_03299_),
    .A(_03677_),
    .Y(_04027_));
 sg13g2_nand2_1 _10079_ (.Y(_04028_),
    .A(_04026_),
    .B(_04027_));
 sg13g2_xnor2_1 _10080_ (.Y(_04029_),
    .A(_04022_),
    .B(_04028_));
 sg13g2_o21ai_1 _10081_ (.B1(_03831_),
    .Y(_04030_),
    .A1(_03819_),
    .A2(_03827_));
 sg13g2_a21oi_1 _10082_ (.A1(_03824_),
    .A2(_03820_),
    .Y(_04032_),
    .B1(_03823_));
 sg13g2_nor2_1 _10083_ (.A(_02783_),
    .B(_04019_),
    .Y(_04033_));
 sg13g2_a22oi_1 _10084_ (.Y(_04034_),
    .B1(_03312_),
    .B2(_03821_),
    .A2(_03815_),
    .A1(_03309_));
 sg13g2_xor2_1 _10085_ (.B(_04034_),
    .A(_04033_),
    .X(_04035_));
 sg13g2_xnor2_1 _10086_ (.Y(_04036_),
    .A(_04032_),
    .B(_04035_));
 sg13g2_nand2b_1 _10087_ (.Y(_04037_),
    .B(_04036_),
    .A_N(_04030_));
 sg13g2_nand2b_1 _10088_ (.Y(_04038_),
    .B(_04030_),
    .A_N(_04036_));
 sg13g2_nand3_1 _10089_ (.B(_03367_),
    .C(_04038_),
    .A(_04037_),
    .Y(_04039_));
 sg13g2_and2_1 _10090_ (.A(_03810_),
    .B(_03802_),
    .X(_04040_));
 sg13g2_xnor2_1 _10091_ (.Y(_04041_),
    .A(_04039_),
    .B(_04040_));
 sg13g2_xor2_1 _10092_ (.B(_04041_),
    .A(_04029_),
    .X(_04043_));
 sg13g2_inv_1 _10093_ (.Y(_04044_),
    .A(_03811_));
 sg13g2_a21oi_1 _10094_ (.A1(_03813_),
    .A2(_03833_),
    .Y(_04045_),
    .B1(_04044_));
 sg13g2_nand2b_1 _10095_ (.Y(_04046_),
    .B(_04045_),
    .A_N(_04043_));
 sg13g2_nand2b_1 _10096_ (.Y(_04047_),
    .B(_04043_),
    .A_N(_04045_));
 sg13g2_nand2_1 _10097_ (.Y(_04048_),
    .A(_02773_),
    .B(_02597_));
 sg13g2_o21ai_1 _10098_ (.B1(_05512_),
    .Y(_04049_),
    .A1(_04048_),
    .A2(_03726_));
 sg13g2_xnor2_1 _10099_ (.Y(_04050_),
    .A(net125),
    .B(_04049_));
 sg13g2_nor2_1 _10100_ (.A(net66),
    .B(_04050_),
    .Y(_04051_));
 sg13g2_a21oi_1 _10101_ (.A1(_04046_),
    .A2(_04047_),
    .Y(_04052_),
    .B1(_04051_));
 sg13g2_nand3_1 _10102_ (.B(_04047_),
    .C(_04051_),
    .A(_04046_),
    .Y(_04054_));
 sg13g2_nand2b_1 _10103_ (.Y(_04055_),
    .B(_04054_),
    .A_N(_04052_));
 sg13g2_xnor2_1 _10104_ (.Y(_04056_),
    .A(_03995_),
    .B(_04055_));
 sg13g2_inv_1 _10105_ (.Y(_04057_),
    .A(_04056_));
 sg13g2_nand2_1 _10106_ (.Y(_04058_),
    .A(_03993_),
    .B(_04057_));
 sg13g2_nand3_1 _10107_ (.B(_03992_),
    .C(_04056_),
    .A(_03948_),
    .Y(_04059_));
 sg13g2_a21oi_1 _10108_ (.A1(_05543_),
    .A2(_03208_),
    .Y(_04060_),
    .B1(_03213_));
 sg13g2_buf_8 _10109_ (.A(_04060_),
    .X(_04061_));
 sg13g2_nand3_1 _10110_ (.B(_04059_),
    .C(net55),
    .A(_04058_),
    .Y(_04062_));
 sg13g2_nor2_1 _10111_ (.A(_04807_),
    .B(_03603_),
    .Y(_04063_));
 sg13g2_nor2_1 _10112_ (.A(_04374_),
    .B(_03350_),
    .Y(_04064_));
 sg13g2_nor2_1 _10113_ (.A(_04335_),
    .B(_03332_),
    .Y(_04065_));
 sg13g2_nor2_1 _10114_ (.A(_04065_),
    .B(_01099_),
    .Y(_04066_));
 sg13g2_xnor2_1 _10115_ (.Y(_04067_),
    .A(_04065_),
    .B(_01099_));
 sg13g2_nand3_1 _10116_ (.B(_02477_),
    .C(_03955_),
    .A(_01005_),
    .Y(_04068_));
 sg13g2_nor3_1 _10117_ (.A(_00061_),
    .B(_03308_),
    .C(_01226_),
    .Y(_04069_));
 sg13g2_inv_1 _10118_ (.Y(_04070_),
    .A(_04069_));
 sg13g2_a21oi_1 _10119_ (.A1(_02477_),
    .A2(_03955_),
    .Y(_04071_),
    .B1(_01005_));
 sg13g2_a21oi_1 _10120_ (.A1(_04068_),
    .A2(_04070_),
    .Y(_04072_),
    .B1(_04071_));
 sg13g2_nor2_1 _10121_ (.A(_04067_),
    .B(_04072_),
    .Y(_04073_));
 sg13g2_xor2_1 _10122_ (.B(_01204_),
    .A(_04064_),
    .X(_04074_));
 sg13g2_o21ai_1 _10123_ (.B1(_04074_),
    .Y(_04075_),
    .A1(_04066_),
    .A2(_04073_));
 sg13g2_o21ai_1 _10124_ (.B1(_04075_),
    .Y(_04076_),
    .A1(_01204_),
    .A2(_04064_));
 sg13g2_nand2_1 _10125_ (.Y(_04077_),
    .A(_03385_),
    .B(_02444_));
 sg13g2_xnor2_1 _10126_ (.Y(_04078_),
    .A(_04077_),
    .B(_01299_));
 sg13g2_nor2b_1 _10127_ (.A(_01299_),
    .B_N(_04077_),
    .Y(_04079_));
 sg13g2_a21o_1 _10128_ (.A2(_04078_),
    .A1(_04076_),
    .B1(_04079_),
    .X(_04080_));
 sg13g2_xor2_1 _10129_ (.B(_01398_),
    .A(_04063_),
    .X(_04081_));
 sg13g2_nand2_1 _10130_ (.Y(_04082_),
    .A(_04080_),
    .B(_04081_));
 sg13g2_o21ai_1 _10131_ (.B1(_04082_),
    .Y(_04083_),
    .A1(_01398_),
    .A2(_04063_));
 sg13g2_nor2_1 _10132_ (.A(_04514_),
    .B(_03729_),
    .Y(_04084_));
 sg13g2_xor2_1 _10133_ (.B(_01652_),
    .A(_04084_),
    .X(_04085_));
 sg13g2_nor2_1 _10134_ (.A(_04084_),
    .B(_01652_),
    .Y(_04086_));
 sg13g2_a21oi_1 _10135_ (.A1(_04083_),
    .A2(_04085_),
    .Y(_04087_),
    .B1(_04086_));
 sg13g2_a21oi_1 _10136_ (.A1(_04087_),
    .A2(_01649_),
    .Y(_04088_),
    .B1(_04061_));
 sg13g2_o21ai_1 _10137_ (.B1(_04088_),
    .Y(_04089_),
    .A1(_01649_),
    .A2(_04087_));
 sg13g2_nand2_2 _10138_ (.Y(_04090_),
    .A(_04062_),
    .B(_04089_));
 sg13g2_nand2_1 _10139_ (.Y(_04091_),
    .A(_03939_),
    .B(_03933_));
 sg13g2_a21oi_1 _10140_ (.A1(_04091_),
    .A2(_03985_),
    .Y(_04092_),
    .B1(_03940_));
 sg13g2_nand2_1 _10141_ (.Y(_04093_),
    .A(_03735_),
    .B(_03609_));
 sg13g2_nand3_1 _10142_ (.B(_03733_),
    .C(_03607_),
    .A(_03732_),
    .Y(_04094_));
 sg13g2_nand2_1 _10143_ (.Y(_04095_),
    .A(_04093_),
    .B(_04094_));
 sg13g2_nand2b_1 _10144_ (.Y(_04096_),
    .B(_03870_),
    .A_N(_03900_));
 sg13g2_nand3_1 _10145_ (.B(_03869_),
    .C(_03900_),
    .A(_03867_),
    .Y(_04097_));
 sg13g2_nand2_1 _10146_ (.Y(_04098_),
    .A(_04096_),
    .B(_04097_));
 sg13g2_nand2_1 _10147_ (.Y(_04099_),
    .A(_04095_),
    .B(_04098_));
 sg13g2_nor2_1 _10148_ (.A(_04092_),
    .B(_04099_),
    .Y(_04100_));
 sg13g2_a21oi_1 _10149_ (.A1(_03736_),
    .A2(_03941_),
    .Y(_04101_),
    .B1(_03945_));
 sg13g2_nor2b_1 _10150_ (.A(_04100_),
    .B_N(_04101_),
    .Y(_04102_));
 sg13g2_nor2_1 _10151_ (.A(_03990_),
    .B(_03737_),
    .Y(_04103_));
 sg13g2_inv_1 _10152_ (.Y(_04104_),
    .A(_03983_));
 sg13g2_xnor2_1 _10153_ (.Y(_04105_),
    .A(_04104_),
    .B(_03981_));
 sg13g2_inv_1 _10154_ (.Y(_04106_),
    .A(_04105_));
 sg13g2_nor2_1 _10155_ (.A(_04106_),
    .B(_03989_),
    .Y(_04107_));
 sg13g2_nand3_1 _10156_ (.B(_03977_),
    .C(_04107_),
    .A(_04103_),
    .Y(_04108_));
 sg13g2_nand2_1 _10157_ (.Y(_04109_),
    .A(_04102_),
    .B(_04108_));
 sg13g2_nand2_1 _10158_ (.Y(_04110_),
    .A(_04109_),
    .B(_03861_));
 sg13g2_inv_1 _10159_ (.Y(_04111_),
    .A(_03861_));
 sg13g2_nand3_1 _10160_ (.B(_04108_),
    .C(_04111_),
    .A(_04102_),
    .Y(_04112_));
 sg13g2_nand3_1 _10161_ (.B(_04112_),
    .C(net55),
    .A(_04110_),
    .Y(_04113_));
 sg13g2_xor2_1 _10162_ (.B(_04083_),
    .A(_04085_),
    .X(_04115_));
 sg13g2_inv_4 _10163_ (.A(_04061_),
    .Y(_04116_));
 sg13g2_nand2b_1 _10164_ (.Y(_04117_),
    .B(_04116_),
    .A_N(_04115_));
 sg13g2_nand2_1 _10165_ (.Y(_04118_),
    .A(_04113_),
    .B(_04117_));
 sg13g2_buf_8 _10166_ (.A(_04118_),
    .X(_04119_));
 sg13g2_xnor2_1 _10167_ (.Y(_04120_),
    .A(net113),
    .B(_05247_));
 sg13g2_inv_1 _10168_ (.Y(_04121_),
    .A(_04120_));
 sg13g2_nor2_1 _10169_ (.A(_02828_),
    .B(_05243_),
    .Y(_04122_));
 sg13g2_inv_1 _10170_ (.Y(_04123_),
    .A(_04122_));
 sg13g2_nand2_1 _10171_ (.Y(_04124_),
    .A(net114),
    .B(_05243_));
 sg13g2_nand2_1 _10172_ (.Y(_04126_),
    .A(_04123_),
    .B(_04124_));
 sg13g2_inv_1 _10173_ (.Y(_04127_),
    .A(_04126_));
 sg13g2_nor2_1 _10174_ (.A(_05201_),
    .B(_03314_),
    .Y(_04128_));
 sg13g2_nand2_1 _10175_ (.Y(_04129_),
    .A(_03314_),
    .B(_05201_));
 sg13g2_inv_1 _10176_ (.Y(_04130_),
    .A(_04129_));
 sg13g2_nor2_1 _10177_ (.A(_04128_),
    .B(_04130_),
    .Y(_04131_));
 sg13g2_xor2_1 _10178_ (.B(_04684_),
    .A(net124),
    .X(_04132_));
 sg13g2_inv_1 _10179_ (.Y(_04133_),
    .A(_04132_));
 sg13g2_inv_1 _10180_ (.Y(_04134_),
    .A(_05239_));
 sg13g2_nor2_1 _10181_ (.A(net103),
    .B(_04134_),
    .Y(_04135_));
 sg13g2_nor2_1 _10182_ (.A(_05239_),
    .B(net112),
    .Y(_04137_));
 sg13g2_nor2_1 _10183_ (.A(_04135_),
    .B(_04137_),
    .Y(_04138_));
 sg13g2_nor2_1 _10184_ (.A(\title_r_pixels_in_scanline[2] ),
    .B(_02970_),
    .Y(_04139_));
 sg13g2_nor2_1 _10185_ (.A(net122),
    .B(_05236_),
    .Y(_04140_));
 sg13g2_nor2_1 _10186_ (.A(_04139_),
    .B(_04140_),
    .Y(_04141_));
 sg13g2_nand4_1 _10187_ (.B(_04133_),
    .C(_04138_),
    .A(_04131_),
    .Y(_04142_),
    .D(_04141_));
 sg13g2_nor4_1 _10188_ (.A(net116),
    .B(_04121_),
    .C(_04127_),
    .D(_04142_),
    .Y(_04143_));
 sg13g2_a21oi_1 _10189_ (.A1(_05244_),
    .A2(net114),
    .Y(_04144_),
    .B1(_05552_));
 sg13g2_nand2_1 _10190_ (.Y(_04145_),
    .A(_04144_),
    .B(_04120_));
 sg13g2_a21oi_1 _10191_ (.A1(net124),
    .A2(_04694_),
    .Y(_04146_),
    .B1(_04128_));
 sg13g2_nor3_1 _10192_ (.A(_04130_),
    .B(_04140_),
    .C(_04146_),
    .Y(_04148_));
 sg13g2_nor3_1 _10193_ (.A(_04137_),
    .B(_04139_),
    .C(_04148_),
    .Y(_04149_));
 sg13g2_a221oi_1 _10194_ (.B2(_05239_),
    .C1(_04149_),
    .B1(net112),
    .A1(_02729_),
    .Y(_04150_),
    .A2(_05243_));
 sg13g2_nand3_1 _10195_ (.B(_05262_),
    .C(_05247_),
    .A(_02751_),
    .Y(_04151_));
 sg13g2_o21ai_1 _10196_ (.B1(_04151_),
    .Y(_04152_),
    .A1(_04145_),
    .A2(_04150_));
 sg13g2_nor2b_1 _10197_ (.A(_04143_),
    .B_N(_04152_),
    .Y(_04153_));
 sg13g2_nand3_1 _10198_ (.B(net125),
    .C(_02806_),
    .A(_02773_),
    .Y(_04154_));
 sg13g2_nand2b_1 _10199_ (.Y(_04155_),
    .B(_02400_),
    .A_N(_04154_));
 sg13g2_nand2_1 _10200_ (.Y(_04156_),
    .A(_04787_),
    .B(_02806_));
 sg13g2_nand4_1 _10201_ (.B(_05504_),
    .C(_04155_),
    .A(_04153_),
    .Y(_04157_),
    .D(_04156_));
 sg13g2_nand3_1 _10202_ (.B(_02608_),
    .C(_04123_),
    .A(_04121_),
    .Y(_04159_));
 sg13g2_a21oi_1 _10203_ (.A1(_04715_),
    .A2(_04694_),
    .Y(_04160_),
    .B1(_04131_));
 sg13g2_nand2_1 _10204_ (.Y(_04161_),
    .A(_02937_),
    .B(_05201_));
 sg13g2_nand2_1 _10205_ (.Y(_04162_),
    .A(net122),
    .B(\title_r_pixels_in_scanline[2] ));
 sg13g2_nand3b_1 _10206_ (.B(_04161_),
    .C(_04162_),
    .Y(_04163_),
    .A_N(_04160_));
 sg13g2_a22oi_1 _10207_ (.Y(_04164_),
    .B1(net112),
    .B2(_04134_),
    .A2(_05236_),
    .A1(_02970_));
 sg13g2_o21ai_1 _10208_ (.B1(_04124_),
    .Y(_04165_),
    .A1(net112),
    .A2(_04134_));
 sg13g2_a21oi_1 _10209_ (.A1(_04163_),
    .A2(_04164_),
    .Y(_04166_),
    .B1(_04165_));
 sg13g2_nand3_1 _10210_ (.B(net113),
    .C(_05247_),
    .A(_05552_),
    .Y(_04167_));
 sg13g2_o21ai_1 _10211_ (.B1(_04167_),
    .Y(_04168_),
    .A1(_04159_),
    .A2(_04166_));
 sg13g2_nor3_1 _10212_ (.A(_02411_),
    .B(_05503_),
    .C(_04154_),
    .Y(_04170_));
 sg13g2_nor4_1 _10213_ (.A(_04138_),
    .B(_04141_),
    .C(_04131_),
    .D(_04133_),
    .Y(_04171_));
 sg13g2_nand4_1 _10214_ (.B(_05552_),
    .C(_04121_),
    .A(_04171_),
    .Y(_04172_),
    .D(_04127_));
 sg13g2_nand3_1 _10215_ (.B(_04170_),
    .C(_04172_),
    .A(_04168_),
    .Y(_04173_));
 sg13g2_o21ai_1 _10216_ (.B1(_00022_),
    .Y(_04174_),
    .A1(_02411_),
    .A2(_04525_));
 sg13g2_o21ai_1 _10217_ (.B1(_05552_),
    .Y(_04175_),
    .A1(_05546_),
    .A2(_04048_));
 sg13g2_nor3_1 _10218_ (.A(_02817_),
    .B(_05503_),
    .C(_04175_),
    .Y(_04176_));
 sg13g2_a21oi_1 _10219_ (.A1(_03102_),
    .A2(net127),
    .Y(_04177_),
    .B1(net129));
 sg13g2_nand2_1 _10220_ (.Y(_04178_),
    .A(_03157_),
    .B(_04177_));
 sg13g2_nand3_1 _10221_ (.B(_04176_),
    .C(_04178_),
    .A(_04174_),
    .Y(_04179_));
 sg13g2_nand3_1 _10222_ (.B(_04173_),
    .C(_04179_),
    .A(_04157_),
    .Y(_04181_));
 sg13g2_nand3b_1 _10223_ (.B(_00204_),
    .C(net86),
    .Y(_04182_),
    .A_N(_00189_));
 sg13g2_nand3_1 _10224_ (.B(_03309_),
    .C(_04182_),
    .A(_04181_),
    .Y(_04183_));
 sg13g2_nand4_1 _10225_ (.B(net17),
    .C(_03221_),
    .A(_04090_),
    .Y(_04184_),
    .D(_04183_));
 sg13g2_inv_2 _10226_ (.Y(_04185_),
    .A(_03363_));
 sg13g2_nor3_1 _10227_ (.A(_05542_),
    .B(_03207_),
    .C(_05543_),
    .Y(_04186_));
 sg13g2_inv_1 _10228_ (.Y(_04187_),
    .A(_04186_));
 sg13g2_nand2_1 _10229_ (.Y(_04188_),
    .A(_04090_),
    .B(_04187_));
 sg13g2_nand3_1 _10230_ (.B(_04185_),
    .C(_04188_),
    .A(_04184_),
    .Y(_04189_));
 sg13g2_a21oi_1 _10231_ (.A1(_03991_),
    .A2(_03988_),
    .Y(_04190_),
    .B1(_03944_));
 sg13g2_xnor2_1 _10232_ (.Y(_04192_),
    .A(_03737_),
    .B(_04190_));
 sg13g2_xnor2_1 _10233_ (.Y(_04193_),
    .A(_04081_),
    .B(_04080_));
 sg13g2_nand2b_1 _10234_ (.Y(_04194_),
    .B(_04116_),
    .A_N(_04193_));
 sg13g2_o21ai_1 _10235_ (.B1(_04194_),
    .Y(_04195_),
    .A1(_04116_),
    .A2(_04192_));
 sg13g2_buf_1 _10236_ (.A(_04195_),
    .X(_04196_));
 sg13g2_nor2_1 _10237_ (.A(_03989_),
    .B(_03986_),
    .Y(_04197_));
 sg13g2_nor3_1 _10238_ (.A(_03940_),
    .B(_04098_),
    .C(_04197_),
    .Y(_04198_));
 sg13g2_o21ai_1 _10239_ (.B1(_04098_),
    .Y(_04199_),
    .A1(_03940_),
    .A2(_04197_));
 sg13g2_nand2_1 _10240_ (.Y(_04200_),
    .A(_04199_),
    .B(net55));
 sg13g2_a21oi_1 _10241_ (.A1(_04076_),
    .A2(_04078_),
    .Y(_04201_),
    .B1(net55));
 sg13g2_o21ai_1 _10242_ (.B1(_04201_),
    .Y(_04203_),
    .A1(_04078_),
    .A2(_04076_));
 sg13g2_o21ai_1 _10243_ (.B1(_04203_),
    .Y(_04204_),
    .A1(_04198_),
    .A2(_04200_));
 sg13g2_buf_8 _10244_ (.A(_04204_),
    .X(_04205_));
 sg13g2_nand2_1 _10245_ (.Y(_04206_),
    .A(_04196_),
    .B(_04205_));
 sg13g2_nor3_1 _10246_ (.A(_04185_),
    .B(net17),
    .C(_04206_),
    .Y(_04207_));
 sg13g2_a21oi_1 _10247_ (.A1(_05529_),
    .A2(_00036_),
    .Y(_04208_),
    .B1(_04207_));
 sg13g2_nand2_1 _10248_ (.Y(_04209_),
    .A(_04189_),
    .B(_04208_));
 sg13g2_nor3_2 _10249_ (.A(_05542_),
    .B(_03207_),
    .C(_05530_),
    .Y(_04210_));
 sg13g2_inv_1 _10250_ (.Y(_04211_),
    .A(_04210_));
 sg13g2_nand2_1 _10251_ (.Y(_04212_),
    .A(_04090_),
    .B(_04118_));
 sg13g2_nor2_1 _10252_ (.A(_04211_),
    .B(_04212_),
    .Y(_04214_));
 sg13g2_nor2_1 _10253_ (.A(_05530_),
    .B(_03225_),
    .Y(_04215_));
 sg13g2_nor2_1 _10254_ (.A(_05533_),
    .B(_04215_),
    .Y(_04216_));
 sg13g2_nand2b_1 _10255_ (.Y(_04217_),
    .B(_04068_),
    .A_N(_04071_));
 sg13g2_xnor2_1 _10256_ (.Y(_04218_),
    .A(_04070_),
    .B(_04217_));
 sg13g2_nand2_1 _10257_ (.Y(_04219_),
    .A(_03975_),
    .B(_03969_));
 sg13g2_nor2_1 _10258_ (.A(_04116_),
    .B(_03977_),
    .Y(_04220_));
 sg13g2_a22oi_1 _10259_ (.Y(_04221_),
    .B1(_04219_),
    .B2(_04220_),
    .A2(_04218_),
    .A1(_04116_));
 sg13g2_nand2_1 _10260_ (.Y(_04222_),
    .A(_04072_),
    .B(_04067_));
 sg13g2_nor2_1 _10261_ (.A(net55),
    .B(_04073_),
    .Y(_04223_));
 sg13g2_xor2_1 _10262_ (.B(_04105_),
    .A(_03977_),
    .X(_04225_));
 sg13g2_a22oi_1 _10263_ (.Y(_04226_),
    .B1(net55),
    .B2(_04225_),
    .A2(_04223_),
    .A1(_04222_));
 sg13g2_nor3_1 _10264_ (.A(_04074_),
    .B(_04066_),
    .C(_04073_),
    .Y(_04227_));
 sg13g2_nor2b_1 _10265_ (.A(_04227_),
    .B_N(_04075_),
    .Y(_04228_));
 sg13g2_nand2_1 _10266_ (.Y(_04229_),
    .A(_03986_),
    .B(_03989_));
 sg13g2_nor2_1 _10267_ (.A(_04116_),
    .B(_04197_),
    .Y(_04230_));
 sg13g2_a22oi_1 _10268_ (.Y(_04231_),
    .B1(_04229_),
    .B2(_04230_),
    .A2(_04228_),
    .A1(_04116_));
 sg13g2_nor2_1 _10269_ (.A(_04226_),
    .B(_04231_),
    .Y(_04232_));
 sg13g2_nand3_1 _10270_ (.B(_04205_),
    .C(_04232_),
    .A(_04196_),
    .Y(_04233_));
 sg13g2_nor3_1 _10271_ (.A(_05533_),
    .B(_04221_),
    .C(_04233_),
    .Y(_04234_));
 sg13g2_nor2_1 _10272_ (.A(_04216_),
    .B(_04234_),
    .Y(_04236_));
 sg13g2_nor2_1 _10273_ (.A(_04214_),
    .B(_04236_),
    .Y(_04237_));
 sg13g2_nand2_1 _10274_ (.Y(_04238_),
    .A(_04209_),
    .B(_04237_));
 sg13g2_nor2_1 _10275_ (.A(_04231_),
    .B(_04206_),
    .Y(_04239_));
 sg13g2_o21ai_1 _10276_ (.B1(_05533_),
    .Y(_04240_),
    .A1(_04181_),
    .A2(_04239_));
 sg13g2_buf_1 _10277_ (.A(_04240_),
    .X(_04241_));
 sg13g2_nand2_2 _10278_ (.Y(_04242_),
    .A(_04836_),
    .B(_02882_));
 sg13g2_a21oi_1 _10279_ (.A1(_04238_),
    .A2(_04241_),
    .Y(_00065_),
    .B1(_04242_));
 sg13g2_o21ai_1 _10280_ (.B1(_04185_),
    .Y(_04243_),
    .A1(_03207_),
    .A2(_05530_));
 sg13g2_inv_1 _10281_ (.Y(_04244_),
    .A(net17));
 sg13g2_nand2_1 _10282_ (.Y(_04246_),
    .A(_04183_),
    .B(_04186_));
 sg13g2_inv_1 _10283_ (.Y(_04247_),
    .A(_04246_));
 sg13g2_nor2_1 _10284_ (.A(_03213_),
    .B(_04247_),
    .Y(_04248_));
 sg13g2_a22oi_1 _10285_ (.Y(_04249_),
    .B1(_04248_),
    .B2(_04188_),
    .A2(_03213_),
    .A1(_04244_));
 sg13g2_nor2_1 _10286_ (.A(net17),
    .B(_04206_),
    .Y(_04250_));
 sg13g2_o21ai_1 _10287_ (.B1(_01226_),
    .Y(_04251_),
    .A1(_00061_),
    .A2(_03308_));
 sg13g2_nor2_1 _10288_ (.A(net55),
    .B(_04069_),
    .Y(_04252_));
 sg13g2_nor2b_1 _10289_ (.A(_03974_),
    .B_N(_03972_),
    .Y(_04253_));
 sg13g2_xnor2_1 _10290_ (.Y(_04254_),
    .A(_03973_),
    .B(_04253_));
 sg13g2_a22oi_1 _10291_ (.Y(_04255_),
    .B1(net55),
    .B2(_04254_),
    .A2(_04252_),
    .A1(_04251_));
 sg13g2_nand2_1 _10292_ (.Y(_04257_),
    .A(_04255_),
    .B(_04215_));
 sg13g2_nor2_1 _10293_ (.A(_04221_),
    .B(_04257_),
    .Y(_04258_));
 sg13g2_nand3_1 _10294_ (.B(_04232_),
    .C(_04258_),
    .A(_04250_),
    .Y(_04259_));
 sg13g2_o21ai_1 _10295_ (.B1(_04259_),
    .Y(_04260_),
    .A1(_04243_),
    .A2(_04249_));
 sg13g2_inv_1 _10296_ (.Y(_04261_),
    .A(_05533_));
 sg13g2_nand2_1 _10297_ (.Y(_04262_),
    .A(_04260_),
    .B(_04261_));
 sg13g2_a21oi_1 _10298_ (.A1(_04262_),
    .A2(_04241_),
    .Y(_00066_),
    .B1(_04242_));
 sg13g2_nand2_1 _10299_ (.Y(_04263_),
    .A(_04212_),
    .B(_02102_));
 sg13g2_nand3_1 _10300_ (.B(net17),
    .C(_04196_),
    .A(_04090_),
    .Y(_04264_));
 sg13g2_nand3_1 _10301_ (.B(_04264_),
    .C(_04247_),
    .A(_04263_),
    .Y(_04265_));
 sg13g2_nand2_1 _10302_ (.Y(_04267_),
    .A(_03783_),
    .B(_03785_));
 sg13g2_nor2_1 _10303_ (.A(_04267_),
    .B(_04188_),
    .Y(_04268_));
 sg13g2_nor2_1 _10304_ (.A(_03209_),
    .B(_04268_),
    .Y(_04269_));
 sg13g2_nand2_1 _10305_ (.Y(_04270_),
    .A(_04265_),
    .B(_04269_));
 sg13g2_nand2_1 _10306_ (.Y(_04271_),
    .A(_02193_),
    .B(_03363_));
 sg13g2_nor4_1 _10307_ (.A(_04231_),
    .B(_04271_),
    .C(_04119_),
    .D(_04206_),
    .Y(_04272_));
 sg13g2_a21oi_1 _10308_ (.A1(_04196_),
    .A2(_03213_),
    .Y(_04273_),
    .B1(_04210_));
 sg13g2_nor2b_1 _10309_ (.A(_04272_),
    .B_N(_04273_),
    .Y(_04274_));
 sg13g2_nand2_1 _10310_ (.Y(_04275_),
    .A(_04270_),
    .B(_04274_));
 sg13g2_a21oi_1 _10311_ (.A1(_04090_),
    .A2(_04119_),
    .Y(_04276_),
    .B1(_02204_));
 sg13g2_nor2b_1 _10312_ (.A(_04276_),
    .B_N(_04264_),
    .Y(_04277_));
 sg13g2_inv_1 _10313_ (.Y(_04278_),
    .A(_04216_));
 sg13g2_a21oi_1 _10314_ (.A1(_04277_),
    .A2(_04210_),
    .Y(_04279_),
    .B1(_04278_));
 sg13g2_nand2_1 _10315_ (.Y(_04280_),
    .A(_04275_),
    .B(_04279_));
 sg13g2_a21oi_1 _10316_ (.A1(_04280_),
    .A2(_04241_),
    .Y(_00067_),
    .B1(_04242_));
 sg13g2_buf_1 _10317_ (.A(_02882_),
    .X(_04281_));
 sg13g2_buf_2 _10318_ (.A(\hvsync_gen.vsync ),
    .X(_04282_));
 sg13g2_buf_1 _10319_ (.A(_04282_),
    .X(_04283_));
 sg13g2_buf_1 _10320_ (.A(net99),
    .X(_04284_));
 sg13g2_nand2_1 _10321_ (.Y(_04285_),
    .A(net117),
    .B(net84));
 sg13g2_inv_1 _10322_ (.Y(_00068_),
    .A(_04285_));
 sg13g2_nand2_1 _10323_ (.Y(_04287_),
    .A(net17),
    .B(_04187_));
 sg13g2_nand3_1 _10324_ (.B(_04185_),
    .C(_04287_),
    .A(_04184_),
    .Y(_04288_));
 sg13g2_nor2_1 _10325_ (.A(_04210_),
    .B(_04207_),
    .Y(_04289_));
 sg13g2_nand2_1 _10326_ (.Y(_04290_),
    .A(_04288_),
    .B(_04289_));
 sg13g2_nor2_1 _10327_ (.A(_04278_),
    .B(_04214_),
    .Y(_04291_));
 sg13g2_nand2_1 _10328_ (.Y(_04292_),
    .A(_04290_),
    .B(_04291_));
 sg13g2_nor2_1 _10329_ (.A(_04257_),
    .B(_04233_),
    .Y(_04293_));
 sg13g2_nor2b_1 _10330_ (.A(_04293_),
    .B_N(_04241_),
    .Y(_04294_));
 sg13g2_a21oi_1 _10331_ (.A1(_04292_),
    .A2(_04294_),
    .Y(_00069_),
    .B1(_04242_));
 sg13g2_a22oi_1 _10332_ (.Y(_04296_),
    .B1(_04248_),
    .B2(_04287_),
    .A2(_04196_),
    .A1(_03213_));
 sg13g2_o21ai_1 _10333_ (.B1(_04259_),
    .Y(_04297_),
    .A1(_04243_),
    .A2(_04296_));
 sg13g2_nand2_1 _10334_ (.Y(_04298_),
    .A(_04297_),
    .B(_04261_));
 sg13g2_a21oi_1 _10335_ (.A1(_04298_),
    .A2(_04241_),
    .Y(_00070_),
    .B1(_04242_));
 sg13g2_nand3_1 _10336_ (.B(_03681_),
    .C(_04187_),
    .A(net17),
    .Y(_04299_));
 sg13g2_nand2_1 _10337_ (.Y(_04300_),
    .A(_04299_),
    .B(_03210_));
 sg13g2_a21oi_1 _10338_ (.A1(_04205_),
    .A2(_03213_),
    .Y(_04301_),
    .B1(_04210_));
 sg13g2_a21oi_1 _10339_ (.A1(_04300_),
    .A2(_04301_),
    .Y(_04302_),
    .B1(_04278_));
 sg13g2_a22oi_1 _10340_ (.Y(_04303_),
    .B1(_01976_),
    .B2(_04212_),
    .A2(_04246_),
    .A1(_04211_));
 sg13g2_nand3_1 _10341_ (.B(net17),
    .C(_04205_),
    .A(_04090_),
    .Y(_04304_));
 sg13g2_nand2_1 _10342_ (.Y(_04306_),
    .A(_04303_),
    .B(_04304_));
 sg13g2_nand2_1 _10343_ (.Y(_04307_),
    .A(_04302_),
    .B(_04306_));
 sg13g2_a21oi_1 _10344_ (.A1(_04307_),
    .A2(_04241_),
    .Y(_00071_),
    .B1(_04242_));
 sg13g2_nand2_1 _10345_ (.Y(_04308_),
    .A(net117),
    .B(hsync));
 sg13g2_inv_1 _10346_ (.Y(_00072_),
    .A(_04308_));
 sg13g2_nor3_1 _10347_ (.A(_05490_),
    .B(_05489_),
    .C(net47),
    .Y(_04309_));
 sg13g2_a21oi_1 _10348_ (.A1(_03355_),
    .A2(_03311_),
    .Y(_04310_),
    .B1(net108));
 sg13g2_nor3_1 _10349_ (.A(net96),
    .B(_04309_),
    .C(_04310_),
    .Y(_00073_));
 sg13g2_nor2_1 _10350_ (.A(net98),
    .B(_04309_),
    .Y(_04311_));
 sg13g2_nand2_1 _10351_ (.Y(_04312_),
    .A(_04309_),
    .B(_03256_));
 sg13g2_inv_1 _10352_ (.Y(_04314_),
    .A(_04312_));
 sg13g2_nor3_1 _10353_ (.A(net96),
    .B(_04311_),
    .C(_04314_),
    .Y(_00074_));
 sg13g2_nor2_1 _10354_ (.A(_05495_),
    .B(_04312_),
    .Y(_04315_));
 sg13g2_nor2_1 _10355_ (.A(_03278_),
    .B(_04314_),
    .Y(_04316_));
 sg13g2_nor3_1 _10356_ (.A(net96),
    .B(_04315_),
    .C(_04316_),
    .Y(_00075_));
 sg13g2_a21oi_1 _10357_ (.A1(net93),
    .A2(net47),
    .Y(_04317_),
    .B1(_03575_));
 sg13g2_nor2_1 _10358_ (.A(net94),
    .B(_04317_),
    .Y(_00076_));
 sg13g2_a21oi_1 _10359_ (.A1(net106),
    .A2(net47),
    .Y(_04318_),
    .B1(_03377_));
 sg13g2_nor2_1 _10360_ (.A(net94),
    .B(_04318_),
    .Y(_00077_));
 sg13g2_a21oi_1 _10361_ (.A1(net100),
    .A2(net47),
    .Y(_04319_),
    .B1(_03476_));
 sg13g2_nor2_1 _10362_ (.A(net94),
    .B(_04319_),
    .Y(_00078_));
 sg13g2_nand2_1 _10363_ (.Y(_04321_),
    .A(net47),
    .B(net118));
 sg13g2_a21oi_1 _10364_ (.A1(_03717_),
    .A2(_04321_),
    .Y(_00079_),
    .B1(net94));
 sg13g2_nand2_1 _10365_ (.Y(_04322_),
    .A(net47),
    .B(_05529_));
 sg13g2_buf_1 _10366_ (.A(net105),
    .X(_04323_));
 sg13g2_a21oi_1 _10367_ (.A1(_04009_),
    .A2(_04322_),
    .Y(_00080_),
    .B1(net83));
 sg13g2_nor2_1 _10368_ (.A(_03207_),
    .B(_03987_),
    .Y(_04324_));
 sg13g2_a21oi_1 _10369_ (.A1(_03355_),
    .A2(_04324_),
    .Y(_04325_),
    .B1(_05528_));
 sg13g2_nor4_1 _10370_ (.A(_05542_),
    .B(_03207_),
    .C(_03987_),
    .D(net47),
    .Y(_04326_));
 sg13g2_nor3_1 _10371_ (.A(net96),
    .B(_04325_),
    .C(_04326_),
    .Y(_00081_));
 sg13g2_xnor2_1 _10372_ (.Y(_04327_),
    .A(\frame_counter[9] ),
    .B(_04326_));
 sg13g2_nor2_1 _10373_ (.A(net94),
    .B(_04327_),
    .Y(_00082_));
 sg13g2_o21ai_1 _10374_ (.B1(net117),
    .Y(_04328_),
    .A1(\envelopeA[0] ),
    .A2(_03553_));
 sg13g2_a21oi_1 _10375_ (.A1(_05489_),
    .A2(_03553_),
    .Y(_00083_),
    .B1(_04328_));
 sg13g2_nor2_1 _10376_ (.A(\noise_counter[1] ),
    .B(\noise_counter[2] ),
    .Y(_04329_));
 sg13g2_xnor2_1 _10377_ (.Y(_04330_),
    .A(_01636_),
    .B(_01747_));
 sg13g2_xnor2_1 _10378_ (.Y(_04331_),
    .A(_05569_),
    .B(_05574_));
 sg13g2_xor2_1 _10379_ (.B(_05587_),
    .A(_00250_),
    .X(_04332_));
 sg13g2_xnor2_1 _10380_ (.Y(_04333_),
    .A(_04331_),
    .B(_04332_));
 sg13g2_xnor2_1 _10381_ (.Y(_04334_),
    .A(_00346_),
    .B(_00292_));
 sg13g2_xnor2_1 _10382_ (.Y(_04336_),
    .A(_00668_),
    .B(_00382_));
 sg13g2_xnor2_1 _10383_ (.Y(_04337_),
    .A(_04334_),
    .B(_04336_));
 sg13g2_xnor2_1 _10384_ (.Y(_04338_),
    .A(_04333_),
    .B(_04337_));
 sg13g2_buf_1 _10385_ (.A(\r1[9] ),
    .X(_04339_));
 sg13g2_xnor2_1 _10386_ (.Y(_04340_),
    .A(_00672_),
    .B(_04339_));
 sg13g2_nand2_1 _10387_ (.Y(_04341_),
    .A(_01070_),
    .B(\r1[10] ));
 sg13g2_nand2_1 _10388_ (.Y(_04342_),
    .A(_01072_),
    .B(_04341_));
 sg13g2_xnor2_1 _10389_ (.Y(_04343_),
    .A(_04340_),
    .B(_04342_));
 sg13g2_nand2_1 _10390_ (.Y(_04344_),
    .A(_01380_),
    .B(_01525_));
 sg13g2_inv_1 _10391_ (.Y(_04345_),
    .A(_04344_));
 sg13g2_nor2_1 _10392_ (.A(_01635_),
    .B(_04345_),
    .Y(_04347_));
 sg13g2_nand2_1 _10393_ (.Y(_04348_),
    .A(\r1[13] ),
    .B(_01179_));
 sg13g2_nor2b_1 _10394_ (.A(_01285_),
    .B_N(_04348_),
    .Y(_04349_));
 sg13g2_xnor2_1 _10395_ (.Y(_04350_),
    .A(_04347_),
    .B(_04349_));
 sg13g2_xnor2_1 _10396_ (.Y(_04351_),
    .A(_04343_),
    .B(_04350_));
 sg13g2_xnor2_1 _10397_ (.Y(_04352_),
    .A(_04338_),
    .B(_04351_));
 sg13g2_xnor2_1 _10398_ (.Y(_04353_),
    .A(_04330_),
    .B(_04352_));
 sg13g2_buf_1 _10399_ (.A(_03058_),
    .X(_04354_));
 sg13g2_nand3b_1 _10400_ (.B(_04353_),
    .C(net54),
    .Y(_04355_),
    .A_N(_04329_));
 sg13g2_o21ai_1 _10401_ (.B1(_04281_),
    .Y(_04356_),
    .A1(_05524_),
    .A2(_04355_));
 sg13g2_a21oi_1 _10402_ (.A1(_05524_),
    .A2(_04355_),
    .Y(_00104_),
    .B1(_04356_));
 sg13g2_nand2b_1 _10403_ (.Y(_04358_),
    .B(_04329_),
    .A_N(\noise_counter[0] ));
 sg13g2_o21ai_1 _10404_ (.B1(net117),
    .Y(_04359_),
    .A1(\noise_counter[0] ),
    .A2(net54));
 sg13g2_a21oi_1 _10405_ (.A1(net54),
    .A2(_04358_),
    .Y(_00105_),
    .B1(_04359_));
 sg13g2_nand3_1 _10406_ (.B(\noise_counter[0] ),
    .C(_04329_),
    .A(net54),
    .Y(_04360_));
 sg13g2_inv_1 _10407_ (.Y(_04361_),
    .A(_03058_));
 sg13g2_nand2_1 _10408_ (.Y(_04362_),
    .A(net53),
    .B(\noise_counter[1] ));
 sg13g2_a21oi_1 _10409_ (.A1(_04360_),
    .A2(_04362_),
    .Y(_00106_),
    .B1(net83));
 sg13g2_and3_1 _10410_ (.X(_00107_),
    .A(net53),
    .B(net117),
    .C(\noise_counter[2] ));
 sg13g2_inv_1 _10411_ (.Y(_04363_),
    .A(\note_counter[7] ));
 sg13g2_inv_1 _10412_ (.Y(_04364_),
    .A(\note_freq[7] ));
 sg13g2_inv_1 _10413_ (.Y(_04365_),
    .A(\note_freq[6] ));
 sg13g2_a22oi_1 _10414_ (.Y(_04366_),
    .B1(\note_counter[6] ),
    .B2(_04365_),
    .A2(\note_counter[7] ),
    .A1(_04364_));
 sg13g2_inv_1 _10415_ (.Y(_04367_),
    .A(\note_freq[4] ));
 sg13g2_nor2_1 _10416_ (.A(\note_counter[4] ),
    .B(_04367_),
    .Y(_04368_));
 sg13g2_inv_1 _10417_ (.Y(_04369_),
    .A(\note_freq[2] ));
 sg13g2_nor2_1 _10418_ (.A(\note_counter[2] ),
    .B(_04369_),
    .Y(_04370_));
 sg13g2_buf_1 _10419_ (.A(\note_freq[1] ),
    .X(_04371_));
 sg13g2_inv_1 _10420_ (.Y(_04372_),
    .A(_04371_));
 sg13g2_inv_1 _10421_ (.Y(_04373_),
    .A(\note_counter[0] ));
 sg13g2_nor2_1 _10422_ (.A(\note_freq[0] ),
    .B(_04373_),
    .Y(_04375_));
 sg13g2_inv_1 _10423_ (.Y(_04376_),
    .A(\note_counter[3] ));
 sg13g2_inv_1 _10424_ (.Y(_04377_),
    .A(\note_counter[1] ));
 sg13g2_o21ai_1 _10425_ (.B1(_04371_),
    .Y(_04378_),
    .A1(_04376_),
    .A2(_04377_));
 sg13g2_a22oi_1 _10426_ (.Y(_04379_),
    .B1(_04375_),
    .B2(_04378_),
    .A2(\note_counter[1] ),
    .A1(_04372_));
 sg13g2_nand2_1 _10427_ (.Y(_04380_),
    .A(_04376_),
    .B(_04371_));
 sg13g2_nand2_1 _10428_ (.Y(_04381_),
    .A(_04369_),
    .B(\note_counter[2] ));
 sg13g2_o21ai_1 _10429_ (.B1(_04381_),
    .Y(_04382_),
    .A1(_04376_),
    .A2(_04371_));
 sg13g2_a22oi_1 _10430_ (.Y(_04383_),
    .B1(_04380_),
    .B2(_04382_),
    .A2(\note_counter[4] ),
    .A1(_04367_));
 sg13g2_o21ai_1 _10431_ (.B1(_04383_),
    .Y(_04384_),
    .A1(_04370_),
    .A2(_04379_));
 sg13g2_buf_1 _10432_ (.A(\note_counter[5] ),
    .X(_04386_));
 sg13g2_nand2b_1 _10433_ (.Y(_04387_),
    .B(\note_freq[5] ),
    .A_N(_04386_));
 sg13g2_nand3b_1 _10434_ (.B(_04384_),
    .C(_04387_),
    .Y(_04388_),
    .A_N(_04368_));
 sg13g2_nand2b_1 _10435_ (.Y(_04389_),
    .B(_04386_),
    .A_N(\note_freq[5] ));
 sg13g2_nand2_1 _10436_ (.Y(_04390_),
    .A(_04388_),
    .B(_04389_));
 sg13g2_o21ai_1 _10437_ (.B1(_04390_),
    .Y(_04391_),
    .A1(\note_counter[6] ),
    .A2(_04365_));
 sg13g2_a22oi_1 _10438_ (.Y(_04392_),
    .B1(_04366_),
    .B2(_04391_),
    .A2(_04363_),
    .A1(\note_freq[7] ));
 sg13g2_nand2_1 _10439_ (.Y(_04393_),
    .A(_04392_),
    .B(net54));
 sg13g2_o21ai_1 _10440_ (.B1(net117),
    .Y(_04394_),
    .A1(_00058_),
    .A2(_04393_));
 sg13g2_a21oi_1 _10441_ (.A1(_05547_),
    .A2(_04393_),
    .Y(_00108_),
    .B1(_04394_));
 sg13g2_inv_1 _10442_ (.Y(_04396_),
    .A(note2));
 sg13g2_inv_1 _10443_ (.Y(_04397_),
    .A(\note2_counter[8] ));
 sg13g2_nor2_1 _10444_ (.A(\note2_freq[8] ),
    .B(_04397_),
    .Y(_04398_));
 sg13g2_inv_1 _10445_ (.Y(_04399_),
    .A(\note2_counter[7] ));
 sg13g2_nor2_1 _10446_ (.A(\note2_freq[7] ),
    .B(_04399_),
    .Y(_04400_));
 sg13g2_nand2_1 _10447_ (.Y(_04401_),
    .A(_04399_),
    .B(\note2_freq[7] ));
 sg13g2_inv_1 _10448_ (.Y(_04402_),
    .A(_04401_));
 sg13g2_nand2_1 _10449_ (.Y(_04403_),
    .A(_04397_),
    .B(\note2_freq[8] ));
 sg13g2_inv_1 _10450_ (.Y(_04404_),
    .A(_04403_));
 sg13g2_nor4_1 _10451_ (.A(_04398_),
    .B(_04400_),
    .C(_04402_),
    .D(_04404_),
    .Y(_04405_));
 sg13g2_inv_1 _10452_ (.Y(_04407_),
    .A(\note2_counter[5] ));
 sg13g2_nand2_1 _10453_ (.Y(_04408_),
    .A(_04407_),
    .B(\note2_freq[5] ));
 sg13g2_inv_1 _10454_ (.Y(_04409_),
    .A(\note2_counter[6] ));
 sg13g2_nor2_1 _10455_ (.A(\note2_freq[6] ),
    .B(_04409_),
    .Y(_04410_));
 sg13g2_nand2_1 _10456_ (.Y(_04411_),
    .A(_04409_),
    .B(\note2_freq[6] ));
 sg13g2_o21ai_1 _10457_ (.B1(_04411_),
    .Y(_04412_),
    .A1(_04408_),
    .A2(_04410_));
 sg13g2_inv_1 _10458_ (.Y(_04413_),
    .A(\note2_counter[2] ));
 sg13g2_inv_1 _10459_ (.Y(_04414_),
    .A(\note2_counter[1] ));
 sg13g2_nand2_1 _10460_ (.Y(_04415_),
    .A(_04414_),
    .B(\note2_freq[1] ));
 sg13g2_inv_1 _10461_ (.Y(_04416_),
    .A(_04415_));
 sg13g2_nor2b_1 _10462_ (.A(\note2_counter[3] ),
    .B_N(\note2_freq[3] ),
    .Y(_04418_));
 sg13g2_inv_1 _10463_ (.Y(_04419_),
    .A(\note2_counter[3] ));
 sg13g2_nor2_1 _10464_ (.A(\note2_freq[3] ),
    .B(_04419_),
    .Y(_04420_));
 sg13g2_buf_1 _10465_ (.A(\note2_counter[4] ),
    .X(_04421_));
 sg13g2_xnor2_1 _10466_ (.Y(_04422_),
    .A(_04421_),
    .B(\note2_freq[4] ));
 sg13g2_inv_1 _10467_ (.Y(_04423_),
    .A(_04422_));
 sg13g2_nor3_1 _10468_ (.A(_04418_),
    .B(_04420_),
    .C(_04423_),
    .Y(_04424_));
 sg13g2_o21ai_1 _10469_ (.B1(_04424_),
    .Y(_04425_),
    .A1(_04413_),
    .A2(_04416_));
 sg13g2_nor2b_1 _10470_ (.A(_04421_),
    .B_N(\note2_freq[4] ),
    .Y(_04426_));
 sg13g2_a21oi_1 _10471_ (.A1(_04422_),
    .A2(_04418_),
    .Y(_04427_),
    .B1(_04426_));
 sg13g2_nand2_1 _10472_ (.Y(_04429_),
    .A(_04425_),
    .B(_04427_));
 sg13g2_inv_1 _10473_ (.Y(_04430_),
    .A(_04410_));
 sg13g2_nand2b_1 _10474_ (.Y(_04431_),
    .B(\note2_counter[5] ),
    .A_N(\note2_freq[5] ));
 sg13g2_nand4_1 _10475_ (.B(_04431_),
    .C(_04411_),
    .A(_04430_),
    .Y(_04432_),
    .D(_04408_));
 sg13g2_nor2b_1 _10476_ (.A(_04432_),
    .B_N(_04405_),
    .Y(_04433_));
 sg13g2_o21ai_1 _10477_ (.B1(_04403_),
    .Y(_04434_),
    .A1(_04401_),
    .A2(_04398_));
 sg13g2_a221oi_1 _10478_ (.B2(_04433_),
    .C1(_04434_),
    .B1(_04429_),
    .A1(_04405_),
    .Y(_04435_),
    .A2(_04412_));
 sg13g2_buf_1 _10479_ (.A(\note2_counter[0] ),
    .X(_04436_));
 sg13g2_nand2b_1 _10480_ (.Y(_04437_),
    .B(_04436_),
    .A_N(\note2_freq[0] ));
 sg13g2_nor2_1 _10481_ (.A(\note2_freq[1] ),
    .B(_04414_),
    .Y(_04438_));
 sg13g2_nor3_1 _10482_ (.A(_04413_),
    .B(_04438_),
    .C(_04416_),
    .Y(_04439_));
 sg13g2_nand4_1 _10483_ (.B(_04437_),
    .C(_04424_),
    .A(_04433_),
    .Y(_04440_),
    .D(_04439_));
 sg13g2_nand3_1 _10484_ (.B(net54),
    .C(_04440_),
    .A(_04435_),
    .Y(_04441_));
 sg13g2_buf_1 _10485_ (.A(_04441_),
    .X(_04442_));
 sg13g2_o21ai_1 _10486_ (.B1(_04281_),
    .Y(_04443_),
    .A1(_00059_),
    .A2(_04442_));
 sg13g2_a21oi_1 _10487_ (.A1(_04396_),
    .A2(_04442_),
    .Y(_00109_),
    .B1(_04443_));
 sg13g2_a21oi_1 _10488_ (.A1(_04435_),
    .A2(_04440_),
    .Y(_04444_),
    .B1(net53));
 sg13g2_o21ai_1 _10489_ (.B1(net117),
    .Y(_04445_),
    .A1(_04436_),
    .A2(_04444_));
 sg13g2_a21oi_1 _10490_ (.A1(_04436_),
    .A2(_04354_),
    .Y(_00110_),
    .B1(_04445_));
 sg13g2_buf_1 _10491_ (.A(net105),
    .X(_04446_));
 sg13g2_a21oi_1 _10492_ (.A1(_04354_),
    .A2(_04436_),
    .Y(_04448_),
    .B1(\note2_counter[1] ));
 sg13g2_nand2_1 _10493_ (.Y(_04449_),
    .A(\note2_counter[1] ),
    .B(_04436_));
 sg13g2_nor2_1 _10494_ (.A(_04449_),
    .B(_04361_),
    .Y(_04450_));
 sg13g2_inv_2 _10495_ (.Y(_04451_),
    .A(_04442_));
 sg13g2_nor4_1 _10496_ (.A(net82),
    .B(_04448_),
    .C(_04450_),
    .D(_04451_),
    .Y(_00111_));
 sg13g2_nor2_1 _10497_ (.A(\note2_counter[2] ),
    .B(_04450_),
    .Y(_04452_));
 sg13g2_inv_1 _10498_ (.Y(_04453_),
    .A(_04436_));
 sg13g2_nor4_2 _10499_ (.A(_04414_),
    .B(_04413_),
    .C(_04453_),
    .Y(_04454_),
    .D(_04361_));
 sg13g2_nor4_1 _10500_ (.A(net82),
    .B(_04452_),
    .C(_04454_),
    .D(_04451_),
    .Y(_00112_));
 sg13g2_nor2_1 _10501_ (.A(\note2_counter[3] ),
    .B(_04454_),
    .Y(_04455_));
 sg13g2_nor2b_1 _10502_ (.A(_04419_),
    .B_N(_04454_),
    .Y(_04457_));
 sg13g2_nor4_1 _10503_ (.A(net82),
    .B(_04455_),
    .C(_04457_),
    .D(_04451_),
    .Y(_00113_));
 sg13g2_nor2_1 _10504_ (.A(_04421_),
    .B(_04457_),
    .Y(_04458_));
 sg13g2_nand2_1 _10505_ (.Y(_04459_),
    .A(_04457_),
    .B(_04421_));
 sg13g2_inv_1 _10506_ (.Y(_04460_),
    .A(_04459_));
 sg13g2_nor4_1 _10507_ (.A(net82),
    .B(_04458_),
    .C(_04460_),
    .D(_04451_),
    .Y(_00114_));
 sg13g2_nor2_1 _10508_ (.A(_04407_),
    .B(_04459_),
    .Y(_04461_));
 sg13g2_nor2_1 _10509_ (.A(\note2_counter[5] ),
    .B(_04460_),
    .Y(_04462_));
 sg13g2_nor4_1 _10510_ (.A(_04446_),
    .B(_04461_),
    .C(_04451_),
    .D(_04462_),
    .Y(_00115_));
 sg13g2_inv_1 _10511_ (.Y(_04463_),
    .A(_04421_));
 sg13g2_nor2_1 _10512_ (.A(_04413_),
    .B(_04449_),
    .Y(_04464_));
 sg13g2_nand3_1 _10513_ (.B(\note2_counter[3] ),
    .C(_04464_),
    .A(_03058_),
    .Y(_04465_));
 sg13g2_nor4_1 _10514_ (.A(_04409_),
    .B(_04407_),
    .C(_04463_),
    .D(_04465_),
    .Y(_04466_));
 sg13g2_inv_1 _10515_ (.Y(_04467_),
    .A(_04466_));
 sg13g2_o21ai_1 _10516_ (.B1(_04467_),
    .Y(_04468_),
    .A1(\note2_counter[6] ),
    .A2(_04461_));
 sg13g2_nor3_1 _10517_ (.A(net96),
    .B(_04451_),
    .C(_04468_),
    .Y(_00116_));
 sg13g2_nor2_1 _10518_ (.A(\note2_counter[7] ),
    .B(_04466_),
    .Y(_04469_));
 sg13g2_nor2_1 _10519_ (.A(_04399_),
    .B(_04467_),
    .Y(_04470_));
 sg13g2_nor4_1 _10520_ (.A(_04446_),
    .B(_04469_),
    .C(_04470_),
    .D(_04451_),
    .Y(_00117_));
 sg13g2_xnor2_1 _10521_ (.Y(_04471_),
    .A(\note2_counter[8] ),
    .B(_04470_));
 sg13g2_nor3_1 _10522_ (.A(net96),
    .B(_04451_),
    .C(_04471_),
    .Y(_00118_));
 sg13g2_nand2_1 _10523_ (.Y(_00119_),
    .A(_04042_),
    .B(_00002_));
 sg13g2_nor3_1 _10524_ (.A(\note_counter[0] ),
    .B(net53),
    .C(_04392_),
    .Y(_04473_));
 sg13g2_a21oi_1 _10525_ (.A1(\note_counter[0] ),
    .A2(net53),
    .Y(_04474_),
    .B1(_04473_));
 sg13g2_nor2_1 _10526_ (.A(net94),
    .B(_04474_),
    .Y(_00122_));
 sg13g2_o21ai_1 _10527_ (.B1(_04377_),
    .Y(_04475_),
    .A1(_04373_),
    .A2(net53));
 sg13g2_nand2_1 _10528_ (.Y(_04476_),
    .A(\note_counter[1] ),
    .B(\note_counter[0] ));
 sg13g2_nand2b_1 _10529_ (.Y(_04477_),
    .B(net54),
    .A_N(_04476_));
 sg13g2_nand3_1 _10530_ (.B(net130),
    .C(_04477_),
    .A(_04475_),
    .Y(_04478_));
 sg13g2_inv_1 _10531_ (.Y(_04479_),
    .A(_04393_));
 sg13g2_nor2_1 _10532_ (.A(_04478_),
    .B(_04479_),
    .Y(_00123_));
 sg13g2_inv_1 _10533_ (.Y(_04481_),
    .A(\note_counter[2] ));
 sg13g2_xnor2_1 _10534_ (.Y(_04482_),
    .A(_04481_),
    .B(_04477_));
 sg13g2_nor3_1 _10535_ (.A(net82),
    .B(_04482_),
    .C(_04479_),
    .Y(_00124_));
 sg13g2_nor2_1 _10536_ (.A(_04481_),
    .B(_04476_),
    .Y(_04483_));
 sg13g2_a21oi_1 _10537_ (.A1(net54),
    .A2(_04483_),
    .Y(_04484_),
    .B1(\note_counter[3] ));
 sg13g2_inv_1 _10538_ (.Y(_04485_),
    .A(_04483_));
 sg13g2_nor3_1 _10539_ (.A(_04376_),
    .B(_04485_),
    .C(net53),
    .Y(_04486_));
 sg13g2_nor4_1 _10540_ (.A(net82),
    .B(_04484_),
    .C(_04486_),
    .D(_04479_),
    .Y(_00125_));
 sg13g2_nor2_1 _10541_ (.A(\note_counter[4] ),
    .B(_04486_),
    .Y(_04487_));
 sg13g2_and2_1 _10542_ (.A(_04486_),
    .B(\note_counter[4] ),
    .X(_04489_));
 sg13g2_buf_1 _10543_ (.A(_04489_),
    .X(_04490_));
 sg13g2_nor4_1 _10544_ (.A(net105),
    .B(_04487_),
    .C(_04490_),
    .D(_04479_),
    .Y(_00126_));
 sg13g2_xnor2_1 _10545_ (.Y(_04491_),
    .A(_04386_),
    .B(_04490_));
 sg13g2_nor3_1 _10546_ (.A(net82),
    .B(_04491_),
    .C(_04479_),
    .Y(_00127_));
 sg13g2_a21oi_1 _10547_ (.A1(_04490_),
    .A2(_04386_),
    .Y(_04492_),
    .B1(\note_counter[6] ));
 sg13g2_and3_1 _10548_ (.X(_04493_),
    .A(_04490_),
    .B(\note_counter[6] ),
    .C(_04386_));
 sg13g2_nor4_1 _10549_ (.A(net105),
    .B(_04492_),
    .C(_04493_),
    .D(_04479_),
    .Y(_00128_));
 sg13g2_xnor2_1 _10550_ (.Y(_04494_),
    .A(\note_counter[7] ),
    .B(_04493_));
 sg13g2_nor3_1 _10551_ (.A(net82),
    .B(_04494_),
    .C(_04479_),
    .Y(_00129_));
 sg13g2_nand2_1 _10552_ (.Y(_00130_),
    .A(_03868_),
    .B(_03793_));
 sg13g2_nand2_1 _10553_ (.Y(_00131_),
    .A(_03846_),
    .B(_03772_));
 sg13g2_inv_1 _10554_ (.Y(_04495_),
    .A(_00031_));
 sg13g2_nor2_1 _10555_ (.A(_04846_),
    .B(net53),
    .Y(_04496_));
 sg13g2_buf_1 _10556_ (.A(_04496_),
    .X(_04497_));
 sg13g2_inv_2 _10557_ (.Y(_04498_),
    .A(_04497_));
 sg13g2_nor2_2 _10558_ (.A(_03179_),
    .B(_04498_),
    .Y(_04499_));
 sg13g2_nor2_1 _10559_ (.A(net113),
    .B(net56),
    .Y(_04500_));
 sg13g2_a22oi_1 _10560_ (.Y(_04501_),
    .B1(net112),
    .B2(net93),
    .A2(_03278_),
    .A1(_02970_));
 sg13g2_xnor2_1 _10561_ (.Y(_04502_),
    .A(net113),
    .B(net61));
 sg13g2_xor2_1 _10562_ (.B(_03443_),
    .A(net114),
    .X(_04504_));
 sg13g2_nand2_1 _10563_ (.Y(_04505_),
    .A(_04502_),
    .B(_04504_));
 sg13g2_inv_1 _10564_ (.Y(_04506_),
    .A(_04505_));
 sg13g2_nand2_1 _10565_ (.Y(_04507_),
    .A(net111),
    .B(_04147_));
 sg13g2_nand3b_1 _10566_ (.B(_04506_),
    .C(_04507_),
    .Y(_04508_),
    .A_N(_04501_));
 sg13g2_nand3_1 _10567_ (.B(net115),
    .C(_02737_),
    .A(_04502_),
    .Y(_04509_));
 sg13g2_nand3b_1 _10568_ (.B(_04508_),
    .C(_04509_),
    .Y(_04510_),
    .A_N(_04500_));
 sg13g2_xnor2_1 _10569_ (.Y(_04511_),
    .A(net126),
    .B(_00228_));
 sg13g2_nor2_1 _10570_ (.A(_00021_),
    .B(_03789_),
    .Y(_04512_));
 sg13g2_nor2_1 _10571_ (.A(_05552_),
    .B(_03790_),
    .Y(_04513_));
 sg13g2_nor3_1 _10572_ (.A(_04511_),
    .B(_04512_),
    .C(_04513_),
    .Y(_04515_));
 sg13g2_nor2_1 _10573_ (.A(_00022_),
    .B(net74),
    .Y(_04516_));
 sg13g2_inv_1 _10574_ (.Y(_04517_),
    .A(net74));
 sg13g2_nor2b_1 _10575_ (.A(_04517_),
    .B_N(_00022_),
    .Y(_04518_));
 sg13g2_nor3_1 _10576_ (.A(_02817_),
    .B(_04516_),
    .C(_04518_),
    .Y(_04519_));
 sg13g2_and2_1 _10577_ (.A(_04515_),
    .B(_04519_),
    .X(_04520_));
 sg13g2_nand2_1 _10578_ (.Y(_04521_),
    .A(_04510_),
    .B(_04520_));
 sg13g2_nand2b_1 _10579_ (.Y(_04522_),
    .B(_04513_),
    .A_N(_04511_));
 sg13g2_o21ai_1 _10580_ (.B1(_04522_),
    .Y(_04523_),
    .A1(_05513_),
    .A2(_00228_));
 sg13g2_a22oi_1 _10581_ (.Y(_04524_),
    .B1(_04519_),
    .B2(_04523_),
    .A2(_00432_),
    .A1(_03014_));
 sg13g2_a22oi_1 _10582_ (.Y(_04526_),
    .B1(_02926_),
    .B2(_05490_),
    .A2(net123),
    .A1(_05486_));
 sg13g2_nand2_1 _10583_ (.Y(_04527_),
    .A(_03314_),
    .B(_03256_));
 sg13g2_nand2b_1 _10584_ (.Y(_04528_),
    .B(_04527_),
    .A_N(_04526_));
 sg13g2_nand2_1 _10585_ (.Y(_04529_),
    .A(_05495_),
    .B(_02959_));
 sg13g2_nand3_1 _10586_ (.B(_04507_),
    .C(_04529_),
    .A(_04501_),
    .Y(_04530_));
 sg13g2_nor2_1 _10587_ (.A(_04530_),
    .B(_04505_),
    .Y(_04531_));
 sg13g2_nand3_1 _10588_ (.B(_04528_),
    .C(_04531_),
    .A(_04520_),
    .Y(_04532_));
 sg13g2_nand3_1 _10589_ (.B(_04524_),
    .C(_04532_),
    .A(_04521_),
    .Y(_04533_));
 sg13g2_nand2_1 _10590_ (.Y(_04534_),
    .A(_04715_),
    .B(net108));
 sg13g2_nand3_1 _10591_ (.B(_04527_),
    .C(_04534_),
    .A(_04526_),
    .Y(_04535_));
 sg13g2_nor2_1 _10592_ (.A(_04530_),
    .B(_04535_),
    .Y(_04537_));
 sg13g2_nand4_1 _10593_ (.B(_04506_),
    .C(_04519_),
    .A(_04515_),
    .Y(_04538_),
    .D(_04537_));
 sg13g2_nand2_1 _10594_ (.Y(_04539_),
    .A(_04533_),
    .B(_04538_));
 sg13g2_buf_2 _10595_ (.A(_04539_),
    .X(_04540_));
 sg13g2_inv_1 _10596_ (.Y(_04541_),
    .A(_04540_));
 sg13g2_buf_1 _10597_ (.A(_04541_),
    .X(_04542_));
 sg13g2_nand2_1 _10598_ (.Y(_04543_),
    .A(_03300_),
    .B(_05574_));
 sg13g2_inv_1 _10599_ (.Y(_04544_),
    .A(_05574_));
 sg13g2_nand2_1 _10600_ (.Y(_04545_),
    .A(_05490_),
    .B(_04544_));
 sg13g2_nand3_1 _10601_ (.B(_04543_),
    .C(_04545_),
    .A(_04542_),
    .Y(_04546_));
 sg13g2_buf_1 _10602_ (.A(_04540_),
    .X(_04548_));
 sg13g2_nor2_1 _10603_ (.A(_04284_),
    .B(_04544_),
    .Y(_04549_));
 sg13g2_nand2_1 _10604_ (.Y(_04550_),
    .A(_04836_),
    .B(_03179_));
 sg13g2_buf_1 _10605_ (.A(_04550_),
    .X(_04551_));
 sg13g2_buf_1 _10606_ (.A(_04551_),
    .X(_04552_));
 sg13g2_a21oi_1 _10607_ (.A1(_04548_),
    .A2(_04549_),
    .Y(_04553_),
    .B1(_04552_));
 sg13g2_inv_1 _10608_ (.Y(_04554_),
    .A(_04551_));
 sg13g2_buf_1 _10609_ (.A(_04554_),
    .X(_04555_));
 sg13g2_nor2_1 _10610_ (.A(_04555_),
    .B(_04497_),
    .Y(_04556_));
 sg13g2_buf_2 _10611_ (.A(_04556_),
    .X(_04557_));
 sg13g2_inv_1 _10612_ (.Y(_04559_),
    .A(_04557_));
 sg13g2_o21ai_1 _10613_ (.B1(net130),
    .Y(_04560_),
    .A1(_04549_),
    .A2(_04559_));
 sg13g2_a221oi_1 _10614_ (.B2(_04553_),
    .C1(_04560_),
    .B1(_04546_),
    .A1(_04495_),
    .Y(_00132_),
    .A2(_04499_));
 sg13g2_nand2_1 _10615_ (.Y(_04561_),
    .A(_03474_),
    .B(_03069_));
 sg13g2_xnor2_1 _10616_ (.Y(_04562_),
    .A(_02543_),
    .B(_04561_));
 sg13g2_nand2_1 _10617_ (.Y(_04563_),
    .A(_03474_),
    .B(_00025_));
 sg13g2_xnor2_1 _10618_ (.Y(_04564_),
    .A(_02389_),
    .B(_04563_));
 sg13g2_nand2_1 _10619_ (.Y(_04565_),
    .A(_04564_),
    .B(_04517_));
 sg13g2_o21ai_1 _10620_ (.B1(_04565_),
    .Y(_04566_),
    .A1(_00025_),
    .A2(_04561_));
 sg13g2_xor2_1 _10621_ (.B(_04566_),
    .A(_04562_),
    .X(_04567_));
 sg13g2_inv_1 _10622_ (.Y(_04568_),
    .A(_04018_));
 sg13g2_a21oi_1 _10623_ (.A1(_04568_),
    .A2(_04013_),
    .Y(_04569_),
    .B1(_04012_));
 sg13g2_nand2_1 _10624_ (.Y(_04570_),
    .A(_04007_),
    .B(_00228_));
 sg13g2_o21ai_1 _10625_ (.B1(_04570_),
    .Y(_04571_),
    .A1(_00023_),
    .A2(_04563_));
 sg13g2_xnor2_1 _10626_ (.Y(_04572_),
    .A(_00432_),
    .B(_04564_));
 sg13g2_nand2_1 _10627_ (.Y(_04573_),
    .A(_04571_),
    .B(_04572_));
 sg13g2_nor2_1 _10628_ (.A(_04572_),
    .B(_04571_),
    .Y(_04574_));
 sg13g2_a21oi_1 _10629_ (.A1(_04569_),
    .A2(_04573_),
    .Y(_04575_),
    .B1(_04574_));
 sg13g2_or2_1 _10630_ (.X(_04576_),
    .B(_04575_),
    .A(_04567_));
 sg13g2_nand2_1 _10631_ (.Y(_04577_),
    .A(_04575_),
    .B(_04567_));
 sg13g2_nand2_1 _10632_ (.Y(_04579_),
    .A(_04576_),
    .B(_04577_));
 sg13g2_buf_1 _10633_ (.A(_04579_),
    .X(_04580_));
 sg13g2_xnor2_1 _10634_ (.Y(_04581_),
    .A(_00978_),
    .B(net21));
 sg13g2_nor2b_1 _10635_ (.A(_04574_),
    .B_N(_04573_),
    .Y(_04582_));
 sg13g2_xnor2_1 _10636_ (.Y(_04583_),
    .A(_04582_),
    .B(_04569_));
 sg13g2_xor2_1 _10637_ (.B(_04583_),
    .A(_04339_),
    .X(_04584_));
 sg13g2_inv_1 _10638_ (.Y(_04585_),
    .A(_04584_));
 sg13g2_inv_1 _10639_ (.Y(_04586_),
    .A(_04019_));
 sg13g2_inv_1 _10640_ (.Y(_04587_),
    .A(_00672_));
 sg13g2_xnor2_1 _10641_ (.Y(_04588_),
    .A(_04587_),
    .B(_04019_));
 sg13g2_inv_1 _10642_ (.Y(_04590_),
    .A(_04588_));
 sg13g2_nor2_1 _10643_ (.A(_00044_),
    .B(_03800_),
    .Y(_04591_));
 sg13g2_xnor2_1 _10644_ (.Y(_04592_),
    .A(_00668_),
    .B(_03800_));
 sg13g2_inv_1 _10645_ (.Y(_04593_),
    .A(_04592_));
 sg13g2_inv_1 _10646_ (.Y(_04594_),
    .A(_00043_));
 sg13g2_inv_1 _10647_ (.Y(_04595_),
    .A(_00032_));
 sg13g2_inv_1 _10648_ (.Y(_04596_),
    .A(_03485_));
 sg13g2_nor2_1 _10649_ (.A(_00286_),
    .B(_03504_),
    .Y(_04597_));
 sg13g2_xnor2_1 _10650_ (.Y(_04598_),
    .A(_00286_),
    .B(_03504_));
 sg13g2_nor2_1 _10651_ (.A(_00253_),
    .B(_03501_),
    .Y(_04599_));
 sg13g2_nand2_1 _10652_ (.Y(_04601_),
    .A(_03519_),
    .B(_05589_));
 sg13g2_nor2_1 _10653_ (.A(_05589_),
    .B(_03519_),
    .Y(_04602_));
 sg13g2_a21oi_1 _10654_ (.A1(_04601_),
    .A2(_05574_),
    .Y(_04603_),
    .B1(_04602_));
 sg13g2_nand2_1 _10655_ (.Y(_04604_),
    .A(_03501_),
    .B(_00253_));
 sg13g2_nor2b_1 _10656_ (.A(_04599_),
    .B_N(_04604_),
    .Y(_04605_));
 sg13g2_nor2b_1 _10657_ (.A(_04603_),
    .B_N(_04605_),
    .Y(_04606_));
 sg13g2_nor2_1 _10658_ (.A(_04599_),
    .B(_04606_),
    .Y(_04607_));
 sg13g2_nor2_1 _10659_ (.A(_04598_),
    .B(_04607_),
    .Y(_04608_));
 sg13g2_nor2_1 _10660_ (.A(_04597_),
    .B(_04608_),
    .Y(_04609_));
 sg13g2_nor2_1 _10661_ (.A(_00340_),
    .B(_03275_),
    .Y(_04610_));
 sg13g2_inv_1 _10662_ (.Y(_04611_),
    .A(_04610_));
 sg13g2_nand2_1 _10663_ (.Y(_04612_),
    .A(_03275_),
    .B(_00340_));
 sg13g2_nand2_1 _10664_ (.Y(_04613_),
    .A(_04611_),
    .B(_04612_));
 sg13g2_or2_1 _10665_ (.X(_04614_),
    .B(_04613_),
    .A(_04609_));
 sg13g2_nand2_1 _10666_ (.Y(_04615_),
    .A(_04614_),
    .B(_04611_));
 sg13g2_inv_1 _10667_ (.Y(_04616_),
    .A(_04615_));
 sg13g2_xnor2_1 _10668_ (.Y(_04617_),
    .A(_00346_),
    .B(_03485_));
 sg13g2_inv_1 _10669_ (.Y(_04618_),
    .A(_04617_));
 sg13g2_nor2_1 _10670_ (.A(_04616_),
    .B(_04618_),
    .Y(_04619_));
 sg13g2_a21oi_1 _10671_ (.A1(_04595_),
    .A2(_04596_),
    .Y(_04620_),
    .B1(_04619_));
 sg13g2_xnor2_1 _10672_ (.Y(_04622_),
    .A(_00382_),
    .B(_03694_));
 sg13g2_inv_1 _10673_ (.Y(_04623_),
    .A(_04622_));
 sg13g2_nor2_1 _10674_ (.A(_04620_),
    .B(_04623_),
    .Y(_04624_));
 sg13g2_a21oi_1 _10675_ (.A1(_04594_),
    .A2(_03815_),
    .Y(_04625_),
    .B1(_04624_));
 sg13g2_nor2_1 _10676_ (.A(_04593_),
    .B(_04625_),
    .Y(_04626_));
 sg13g2_nor2_1 _10677_ (.A(_04591_),
    .B(_04626_),
    .Y(_04627_));
 sg13g2_inv_1 _10678_ (.Y(_04628_),
    .A(_04627_));
 sg13g2_a22oi_1 _10679_ (.Y(_04629_),
    .B1(_04590_),
    .B2(_04628_),
    .A2(_04586_),
    .A1(_00776_));
 sg13g2_nand2_1 _10680_ (.Y(_04630_),
    .A(_04583_),
    .B(_00784_));
 sg13g2_o21ai_1 _10681_ (.B1(_04630_),
    .Y(_04631_),
    .A1(_04585_),
    .A2(_04629_));
 sg13g2_inv_1 _10682_ (.Y(_04633_),
    .A(_04631_));
 sg13g2_nor2_1 _10683_ (.A(_04581_),
    .B(_04633_),
    .Y(_04634_));
 sg13g2_nand2_1 _10684_ (.Y(_04635_),
    .A(_04633_),
    .B(_04581_));
 sg13g2_nand3b_1 _10685_ (.B(_04499_),
    .C(_04635_),
    .Y(_04636_),
    .A_N(_04634_));
 sg13g2_nor2_1 _10686_ (.A(net99),
    .B(_00978_),
    .Y(_04637_));
 sg13g2_buf_1 _10687_ (.A(_04555_),
    .X(_04638_));
 sg13g2_buf_1 _10688_ (.A(_04540_),
    .X(_04639_));
 sg13g2_xnor2_1 _10689_ (.Y(_04640_),
    .A(_00672_),
    .B(net74));
 sg13g2_xnor2_1 _10690_ (.Y(_04641_),
    .A(_00430_),
    .B(_00228_));
 sg13g2_nor2_1 _10691_ (.A(_00043_),
    .B(_03790_),
    .Y(_04642_));
 sg13g2_inv_1 _10692_ (.Y(_04643_),
    .A(_00346_));
 sg13g2_xnor2_1 _10693_ (.Y(_04644_),
    .A(_04643_),
    .B(net61));
 sg13g2_nor2_1 _10694_ (.A(net106),
    .B(_00340_),
    .Y(_04645_));
 sg13g2_nor2_1 _10695_ (.A(_00292_),
    .B(net86),
    .Y(_04646_));
 sg13g2_xor2_1 _10696_ (.B(_05569_),
    .A(net98),
    .X(_04647_));
 sg13g2_inv_1 _10697_ (.Y(_04648_),
    .A(_04647_));
 sg13g2_nand2_1 _10698_ (.Y(_04649_),
    .A(net98),
    .B(_05569_));
 sg13g2_o21ai_1 _10699_ (.B1(_04649_),
    .Y(_04650_),
    .A1(_04543_),
    .A2(_04648_));
 sg13g2_xor2_1 _10700_ (.B(_05587_),
    .A(net109),
    .X(_04651_));
 sg13g2_and2_1 _10701_ (.A(_04650_),
    .B(_04651_),
    .X(_04652_));
 sg13g2_a21oi_1 _10702_ (.A1(net109),
    .A2(_05587_),
    .Y(_04654_),
    .B1(_04652_));
 sg13g2_nand2_1 _10703_ (.Y(_04655_),
    .A(net93),
    .B(_00250_));
 sg13g2_nor2_1 _10704_ (.A(net93),
    .B(_00250_),
    .Y(_04656_));
 sg13g2_a21oi_1 _10705_ (.A1(_04654_),
    .A2(_04655_),
    .Y(_04657_),
    .B1(_04656_));
 sg13g2_nand2b_1 _10706_ (.Y(_04658_),
    .B(_04657_),
    .A_N(_04646_));
 sg13g2_nand2b_1 _10707_ (.Y(_04659_),
    .B(_04658_),
    .A_N(_04645_));
 sg13g2_a22oi_1 _10708_ (.Y(_04660_),
    .B1(_04644_),
    .B2(_04659_),
    .A2(net61),
    .A1(_04595_));
 sg13g2_inv_1 _10709_ (.Y(_04661_),
    .A(_04641_));
 sg13g2_xnor2_1 _10710_ (.Y(_04662_),
    .A(_00383_),
    .B(_03789_));
 sg13g2_inv_1 _10711_ (.Y(_04663_),
    .A(_04662_));
 sg13g2_nor2_1 _10712_ (.A(_04661_),
    .B(_04663_),
    .Y(_04665_));
 sg13g2_nor2b_1 _10713_ (.A(_04660_),
    .B_N(_04665_),
    .Y(_04666_));
 sg13g2_a221oi_1 _10714_ (.B2(_04642_),
    .C1(_04666_),
    .B1(_04641_),
    .A1(_00668_),
    .Y(_04667_),
    .A2(_04005_));
 sg13g2_nor2_1 _10715_ (.A(_04640_),
    .B(_04667_),
    .Y(_04668_));
 sg13g2_a21oi_1 _10716_ (.A1(_00776_),
    .A2(net74),
    .Y(_04669_),
    .B1(_04668_));
 sg13g2_nor2_1 _10717_ (.A(_00040_),
    .B(_04669_),
    .Y(_04670_));
 sg13g2_xnor2_1 _10718_ (.Y(_04671_),
    .A(_00877_),
    .B(_04670_));
 sg13g2_nand2_1 _10719_ (.Y(_04672_),
    .A(net24),
    .B(_04637_));
 sg13g2_o21ai_1 _10720_ (.B1(_04672_),
    .Y(_04673_),
    .A1(net24),
    .A2(_04671_));
 sg13g2_a22oi_1 _10721_ (.Y(_04674_),
    .B1(net36),
    .B2(_04673_),
    .A2(_04637_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10722_ (.A1(_04636_),
    .A2(_04674_),
    .Y(_00133_),
    .B1(net83));
 sg13g2_inv_1 _10723_ (.Y(_04675_),
    .A(_01070_));
 sg13g2_xnor2_1 _10724_ (.Y(_04676_),
    .A(_04675_),
    .B(net21));
 sg13g2_inv_1 _10725_ (.Y(_04677_),
    .A(net21));
 sg13g2_a21oi_1 _10726_ (.A1(_00877_),
    .A2(_04677_),
    .Y(_04678_),
    .B1(_04634_));
 sg13g2_nor2_1 _10727_ (.A(_04676_),
    .B(_04678_),
    .Y(_04679_));
 sg13g2_nand2_1 _10728_ (.Y(_04680_),
    .A(_04678_),
    .B(_04676_));
 sg13g2_nand3b_1 _10729_ (.B(_04499_),
    .C(_04680_),
    .Y(_04681_),
    .A_N(_04679_));
 sg13g2_nor2_1 _10730_ (.A(net99),
    .B(_04675_),
    .Y(_04682_));
 sg13g2_inv_1 _10731_ (.Y(_04683_),
    .A(_04339_));
 sg13g2_nor3_1 _10732_ (.A(_00978_),
    .B(_04683_),
    .C(_04669_),
    .Y(_04685_));
 sg13g2_xnor2_1 _10733_ (.Y(_04686_),
    .A(_00983_),
    .B(_04685_));
 sg13g2_nand2_1 _10734_ (.Y(_04687_),
    .A(net24),
    .B(_04682_));
 sg13g2_o21ai_1 _10735_ (.B1(_04687_),
    .Y(_04688_),
    .A1(net24),
    .A2(_04686_));
 sg13g2_a22oi_1 _10736_ (.Y(_04689_),
    .B1(net36),
    .B2(_04688_),
    .A2(_04682_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10737_ (.A1(_04681_),
    .A2(_04689_),
    .Y(_00134_),
    .B1(net83));
 sg13g2_buf_1 _10738_ (.A(_04555_),
    .X(_04690_));
 sg13g2_buf_1 _10739_ (.A(net35),
    .X(_04691_));
 sg13g2_inv_1 _10740_ (.Y(_04692_),
    .A(_01179_));
 sg13g2_nor2_1 _10741_ (.A(net84),
    .B(_04692_),
    .Y(_04693_));
 sg13g2_inv_1 _10742_ (.Y(_04695_),
    .A(_04670_));
 sg13g2_nor2_1 _10743_ (.A(_04341_),
    .B(_04695_),
    .Y(_04696_));
 sg13g2_xnor2_1 _10744_ (.Y(_04697_),
    .A(_01077_),
    .B(_04696_));
 sg13g2_nor2_1 _10745_ (.A(net24),
    .B(_04697_),
    .Y(_04698_));
 sg13g2_a21oi_1 _10746_ (.A1(net25),
    .A2(_04693_),
    .Y(_04699_),
    .B1(_04698_));
 sg13g2_xnor2_1 _10747_ (.Y(_04700_),
    .A(_04692_),
    .B(net21));
 sg13g2_a21oi_1 _10748_ (.A1(_00983_),
    .A2(_04677_),
    .Y(_04701_),
    .B1(_04679_));
 sg13g2_nor2_1 _10749_ (.A(_04700_),
    .B(_04701_),
    .Y(_04702_));
 sg13g2_buf_1 _10750_ (.A(_04497_),
    .X(_04703_));
 sg13g2_nand2_1 _10751_ (.Y(_04704_),
    .A(_04701_),
    .B(_04700_));
 sg13g2_nand3b_1 _10752_ (.B(net39),
    .C(_04704_),
    .Y(_04706_),
    .A_N(_04702_));
 sg13g2_buf_1 _10753_ (.A(_04498_),
    .X(_04707_));
 sg13g2_buf_1 _10754_ (.A(_04555_),
    .X(_04708_));
 sg13g2_a21oi_1 _10755_ (.A1(net34),
    .A2(_04693_),
    .Y(_04709_),
    .B1(net33));
 sg13g2_buf_1 _10756_ (.A(net105),
    .X(_04710_));
 sg13g2_a221oi_1 _10757_ (.B2(_04709_),
    .C1(net81),
    .B1(_04706_),
    .A1(net30),
    .Y(_00135_),
    .A2(_04699_));
 sg13g2_xnor2_1 _10758_ (.Y(_04711_),
    .A(_01382_),
    .B(net21));
 sg13g2_a21oi_1 _10759_ (.A1(_01077_),
    .A2(_04677_),
    .Y(_04712_),
    .B1(_04702_));
 sg13g2_nor2_1 _10760_ (.A(_04711_),
    .B(_04712_),
    .Y(_04713_));
 sg13g2_nand2_1 _10761_ (.Y(_04714_),
    .A(_04712_),
    .B(_04711_));
 sg13g2_nand3b_1 _10762_ (.B(_04499_),
    .C(_04714_),
    .Y(_04716_),
    .A_N(_04713_));
 sg13g2_nor2_1 _10763_ (.A(net99),
    .B(_01382_),
    .Y(_04717_));
 sg13g2_nand3_1 _10764_ (.B(_01070_),
    .C(_01179_),
    .A(_04685_),
    .Y(_04718_));
 sg13g2_xnor2_1 _10765_ (.Y(_04719_),
    .A(_01187_),
    .B(_04718_));
 sg13g2_nand2_1 _10766_ (.Y(_04720_),
    .A(_04540_),
    .B(_04717_));
 sg13g2_o21ai_1 _10767_ (.B1(_04720_),
    .Y(_04721_),
    .A1(_04639_),
    .A2(_04719_));
 sg13g2_a22oi_1 _10768_ (.Y(_04722_),
    .B1(net36),
    .B2(_04721_),
    .A2(_04717_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10769_ (.A1(_04716_),
    .A2(_04722_),
    .Y(_00136_),
    .B1(net83));
 sg13g2_xnor2_1 _10770_ (.Y(_04723_),
    .A(_01381_),
    .B(net21));
 sg13g2_inv_1 _10771_ (.Y(_04724_),
    .A(_04723_));
 sg13g2_nor2_1 _10772_ (.A(_01187_),
    .B(net21),
    .Y(_04726_));
 sg13g2_nor2_1 _10773_ (.A(_04726_),
    .B(_04713_),
    .Y(_04727_));
 sg13g2_xnor2_1 _10774_ (.Y(_04728_),
    .A(_04724_),
    .B(_04727_));
 sg13g2_inv_2 _10775_ (.Y(_04729_),
    .A(_04282_));
 sg13g2_buf_1 _10776_ (.A(_04729_),
    .X(_04730_));
 sg13g2_nand2_1 _10777_ (.Y(_04731_),
    .A(net80),
    .B(_01380_));
 sg13g2_a21oi_1 _10778_ (.A1(net34),
    .A2(_04731_),
    .Y(_04732_),
    .B1(net35));
 sg13g2_o21ai_1 _10779_ (.B1(_04732_),
    .Y(_04733_),
    .A1(net34),
    .A2(_04728_));
 sg13g2_nor3_2 _10780_ (.A(_04341_),
    .B(_04348_),
    .C(_04695_),
    .Y(_04734_));
 sg13g2_xnor2_1 _10781_ (.Y(_04735_),
    .A(_00045_),
    .B(_04734_));
 sg13g2_a21oi_1 _10782_ (.A1(net25),
    .A2(_04731_),
    .Y(_04737_),
    .B1(net43));
 sg13g2_o21ai_1 _10783_ (.B1(_04737_),
    .Y(_04738_),
    .A1(net25),
    .A2(_04735_));
 sg13g2_a21oi_1 _10784_ (.A1(_04733_),
    .A2(_04738_),
    .Y(_00137_),
    .B1(net83));
 sg13g2_xor2_1 _10785_ (.B(net21),
    .A(_01525_),
    .X(_04739_));
 sg13g2_inv_1 _10786_ (.Y(_04740_),
    .A(_04727_));
 sg13g2_a22oi_1 _10787_ (.Y(_04741_),
    .B1(_04724_),
    .B2(_04740_),
    .A2(_04677_),
    .A1(_01284_));
 sg13g2_xor2_1 _10788_ (.B(_04741_),
    .A(_04739_),
    .X(_04742_));
 sg13g2_nand2_1 _10789_ (.Y(_04743_),
    .A(net80),
    .B(_01525_));
 sg13g2_a21oi_1 _10790_ (.A1(_04498_),
    .A2(_04743_),
    .Y(_04744_),
    .B1(net35));
 sg13g2_o21ai_1 _10791_ (.B1(_04744_),
    .Y(_04745_),
    .A1(_04707_),
    .A2(_04742_));
 sg13g2_nor3_1 _10792_ (.A(_01381_),
    .B(_01382_),
    .C(_04718_),
    .Y(_04747_));
 sg13g2_xnor2_1 _10793_ (.Y(_04748_),
    .A(_00039_),
    .B(_04747_));
 sg13g2_a21oi_1 _10794_ (.A1(_04639_),
    .A2(_04743_),
    .Y(_04749_),
    .B1(net43));
 sg13g2_o21ai_1 _10795_ (.B1(_04749_),
    .Y(_04750_),
    .A1(net25),
    .A2(_04748_));
 sg13g2_a21oi_1 _10796_ (.A1(_04745_),
    .A2(_04750_),
    .Y(_00138_),
    .B1(net83));
 sg13g2_xnor2_1 _10797_ (.Y(_04751_),
    .A(_01637_),
    .B(_04580_));
 sg13g2_nor2_1 _10798_ (.A(_04739_),
    .B(_04741_),
    .Y(_04752_));
 sg13g2_a21oi_1 _10799_ (.A1(_01389_),
    .A2(_04677_),
    .Y(_04753_),
    .B1(_04752_));
 sg13g2_nor2_1 _10800_ (.A(_04751_),
    .B(_04753_),
    .Y(_04754_));
 sg13g2_nor2_1 _10801_ (.A(_04707_),
    .B(_04754_),
    .Y(_04755_));
 sg13g2_nand2_1 _10802_ (.Y(_04757_),
    .A(_04753_),
    .B(_04751_));
 sg13g2_nand2_1 _10803_ (.Y(_04758_),
    .A(net80),
    .B(_01636_));
 sg13g2_nor2_1 _10804_ (.A(_04758_),
    .B(net39),
    .Y(_04759_));
 sg13g2_a21oi_1 _10805_ (.A1(_04755_),
    .A2(_04757_),
    .Y(_04760_),
    .B1(_04759_));
 sg13g2_buf_1 _10806_ (.A(_04551_),
    .X(_04761_));
 sg13g2_a21oi_1 _10807_ (.A1(_04734_),
    .A2(_04345_),
    .Y(_04762_),
    .B1(_01529_));
 sg13g2_nand3_1 _10808_ (.B(_01529_),
    .C(_04345_),
    .A(_04734_),
    .Y(_04763_));
 sg13g2_nand3b_1 _10809_ (.B(net23),
    .C(_04763_),
    .Y(_04764_),
    .A_N(_04762_));
 sg13g2_o21ai_1 _10810_ (.B1(_04764_),
    .Y(_04765_),
    .A1(net23),
    .A2(_04758_));
 sg13g2_o21ai_1 _10811_ (.B1(net117),
    .Y(_04766_),
    .A1(net43),
    .A2(_04765_));
 sg13g2_a21oi_1 _10812_ (.A1(_04760_),
    .A2(net42),
    .Y(_00139_),
    .B1(_04766_));
 sg13g2_nor3_1 _10813_ (.A(_01637_),
    .B(_04677_),
    .C(_04753_),
    .Y(_04768_));
 sg13g2_nor3_1 _10814_ (.A(_01529_),
    .B(_04580_),
    .C(_04754_),
    .Y(_04769_));
 sg13g2_o21ai_1 _10815_ (.B1(_04497_),
    .Y(_04770_),
    .A1(_04768_),
    .A2(_04769_));
 sg13g2_o21ai_1 _10816_ (.B1(_01747_),
    .Y(_04771_),
    .A1(net80),
    .A2(_04497_));
 sg13g2_inv_1 _10817_ (.Y(_04772_),
    .A(_01747_));
 sg13g2_nor2_1 _10818_ (.A(_04772_),
    .B(_04770_),
    .Y(_04773_));
 sg13g2_a21oi_1 _10819_ (.A1(_04770_),
    .A2(_04771_),
    .Y(_04774_),
    .B1(_04773_));
 sg13g2_nand2_1 _10820_ (.Y(_04775_),
    .A(_04774_),
    .B(_04761_));
 sg13g2_nor4_1 _10821_ (.A(_01382_),
    .B(_01637_),
    .C(_04344_),
    .D(_04718_),
    .Y(_04776_));
 sg13g2_a21oi_1 _10822_ (.A1(_04776_),
    .A2(_01633_),
    .Y(_04778_),
    .B1(_04540_));
 sg13g2_o21ai_1 _10823_ (.B1(_04778_),
    .Y(_04779_),
    .A1(_01633_),
    .A2(_04776_));
 sg13g2_o21ai_1 _10824_ (.B1(_04548_),
    .Y(_04780_),
    .A1(_04772_),
    .A2(_04284_));
 sg13g2_nand3_1 _10825_ (.B(net33),
    .C(_04780_),
    .A(_04779_),
    .Y(_04781_));
 sg13g2_a21oi_1 _10826_ (.A1(_04775_),
    .A2(_04781_),
    .Y(_00140_),
    .B1(_04323_));
 sg13g2_nor2_1 _10827_ (.A(net84),
    .B(_05589_),
    .Y(_04782_));
 sg13g2_nand2b_1 _10828_ (.Y(_04783_),
    .B(_04601_),
    .A_N(_04602_));
 sg13g2_xnor2_1 _10829_ (.Y(_04784_),
    .A(_04495_),
    .B(_04783_));
 sg13g2_a22oi_1 _10830_ (.Y(_04785_),
    .B1(_04499_),
    .B2(_04784_),
    .A2(_04782_),
    .A1(_04557_));
 sg13g2_xor2_1 _10831_ (.B(_04647_),
    .A(_04543_),
    .X(_04786_));
 sg13g2_a21oi_1 _10832_ (.A1(net23),
    .A2(_04786_),
    .Y(_04788_),
    .B1(_04551_));
 sg13g2_o21ai_1 _10833_ (.B1(_04788_),
    .Y(_04789_),
    .A1(_04542_),
    .A2(_04782_));
 sg13g2_a21oi_1 _10834_ (.A1(_04785_),
    .A2(_04789_),
    .Y(_00141_),
    .B1(_04323_));
 sg13g2_inv_1 _10835_ (.Y(_04790_),
    .A(_04603_));
 sg13g2_nor3_1 _10836_ (.A(_04555_),
    .B(_04498_),
    .C(_04606_),
    .Y(_04791_));
 sg13g2_o21ai_1 _10837_ (.B1(_04791_),
    .Y(_04792_),
    .A1(_04790_),
    .A2(_04605_));
 sg13g2_nor2_1 _10838_ (.A(net99),
    .B(_00253_),
    .Y(_04793_));
 sg13g2_xnor2_1 _10839_ (.Y(_04794_),
    .A(_04651_),
    .B(_04650_));
 sg13g2_nand2_1 _10840_ (.Y(_04795_),
    .A(_04540_),
    .B(_04793_));
 sg13g2_o21ai_1 _10841_ (.B1(_04795_),
    .Y(_04796_),
    .A1(net24),
    .A2(_04794_));
 sg13g2_a22oi_1 _10842_ (.Y(_04798_),
    .B1(net36),
    .B2(_04796_),
    .A2(_04793_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10843_ (.A1(_04792_),
    .A2(_04798_),
    .Y(_00142_),
    .B1(net83));
 sg13g2_nor3_1 _10844_ (.A(_04555_),
    .B(net34),
    .C(_04608_),
    .Y(_04799_));
 sg13g2_nand2_1 _10845_ (.Y(_04800_),
    .A(_04607_),
    .B(_04598_));
 sg13g2_nand2_1 _10846_ (.Y(_04801_),
    .A(_04799_),
    .B(_04800_));
 sg13g2_nor2_1 _10847_ (.A(net99),
    .B(_00286_),
    .Y(_04802_));
 sg13g2_nor2b_1 _10848_ (.A(_04656_),
    .B_N(_04655_),
    .Y(_04803_));
 sg13g2_xnor2_1 _10849_ (.Y(_04804_),
    .A(_04803_),
    .B(_04654_));
 sg13g2_mux2_1 _10850_ (.A0(_04804_),
    .A1(_04802_),
    .S(net24),
    .X(_04805_));
 sg13g2_a22oi_1 _10851_ (.Y(_04806_),
    .B1(net33),
    .B2(_04805_),
    .A2(_04802_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10852_ (.A1(_04801_),
    .A2(_04806_),
    .Y(_00143_),
    .B1(net81));
 sg13g2_nor2_1 _10853_ (.A(net84),
    .B(_00340_),
    .Y(_04808_));
 sg13g2_nand2_1 _10854_ (.Y(_04809_),
    .A(net25),
    .B(_04808_));
 sg13g2_nor2_1 _10855_ (.A(_04645_),
    .B(_04646_),
    .Y(_04810_));
 sg13g2_xor2_1 _10856_ (.B(_04657_),
    .A(_04810_),
    .X(_04811_));
 sg13g2_a21oi_1 _10857_ (.A1(net23),
    .A2(_04811_),
    .Y(_04812_),
    .B1(net43));
 sg13g2_nand2_1 _10858_ (.Y(_04813_),
    .A(_04613_),
    .B(_04609_));
 sg13g2_nand3_1 _10859_ (.B(net39),
    .C(_04813_),
    .A(_04614_),
    .Y(_04814_));
 sg13g2_a21oi_1 _10860_ (.A1(net34),
    .A2(_04808_),
    .Y(_04815_),
    .B1(net33));
 sg13g2_a221oi_1 _10861_ (.B2(_04815_),
    .C1(net81),
    .B1(_04814_),
    .A1(_04809_),
    .Y(_00144_),
    .A2(_04812_));
 sg13g2_xor2_1 _10862_ (.B(_04659_),
    .A(_04644_),
    .X(_04817_));
 sg13g2_nand2_1 _10863_ (.Y(_04818_),
    .A(_04817_),
    .B(net23));
 sg13g2_nor2_1 _10864_ (.A(net84),
    .B(_04643_),
    .Y(_04819_));
 sg13g2_a21oi_1 _10865_ (.A1(net25),
    .A2(_04819_),
    .Y(_04820_),
    .B1(net43));
 sg13g2_nand2_1 _10866_ (.Y(_04821_),
    .A(_04618_),
    .B(_04616_));
 sg13g2_nor2_1 _10867_ (.A(_04498_),
    .B(_04619_),
    .Y(_04822_));
 sg13g2_a22oi_1 _10868_ (.Y(_04823_),
    .B1(_04821_),
    .B2(_04822_),
    .A2(_04819_),
    .A1(net34));
 sg13g2_a221oi_1 _10869_ (.B2(net42),
    .C1(net81),
    .B1(_04823_),
    .A1(_04818_),
    .Y(_00145_),
    .A2(_04820_));
 sg13g2_nor2_1 _10870_ (.A(_04663_),
    .B(_04660_),
    .Y(_04824_));
 sg13g2_nand2_1 _10871_ (.Y(_04825_),
    .A(_04660_),
    .B(_04663_));
 sg13g2_nand3b_1 _10872_ (.B(net23),
    .C(_04825_),
    .Y(_04827_),
    .A_N(_04824_));
 sg13g2_nor2_1 _10873_ (.A(net84),
    .B(_00383_),
    .Y(_04828_));
 sg13g2_a21oi_1 _10874_ (.A1(net25),
    .A2(_04828_),
    .Y(_04829_),
    .B1(net43));
 sg13g2_nand2_1 _10875_ (.Y(_04830_),
    .A(_04623_),
    .B(_04620_));
 sg13g2_nor2_1 _10876_ (.A(_04498_),
    .B(_04624_),
    .Y(_04831_));
 sg13g2_a22oi_1 _10877_ (.Y(_04832_),
    .B1(_04830_),
    .B2(_04831_),
    .A2(_04828_),
    .A1(net34));
 sg13g2_a221oi_1 _10878_ (.B2(net42),
    .C1(net81),
    .B1(_04832_),
    .A1(_04827_),
    .Y(_00146_),
    .A2(_04829_));
 sg13g2_nor2b_1 _10879_ (.A(net84),
    .B_N(_00668_),
    .Y(_04833_));
 sg13g2_nor2_1 _10880_ (.A(_04642_),
    .B(_04824_),
    .Y(_04834_));
 sg13g2_o21ai_1 _10881_ (.B1(_04541_),
    .Y(_04835_),
    .A1(_04661_),
    .A2(_04834_));
 sg13g2_a21oi_1 _10882_ (.A1(_04661_),
    .A2(_04834_),
    .Y(_04837_),
    .B1(_04835_));
 sg13g2_a21oi_1 _10883_ (.A1(net25),
    .A2(_04833_),
    .Y(_04838_),
    .B1(_04837_));
 sg13g2_nand2_1 _10884_ (.Y(_04839_),
    .A(_04625_),
    .B(_04593_));
 sg13g2_nand3b_1 _10885_ (.B(net39),
    .C(_04839_),
    .Y(_04840_),
    .A_N(_04626_));
 sg13g2_a21oi_1 _10886_ (.A1(net34),
    .A2(_04833_),
    .Y(_04841_),
    .B1(net33));
 sg13g2_a221oi_1 _10887_ (.B2(_04841_),
    .C1(net81),
    .B1(_04840_),
    .A1(net30),
    .Y(_00147_),
    .A2(_04838_));
 sg13g2_nand2_1 _10888_ (.Y(_04842_),
    .A(_04628_),
    .B(_04590_));
 sg13g2_nand2_1 _10889_ (.Y(_04843_),
    .A(_04627_),
    .B(_04588_));
 sg13g2_nand3_1 _10890_ (.B(_04499_),
    .C(_04843_),
    .A(_04842_),
    .Y(_04844_));
 sg13g2_nor2_1 _10891_ (.A(net99),
    .B(_04587_),
    .Y(_04845_));
 sg13g2_xnor2_1 _10892_ (.Y(_04847_),
    .A(_04640_),
    .B(_04667_));
 sg13g2_nand2_1 _10893_ (.Y(_04848_),
    .A(_04540_),
    .B(_04845_));
 sg13g2_o21ai_1 _10894_ (.B1(_04848_),
    .Y(_04849_),
    .A1(net24),
    .A2(_04847_));
 sg13g2_a22oi_1 _10895_ (.Y(_04850_),
    .B1(net33),
    .B2(_04849_),
    .A2(_04845_),
    .A1(_04557_));
 sg13g2_a21oi_1 _10896_ (.A1(_04844_),
    .A2(_04850_),
    .Y(_00148_),
    .B1(net81));
 sg13g2_xnor2_1 _10897_ (.Y(_04851_),
    .A(_04584_),
    .B(_04629_));
 sg13g2_nand2_1 _10898_ (.Y(_04852_),
    .A(net80),
    .B(_04339_));
 sg13g2_nor2_1 _10899_ (.A(_04852_),
    .B(net39),
    .Y(_04853_));
 sg13g2_a21oi_1 _10900_ (.A1(_04851_),
    .A2(net39),
    .Y(_04854_),
    .B1(_04853_));
 sg13g2_nand2_1 _10901_ (.Y(_04855_),
    .A(_04669_),
    .B(_00040_));
 sg13g2_nand3_1 _10902_ (.B(_04855_),
    .C(net23),
    .A(_04695_),
    .Y(_04857_));
 sg13g2_o21ai_1 _10903_ (.B1(_04857_),
    .Y(_04858_),
    .A1(net23),
    .A2(_04852_));
 sg13g2_o21ai_1 _10904_ (.B1(net130),
    .Y(_04859_),
    .A1(net43),
    .A2(_04858_));
 sg13g2_a21oi_1 _10905_ (.A1(_04854_),
    .A2(net42),
    .Y(_00149_),
    .B1(_04859_));
 sg13g2_nand2_1 _10906_ (.Y(_04860_),
    .A(net80),
    .B(_00217_));
 sg13g2_inv_1 _10907_ (.Y(_04861_),
    .A(_03306_));
 sg13g2_o21ai_1 _10908_ (.B1(_03347_),
    .Y(_04862_),
    .A1(_03316_),
    .A2(_04861_));
 sg13g2_nand3b_1 _10909_ (.B(_04862_),
    .C(_03378_),
    .Y(_04863_),
    .A_N(_03326_));
 sg13g2_nand3b_1 _10910_ (.B(_04863_),
    .C(_03598_),
    .Y(_04864_),
    .A_N(_03345_));
 sg13g2_nor2_1 _10911_ (.A(_03381_),
    .B(_03594_),
    .Y(_04865_));
 sg13g2_nand2_1 _10912_ (.Y(_04867_),
    .A(_04864_),
    .B(_04865_));
 sg13g2_nor2_1 _10913_ (.A(net125),
    .B(_05513_),
    .Y(_04868_));
 sg13g2_nand2_1 _10914_ (.Y(_04869_),
    .A(_02674_),
    .B(_02817_));
 sg13g2_nor4_1 _10915_ (.A(_03595_),
    .B(_04868_),
    .C(_04705_),
    .D(_04869_),
    .Y(_04870_));
 sg13g2_nand2_1 _10916_ (.Y(_04871_),
    .A(_04867_),
    .B(_04870_));
 sg13g2_buf_1 _10917_ (.A(_04871_),
    .X(_04872_));
 sg13g2_buf_1 _10918_ (.A(_04872_),
    .X(_04873_));
 sg13g2_buf_1 _10919_ (.A(net29),
    .X(_04874_));
 sg13g2_buf_1 _10920_ (.A(_05132_),
    .X(_04875_));
 sg13g2_a21oi_1 _10921_ (.A1(net27),
    .A2(_04860_),
    .Y(_04876_),
    .B1(net41));
 sg13g2_inv_1 _10922_ (.Y(_04878_),
    .A(_04872_));
 sg13g2_buf_1 _10923_ (.A(_04878_),
    .X(_04879_));
 sg13g2_nand2_1 _10924_ (.Y(_04880_),
    .A(net26),
    .B(_00218_));
 sg13g2_nand2_1 _10925_ (.Y(_04881_),
    .A(_04876_),
    .B(_04880_));
 sg13g2_nor2_1 _10926_ (.A(_03058_),
    .B(_04846_),
    .Y(_04882_));
 sg13g2_buf_2 _10927_ (.A(_04882_),
    .X(_04883_));
 sg13g2_nor2_2 _10928_ (.A(_04797_),
    .B(_04767_),
    .Y(_04884_));
 sg13g2_inv_1 _10929_ (.Y(_04885_),
    .A(_04884_));
 sg13g2_buf_1 _10930_ (.A(_04885_),
    .X(_04886_));
 sg13g2_a21oi_1 _10931_ (.A1(_04883_),
    .A2(_00217_),
    .Y(_04887_),
    .B1(net40));
 sg13g2_inv_1 _10932_ (.Y(_04889_),
    .A(_04883_));
 sg13g2_nand2_1 _10933_ (.Y(_04890_),
    .A(net38),
    .B(_04860_));
 sg13g2_a21oi_1 _10934_ (.A1(_04887_),
    .A2(_04890_),
    .Y(_04891_),
    .B1(_04708_));
 sg13g2_a221oi_1 _10935_ (.B2(_04891_),
    .C1(_04710_),
    .B1(_04881_),
    .A1(net30),
    .Y(_00150_),
    .A2(_04860_));
 sg13g2_nand2_1 _10936_ (.Y(_04892_),
    .A(_04729_),
    .B(_00792_));
 sg13g2_inv_1 _10937_ (.Y(_04893_),
    .A(_00053_));
 sg13g2_xnor2_1 _10938_ (.Y(_04894_),
    .A(_00299_),
    .B(_03385_));
 sg13g2_inv_1 _10939_ (.Y(_04895_),
    .A(_00055_));
 sg13g2_xnor2_1 _10940_ (.Y(_04896_),
    .A(_05596_),
    .B(_03332_));
 sg13g2_nor2_1 _10941_ (.A(_00057_),
    .B(_03323_),
    .Y(_04897_));
 sg13g2_xnor2_1 _10942_ (.Y(_04899_),
    .A(_05583_),
    .B(_03323_));
 sg13g2_inv_1 _10943_ (.Y(_04900_),
    .A(_04899_));
 sg13g2_xnor2_1 _10944_ (.Y(_04901_),
    .A(_05573_),
    .B(_03308_));
 sg13g2_and2_1 _10945_ (.A(_04901_),
    .B(_00217_),
    .X(_04902_));
 sg13g2_a21oi_1 _10946_ (.A1(_05573_),
    .A2(_03953_),
    .Y(_04903_),
    .B1(_04902_));
 sg13g2_nor2_1 _10947_ (.A(_04900_),
    .B(_04903_),
    .Y(_04904_));
 sg13g2_nor2_1 _10948_ (.A(_04897_),
    .B(_04904_),
    .Y(_04905_));
 sg13g2_inv_1 _10949_ (.Y(_04906_),
    .A(_04905_));
 sg13g2_a22oi_1 _10950_ (.Y(_04907_),
    .B1(_04896_),
    .B2(_04906_),
    .A2(_03334_),
    .A1(_04895_));
 sg13g2_xnor2_1 _10951_ (.Y(_04908_),
    .A(_00258_),
    .B(_03350_));
 sg13g2_nand2b_1 _10952_ (.Y(_04910_),
    .B(_04908_),
    .A_N(_04907_));
 sg13g2_o21ai_1 _10953_ (.B1(_04910_),
    .Y(_04911_),
    .A1(_00054_),
    .A2(_03350_));
 sg13g2_a22oi_1 _10954_ (.Y(_04912_),
    .B1(_04894_),
    .B2(_04911_),
    .A2(_03385_),
    .A1(_04893_));
 sg13g2_xnor2_1 _10955_ (.Y(_04913_),
    .A(_00354_),
    .B(_03603_));
 sg13g2_nand2b_1 _10956_ (.Y(_04914_),
    .B(_04913_),
    .A_N(_04912_));
 sg13g2_o21ai_1 _10957_ (.B1(_04914_),
    .Y(_04915_),
    .A1(_00052_),
    .A2(_03603_));
 sg13g2_xnor2_1 _10958_ (.Y(_04916_),
    .A(_00451_),
    .B(_03727_));
 sg13g2_nand2_1 _10959_ (.Y(_04917_),
    .A(_04915_),
    .B(_04916_));
 sg13g2_o21ai_1 _10960_ (.B1(_04917_),
    .Y(_04918_),
    .A1(_00051_),
    .A2(_03729_));
 sg13g2_xnor2_1 _10961_ (.Y(_04919_),
    .A(_00447_),
    .B(_03850_));
 sg13g2_nand2_1 _10962_ (.Y(_04921_),
    .A(_04918_),
    .B(_04919_));
 sg13g2_o21ai_1 _10963_ (.B1(_04921_),
    .Y(_04922_),
    .A1(_00050_),
    .A2(_03850_));
 sg13g2_xnor2_1 _10964_ (.Y(_04923_),
    .A(_00678_),
    .B(_04050_));
 sg13g2_nand2_1 _10965_ (.Y(_04924_),
    .A(_04922_),
    .B(_04923_));
 sg13g2_o21ai_1 _10966_ (.B1(_04924_),
    .Y(_04925_),
    .A1(_00028_),
    .A2(_04050_));
 sg13g2_a21oi_1 _10967_ (.A1(_03847_),
    .A2(_02773_),
    .Y(_04926_),
    .B1(_05546_));
 sg13g2_nand2b_1 _10968_ (.Y(_04927_),
    .B(_02817_),
    .A_N(_04926_));
 sg13g2_nand2_1 _10969_ (.Y(_04928_),
    .A(_04926_),
    .B(_02806_));
 sg13g2_nand2_1 _10970_ (.Y(_04929_),
    .A(_04927_),
    .B(_04928_));
 sg13g2_buf_1 _10971_ (.A(_04929_),
    .X(_04930_));
 sg13g2_nor2_1 _10972_ (.A(_00793_),
    .B(net22),
    .Y(_04932_));
 sg13g2_inv_2 _10973_ (.Y(_04933_),
    .A(net22));
 sg13g2_nor2_1 _10974_ (.A(_00792_),
    .B(_04933_),
    .Y(_04934_));
 sg13g2_nor2_1 _10975_ (.A(_04932_),
    .B(_04934_),
    .Y(_04935_));
 sg13g2_nor2_1 _10976_ (.A(_04885_),
    .B(net38),
    .Y(_04936_));
 sg13g2_o21ai_1 _10977_ (.B1(_04936_),
    .Y(_04937_),
    .A1(_04935_),
    .A2(_04925_));
 sg13g2_a21o_1 _10978_ (.A2(_04935_),
    .A1(_04925_),
    .B1(_04937_),
    .X(_04938_));
 sg13g2_nor2_1 _10979_ (.A(net118),
    .B(_00298_),
    .Y(_04939_));
 sg13g2_nor2_1 _10980_ (.A(_05484_),
    .B(_05583_),
    .Y(_04940_));
 sg13g2_nand2_1 _10981_ (.Y(_04941_),
    .A(net98),
    .B(_00217_));
 sg13g2_xor2_1 _10982_ (.B(_05573_),
    .A(net109),
    .X(_04943_));
 sg13g2_nor2b_1 _10983_ (.A(_04941_),
    .B_N(_04943_),
    .Y(_04944_));
 sg13g2_a21oi_1 _10984_ (.A1(net109),
    .A2(_05573_),
    .Y(_04945_),
    .B1(_04944_));
 sg13g2_nand2_1 _10985_ (.Y(_04946_),
    .A(_05484_),
    .B(_05583_));
 sg13g2_o21ai_1 _10986_ (.B1(_04946_),
    .Y(_04947_),
    .A1(_04940_),
    .A2(_04945_));
 sg13g2_inv_1 _10987_ (.Y(_04948_),
    .A(_04947_));
 sg13g2_nand2_1 _10988_ (.Y(_04949_),
    .A(net106),
    .B(_05596_));
 sg13g2_nor2_1 _10989_ (.A(net106),
    .B(_05596_),
    .Y(_04950_));
 sg13g2_a21oi_1 _10990_ (.A1(_04948_),
    .A2(_04949_),
    .Y(_04951_),
    .B1(_04950_));
 sg13g2_xor2_1 _10991_ (.B(_00258_),
    .A(net100),
    .X(_04952_));
 sg13g2_nand2_1 _10992_ (.Y(_04954_),
    .A(net100),
    .B(_00258_));
 sg13g2_inv_1 _10993_ (.Y(_04955_),
    .A(_04954_));
 sg13g2_a221oi_1 _10994_ (.B2(_04952_),
    .C1(_04955_),
    .B1(_04951_),
    .A1(net118),
    .Y(_04956_),
    .A2(_00298_));
 sg13g2_nor2_1 _10995_ (.A(_04939_),
    .B(_04956_),
    .Y(_04957_));
 sg13g2_nand2_1 _10996_ (.Y(_04958_),
    .A(_04957_),
    .B(_00354_));
 sg13g2_inv_1 _10997_ (.Y(_04959_),
    .A(_04958_));
 sg13g2_nor2_1 _10998_ (.A(\r2[7] ),
    .B(_04959_),
    .Y(_04960_));
 sg13g2_inv_1 _10999_ (.Y(_04961_),
    .A(_04960_));
 sg13g2_nor2_1 _11000_ (.A(_00678_),
    .B(_00449_),
    .Y(_04962_));
 sg13g2_inv_1 _11001_ (.Y(_04963_),
    .A(_00028_));
 sg13g2_a21oi_2 _11002_ (.B1(_04963_),
    .Y(_04965_),
    .A2(_04962_),
    .A1(_04961_));
 sg13g2_inv_1 _11003_ (.Y(_04966_),
    .A(_04965_));
 sg13g2_nand2_1 _11004_ (.Y(_04967_),
    .A(_04966_),
    .B(_00793_));
 sg13g2_nand2_1 _11005_ (.Y(_04968_),
    .A(_04965_),
    .B(_00792_));
 sg13g2_nand3_1 _11006_ (.B(net26),
    .C(_04968_),
    .A(_04967_),
    .Y(_04969_));
 sg13g2_a21oi_1 _11007_ (.A1(net27),
    .A2(_04892_),
    .Y(_04970_),
    .B1(net41));
 sg13g2_nor2_1 _11008_ (.A(_04885_),
    .B(_04883_),
    .Y(_04971_));
 sg13g2_inv_1 _11009_ (.Y(_04972_),
    .A(_04971_));
 sg13g2_o21ai_1 _11010_ (.B1(_04551_),
    .Y(_04973_),
    .A1(_04892_),
    .A2(_04972_));
 sg13g2_a21oi_1 _11011_ (.A1(_04969_),
    .A2(_04970_),
    .Y(_04974_),
    .B1(_04973_));
 sg13g2_buf_1 _11012_ (.A(_03520_),
    .X(_04976_));
 sg13g2_a221oi_1 _11013_ (.B2(_04974_),
    .C1(net79),
    .B1(_04938_),
    .A1(net30),
    .Y(_00151_),
    .A2(_04892_));
 sg13g2_nor2_1 _11014_ (.A(_04282_),
    .B(_00881_),
    .Y(_04977_));
 sg13g2_nand2_1 _11015_ (.Y(_04978_),
    .A(_04498_),
    .B(_04884_));
 sg13g2_nor2_1 _11016_ (.A(_00881_),
    .B(net22),
    .Y(_04979_));
 sg13g2_nor2_1 _11017_ (.A(_00880_),
    .B(_04933_),
    .Y(_04980_));
 sg13g2_nor2_1 _11018_ (.A(_04979_),
    .B(_04980_),
    .Y(_04981_));
 sg13g2_inv_1 _11019_ (.Y(_04982_),
    .A(_04981_));
 sg13g2_inv_1 _11020_ (.Y(_04983_),
    .A(_04934_));
 sg13g2_a21oi_2 _11021_ (.B1(_04932_),
    .Y(_04984_),
    .A2(_04983_),
    .A1(_04925_));
 sg13g2_xnor2_1 _11022_ (.Y(_04986_),
    .A(_04982_),
    .B(_04984_));
 sg13g2_nand2_1 _11023_ (.Y(_04987_),
    .A(_04986_),
    .B(_04836_));
 sg13g2_o21ai_1 _11024_ (.B1(_04987_),
    .Y(_04988_),
    .A1(_04836_),
    .A2(_04977_));
 sg13g2_o21ai_1 _11025_ (.B1(_05122_),
    .Y(_04989_),
    .A1(_04977_),
    .A2(_04878_));
 sg13g2_nand2_1 _11026_ (.Y(_04990_),
    .A(net118),
    .B(_00298_));
 sg13g2_inv_1 _11027_ (.Y(_04991_),
    .A(_04990_));
 sg13g2_inv_1 _11028_ (.Y(_04992_),
    .A(_04949_));
 sg13g2_nor2_1 _11029_ (.A(_04950_),
    .B(_04992_),
    .Y(_04993_));
 sg13g2_nand2_1 _11030_ (.Y(_04994_),
    .A(_04993_),
    .B(_04952_));
 sg13g2_a21oi_1 _11031_ (.A1(_04952_),
    .A2(_04992_),
    .Y(_04995_),
    .B1(_04955_));
 sg13g2_o21ai_1 _11032_ (.B1(_04995_),
    .Y(_04997_),
    .A1(_04994_),
    .A2(_04948_));
 sg13g2_nor2_1 _11033_ (.A(_04939_),
    .B(_04991_),
    .Y(_04998_));
 sg13g2_nand2_1 _11034_ (.Y(_04999_),
    .A(_04997_),
    .B(_04998_));
 sg13g2_inv_1 _11035_ (.Y(_05000_),
    .A(_04999_));
 sg13g2_a22oi_1 _11036_ (.Y(_05001_),
    .B1(_00396_),
    .B2(_05000_),
    .A2(_04991_),
    .A1(_00354_));
 sg13g2_a21oi_1 _11037_ (.A1(_05001_),
    .A2(_00451_),
    .Y(_05002_),
    .B1(_00449_));
 sg13g2_nor2_1 _11038_ (.A(_00678_),
    .B(_05002_),
    .Y(_05003_));
 sg13g2_nor2_1 _11039_ (.A(_00793_),
    .B(_05003_),
    .Y(_05004_));
 sg13g2_a21oi_1 _11040_ (.A1(_05004_),
    .A2(_00881_),
    .Y(_05005_),
    .B1(_04872_));
 sg13g2_o21ai_1 _11041_ (.B1(_05005_),
    .Y(_05006_),
    .A1(_00881_),
    .A2(_05004_));
 sg13g2_nand2b_1 _11042_ (.Y(_05008_),
    .B(_05006_),
    .A_N(_04989_));
 sg13g2_o21ai_1 _11043_ (.B1(_05008_),
    .Y(_05009_),
    .A1(_04978_),
    .A2(_04988_));
 sg13g2_a22oi_1 _11044_ (.Y(_05010_),
    .B1(net42),
    .B2(_05009_),
    .A2(_04977_),
    .A1(_04559_));
 sg13g2_nor2_1 _11045_ (.A(net94),
    .B(_05010_),
    .Y(_00152_));
 sg13g2_xnor2_1 _11046_ (.Y(_05011_),
    .A(_00986_),
    .B(net22));
 sg13g2_inv_1 _11047_ (.Y(_05012_),
    .A(_05011_));
 sg13g2_inv_1 _11048_ (.Y(_05013_),
    .A(_04979_));
 sg13g2_o21ai_1 _11049_ (.B1(_05013_),
    .Y(_05014_),
    .A1(_04980_),
    .A2(_04984_));
 sg13g2_nor2_1 _11050_ (.A(_05012_),
    .B(_05014_),
    .Y(_05015_));
 sg13g2_nand2_1 _11051_ (.Y(_05016_),
    .A(_05014_),
    .B(_05012_));
 sg13g2_nand2_1 _11052_ (.Y(_05018_),
    .A(_05016_),
    .B(_04883_));
 sg13g2_nor2_1 _11053_ (.A(_04283_),
    .B(_00986_),
    .Y(_05019_));
 sg13g2_a21oi_1 _11054_ (.A1(net38),
    .A2(_05019_),
    .Y(_05020_),
    .B1(net40));
 sg13g2_o21ai_1 _11055_ (.B1(_05020_),
    .Y(_05021_),
    .A1(_05015_),
    .A2(_05018_));
 sg13g2_inv_1 _11056_ (.Y(_05022_),
    .A(_00030_));
 sg13g2_nand2_1 _11057_ (.Y(_05023_),
    .A(_00880_),
    .B(_00792_));
 sg13g2_nor2_1 _11058_ (.A(_05023_),
    .B(_04965_),
    .Y(_05024_));
 sg13g2_xnor2_1 _11059_ (.Y(_05025_),
    .A(_05022_),
    .B(_05024_));
 sg13g2_a21oi_1 _11060_ (.A1(net29),
    .A2(_05019_),
    .Y(_05026_),
    .B1(_05132_));
 sg13g2_o21ai_1 _11061_ (.B1(_05026_),
    .Y(_05027_),
    .A1(net27),
    .A2(_05025_));
 sg13g2_nand2_1 _11062_ (.Y(_05029_),
    .A(_05021_),
    .B(_05027_));
 sg13g2_o21ai_1 _11063_ (.B1(net130),
    .Y(_05030_),
    .A1(_05019_),
    .A2(_04552_));
 sg13g2_a21oi_1 _11064_ (.A1(_05029_),
    .A2(_04761_),
    .Y(_00153_),
    .B1(_05030_));
 sg13g2_nor2_1 _11065_ (.A(_04282_),
    .B(_01083_),
    .Y(_05031_));
 sg13g2_inv_1 _11066_ (.Y(_05032_),
    .A(_05031_));
 sg13g2_nor3_1 _11067_ (.A(_04982_),
    .B(_05011_),
    .C(_04984_),
    .Y(_05033_));
 sg13g2_a221oi_1 _11068_ (.B2(_04933_),
    .C1(_05033_),
    .B1(_05022_),
    .A1(_00986_),
    .Y(_05034_),
    .A2(_04979_));
 sg13g2_xnor2_1 _11069_ (.Y(_05035_),
    .A(_01081_),
    .B(net22));
 sg13g2_nand2b_1 _11070_ (.Y(_05036_),
    .B(_05035_),
    .A_N(_05034_));
 sg13g2_inv_1 _11071_ (.Y(_05037_),
    .A(_05035_));
 sg13g2_nand2_1 _11072_ (.Y(_05039_),
    .A(_05034_),
    .B(_05037_));
 sg13g2_a21oi_1 _11073_ (.A1(_05036_),
    .A2(_05039_),
    .Y(_05040_),
    .B1(_04846_));
 sg13g2_a21oi_1 _11074_ (.A1(_04846_),
    .A2(_05032_),
    .Y(_05041_),
    .B1(_05040_));
 sg13g2_a21oi_1 _11075_ (.A1(net39),
    .A2(_05032_),
    .Y(_05042_),
    .B1(_04886_));
 sg13g2_o21ai_1 _11076_ (.B1(_05042_),
    .Y(_05043_),
    .A1(net39),
    .A2(_05041_));
 sg13g2_nand2_1 _11077_ (.Y(_05044_),
    .A(_04872_),
    .B(_04283_));
 sg13g2_nor2_1 _11078_ (.A(_00986_),
    .B(_05023_),
    .Y(_05045_));
 sg13g2_nor2b_1 _11079_ (.A(_05003_),
    .B_N(_05045_),
    .Y(_05046_));
 sg13g2_a22oi_1 _11080_ (.Y(_05047_),
    .B1(net26),
    .B2(_05046_),
    .A2(_05044_),
    .A1(_01081_));
 sg13g2_nor2_1 _11081_ (.A(_04875_),
    .B(_05047_),
    .Y(_05048_));
 sg13g2_nand3_1 _11082_ (.B(_01081_),
    .C(net26),
    .A(_05046_),
    .Y(_05050_));
 sg13g2_a21oi_1 _11083_ (.A1(_05048_),
    .A2(_05050_),
    .Y(_05051_),
    .B1(net33));
 sg13g2_a221oi_1 _11084_ (.B2(_05051_),
    .C1(_04976_),
    .B1(_05043_),
    .A1(_04691_),
    .Y(_00154_),
    .A2(_05032_));
 sg13g2_nor2_1 _11085_ (.A(_04282_),
    .B(_01193_),
    .Y(_05052_));
 sg13g2_inv_1 _11086_ (.Y(_05053_),
    .A(_05052_));
 sg13g2_o21ai_1 _11087_ (.B1(_04933_),
    .Y(_05054_),
    .A1(_01081_),
    .A2(_05022_));
 sg13g2_o21ai_1 _11088_ (.B1(_05054_),
    .Y(_05055_),
    .A1(_05037_),
    .A2(_05016_));
 sg13g2_xnor2_1 _11089_ (.Y(_05056_),
    .A(_01192_),
    .B(net22));
 sg13g2_a21oi_1 _11090_ (.A1(_05055_),
    .A2(_05056_),
    .Y(_05057_),
    .B1(_04846_));
 sg13g2_o21ai_1 _11091_ (.B1(_05057_),
    .Y(_05058_),
    .A1(_05055_),
    .A2(_05056_));
 sg13g2_a21oi_1 _11092_ (.A1(_04846_),
    .A2(_05052_),
    .Y(_05060_),
    .B1(_04703_));
 sg13g2_o21ai_1 _11093_ (.B1(_04884_),
    .Y(_05061_),
    .A1(_05052_),
    .A2(_04498_));
 sg13g2_a21o_1 _11094_ (.A2(_05060_),
    .A1(_05058_),
    .B1(_05061_),
    .X(_05062_));
 sg13g2_nand2_1 _11095_ (.Y(_05063_),
    .A(_01081_),
    .B(\r2[12] ));
 sg13g2_nor3_1 _11096_ (.A(_05023_),
    .B(_05063_),
    .C(_04965_),
    .Y(_05064_));
 sg13g2_a21oi_1 _11097_ (.A1(_05064_),
    .A2(_01193_),
    .Y(_05065_),
    .B1(_04873_));
 sg13g2_o21ai_1 _11098_ (.B1(_05065_),
    .Y(_05066_),
    .A1(_01193_),
    .A2(_05064_));
 sg13g2_a21oi_1 _11099_ (.A1(_04874_),
    .A2(_05053_),
    .Y(_05067_),
    .B1(_04875_));
 sg13g2_a21oi_1 _11100_ (.A1(_05066_),
    .A2(_05067_),
    .Y(_05068_),
    .B1(_04708_));
 sg13g2_a221oi_1 _11101_ (.B2(_05068_),
    .C1(_04976_),
    .B1(_05062_),
    .A1(net30),
    .Y(_00155_),
    .A2(_05053_));
 sg13g2_xnor2_1 _11102_ (.Y(_05070_),
    .A(_01377_),
    .B(net22));
 sg13g2_inv_1 _11103_ (.Y(_05071_),
    .A(_05056_));
 sg13g2_o21ai_1 _11104_ (.B1(_04933_),
    .Y(_05072_),
    .A1(_01192_),
    .A2(_01081_));
 sg13g2_o21ai_1 _11105_ (.B1(_05072_),
    .Y(_05073_),
    .A1(_05071_),
    .A2(_05036_));
 sg13g2_inv_1 _11106_ (.Y(_05074_),
    .A(_05073_));
 sg13g2_nor2_1 _11107_ (.A(_05070_),
    .B(_05074_),
    .Y(_05075_));
 sg13g2_a21o_1 _11108_ (.A2(_05070_),
    .A1(_05074_),
    .B1(net38),
    .X(_05076_));
 sg13g2_nor2_1 _11109_ (.A(_04282_),
    .B(_01377_),
    .Y(_05077_));
 sg13g2_a21oi_1 _11110_ (.A1(net38),
    .A2(_05077_),
    .Y(_05078_),
    .B1(_04885_));
 sg13g2_o21ai_1 _11111_ (.B1(_05078_),
    .Y(_05079_),
    .A1(_05075_),
    .A2(_05076_));
 sg13g2_nor3_1 _11112_ (.A(_01193_),
    .B(_00881_),
    .C(_05063_),
    .Y(_05081_));
 sg13g2_a21oi_1 _11113_ (.A1(_05004_),
    .A2(_05081_),
    .Y(_05082_),
    .B1(_01283_));
 sg13g2_nand3_1 _11114_ (.B(_01283_),
    .C(_05081_),
    .A(_05004_),
    .Y(_05083_));
 sg13g2_nand2b_1 _11115_ (.Y(_05084_),
    .B(_05083_),
    .A_N(_05082_));
 sg13g2_a21oi_1 _11116_ (.A1(net29),
    .A2(_05077_),
    .Y(_05085_),
    .B1(_05132_));
 sg13g2_o21ai_1 _11117_ (.B1(_05085_),
    .Y(_05086_),
    .A1(_04874_),
    .A2(_05084_));
 sg13g2_nand2_1 _11118_ (.Y(_05087_),
    .A(_05079_),
    .B(_05086_));
 sg13g2_o21ai_1 _11119_ (.B1(net130),
    .Y(_05088_),
    .A1(_05077_),
    .A2(net43));
 sg13g2_a21oi_1 _11120_ (.A1(_05087_),
    .A2(net42),
    .Y(_00156_),
    .B1(_05088_));
 sg13g2_nor2_1 _11121_ (.A(net99),
    .B(_01523_),
    .Y(_05089_));
 sg13g2_nand2_1 _11122_ (.Y(_05091_),
    .A(\r2[15] ),
    .B(_01192_));
 sg13g2_nand2b_1 _11123_ (.Y(_05092_),
    .B(_05064_),
    .A_N(_05091_));
 sg13g2_a21oi_1 _11124_ (.A1(_05092_),
    .A2(_01379_),
    .Y(_05093_),
    .B1(net29));
 sg13g2_o21ai_1 _11125_ (.B1(_05093_),
    .Y(_05094_),
    .A1(_01379_),
    .A2(_05092_));
 sg13g2_a21oi_1 _11126_ (.A1(net29),
    .A2(_05089_),
    .Y(_05095_),
    .B1(_05132_));
 sg13g2_a21oi_1 _11127_ (.A1(_05094_),
    .A2(_05095_),
    .Y(_05096_),
    .B1(net35));
 sg13g2_a21oi_1 _11128_ (.A1(_01283_),
    .A2(_04933_),
    .Y(_05097_),
    .B1(_05075_));
 sg13g2_xnor2_1 _11129_ (.Y(_05098_),
    .A(_01523_),
    .B(_04930_));
 sg13g2_a21oi_1 _11130_ (.A1(_05097_),
    .A2(_05098_),
    .Y(_05099_),
    .B1(net38));
 sg13g2_or2_1 _11131_ (.X(_05100_),
    .B(_05097_),
    .A(_05098_));
 sg13g2_nand2_1 _11132_ (.Y(_05102_),
    .A(_05099_),
    .B(_05100_));
 sg13g2_nand2_1 _11133_ (.Y(_05103_),
    .A(_04703_),
    .B(_05089_));
 sg13g2_a21oi_1 _11134_ (.A1(_04846_),
    .A2(_05089_),
    .Y(_05104_),
    .B1(_04885_));
 sg13g2_nand3_1 _11135_ (.B(_05103_),
    .C(_05104_),
    .A(_05102_),
    .Y(_05105_));
 sg13g2_a22oi_1 _11136_ (.Y(_05106_),
    .B1(_05096_),
    .B2(_05105_),
    .A2(_05089_),
    .A1(net36));
 sg13g2_nor2_1 _11137_ (.A(_05482_),
    .B(_05106_),
    .Y(_00157_));
 sg13g2_nand2_1 _11138_ (.Y(_05107_),
    .A(_04730_),
    .B(\r2[17] ));
 sg13g2_o21ai_1 _11139_ (.B1(_05100_),
    .Y(_05108_),
    .A1(_01379_),
    .A2(_04930_));
 sg13g2_xnor2_1 _11140_ (.Y(_05109_),
    .A(_01631_),
    .B(net22));
 sg13g2_a21oi_1 _11141_ (.A1(_05108_),
    .A2(_05109_),
    .Y(_05110_),
    .B1(net38));
 sg13g2_o21ai_1 _11142_ (.B1(_05110_),
    .Y(_05112_),
    .A1(_05108_),
    .A2(_05109_));
 sg13g2_buf_1 _11143_ (.A(net38),
    .X(_05113_));
 sg13g2_a21oi_1 _11144_ (.A1(net32),
    .A2(_05107_),
    .Y(_05114_),
    .B1(net40));
 sg13g2_nand2_1 _11145_ (.Y(_05115_),
    .A(_05112_),
    .B(_05114_));
 sg13g2_nor3_1 _11146_ (.A(_01083_),
    .B(_01523_),
    .C(_05091_),
    .Y(_05116_));
 sg13g2_a21oi_1 _11147_ (.A1(_05046_),
    .A2(_05116_),
    .Y(_05117_),
    .B1(_01631_));
 sg13g2_nand3_1 _11148_ (.B(_01631_),
    .C(_05116_),
    .A(_05046_),
    .Y(_05118_));
 sg13g2_nand3b_1 _11149_ (.B(net26),
    .C(_05118_),
    .Y(_05119_),
    .A_N(_05117_));
 sg13g2_a21oi_1 _11150_ (.A1(net27),
    .A2(_05107_),
    .Y(_05120_),
    .B1(net41));
 sg13g2_a21oi_1 _11151_ (.A1(_05119_),
    .A2(_05120_),
    .Y(_05121_),
    .B1(net33));
 sg13g2_a221oi_1 _11152_ (.B2(_05121_),
    .C1(net79),
    .B1(_05115_),
    .A1(net30),
    .Y(_00158_),
    .A2(_05107_));
 sg13g2_nand2_1 _11153_ (.Y(_05123_),
    .A(_04729_),
    .B(\r2[18] ));
 sg13g2_nand2b_1 _11154_ (.Y(_05124_),
    .B(_05108_),
    .A_N(_05109_));
 sg13g2_nand3_1 _11155_ (.B(_00013_),
    .C(_04933_),
    .A(_05124_),
    .Y(_05125_));
 sg13g2_o21ai_1 _11156_ (.B1(_05125_),
    .Y(_05126_),
    .A1(_04933_),
    .A2(_05124_));
 sg13g2_xnor2_1 _11157_ (.Y(_05127_),
    .A(_00015_),
    .B(_05126_));
 sg13g2_a21oi_1 _11158_ (.A1(net32),
    .A2(_05123_),
    .Y(_05128_),
    .B1(net40));
 sg13g2_o21ai_1 _11159_ (.B1(_05128_),
    .Y(_05129_),
    .A1(net32),
    .A2(_05127_));
 sg13g2_nand4_1 _11160_ (.B(\r2[17] ),
    .C(_05045_),
    .A(_04966_),
    .Y(_05130_),
    .D(_05116_));
 sg13g2_a21oi_1 _11161_ (.A1(_05130_),
    .A2(\r2[18] ),
    .Y(_05131_),
    .B1(net29));
 sg13g2_o21ai_1 _11162_ (.B1(_05131_),
    .Y(_05133_),
    .A1(\r2[18] ),
    .A2(_05130_));
 sg13g2_a21oi_1 _11163_ (.A1(net27),
    .A2(_05123_),
    .Y(_05134_),
    .B1(net41));
 sg13g2_a21oi_1 _11164_ (.A1(_05133_),
    .A2(_05134_),
    .Y(_05135_),
    .B1(net35));
 sg13g2_a221oi_1 _11165_ (.B2(_05135_),
    .C1(net79),
    .B1(_05129_),
    .A1(net30),
    .Y(_00159_),
    .A2(_05123_));
 sg13g2_nand2_1 _11166_ (.Y(_05136_),
    .A(net80),
    .B(_05573_));
 sg13g2_xnor2_1 _11167_ (.Y(_05137_),
    .A(_04941_),
    .B(_04943_));
 sg13g2_a21oi_1 _11168_ (.A1(net27),
    .A2(_05136_),
    .Y(_05138_),
    .B1(net41));
 sg13g2_o21ai_1 _11169_ (.B1(_05138_),
    .Y(_05139_),
    .A1(net27),
    .A2(_05137_));
 sg13g2_a21oi_1 _11170_ (.A1(_04889_),
    .A2(_05136_),
    .Y(_05140_),
    .B1(net40));
 sg13g2_nor2_1 _11171_ (.A(_00217_),
    .B(_04901_),
    .Y(_05141_));
 sg13g2_o21ai_1 _11172_ (.B1(_04883_),
    .Y(_05143_),
    .A1(_04902_),
    .A2(_05141_));
 sg13g2_a21oi_1 _11173_ (.A1(_05140_),
    .A2(_05143_),
    .Y(_05144_),
    .B1(net35));
 sg13g2_a221oi_1 _11174_ (.B2(_05144_),
    .C1(net79),
    .B1(_05139_),
    .A1(_04691_),
    .Y(_00160_),
    .A2(_05136_));
 sg13g2_nand2b_1 _11175_ (.Y(_05145_),
    .B(_04946_),
    .A_N(_04940_));
 sg13g2_xnor2_1 _11176_ (.Y(_05146_),
    .A(_05145_),
    .B(_04945_));
 sg13g2_nand2_1 _11177_ (.Y(_05147_),
    .A(_04879_),
    .B(_05122_));
 sg13g2_nand2_1 _11178_ (.Y(_05148_),
    .A(_04903_),
    .B(_04900_));
 sg13g2_nand3b_1 _11179_ (.B(_04936_),
    .C(_05148_),
    .Y(_05149_),
    .A_N(_04904_));
 sg13g2_o21ai_1 _11180_ (.B1(_05149_),
    .Y(_05150_),
    .A1(_05146_),
    .A2(_05147_));
 sg13g2_nand2_1 _11181_ (.Y(_05151_),
    .A(_05150_),
    .B(net42));
 sg13g2_nand2_1 _11182_ (.Y(_05153_),
    .A(_04872_),
    .B(_05122_));
 sg13g2_nand3_1 _11183_ (.B(_04551_),
    .C(_04972_),
    .A(_05153_),
    .Y(_05154_));
 sg13g2_nand3_1 _11184_ (.B(_05583_),
    .C(_04730_),
    .A(_05154_),
    .Y(_05155_));
 sg13g2_a21oi_1 _11185_ (.A1(_05151_),
    .A2(_05155_),
    .Y(_00161_),
    .B1(net81));
 sg13g2_nor2_1 _11186_ (.A(net84),
    .B(_05598_),
    .Y(_05156_));
 sg13g2_xnor2_1 _11187_ (.Y(_05157_),
    .A(_04993_),
    .B(_04947_));
 sg13g2_nand2_1 _11188_ (.Y(_05158_),
    .A(_04906_),
    .B(_04896_));
 sg13g2_nand2b_1 _11189_ (.Y(_05159_),
    .B(_04905_),
    .A_N(_04896_));
 sg13g2_nand3_1 _11190_ (.B(_05159_),
    .C(_04936_),
    .A(_05158_),
    .Y(_05160_));
 sg13g2_o21ai_1 _11191_ (.B1(_05160_),
    .Y(_05161_),
    .A1(_05147_),
    .A2(_05157_));
 sg13g2_a22oi_1 _11192_ (.Y(_05163_),
    .B1(net42),
    .B2(_05161_),
    .A2(_05156_),
    .A1(_05154_));
 sg13g2_nor2_1 _11193_ (.A(net94),
    .B(_05163_),
    .Y(_00162_));
 sg13g2_nand2_1 _11194_ (.Y(_05164_),
    .A(_04729_),
    .B(_00258_));
 sg13g2_nand2b_1 _11195_ (.Y(_05165_),
    .B(_04907_),
    .A_N(_04908_));
 sg13g2_nand3_1 _11196_ (.B(_05165_),
    .C(_04883_),
    .A(_04910_),
    .Y(_05166_));
 sg13g2_o21ai_1 _11197_ (.B1(_05166_),
    .Y(_05167_),
    .A1(_04883_),
    .A2(_05164_));
 sg13g2_nand2_1 _11198_ (.Y(_05168_),
    .A(_05167_),
    .B(_04884_));
 sg13g2_xnor2_1 _11199_ (.Y(_05169_),
    .A(_04952_),
    .B(_04951_));
 sg13g2_nand2_1 _11200_ (.Y(_05170_),
    .A(_05169_),
    .B(_04879_));
 sg13g2_a21oi_1 _11201_ (.A1(net27),
    .A2(_05164_),
    .Y(_05171_),
    .B1(net41));
 sg13g2_a21oi_1 _11202_ (.A1(_05170_),
    .A2(_05171_),
    .Y(_05173_),
    .B1(net35));
 sg13g2_a221oi_1 _11203_ (.B2(_05173_),
    .C1(net79),
    .B1(_05168_),
    .A1(net30),
    .Y(_00163_),
    .A2(_05164_));
 sg13g2_nand2_1 _11204_ (.Y(_05174_),
    .A(net80),
    .B(_00298_));
 sg13g2_xor2_1 _11205_ (.B(_04911_),
    .A(_04894_),
    .X(_05175_));
 sg13g2_a21oi_1 _11206_ (.A1(net32),
    .A2(_05174_),
    .Y(_05176_),
    .B1(net40));
 sg13g2_o21ai_1 _11207_ (.B1(_05176_),
    .Y(_05177_),
    .A1(net32),
    .A2(_05175_));
 sg13g2_o21ai_1 _11208_ (.B1(_04551_),
    .Y(_05178_),
    .A1(_05174_),
    .A2(_05153_));
 sg13g2_nor2_1 _11209_ (.A(_04998_),
    .B(_04997_),
    .Y(_05179_));
 sg13g2_nor3_1 _11210_ (.A(_05147_),
    .B(_05179_),
    .C(_05000_),
    .Y(_05180_));
 sg13g2_nor2_1 _11211_ (.A(_05178_),
    .B(_05180_),
    .Y(_05181_));
 sg13g2_a221oi_1 _11212_ (.B2(_05181_),
    .C1(net79),
    .B1(_05177_),
    .A1(net36),
    .Y(_00164_),
    .A2(_05174_));
 sg13g2_nor2_1 _11213_ (.A(_04282_),
    .B(_00356_),
    .Y(_05183_));
 sg13g2_inv_1 _11214_ (.Y(_05184_),
    .A(_05183_));
 sg13g2_nand2b_1 _11215_ (.Y(_05185_),
    .B(_04912_),
    .A_N(_04913_));
 sg13g2_nand3_1 _11216_ (.B(_04936_),
    .C(_05185_),
    .A(_04914_),
    .Y(_05186_));
 sg13g2_a21oi_1 _11217_ (.A1(_04971_),
    .A2(_05183_),
    .Y(_05187_),
    .B1(_04555_));
 sg13g2_o21ai_1 _11218_ (.B1(_05187_),
    .Y(_05188_),
    .A1(_05184_),
    .A2(_05153_));
 sg13g2_nor2_1 _11219_ (.A(_00354_),
    .B(_04957_),
    .Y(_05189_));
 sg13g2_nor3_1 _11220_ (.A(_05147_),
    .B(_05189_),
    .C(_04959_),
    .Y(_05190_));
 sg13g2_nor2_1 _11221_ (.A(_05188_),
    .B(_05190_),
    .Y(_05191_));
 sg13g2_a221oi_1 _11222_ (.B2(_05191_),
    .C1(net79),
    .B1(_05186_),
    .A1(net36),
    .Y(_00165_),
    .A2(_05184_));
 sg13g2_nand2_1 _11223_ (.Y(_05192_),
    .A(_04729_),
    .B(\r2[7] ));
 sg13g2_xor2_1 _11224_ (.B(_04915_),
    .A(_04916_),
    .X(_05193_));
 sg13g2_a21oi_1 _11225_ (.A1(net32),
    .A2(_05192_),
    .Y(_05194_),
    .B1(net40));
 sg13g2_o21ai_1 _11226_ (.B1(_05194_),
    .Y(_05195_),
    .A1(net32),
    .A2(_05193_));
 sg13g2_nand2b_1 _11227_ (.Y(_05196_),
    .B(_00392_),
    .A_N(_05001_));
 sg13g2_nand2_1 _11228_ (.Y(_05197_),
    .A(_05001_),
    .B(_00051_));
 sg13g2_nand3_1 _11229_ (.B(net26),
    .C(_05197_),
    .A(_05196_),
    .Y(_05198_));
 sg13g2_a21oi_1 _11230_ (.A1(_04873_),
    .A2(_05192_),
    .Y(_05199_),
    .B1(net41));
 sg13g2_a21oi_1 _11231_ (.A1(_05198_),
    .A2(_05199_),
    .Y(_05200_),
    .B1(net35));
 sg13g2_a221oi_1 _11232_ (.B2(_05200_),
    .C1(net79),
    .B1(_05195_),
    .A1(net36),
    .Y(_00166_),
    .A2(_05192_));
 sg13g2_nand2_1 _11233_ (.Y(_05202_),
    .A(_04729_),
    .B(_00447_));
 sg13g2_xor2_1 _11234_ (.B(_04918_),
    .A(_04919_),
    .X(_05203_));
 sg13g2_a21oi_1 _11235_ (.A1(_05113_),
    .A2(_05202_),
    .Y(_05204_),
    .B1(net40));
 sg13g2_o21ai_1 _11236_ (.B1(_05204_),
    .Y(_05205_),
    .A1(net32),
    .A2(_05203_));
 sg13g2_nand2_1 _11237_ (.Y(_05206_),
    .A(_04961_),
    .B(_00449_));
 sg13g2_nand2_1 _11238_ (.Y(_05207_),
    .A(_04960_),
    .B(_00447_));
 sg13g2_nand3_1 _11239_ (.B(net26),
    .C(_05207_),
    .A(_05206_),
    .Y(_05208_));
 sg13g2_a21oi_1 _11240_ (.A1(net29),
    .A2(_05202_),
    .Y(_05209_),
    .B1(net41));
 sg13g2_a21oi_1 _11241_ (.A1(_05208_),
    .A2(_05209_),
    .Y(_05210_),
    .B1(_04690_));
 sg13g2_a221oi_1 _11242_ (.B2(_05210_),
    .C1(net96),
    .B1(_05205_),
    .A1(_04638_),
    .Y(_00167_),
    .A2(_05202_));
 sg13g2_nand2_1 _11243_ (.Y(_05212_),
    .A(_04729_),
    .B(_00678_));
 sg13g2_xor2_1 _11244_ (.B(_04922_),
    .A(_04923_),
    .X(_05213_));
 sg13g2_a21oi_1 _11245_ (.A1(_04889_),
    .A2(_05212_),
    .Y(_05214_),
    .B1(_04886_));
 sg13g2_o21ai_1 _11246_ (.B1(_05214_),
    .Y(_05215_),
    .A1(_05113_),
    .A2(_05213_));
 sg13g2_nand2b_1 _11247_ (.Y(_05216_),
    .B(_00028_),
    .A_N(_05002_));
 sg13g2_nand2_1 _11248_ (.Y(_05217_),
    .A(_05002_),
    .B(_04963_));
 sg13g2_nand3_1 _11249_ (.B(net26),
    .C(_05217_),
    .A(_05216_),
    .Y(_05218_));
 sg13g2_a21oi_1 _11250_ (.A1(net29),
    .A2(_05212_),
    .Y(_05219_),
    .B1(_05132_));
 sg13g2_a21oi_1 _11251_ (.A1(_05218_),
    .A2(_05219_),
    .Y(_05220_),
    .B1(_04690_));
 sg13g2_a221oi_1 _11252_ (.B2(_05220_),
    .C1(net96),
    .B1(_05215_),
    .A1(_04638_),
    .Y(_00168_),
    .A2(_05212_));
 sg13g2_xor2_1 _11253_ (.B(_05069_),
    .A(net95),
    .X(_05222_));
 sg13g2_inv_1 _11254_ (.Y(_05223_),
    .A(_05400_));
 sg13g2_a21oi_1 _11255_ (.A1(_05059_),
    .A2(_05386_),
    .Y(_05224_),
    .B1(net95));
 sg13g2_a21oi_1 _11256_ (.A1(_05223_),
    .A2(_05421_),
    .Y(_05225_),
    .B1(_05224_));
 sg13g2_xnor2_1 _11257_ (.Y(_05226_),
    .A(_05222_),
    .B(_05225_));
 sg13g2_a21oi_1 _11258_ (.A1(_05433_),
    .A2(_05404_),
    .Y(_05227_),
    .B1(_05432_));
 sg13g2_o21ai_1 _11259_ (.B1(_05227_),
    .Y(_05228_),
    .A1(_05430_),
    .A2(_05419_));
 sg13g2_xor2_1 _11260_ (.B(_05429_),
    .A(_05069_),
    .X(_05229_));
 sg13g2_a21oi_1 _11261_ (.A1(_05228_),
    .A2(_05229_),
    .Y(_05230_),
    .B1(_04777_));
 sg13g2_o21ai_1 _11262_ (.B1(_05230_),
    .Y(_05232_),
    .A1(_05228_),
    .A2(_05229_));
 sg13g2_o21ai_1 _11263_ (.B1(_05232_),
    .Y(_05233_),
    .A1(net58),
    .A2(_05226_));
 sg13g2_nand2_1 _11264_ (.Y(_05234_),
    .A(_05233_),
    .B(net28));
 sg13g2_a21oi_1 _11265_ (.A1(net31),
    .A2(_05069_),
    .Y(_05235_),
    .B1(_04866_));
 sg13g2_a21oi_1 _11266_ (.A1(_05234_),
    .A2(_05235_),
    .Y(_00173_),
    .B1(_04710_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _11268_ (.A(net140),
    .X(uio_oe[0]));
 sg13g2_buf_1 _11269_ (.A(net141),
    .X(uio_oe[1]));
 sg13g2_buf_1 _11270_ (.A(net142),
    .X(uio_oe[2]));
 sg13g2_buf_1 _11271_ (.A(net143),
    .X(uio_oe[3]));
 sg13g2_buf_1 _11272_ (.A(net144),
    .X(uio_oe[4]));
 sg13g2_buf_1 _11273_ (.A(net145),
    .X(uio_oe[5]));
 sg13g2_buf_1 _11274_ (.A(net146),
    .X(uio_oe[6]));
 sg13g2_buf_1 _11275_ (.A(net147),
    .X(uio_oe[7]));
 sg13g2_buf_1 _11276_ (.A(net8),
    .X(net1));
 sg13g2_buf_1 _11277_ (.A(net8),
    .X(net2));
 sg13g2_buf_1 _11278_ (.A(net8),
    .X(net3));
 sg13g2_buf_1 _11279_ (.A(net8),
    .X(net4));
 sg13g2_buf_1 _11280_ (.A(net8),
    .X(net5));
 sg13g2_buf_1 _11281_ (.A(net8),
    .X(net6));
 sg13g2_buf_1 _11282_ (.A(net8),
    .X(net7));
 sg13g2_dfrbp_1 \frame_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net148),
    .D(_00073_),
    .Q_N(_00037_),
    .Q(\center_y[0] ));
 sg13g2_dfrbp_1 \frame_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net149),
    .D(_00074_),
    .Q_N(_00012_),
    .Q(\center_x[0] ));
 sg13g2_dfrbp_1 \frame_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net150),
    .D(_00075_),
    .Q_N(_00056_),
    .Q(\center_x[1] ));
 sg13g2_dfrbp_1 \frame_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net151),
    .D(_00076_),
    .Q_N(_00035_),
    .Q(\center_x[2] ));
 sg13g2_dfrbp_1 \frame_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net152),
    .D(_00077_),
    .Q_N(_00033_),
    .Q(\center_x[3] ));
 sg13g2_dfrbp_1 \frame_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net153),
    .D(_00078_),
    .Q_N(_00029_),
    .Q(\center_x[4] ));
 sg13g2_dfrbp_1 \frame_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net154),
    .D(_00079_),
    .Q_N(_00027_),
    .Q(\center_x[5] ));
 sg13g2_dfrbp_1 \frame_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net155),
    .D(_00080_),
    .Q_N(_00026_),
    .Q(\frame_counter[7] ));
 sg13g2_dfrbp_1 \frame_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_30__leaf_clk),
    .RESET_B(net156),
    .D(_00081_),
    .Q_N(_00018_),
    .Q(\frame_counter[8] ));
 sg13g2_dfrbp_1 \frame_counter[9]$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net157),
    .D(_00082_),
    .Q_N(_00036_),
    .Q(\frame_counter[9] ));
 sg13g2_dfrbp_1 \frame_counter_frac$_SDFFE_PN0P_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net158),
    .D(_00083_),
    .Q_N(\envelopeA[0] ),
    .Q(frame_counter_frac));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[0]$_SDFF_PP0_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net159),
    .D(_00084_),
    .Q_N(_00060_),
    .Q(\hvsync_gen.hpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[1]$_SDFF_PP0_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net160),
    .D(_00085_),
    .Q_N(_05680_),
    .Q(\hvsync_gen.hpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[2]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net161),
    .D(_00086_),
    .Q_N(_00034_),
    .Q(\hvsync_gen.hpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[3]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net162),
    .D(_00087_),
    .Q_N(_05679_),
    .Q(\hvsync_gen.hpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[4]$_SDFF_PP0_  (.CLK(clknet_5_28__leaf_clk),
    .RESET_B(net163),
    .D(_00088_),
    .Q_N(_05678_),
    .Q(\hvsync_gen.hpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[5]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net164),
    .D(_00089_),
    .Q_N(_05677_),
    .Q(\hvsync_gen.hpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[6]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net165),
    .D(_00090_),
    .Q_N(_00021_),
    .Q(\hvsync_gen.hpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[7]$_SDFF_PP0_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net166),
    .D(_00091_),
    .Q_N(_00024_),
    .Q(\hvsync_gen.hpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[8]$_SDFF_PP0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net167),
    .D(_00092_),
    .Q_N(_00022_),
    .Q(\hvsync_gen.hpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.hpos[9]$_SDFF_PP0_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net168),
    .D(_00093_),
    .Q_N(_00017_),
    .Q(\hvsync_gen.hpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.hsync$_DFF_P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net169),
    .D(_00010_),
    .Q_N(_05676_),
    .Q(hsync));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net170),
    .D(_00094_),
    .Q_N(_00061_),
    .Q(\hvsync_gen.vpos[0] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_25__leaf_clk),
    .RESET_B(net171),
    .D(_00095_),
    .Q_N(_05675_),
    .Q(\hvsync_gen.vpos[1] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[2]$_SDFFCE_PP0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net172),
    .D(_00096_),
    .Q_N(_05674_),
    .Q(\hvsync_gen.vpos[2] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net173),
    .D(_00097_),
    .Q_N(_05673_),
    .Q(\hvsync_gen.vpos[3] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net174),
    .D(_00098_),
    .Q_N(_00019_),
    .Q(\hvsync_gen.vpos[4] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[5]$_SDFFCE_PP0P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net175),
    .D(_00099_),
    .Q_N(_00020_),
    .Q(\hvsync_gen.vpos[5] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[6]$_SDFFCE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net176),
    .D(_00100_),
    .Q_N(_00023_),
    .Q(\hvsync_gen.vpos[6] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[7]$_SDFFCE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net177),
    .D(_00101_),
    .Q_N(_00025_),
    .Q(\hvsync_gen.vpos[7] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[8]$_SDFFCE_PP0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net178),
    .D(_00102_),
    .Q_N(_05672_),
    .Q(\hvsync_gen.vpos[8] ));
 sg13g2_dfrbp_1 \hvsync_gen.vpos[9]$_SDFFCE_PP0P_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net179),
    .D(_00103_),
    .Q_N(_05690_),
    .Q(\hvsync_gen.vpos[9] ));
 sg13g2_dfrbp_1 \hvsync_gen.vsync$_DFF_P_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net180),
    .D(_00011_),
    .Q_N(_05671_),
    .Q(\hvsync_gen.vsync ));
 sg13g2_dfrbp_1 \noise$_SDFFE_PN0P_  (.CLK(clknet_5_19__leaf_clk),
    .RESET_B(net181),
    .D(_00104_),
    .Q_N(_05670_),
    .Q(noise));
 sg13g2_dfrbp_1 \noise_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net182),
    .D(_00105_),
    .Q_N(_05669_),
    .Q(\noise_counter[0] ));
 sg13g2_dfrbp_1 \noise_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net183),
    .D(_00106_),
    .Q_N(_05668_),
    .Q(\noise_counter[1] ));
 sg13g2_dfrbp_1 \noise_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net184),
    .D(_00107_),
    .Q_N(_05667_),
    .Q(\noise_counter[2] ));
 sg13g2_dfrbp_1 \note$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net185),
    .D(_00108_),
    .Q_N(_00058_),
    .Q(note));
 sg13g2_dfrbp_1 \note2$_SDFFE_PN0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net186),
    .D(_00109_),
    .Q_N(_00059_),
    .Q(note2));
 sg13g2_dfrbp_1 \note2_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net187),
    .D(_00110_),
    .Q_N(_05666_),
    .Q(\note2_counter[0] ));
 sg13g2_dfrbp_1 \note2_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net188),
    .D(_00111_),
    .Q_N(_05665_),
    .Q(\note2_counter[1] ));
 sg13g2_dfrbp_1 \note2_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net189),
    .D(_00112_),
    .Q_N(_05664_),
    .Q(\note2_counter[2] ));
 sg13g2_dfrbp_1 \note2_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net190),
    .D(_00113_),
    .Q_N(_05663_),
    .Q(\note2_counter[3] ));
 sg13g2_dfrbp_1 \note2_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net191),
    .D(_00114_),
    .Q_N(_05662_),
    .Q(\note2_counter[4] ));
 sg13g2_dfrbp_1 \note2_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net192),
    .D(_00115_),
    .Q_N(_05661_),
    .Q(\note2_counter[5] ));
 sg13g2_dfrbp_1 \note2_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net193),
    .D(_00116_),
    .Q_N(_05660_),
    .Q(\note2_counter[6] ));
 sg13g2_dfrbp_1 \note2_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net194),
    .D(_00117_),
    .Q_N(_05659_),
    .Q(\note2_counter[7] ));
 sg13g2_dfrbp_1 \note2_counter[8]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net195),
    .D(_00118_),
    .Q_N(_05691_),
    .Q(\note2_counter[8] ));
 sg13g2_dfrbp_1 \note2_freq[0]$_DFF_P_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net196),
    .D(_00000_),
    .Q_N(_05658_),
    .Q(\note2_freq[0] ));
 sg13g2_dfrbp_1 \note2_freq[1]$_SDFF_PN1_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net197),
    .D(_00119_),
    .Q_N(_05657_),
    .Q(\note2_freq[1] ));
 sg13g2_dfrbp_1 \note2_freq[3]$_SDFF_PN1_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net198),
    .D(_00120_),
    .Q_N(_05692_),
    .Q(\note2_freq[3] ));
 sg13g2_dfrbp_1 \note2_freq[4]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net199),
    .D(_00001_),
    .Q_N(_05693_),
    .Q(\note2_freq[4] ));
 sg13g2_dfrbp_1 \note2_freq[5]$_DFF_P_  (.CLK(clknet_5_9__leaf_clk),
    .RESET_B(net200),
    .D(_00002_),
    .Q_N(_05694_),
    .Q(\note2_freq[5] ));
 sg13g2_dfrbp_1 \note2_freq[6]$_DFF_P_  (.CLK(clknet_5_4__leaf_clk),
    .RESET_B(net201),
    .D(_00003_),
    .Q_N(_05656_),
    .Q(\note2_freq[6] ));
 sg13g2_dfrbp_1 \note2_freq[7]$_SDFF_PP1_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net202),
    .D(_00121_),
    .Q_N(_05695_),
    .Q(\note2_freq[7] ));
 sg13g2_dfrbp_1 \note2_freq[8]$_DFF_P_  (.CLK(clknet_5_7__leaf_clk),
    .RESET_B(net203),
    .D(_00004_),
    .Q_N(_05655_),
    .Q(\note2_freq[8] ));
 sg13g2_dfrbp_1 \note_counter[0]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net204),
    .D(_00122_),
    .Q_N(_05654_),
    .Q(\note_counter[0] ));
 sg13g2_dfrbp_1 \note_counter[1]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net205),
    .D(_00123_),
    .Q_N(_05653_),
    .Q(\note_counter[1] ));
 sg13g2_dfrbp_1 \note_counter[2]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net206),
    .D(_00124_),
    .Q_N(_05652_),
    .Q(\note_counter[2] ));
 sg13g2_dfrbp_1 \note_counter[3]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net207),
    .D(_00125_),
    .Q_N(_05651_),
    .Q(\note_counter[3] ));
 sg13g2_dfrbp_1 \note_counter[4]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net208),
    .D(_00126_),
    .Q_N(_05650_),
    .Q(\note_counter[4] ));
 sg13g2_dfrbp_1 \note_counter[5]$_SDFFE_PN0P_  (.CLK(clknet_5_0__leaf_clk),
    .RESET_B(net209),
    .D(_00127_),
    .Q_N(_05649_),
    .Q(\note_counter[5] ));
 sg13g2_dfrbp_1 \note_counter[6]$_SDFFE_PN0P_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net210),
    .D(_00128_),
    .Q_N(_05648_),
    .Q(\note_counter[6] ));
 sg13g2_dfrbp_1 \note_counter[7]$_SDFFE_PN0P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net211),
    .D(_00129_),
    .Q_N(_05647_),
    .Q(\note_counter[7] ));
 sg13g2_dfrbp_1 \note_freq[0]$_SDFF_PN1_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net212),
    .D(_00130_),
    .Q_N(_05696_),
    .Q(\note_freq[0] ));
 sg13g2_dfrbp_1 \note_freq[2]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net213),
    .D(_00005_),
    .Q_N(_05646_),
    .Q(\note_freq[2] ));
 sg13g2_dfrbp_1 \note_freq[3]$_SDFF_PN1_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net214),
    .D(_00131_),
    .Q_N(_05697_),
    .Q(\note_freq[1] ));
 sg13g2_dfrbp_1 \note_freq[4]$_DFF_P_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net215),
    .D(_00006_),
    .Q_N(_05698_),
    .Q(\note_freq[4] ));
 sg13g2_dfrbp_1 \note_freq[5]$_DFF_P_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net216),
    .D(_00007_),
    .Q_N(_05699_),
    .Q(\note_freq[5] ));
 sg13g2_dfrbp_1 \note_freq[6]$_DFF_P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net217),
    .D(_00008_),
    .Q_N(_05700_),
    .Q(\note_freq[6] ));
 sg13g2_dfrbp_1 \note_freq[7]$_DFF_P_  (.CLK(clknet_5_1__leaf_clk),
    .RESET_B(net218),
    .D(_00009_),
    .Q_N(_05645_),
    .Q(\note_freq[7] ));
 sg13g2_dfrbp_1 \r1[0]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net219),
    .D(_00132_),
    .Q_N(_00031_),
    .Q(\r1[0] ));
 sg13g2_dfrbp_1 \r1[10]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net220),
    .D(_00133_),
    .Q_N(_00041_),
    .Q(\r1[10] ));
 sg13g2_dfrbp_1 \r1[11]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net221),
    .D(_00134_),
    .Q_N(_00049_),
    .Q(\r1[11] ));
 sg13g2_dfrbp_1 \r1[12]$_SDFF_PN0_  (.CLK(clknet_5_3__leaf_clk),
    .RESET_B(net222),
    .D(_00135_),
    .Q_N(_00048_),
    .Q(\r1[12] ));
 sg13g2_dfrbp_1 \r1[13]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net223),
    .D(_00136_),
    .Q_N(_00047_),
    .Q(\r1[13] ));
 sg13g2_dfrbp_1 \r1[14]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net224),
    .D(_00137_),
    .Q_N(_00045_),
    .Q(\r1[14] ));
 sg13g2_dfrbp_1 \r1[15]$_SDFF_PN0_  (.CLK(clknet_5_6__leaf_clk),
    .RESET_B(net225),
    .D(_00138_),
    .Q_N(_00039_),
    .Q(\r1[15] ));
 sg13g2_dfrbp_1 \r1[16]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net226),
    .D(_00139_),
    .Q_N(_00014_),
    .Q(\r1[16] ));
 sg13g2_dfrbp_1 \r1[17]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net227),
    .D(_00140_),
    .Q_N(_00016_),
    .Q(\r1[17] ));
 sg13g2_dfrbp_1 \r1[1]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net228),
    .D(_00141_),
    .Q_N(_05644_),
    .Q(\r1[1] ));
 sg13g2_dfrbp_1 \r1[2]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net229),
    .D(_00142_),
    .Q_N(_05643_),
    .Q(\r1[2] ));
 sg13g2_dfrbp_1 \r1[3]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net230),
    .D(_00143_),
    .Q_N(_05642_),
    .Q(\r1[3] ));
 sg13g2_dfrbp_1 \r1[4]$_SDFF_PN0_  (.CLK(clknet_5_11__leaf_clk),
    .RESET_B(net231),
    .D(_00144_),
    .Q_N(_05641_),
    .Q(\r1[4] ));
 sg13g2_dfrbp_1 \r1[5]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net232),
    .D(_00145_),
    .Q_N(_00032_),
    .Q(\r1[5] ));
 sg13g2_dfrbp_1 \r1[6]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net233),
    .D(_00146_),
    .Q_N(_00043_),
    .Q(\r1[6] ));
 sg13g2_dfrbp_1 \r1[7]$_SDFF_PN0_  (.CLK(clknet_5_10__leaf_clk),
    .RESET_B(net234),
    .D(_00147_),
    .Q_N(_00044_),
    .Q(\r1[7] ));
 sg13g2_dfrbp_1 \r1[8]$_SDFF_PN0_  (.CLK(clknet_5_8__leaf_clk),
    .RESET_B(net235),
    .D(_00148_),
    .Q_N(_00042_),
    .Q(\r1[8] ));
 sg13g2_dfrbp_1 \r1[9]$_SDFF_PN0_  (.CLK(clknet_5_2__leaf_clk),
    .RESET_B(net236),
    .D(_00149_),
    .Q_N(_00040_),
    .Q(\r1[9] ));
 sg13g2_dfrbp_1 \r2[0]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net237),
    .D(_00150_),
    .Q_N(_05640_),
    .Q(\r2[0] ));
 sg13g2_dfrbp_1 \r2[10]$_SDFF_PN0_  (.CLK(clknet_5_13__leaf_clk),
    .RESET_B(net238),
    .D(_00151_),
    .Q_N(_05639_),
    .Q(\r2[10] ));
 sg13g2_dfrbp_1 \r2[11]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net239),
    .D(_00152_),
    .Q_N(_05638_),
    .Q(\r2[11] ));
 sg13g2_dfrbp_1 \r2[12]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net240),
    .D(_00153_),
    .Q_N(_00030_),
    .Q(\r2[12] ));
 sg13g2_dfrbp_1 \r2[13]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net241),
    .D(_00154_),
    .Q_N(_05637_),
    .Q(\r2[13] ));
 sg13g2_dfrbp_1 \r2[14]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net242),
    .D(_00155_),
    .Q_N(_05636_),
    .Q(\r2[14] ));
 sg13g2_dfrbp_1 \r2[15]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net243),
    .D(_00156_),
    .Q_N(_00046_),
    .Q(\r2[15] ));
 sg13g2_dfrbp_1 \r2[16]$_SDFF_PN0_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net244),
    .D(_00157_),
    .Q_N(_00038_),
    .Q(\r2[16] ));
 sg13g2_dfrbp_1 \r2[17]$_SDFF_PN0_  (.CLK(clknet_5_5__leaf_clk),
    .RESET_B(net245),
    .D(_00158_),
    .Q_N(_00013_),
    .Q(\r2[17] ));
 sg13g2_dfrbp_1 \r2[18]$_SDFF_PN0_  (.CLK(clknet_5_12__leaf_clk),
    .RESET_B(net246),
    .D(_00159_),
    .Q_N(_00015_),
    .Q(\r2[18] ));
 sg13g2_dfrbp_1 \r2[1]$_SDFF_PN0_  (.CLK(clknet_5_26__leaf_clk),
    .RESET_B(net247),
    .D(_00160_),
    .Q_N(_05635_),
    .Q(\r2[1] ));
 sg13g2_dfrbp_1 \r2[2]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net248),
    .D(_00161_),
    .Q_N(_00057_),
    .Q(\r2[2] ));
 sg13g2_dfrbp_1 \r2[3]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net249),
    .D(_00162_),
    .Q_N(_00055_),
    .Q(\r2[3] ));
 sg13g2_dfrbp_1 \r2[4]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net250),
    .D(_00163_),
    .Q_N(_00054_),
    .Q(\r2[4] ));
 sg13g2_dfrbp_1 \r2[5]$_SDFF_PN0_  (.CLK(clknet_5_14__leaf_clk),
    .RESET_B(net251),
    .D(_00164_),
    .Q_N(_00053_),
    .Q(\r2[5] ));
 sg13g2_dfrbp_1 \r2[6]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net252),
    .D(_00165_),
    .Q_N(_00052_),
    .Q(\r2[6] ));
 sg13g2_dfrbp_1 \r2[7]$_SDFF_PN0_  (.CLK(clknet_5_15__leaf_clk),
    .RESET_B(net253),
    .D(_00166_),
    .Q_N(_00051_),
    .Q(\r2[7] ));
 sg13g2_dfrbp_1 \r2[8]$_SDFF_PN0_  (.CLK(clknet_5_27__leaf_clk),
    .RESET_B(net254),
    .D(_00167_),
    .Q_N(_00050_),
    .Q(\r2[8] ));
 sg13g2_dfrbp_1 \r2[9]$_SDFF_PN0_  (.CLK(clknet_5_18__leaf_clk),
    .RESET_B(net255),
    .D(_00168_),
    .Q_N(_00028_),
    .Q(\r2[9] ));
 sg13g2_dfrbp_1 \title_r[0]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net256),
    .D(_00169_),
    .Q_N(_00062_),
    .Q(\title_r[0] ));
 sg13g2_dfrbp_1 \title_r[10]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net257),
    .D(_00170_),
    .Q_N(_05634_),
    .Q(\title_r[10] ));
 sg13g2_dfrbp_1 \title_r[11]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net258),
    .D(_00171_),
    .Q_N(_05633_),
    .Q(\title_r[11] ));
 sg13g2_dfrbp_1 \title_r[12]$_SDFFE_PP0P_  (.CLK(clknet_5_17__leaf_clk),
    .RESET_B(net259),
    .D(_00172_),
    .Q_N(_05632_),
    .Q(\title_r[12] ));
 sg13g2_dfrbp_1 \title_r[13]$_SDFFE_PN0P_  (.CLK(clknet_5_16__leaf_clk),
    .RESET_B(net260),
    .D(_00173_),
    .Q_N(_05631_),
    .Q(\title_r[13] ));
 sg13g2_dfrbp_1 \title_r[1]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net261),
    .D(_00174_),
    .Q_N(_05630_),
    .Q(\title_r[1] ));
 sg13g2_dfrbp_1 \title_r[2]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net262),
    .D(_00175_),
    .Q_N(_05629_),
    .Q(\title_r[2] ));
 sg13g2_dfrbp_1 \title_r[3]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net263),
    .D(_00176_),
    .Q_N(_05628_),
    .Q(\title_r[3] ));
 sg13g2_dfrbp_1 \title_r[4]$_SDFFE_PP0P_  (.CLK(clknet_5_21__leaf_clk),
    .RESET_B(net264),
    .D(_00177_),
    .Q_N(_05627_),
    .Q(\title_r[4] ));
 sg13g2_dfrbp_1 \title_r[5]$_SDFFE_PP0P_  (.CLK(clknet_5_22__leaf_clk),
    .RESET_B(net265),
    .D(_00178_),
    .Q_N(_05626_),
    .Q(\title_r[5] ));
 sg13g2_dfrbp_1 \title_r[6]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net266),
    .D(_00179_),
    .Q_N(_05625_),
    .Q(\title_r[6] ));
 sg13g2_dfrbp_1 \title_r[7]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net267),
    .D(_00180_),
    .Q_N(_05624_),
    .Q(\title_r[7] ));
 sg13g2_dfrbp_1 \title_r[8]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net268),
    .D(_00181_),
    .Q_N(_05623_),
    .Q(\title_r[8] ));
 sg13g2_dfrbp_1 \title_r[9]$_SDFFE_PP0P_  (.CLK(clknet_5_20__leaf_clk),
    .RESET_B(net269),
    .D(_00182_),
    .Q_N(_05622_),
    .Q(\title_r[9] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[0]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net270),
    .D(_00183_),
    .Q_N(_00063_),
    .Q(\title_r_pixels_in_scanline[0] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[1]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net271),
    .D(_00184_),
    .Q_N(_05621_),
    .Q(\title_r_pixels_in_scanline[1] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[2]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net272),
    .D(_00185_),
    .Q_N(_05620_),
    .Q(\title_r_pixels_in_scanline[2] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[3]$_SDFFCE_PP0P_  (.CLK(clknet_5_29__leaf_clk),
    .RESET_B(net273),
    .D(_00186_),
    .Q_N(_05619_),
    .Q(\title_r_pixels_in_scanline[3] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[4]$_SDFFCE_PP0P_  (.CLK(clknet_5_24__leaf_clk),
    .RESET_B(net274),
    .D(_00187_),
    .Q_N(_05618_),
    .Q(\title_r_pixels_in_scanline[4] ));
 sg13g2_dfrbp_1 \title_r_pixels_in_scanline[5]$_SDFFCE_PP0P_  (.CLK(clknet_5_23__leaf_clk),
    .RESET_B(net275),
    .D(_00188_),
    .Q_N(_05617_),
    .Q(\title_r_pixels_in_scanline[5] ));
 sg13g2_buf_1 output1 (.A(net1),
    .X(uio_out[0]));
 sg13g2_buf_1 output2 (.A(net2),
    .X(uio_out[1]));
 sg13g2_buf_1 output3 (.A(net3),
    .X(uio_out[2]));
 sg13g2_buf_1 output4 (.A(net4),
    .X(uio_out[3]));
 sg13g2_buf_1 output5 (.A(net5),
    .X(uio_out[4]));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uio_out[5]));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uio_out[6]));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uio_out[7]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[0]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[1]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[2]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[3]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[4]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[5]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[6]));
 sg13g2_buf_1 output16 (.A(net16),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout17 (.A(_04119_),
    .X(net17));
 sg13g2_buf_4 fanout18 (.X(net18),
    .A(_02102_));
 sg13g2_buf_2 fanout19 (.A(_02018_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_01976_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_04580_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_04930_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_04542_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_04639_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_04548_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_04879_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_04874_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_05384_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_04873_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_04691_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_05273_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_05113_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_04708_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_04707_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_04690_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_04638_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_05274_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_04889_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_04703_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_04886_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_04875_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_04761_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_04552_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_01112_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_00232_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_04385_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_03553_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_03216_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_00649_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_00231_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_00207_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_05172_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_04361_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_04354_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_04061_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_01502_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_05567_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_05380_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_03365_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_03313_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_01817_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_00551_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_00325_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_00202_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_00193_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_03593_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_01487_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_00610_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_00555_),
    .X(net69));
 sg13g2_buf_4 fanout70 (.X(net70),
    .A(_00201_));
 sg13g2_buf_2 fanout71 (.A(_05565_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_03976_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_02369_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_00432_),
    .X(net74));
 sg13g2_buf_2 fanout75 (.A(_00333_),
    .X(net75));
 sg13g2_buf_2 fanout76 (.A(_05495_),
    .X(net76));
 sg13g2_buf_2 fanout77 (.A(_05262_),
    .X(net77));
 sg13g2_buf_2 fanout78 (.A(_03684_),
    .X(net78));
 sg13g2_buf_2 fanout79 (.A(_04976_),
    .X(net79));
 sg13g2_buf_2 fanout80 (.A(_04730_),
    .X(net80));
 sg13g2_buf_2 fanout81 (.A(_04710_),
    .X(net81));
 sg13g2_buf_2 fanout82 (.A(_04446_),
    .X(net82));
 sg13g2_buf_2 fanout83 (.A(_04323_),
    .X(net83));
 sg13g2_buf_2 fanout84 (.A(_04284_),
    .X(net84));
 sg13g2_buf_2 fanout85 (.A(_03304_),
    .X(net85));
 sg13g2_buf_2 fanout86 (.A(_02737_),
    .X(net86));
 sg13g2_buf_2 fanout87 (.A(_02562_),
    .X(net87));
 sg13g2_buf_2 fanout88 (.A(_02467_),
    .X(net88));
 sg13g2_buf_2 fanout89 (.A(_02458_),
    .X(net89));
 sg13g2_buf_2 fanout90 (.A(_01009_),
    .X(net90));
 sg13g2_buf_2 fanout91 (.A(_05494_),
    .X(net91));
 sg13g2_buf_2 fanout92 (.A(_05486_),
    .X(net92));
 sg13g2_buf_2 fanout93 (.A(_05484_),
    .X(net93));
 sg13g2_buf_2 fanout94 (.A(_05482_),
    .X(net94));
 sg13g2_buf_2 fanout95 (.A(_05259_),
    .X(net95));
 sg13g2_buf_2 fanout96 (.A(_05252_),
    .X(net96));
 sg13g2_buf_2 fanout97 (.A(_04514_),
    .X(net97));
 sg13g2_buf_2 fanout98 (.A(_03256_),
    .X(net98));
 sg13g2_buf_2 fanout99 (.A(_04283_),
    .X(net99));
 sg13g2_buf_2 fanout100 (.A(_02783_),
    .X(net100));
 sg13g2_buf_2 fanout101 (.A(_00412_),
    .X(net101));
 sg13g2_buf_2 fanout102 (.A(_05483_),
    .X(net102));
 sg13g2_buf_2 fanout103 (.A(_04147_),
    .X(net103));
 sg13g2_buf_2 fanout104 (.A(_03921_),
    .X(net104));
 sg13g2_buf_2 fanout105 (.A(_03520_),
    .X(net105));
 sg13g2_buf_2 fanout106 (.A(_03443_),
    .X(net106));
 sg13g2_buf_2 fanout107 (.A(_03421_),
    .X(net107));
 sg13g2_buf_2 fanout108 (.A(_03300_),
    .X(net108));
 sg13g2_buf_2 fanout109 (.A(_03278_),
    .X(net109));
 sg13g2_buf_2 fanout110 (.A(_03245_),
    .X(net110));
 sg13g2_buf_2 fanout111 (.A(_03223_),
    .X(net111));
 sg13g2_buf_2 fanout112 (.A(_02992_),
    .X(net112));
 sg13g2_buf_2 fanout113 (.A(_02839_),
    .X(net113));
 sg13g2_buf_2 fanout114 (.A(_02828_),
    .X(net114));
 sg13g2_buf_2 fanout115 (.A(_02729_),
    .X(net115));
 sg13g2_buf_2 fanout116 (.A(_02608_),
    .X(net116));
 sg13g2_buf_2 fanout117 (.A(_04281_),
    .X(net117));
 sg13g2_buf_2 fanout118 (.A(_03932_),
    .X(net118));
 sg13g2_buf_2 fanout119 (.A(_03432_),
    .X(net119));
 sg13g2_buf_4 fanout120 (.X(net120),
    .A(_03267_));
 sg13g2_buf_2 fanout121 (.A(_03234_),
    .X(net121));
 sg13g2_buf_2 fanout122 (.A(_02959_),
    .X(net122));
 sg13g2_buf_2 fanout123 (.A(_02937_),
    .X(net123));
 sg13g2_buf_2 fanout124 (.A(_02926_),
    .X(net124));
 sg13g2_buf_2 fanout125 (.A(_02641_),
    .X(net125));
 sg13g2_buf_2 fanout126 (.A(_02586_),
    .X(net126));
 sg13g2_buf_2 fanout127 (.A(_02510_),
    .X(net127));
 sg13g2_buf_2 fanout128 (.A(_02477_),
    .X(net128));
 sg13g2_buf_2 fanout129 (.A(_02466_),
    .X(net129));
 sg13g2_buf_2 fanout130 (.A(_02882_),
    .X(net130));
 sg13g2_tiehi \AUDIO_OUT[0]$_SDFF_PN0__131  (.L_HI(net131));
 sg13g2_tiehi \VIDEO_OUT[0]$_SDFF_PN0__132  (.L_HI(net132));
 sg13g2_tiehi \VIDEO_OUT[1]$_SDFF_PN0__133  (.L_HI(net133));
 sg13g2_tiehi \VIDEO_OUT[2]$_SDFF_PN0__134  (.L_HI(net134));
 sg13g2_tiehi \VIDEO_OUT[3]$_SDFF_PN0__135  (.L_HI(net135));
 sg13g2_tiehi \VIDEO_OUT[4]$_SDFF_PN0__136  (.L_HI(net136));
 sg13g2_tiehi \VIDEO_OUT[5]$_SDFF_PN0__137  (.L_HI(net137));
 sg13g2_tiehi \VIDEO_OUT[6]$_SDFF_PN0__138  (.L_HI(net138));
 sg13g2_tiehi \VIDEO_OUT[7]$_SDFF_PN0__139  (.L_HI(net139));
 sg13g2_tiehi _11268__140 (.L_HI(net140));
 sg13g2_tiehi _11269__141 (.L_HI(net141));
 sg13g2_tiehi _11270__142 (.L_HI(net142));
 sg13g2_tiehi _11271__143 (.L_HI(net143));
 sg13g2_tiehi _11272__144 (.L_HI(net144));
 sg13g2_tiehi _11273__145 (.L_HI(net145));
 sg13g2_tiehi _11274__146 (.L_HI(net146));
 sg13g2_tiehi _11275__147 (.L_HI(net147));
 sg13g2_tiehi \frame_counter[0]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \frame_counter[1]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \frame_counter[2]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \frame_counter[3]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \frame_counter[4]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \frame_counter[5]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \frame_counter[6]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \frame_counter[7]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \frame_counter[8]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \frame_counter[9]$_SDFFE_PN0P__157  (.L_HI(net157));
 sg13g2_tiehi \frame_counter_frac$_SDFFE_PN0P__158  (.L_HI(net158));
 sg13g2_tiehi \hvsync_gen.hpos[0]$_SDFF_PP0__159  (.L_HI(net159));
 sg13g2_tiehi \hvsync_gen.hpos[1]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \hvsync_gen.hpos[2]$_SDFF_PP0__161  (.L_HI(net161));
 sg13g2_tiehi \hvsync_gen.hpos[3]$_SDFF_PP0__162  (.L_HI(net162));
 sg13g2_tiehi \hvsync_gen.hpos[4]$_SDFF_PP0__163  (.L_HI(net163));
 sg13g2_tiehi \hvsync_gen.hpos[5]$_SDFF_PP0__164  (.L_HI(net164));
 sg13g2_tiehi \hvsync_gen.hpos[6]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \hvsync_gen.hpos[7]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \hvsync_gen.hpos[8]$_SDFF_PP0__167  (.L_HI(net167));
 sg13g2_tiehi \hvsync_gen.hpos[9]$_SDFF_PP0__168  (.L_HI(net168));
 sg13g2_tiehi \hvsync_gen.hsync$_DFF_P__169  (.L_HI(net169));
 sg13g2_tiehi \hvsync_gen.vpos[0]$_SDFFCE_PP0P__170  (.L_HI(net170));
 sg13g2_tiehi \hvsync_gen.vpos[1]$_SDFFCE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \hvsync_gen.vpos[2]$_SDFFCE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \hvsync_gen.vpos[3]$_SDFFCE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \hvsync_gen.vpos[4]$_SDFFCE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \hvsync_gen.vpos[5]$_SDFFCE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \hvsync_gen.vpos[6]$_SDFFCE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \hvsync_gen.vpos[7]$_SDFFCE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \hvsync_gen.vpos[8]$_SDFFCE_PP0P__178  (.L_HI(net178));
 sg13g2_tiehi \hvsync_gen.vpos[9]$_SDFFCE_PP0P__179  (.L_HI(net179));
 sg13g2_tiehi \hvsync_gen.vsync$_DFF_P__180  (.L_HI(net180));
 sg13g2_tiehi \noise$_SDFFE_PN0P__181  (.L_HI(net181));
 sg13g2_tiehi \noise_counter[0]$_SDFFE_PN0P__182  (.L_HI(net182));
 sg13g2_tiehi \noise_counter[1]$_SDFFE_PN0P__183  (.L_HI(net183));
 sg13g2_tiehi \noise_counter[2]$_SDFFE_PN0P__184  (.L_HI(net184));
 sg13g2_tiehi \note$_SDFFE_PN0P__185  (.L_HI(net185));
 sg13g2_tiehi \note2$_SDFFE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \note2_counter[0]$_SDFFE_PN0P__187  (.L_HI(net187));
 sg13g2_tiehi \note2_counter[1]$_SDFFE_PN0P__188  (.L_HI(net188));
 sg13g2_tiehi \note2_counter[2]$_SDFFE_PN0P__189  (.L_HI(net189));
 sg13g2_tiehi \note2_counter[3]$_SDFFE_PN0P__190  (.L_HI(net190));
 sg13g2_tiehi \note2_counter[4]$_SDFFE_PN0P__191  (.L_HI(net191));
 sg13g2_tiehi \note2_counter[5]$_SDFFE_PN0P__192  (.L_HI(net192));
 sg13g2_tiehi \note2_counter[6]$_SDFFE_PN0P__193  (.L_HI(net193));
 sg13g2_tiehi \note2_counter[7]$_SDFFE_PN0P__194  (.L_HI(net194));
 sg13g2_tiehi \note2_counter[8]$_SDFFE_PN0P__195  (.L_HI(net195));
 sg13g2_tiehi \note2_freq[0]$_DFF_P__196  (.L_HI(net196));
 sg13g2_tiehi \note2_freq[1]$_SDFF_PN1__197  (.L_HI(net197));
 sg13g2_tiehi \note2_freq[3]$_SDFF_PN1__198  (.L_HI(net198));
 sg13g2_tiehi \note2_freq[4]$_DFF_P__199  (.L_HI(net199));
 sg13g2_tiehi \note2_freq[5]$_DFF_P__200  (.L_HI(net200));
 sg13g2_tiehi \note2_freq[6]$_DFF_P__201  (.L_HI(net201));
 sg13g2_tiehi \note2_freq[7]$_SDFF_PP1__202  (.L_HI(net202));
 sg13g2_tiehi \note2_freq[8]$_DFF_P__203  (.L_HI(net203));
 sg13g2_tiehi \note_counter[0]$_SDFFE_PN0P__204  (.L_HI(net204));
 sg13g2_tiehi \note_counter[1]$_SDFFE_PN0P__205  (.L_HI(net205));
 sg13g2_tiehi \note_counter[2]$_SDFFE_PN0P__206  (.L_HI(net206));
 sg13g2_tiehi \note_counter[3]$_SDFFE_PN0P__207  (.L_HI(net207));
 sg13g2_tiehi \note_counter[4]$_SDFFE_PN0P__208  (.L_HI(net208));
 sg13g2_tiehi \note_counter[5]$_SDFFE_PN0P__209  (.L_HI(net209));
 sg13g2_tiehi \note_counter[6]$_SDFFE_PN0P__210  (.L_HI(net210));
 sg13g2_tiehi \note_counter[7]$_SDFFE_PN0P__211  (.L_HI(net211));
 sg13g2_tiehi \note_freq[0]$_SDFF_PN1__212  (.L_HI(net212));
 sg13g2_tiehi \note_freq[2]$_DFF_P__213  (.L_HI(net213));
 sg13g2_tiehi \note_freq[3]$_SDFF_PN1__214  (.L_HI(net214));
 sg13g2_tiehi \note_freq[4]$_DFF_P__215  (.L_HI(net215));
 sg13g2_tiehi \note_freq[5]$_DFF_P__216  (.L_HI(net216));
 sg13g2_tiehi \note_freq[6]$_DFF_P__217  (.L_HI(net217));
 sg13g2_tiehi \note_freq[7]$_DFF_P__218  (.L_HI(net218));
 sg13g2_tiehi \r1[0]$_SDFF_PN0__219  (.L_HI(net219));
 sg13g2_tiehi \r1[10]$_SDFF_PN0__220  (.L_HI(net220));
 sg13g2_tiehi \r1[11]$_SDFF_PN0__221  (.L_HI(net221));
 sg13g2_tiehi \r1[12]$_SDFF_PN0__222  (.L_HI(net222));
 sg13g2_tiehi \r1[13]$_SDFF_PN0__223  (.L_HI(net223));
 sg13g2_tiehi \r1[14]$_SDFF_PN0__224  (.L_HI(net224));
 sg13g2_tiehi \r1[15]$_SDFF_PN0__225  (.L_HI(net225));
 sg13g2_tiehi \r1[16]$_SDFF_PN0__226  (.L_HI(net226));
 sg13g2_tiehi \r1[17]$_SDFF_PN0__227  (.L_HI(net227));
 sg13g2_tiehi \r1[1]$_SDFF_PN0__228  (.L_HI(net228));
 sg13g2_tiehi \r1[2]$_SDFF_PN0__229  (.L_HI(net229));
 sg13g2_tiehi \r1[3]$_SDFF_PN0__230  (.L_HI(net230));
 sg13g2_tiehi \r1[4]$_SDFF_PN0__231  (.L_HI(net231));
 sg13g2_tiehi \r1[5]$_SDFF_PN0__232  (.L_HI(net232));
 sg13g2_tiehi \r1[6]$_SDFF_PN0__233  (.L_HI(net233));
 sg13g2_tiehi \r1[7]$_SDFF_PN0__234  (.L_HI(net234));
 sg13g2_tiehi \r1[8]$_SDFF_PN0__235  (.L_HI(net235));
 sg13g2_tiehi \r1[9]$_SDFF_PN0__236  (.L_HI(net236));
 sg13g2_tiehi \r2[0]$_SDFF_PN0__237  (.L_HI(net237));
 sg13g2_tiehi \r2[10]$_SDFF_PN0__238  (.L_HI(net238));
 sg13g2_tiehi \r2[11]$_SDFF_PN0__239  (.L_HI(net239));
 sg13g2_tiehi \r2[12]$_SDFF_PN0__240  (.L_HI(net240));
 sg13g2_tiehi \r2[13]$_SDFF_PN0__241  (.L_HI(net241));
 sg13g2_tiehi \r2[14]$_SDFF_PN0__242  (.L_HI(net242));
 sg13g2_tiehi \r2[15]$_SDFF_PN0__243  (.L_HI(net243));
 sg13g2_tiehi \r2[16]$_SDFF_PN0__244  (.L_HI(net244));
 sg13g2_tiehi \r2[17]$_SDFF_PN0__245  (.L_HI(net245));
 sg13g2_tiehi \r2[18]$_SDFF_PN0__246  (.L_HI(net246));
 sg13g2_tiehi \r2[1]$_SDFF_PN0__247  (.L_HI(net247));
 sg13g2_tiehi \r2[2]$_SDFF_PN0__248  (.L_HI(net248));
 sg13g2_tiehi \r2[3]$_SDFF_PN0__249  (.L_HI(net249));
 sg13g2_tiehi \r2[4]$_SDFF_PN0__250  (.L_HI(net250));
 sg13g2_tiehi \r2[5]$_SDFF_PN0__251  (.L_HI(net251));
 sg13g2_tiehi \r2[6]$_SDFF_PN0__252  (.L_HI(net252));
 sg13g2_tiehi \r2[7]$_SDFF_PN0__253  (.L_HI(net253));
 sg13g2_tiehi \r2[8]$_SDFF_PN0__254  (.L_HI(net254));
 sg13g2_tiehi \r2[9]$_SDFF_PN0__255  (.L_HI(net255));
 sg13g2_tiehi \title_r[0]$_SDFFE_PP0P__256  (.L_HI(net256));
 sg13g2_tiehi \title_r[10]$_SDFFE_PP0P__257  (.L_HI(net257));
 sg13g2_tiehi \title_r[11]$_SDFFE_PP0P__258  (.L_HI(net258));
 sg13g2_tiehi \title_r[12]$_SDFFE_PP0P__259  (.L_HI(net259));
 sg13g2_tiehi \title_r[13]$_SDFFE_PN0P__260  (.L_HI(net260));
 sg13g2_tiehi \title_r[1]$_SDFFE_PP0P__261  (.L_HI(net261));
 sg13g2_tiehi \title_r[2]$_SDFFE_PP0P__262  (.L_HI(net262));
 sg13g2_tiehi \title_r[3]$_SDFFE_PP0P__263  (.L_HI(net263));
 sg13g2_tiehi \title_r[4]$_SDFFE_PP0P__264  (.L_HI(net264));
 sg13g2_tiehi \title_r[5]$_SDFFE_PP0P__265  (.L_HI(net265));
 sg13g2_tiehi \title_r[6]$_SDFFE_PP0P__266  (.L_HI(net266));
 sg13g2_tiehi \title_r[7]$_SDFFE_PP0P__267  (.L_HI(net267));
 sg13g2_tiehi \title_r[8]$_SDFFE_PP0P__268  (.L_HI(net268));
 sg13g2_tiehi \title_r[9]$_SDFFE_PP0P__269  (.L_HI(net269));
 sg13g2_tiehi \title_r_pixels_in_scanline[0]$_SDFFCE_PP0P__270  (.L_HI(net270));
 sg13g2_tiehi \title_r_pixels_in_scanline[1]$_SDFFCE_PP0P__271  (.L_HI(net271));
 sg13g2_tiehi \title_r_pixels_in_scanline[2]$_SDFFCE_PP0P__272  (.L_HI(net272));
 sg13g2_tiehi \title_r_pixels_in_scanline[3]$_SDFFCE_PP0P__273  (.L_HI(net273));
 sg13g2_tiehi \title_r_pixels_in_scanline[4]$_SDFFCE_PP0P__274  (.L_HI(net274));
 sg13g2_tiehi \title_r_pixels_in_scanline[5]$_SDFFCE_PP0P__275  (.L_HI(net275));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sg13g2_buf_1 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sg13g2_buf_1 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sg13g2_buf_1 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sg13g2_buf_1 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sg13g2_buf_1 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sg13g2_buf_1 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sg13g2_buf_1 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sg13g2_buf_1 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sg13g2_buf_1 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sg13g2_buf_1 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sg13g2_buf_1 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sg13g2_buf_1 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sg13g2_buf_1 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sg13g2_buf_1 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sg13g2_buf_1 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sg13g2_buf_1 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sg13g2_buf_1 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sg13g2_buf_1 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sg13g2_buf_1 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sg13g2_buf_1 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sg13g2_buf_1 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sg13g2_buf_1 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sg13g2_buf_1 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sg13g2_buf_1 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sg13g2_buf_1 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sg13g2_buf_1 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sg13g2_buf_1 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sg13g2_buf_1 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sg13g2_buf_1 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sg13g2_buf_1 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sg13g2_buf_1 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_5_1__leaf_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_5_3__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_5_5__leaf_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_5_9__leaf_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_5_13__leaf_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_5_17__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_5_21__leaf_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_5_25__leaf_clk));
 sg13g2_inv_1 clkload8 (.A(clknet_5_29__leaf_clk));
 sg13g2_antennanp ANTENNA_1 (.A(clk));
 sg13g2_antennanp ANTENNA_2 (.A(clk));
 sg13g2_antennanp ANTENNA_3 (.A(clk));
 sg13g2_fill_2 FILLER_0_0 ();
 sg13g2_fill_1 FILLER_0_14 ();
 sg13g2_fill_1 FILLER_0_49 ();
 sg13g2_fill_2 FILLER_0_163 ();
 sg13g2_fill_2 FILLER_0_195 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_220 ();
 sg13g2_fill_1 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_288 ();
 sg13g2_fill_1 FILLER_0_308 ();
 sg13g2_fill_1 FILLER_0_333 ();
 sg13g2_decap_8 FILLER_0_359 ();
 sg13g2_fill_2 FILLER_0_366 ();
 sg13g2_fill_1 FILLER_0_368 ();
 sg13g2_fill_2 FILLER_0_386 ();
 sg13g2_fill_1 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_410 ();
 sg13g2_decap_8 FILLER_0_417 ();
 sg13g2_decap_4 FILLER_0_424 ();
 sg13g2_fill_2 FILLER_0_428 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_55 ();
 sg13g2_fill_1 FILLER_1_193 ();
 sg13g2_fill_1 FILLER_1_208 ();
 sg13g2_fill_1 FILLER_1_228 ();
 sg13g2_fill_1 FILLER_1_256 ();
 sg13g2_fill_1 FILLER_1_261 ();
 sg13g2_fill_2 FILLER_1_284 ();
 sg13g2_fill_1 FILLER_1_291 ();
 sg13g2_fill_2 FILLER_1_299 ();
 sg13g2_fill_2 FILLER_1_310 ();
 sg13g2_fill_1 FILLER_1_316 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_1 FILLER_1_328 ();
 sg13g2_fill_1 FILLER_1_335 ();
 sg13g2_fill_1 FILLER_1_341 ();
 sg13g2_fill_1 FILLER_1_360 ();
 sg13g2_fill_2 FILLER_1_365 ();
 sg13g2_fill_1 FILLER_1_367 ();
 sg13g2_fill_1 FILLER_1_376 ();
 sg13g2_fill_1 FILLER_1_381 ();
 sg13g2_fill_2 FILLER_1_385 ();
 sg13g2_fill_1 FILLER_1_391 ();
 sg13g2_fill_1 FILLER_1_397 ();
 sg13g2_fill_2 FILLER_1_402 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_fill_2 FILLER_1_427 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_fill_1 FILLER_2_214 ();
 sg13g2_fill_2 FILLER_2_227 ();
 sg13g2_fill_1 FILLER_2_263 ();
 sg13g2_fill_1 FILLER_2_272 ();
 sg13g2_fill_1 FILLER_2_277 ();
 sg13g2_fill_1 FILLER_2_283 ();
 sg13g2_fill_1 FILLER_2_311 ();
 sg13g2_fill_1 FILLER_2_317 ();
 sg13g2_fill_1 FILLER_2_348 ();
 sg13g2_fill_2 FILLER_2_356 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_fill_2 FILLER_2_395 ();
 sg13g2_fill_1 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_421 ();
 sg13g2_fill_2 FILLER_2_428 ();
 sg13g2_fill_1 FILLER_3_22 ();
 sg13g2_fill_1 FILLER_3_168 ();
 sg13g2_fill_1 FILLER_3_173 ();
 sg13g2_fill_1 FILLER_3_183 ();
 sg13g2_fill_2 FILLER_3_208 ();
 sg13g2_fill_2 FILLER_3_240 ();
 sg13g2_fill_2 FILLER_3_257 ();
 sg13g2_fill_1 FILLER_3_322 ();
 sg13g2_fill_1 FILLER_3_327 ();
 sg13g2_fill_1 FILLER_3_337 ();
 sg13g2_fill_2 FILLER_3_343 ();
 sg13g2_fill_2 FILLER_3_363 ();
 sg13g2_fill_1 FILLER_3_369 ();
 sg13g2_fill_2 FILLER_3_374 ();
 sg13g2_decap_4 FILLER_3_387 ();
 sg13g2_fill_2 FILLER_3_427 ();
 sg13g2_fill_1 FILLER_3_429 ();
 sg13g2_fill_1 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_50 ();
 sg13g2_fill_1 FILLER_4_59 ();
 sg13g2_fill_1 FILLER_4_65 ();
 sg13g2_fill_1 FILLER_4_71 ();
 sg13g2_fill_1 FILLER_4_76 ();
 sg13g2_fill_2 FILLER_4_114 ();
 sg13g2_fill_1 FILLER_4_200 ();
 sg13g2_fill_2 FILLER_4_215 ();
 sg13g2_fill_1 FILLER_4_221 ();
 sg13g2_fill_1 FILLER_4_233 ();
 sg13g2_fill_1 FILLER_4_239 ();
 sg13g2_fill_2 FILLER_4_248 ();
 sg13g2_fill_2 FILLER_4_269 ();
 sg13g2_fill_1 FILLER_4_284 ();
 sg13g2_fill_1 FILLER_4_289 ();
 sg13g2_fill_1 FILLER_4_338 ();
 sg13g2_fill_1 FILLER_4_356 ();
 sg13g2_fill_1 FILLER_4_361 ();
 sg13g2_fill_1 FILLER_4_366 ();
 sg13g2_fill_1 FILLER_4_376 ();
 sg13g2_fill_1 FILLER_4_381 ();
 sg13g2_fill_1 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_404 ();
 sg13g2_fill_1 FILLER_4_411 ();
 sg13g2_fill_1 FILLER_4_417 ();
 sg13g2_fill_1 FILLER_4_422 ();
 sg13g2_fill_2 FILLER_4_427 ();
 sg13g2_fill_1 FILLER_4_429 ();
 sg13g2_fill_1 FILLER_5_0 ();
 sg13g2_fill_2 FILLER_5_50 ();
 sg13g2_fill_2 FILLER_5_92 ();
 sg13g2_fill_1 FILLER_5_107 ();
 sg13g2_fill_1 FILLER_5_127 ();
 sg13g2_fill_2 FILLER_5_139 ();
 sg13g2_fill_1 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_163 ();
 sg13g2_fill_1 FILLER_5_172 ();
 sg13g2_fill_1 FILLER_5_182 ();
 sg13g2_fill_2 FILLER_5_225 ();
 sg13g2_fill_2 FILLER_5_256 ();
 sg13g2_fill_2 FILLER_5_297 ();
 sg13g2_fill_1 FILLER_5_326 ();
 sg13g2_fill_1 FILLER_5_335 ();
 sg13g2_fill_1 FILLER_5_341 ();
 sg13g2_fill_1 FILLER_5_380 ();
 sg13g2_fill_2 FILLER_5_384 ();
 sg13g2_fill_1 FILLER_5_386 ();
 sg13g2_fill_1 FILLER_5_391 ();
 sg13g2_decap_4 FILLER_5_400 ();
 sg13g2_fill_1 FILLER_5_404 ();
 sg13g2_decap_4 FILLER_5_413 ();
 sg13g2_fill_2 FILLER_6_63 ();
 sg13g2_fill_1 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_99 ();
 sg13g2_fill_1 FILLER_6_111 ();
 sg13g2_fill_1 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_163 ();
 sg13g2_fill_1 FILLER_6_167 ();
 sg13g2_fill_1 FILLER_6_181 ();
 sg13g2_fill_1 FILLER_6_207 ();
 sg13g2_fill_1 FILLER_6_223 ();
 sg13g2_fill_2 FILLER_6_242 ();
 sg13g2_fill_1 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_320 ();
 sg13g2_fill_1 FILLER_6_332 ();
 sg13g2_fill_2 FILLER_6_349 ();
 sg13g2_fill_1 FILLER_6_355 ();
 sg13g2_fill_1 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_365 ();
 sg13g2_fill_1 FILLER_6_371 ();
 sg13g2_fill_2 FILLER_6_376 ();
 sg13g2_fill_1 FILLER_6_382 ();
 sg13g2_fill_1 FILLER_6_395 ();
 sg13g2_fill_2 FILLER_6_399 ();
 sg13g2_fill_2 FILLER_6_409 ();
 sg13g2_fill_1 FILLER_6_411 ();
 sg13g2_fill_2 FILLER_6_418 ();
 sg13g2_fill_1 FILLER_7_30 ();
 sg13g2_fill_1 FILLER_7_35 ();
 sg13g2_fill_1 FILLER_7_160 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_fill_1 FILLER_7_192 ();
 sg13g2_fill_1 FILLER_7_197 ();
 sg13g2_fill_1 FILLER_7_206 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_fill_1 FILLER_7_236 ();
 sg13g2_fill_2 FILLER_7_252 ();
 sg13g2_fill_2 FILLER_7_284 ();
 sg13g2_fill_1 FILLER_7_319 ();
 sg13g2_fill_1 FILLER_7_338 ();
 sg13g2_fill_2 FILLER_7_347 ();
 sg13g2_fill_2 FILLER_7_362 ();
 sg13g2_fill_2 FILLER_7_383 ();
 sg13g2_fill_1 FILLER_7_389 ();
 sg13g2_fill_1 FILLER_7_411 ();
 sg13g2_fill_1 FILLER_7_424 ();
 sg13g2_fill_2 FILLER_8_21 ();
 sg13g2_fill_1 FILLER_8_104 ();
 sg13g2_fill_2 FILLER_8_146 ();
 sg13g2_fill_1 FILLER_8_191 ();
 sg13g2_fill_1 FILLER_8_196 ();
 sg13g2_fill_1 FILLER_8_208 ();
 sg13g2_fill_1 FILLER_8_217 ();
 sg13g2_fill_1 FILLER_8_240 ();
 sg13g2_fill_2 FILLER_8_254 ();
 sg13g2_fill_1 FILLER_8_261 ();
 sg13g2_fill_1 FILLER_8_267 ();
 sg13g2_fill_1 FILLER_8_295 ();
 sg13g2_fill_2 FILLER_8_314 ();
 sg13g2_fill_2 FILLER_8_330 ();
 sg13g2_decap_4 FILLER_8_355 ();
 sg13g2_fill_2 FILLER_8_359 ();
 sg13g2_decap_4 FILLER_8_366 ();
 sg13g2_decap_8 FILLER_8_374 ();
 sg13g2_fill_2 FILLER_8_388 ();
 sg13g2_fill_1 FILLER_8_409 ();
 sg13g2_fill_1 FILLER_8_415 ();
 sg13g2_fill_1 FILLER_8_419 ();
 sg13g2_fill_1 FILLER_8_425 ();
 sg13g2_fill_1 FILLER_9_26 ();
 sg13g2_fill_1 FILLER_9_33 ();
 sg13g2_fill_1 FILLER_9_44 ();
 sg13g2_fill_1 FILLER_9_80 ();
 sg13g2_fill_1 FILLER_9_85 ();
 sg13g2_fill_1 FILLER_9_114 ();
 sg13g2_fill_2 FILLER_9_120 ();
 sg13g2_fill_1 FILLER_9_142 ();
 sg13g2_fill_1 FILLER_9_181 ();
 sg13g2_fill_2 FILLER_9_217 ();
 sg13g2_fill_1 FILLER_9_224 ();
 sg13g2_fill_1 FILLER_9_233 ();
 sg13g2_fill_1 FILLER_9_275 ();
 sg13g2_decap_4 FILLER_9_284 ();
 sg13g2_fill_1 FILLER_9_288 ();
 sg13g2_fill_1 FILLER_9_302 ();
 sg13g2_fill_2 FILLER_9_318 ();
 sg13g2_fill_2 FILLER_9_329 ();
 sg13g2_fill_2 FILLER_9_355 ();
 sg13g2_fill_1 FILLER_9_365 ();
 sg13g2_fill_1 FILLER_9_371 ();
 sg13g2_fill_1 FILLER_9_401 ();
 sg13g2_fill_2 FILLER_9_406 ();
 sg13g2_decap_4 FILLER_9_425 ();
 sg13g2_fill_1 FILLER_9_429 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_fill_2 FILLER_10_123 ();
 sg13g2_fill_1 FILLER_10_130 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_fill_1 FILLER_10_148 ();
 sg13g2_fill_2 FILLER_10_154 ();
 sg13g2_fill_1 FILLER_10_160 ();
 sg13g2_fill_1 FILLER_10_187 ();
 sg13g2_fill_1 FILLER_10_193 ();
 sg13g2_fill_1 FILLER_10_202 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_222 ();
 sg13g2_fill_2 FILLER_10_264 ();
 sg13g2_fill_1 FILLER_10_271 ();
 sg13g2_decap_4 FILLER_10_277 ();
 sg13g2_fill_2 FILLER_10_286 ();
 sg13g2_fill_1 FILLER_10_313 ();
 sg13g2_fill_1 FILLER_10_318 ();
 sg13g2_fill_1 FILLER_10_324 ();
 sg13g2_decap_4 FILLER_10_340 ();
 sg13g2_fill_1 FILLER_10_348 ();
 sg13g2_fill_2 FILLER_10_356 ();
 sg13g2_fill_1 FILLER_10_361 ();
 sg13g2_fill_1 FILLER_10_365 ();
 sg13g2_fill_1 FILLER_10_422 ();
 sg13g2_fill_1 FILLER_11_74 ();
 sg13g2_fill_2 FILLER_11_115 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_fill_1 FILLER_11_172 ();
 sg13g2_fill_1 FILLER_11_177 ();
 sg13g2_fill_1 FILLER_11_191 ();
 sg13g2_fill_1 FILLER_11_196 ();
 sg13g2_fill_1 FILLER_11_202 ();
 sg13g2_fill_1 FILLER_11_211 ();
 sg13g2_fill_1 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_225 ();
 sg13g2_fill_1 FILLER_11_230 ();
 sg13g2_fill_1 FILLER_11_235 ();
 sg13g2_decap_4 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_254 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_1 FILLER_11_332 ();
 sg13g2_fill_1 FILLER_11_342 ();
 sg13g2_fill_1 FILLER_11_352 ();
 sg13g2_fill_2 FILLER_11_363 ();
 sg13g2_fill_1 FILLER_11_369 ();
 sg13g2_fill_1 FILLER_12_8 ();
 sg13g2_fill_1 FILLER_12_76 ();
 sg13g2_fill_2 FILLER_12_102 ();
 sg13g2_fill_2 FILLER_12_112 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_164 ();
 sg13g2_fill_1 FILLER_12_226 ();
 sg13g2_fill_1 FILLER_12_246 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_279 ();
 sg13g2_fill_2 FILLER_12_284 ();
 sg13g2_fill_2 FILLER_12_291 ();
 sg13g2_fill_2 FILLER_12_297 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_337 ();
 sg13g2_fill_1 FILLER_12_343 ();
 sg13g2_fill_1 FILLER_12_364 ();
 sg13g2_fill_1 FILLER_12_369 ();
 sg13g2_fill_1 FILLER_12_374 ();
 sg13g2_fill_1 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_389 ();
 sg13g2_fill_2 FILLER_12_394 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_1 FILLER_13_35 ();
 sg13g2_fill_2 FILLER_13_62 ();
 sg13g2_fill_2 FILLER_13_80 ();
 sg13g2_fill_1 FILLER_13_132 ();
 sg13g2_fill_2 FILLER_13_178 ();
 sg13g2_fill_1 FILLER_13_193 ();
 sg13g2_decap_8 FILLER_13_237 ();
 sg13g2_fill_1 FILLER_13_248 ();
 sg13g2_fill_1 FILLER_13_261 ();
 sg13g2_fill_1 FILLER_13_265 ();
 sg13g2_fill_1 FILLER_13_290 ();
 sg13g2_fill_1 FILLER_13_295 ();
 sg13g2_fill_2 FILLER_13_360 ();
 sg13g2_fill_1 FILLER_13_375 ();
 sg13g2_decap_4 FILLER_13_388 ();
 sg13g2_fill_1 FILLER_13_400 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_94 ();
 sg13g2_fill_1 FILLER_14_178 ();
 sg13g2_fill_2 FILLER_14_203 ();
 sg13g2_decap_4 FILLER_14_226 ();
 sg13g2_fill_2 FILLER_14_230 ();
 sg13g2_fill_1 FILLER_14_237 ();
 sg13g2_fill_2 FILLER_14_243 ();
 sg13g2_fill_1 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_250 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_fill_2 FILLER_14_285 ();
 sg13g2_decap_4 FILLER_14_299 ();
 sg13g2_fill_1 FILLER_14_332 ();
 sg13g2_fill_2 FILLER_14_376 ();
 sg13g2_fill_1 FILLER_14_378 ();
 sg13g2_decap_4 FILLER_14_388 ();
 sg13g2_fill_1 FILLER_14_392 ();
 sg13g2_fill_2 FILLER_14_410 ();
 sg13g2_fill_2 FILLER_14_417 ();
 sg13g2_fill_1 FILLER_14_419 ();
 sg13g2_fill_1 FILLER_14_423 ();
 sg13g2_fill_2 FILLER_14_428 ();
 sg13g2_fill_1 FILLER_15_9 ();
 sg13g2_fill_2 FILLER_15_76 ();
 sg13g2_fill_1 FILLER_15_86 ();
 sg13g2_fill_1 FILLER_15_127 ();
 sg13g2_fill_1 FILLER_15_141 ();
 sg13g2_fill_1 FILLER_15_150 ();
 sg13g2_fill_1 FILLER_15_155 ();
 sg13g2_fill_2 FILLER_15_213 ();
 sg13g2_fill_1 FILLER_15_215 ();
 sg13g2_fill_1 FILLER_15_219 ();
 sg13g2_fill_2 FILLER_15_224 ();
 sg13g2_decap_4 FILLER_15_229 ();
 sg13g2_fill_2 FILLER_15_238 ();
 sg13g2_fill_1 FILLER_15_243 ();
 sg13g2_fill_2 FILLER_15_249 ();
 sg13g2_fill_1 FILLER_15_251 ();
 sg13g2_fill_2 FILLER_15_277 ();
 sg13g2_fill_1 FILLER_15_279 ();
 sg13g2_decap_4 FILLER_15_284 ();
 sg13g2_fill_1 FILLER_15_288 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_fill_2 FILLER_15_335 ();
 sg13g2_fill_1 FILLER_15_337 ();
 sg13g2_fill_1 FILLER_15_349 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_365 ();
 sg13g2_fill_1 FILLER_15_367 ();
 sg13g2_fill_1 FILLER_15_388 ();
 sg13g2_fill_2 FILLER_15_405 ();
 sg13g2_fill_1 FILLER_15_407 ();
 sg13g2_decap_4 FILLER_15_417 ();
 sg13g2_fill_1 FILLER_15_429 ();
 sg13g2_fill_2 FILLER_16_8 ();
 sg13g2_fill_2 FILLER_16_41 ();
 sg13g2_fill_1 FILLER_16_89 ();
 sg13g2_fill_1 FILLER_16_115 ();
 sg13g2_fill_2 FILLER_16_190 ();
 sg13g2_fill_2 FILLER_16_206 ();
 sg13g2_fill_2 FILLER_16_213 ();
 sg13g2_decap_4 FILLER_16_219 ();
 sg13g2_fill_1 FILLER_16_223 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_1 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_284 ();
 sg13g2_fill_1 FILLER_16_319 ();
 sg13g2_fill_1 FILLER_16_329 ();
 sg13g2_fill_1 FILLER_16_338 ();
 sg13g2_fill_2 FILLER_16_383 ();
 sg13g2_fill_1 FILLER_16_385 ();
 sg13g2_fill_1 FILLER_16_394 ();
 sg13g2_fill_1 FILLER_16_399 ();
 sg13g2_fill_1 FILLER_16_405 ();
 sg13g2_fill_1 FILLER_16_419 ();
 sg13g2_fill_2 FILLER_16_428 ();
 sg13g2_fill_1 FILLER_17_38 ();
 sg13g2_fill_2 FILLER_17_59 ();
 sg13g2_fill_1 FILLER_17_70 ();
 sg13g2_fill_2 FILLER_17_75 ();
 sg13g2_fill_1 FILLER_17_88 ();
 sg13g2_fill_1 FILLER_17_96 ();
 sg13g2_fill_1 FILLER_17_119 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_2 FILLER_17_172 ();
 sg13g2_fill_2 FILLER_17_232 ();
 sg13g2_fill_1 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_276 ();
 sg13g2_fill_2 FILLER_17_280 ();
 sg13g2_fill_2 FILLER_17_308 ();
 sg13g2_fill_1 FILLER_17_310 ();
 sg13g2_decap_4 FILLER_17_330 ();
 sg13g2_fill_2 FILLER_17_428 ();
 sg13g2_fill_1 FILLER_18_13 ();
 sg13g2_fill_1 FILLER_18_44 ();
 sg13g2_fill_1 FILLER_18_50 ();
 sg13g2_fill_1 FILLER_18_56 ();
 sg13g2_fill_1 FILLER_18_62 ();
 sg13g2_fill_1 FILLER_18_68 ();
 sg13g2_fill_1 FILLER_18_75 ();
 sg13g2_fill_2 FILLER_18_107 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_1 FILLER_18_127 ();
 sg13g2_fill_1 FILLER_18_132 ();
 sg13g2_fill_2 FILLER_18_146 ();
 sg13g2_fill_2 FILLER_18_204 ();
 sg13g2_fill_2 FILLER_18_219 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_fill_1 FILLER_18_231 ();
 sg13g2_fill_2 FILLER_18_236 ();
 sg13g2_fill_2 FILLER_18_242 ();
 sg13g2_fill_2 FILLER_18_249 ();
 sg13g2_fill_1 FILLER_18_266 ();
 sg13g2_fill_1 FILLER_18_287 ();
 sg13g2_fill_2 FILLER_18_292 ();
 sg13g2_fill_2 FILLER_18_298 ();
 sg13g2_fill_2 FILLER_18_304 ();
 sg13g2_fill_1 FILLER_18_306 ();
 sg13g2_fill_1 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_349 ();
 sg13g2_fill_1 FILLER_18_354 ();
 sg13g2_fill_1 FILLER_18_376 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_1 FILLER_18_392 ();
 sg13g2_fill_1 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_406 ();
 sg13g2_fill_1 FILLER_18_429 ();
 sg13g2_fill_2 FILLER_19_0 ();
 sg13g2_fill_1 FILLER_19_75 ();
 sg13g2_fill_1 FILLER_19_96 ();
 sg13g2_fill_1 FILLER_19_135 ();
 sg13g2_fill_2 FILLER_19_140 ();
 sg13g2_fill_2 FILLER_19_216 ();
 sg13g2_fill_2 FILLER_19_223 ();
 sg13g2_fill_2 FILLER_19_261 ();
 sg13g2_fill_1 FILLER_19_297 ();
 sg13g2_fill_2 FILLER_19_304 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_315 ();
 sg13g2_fill_2 FILLER_19_367 ();
 sg13g2_fill_1 FILLER_19_396 ();
 sg13g2_fill_2 FILLER_19_424 ();
 sg13g2_fill_1 FILLER_20_34 ();
 sg13g2_fill_1 FILLER_20_51 ();
 sg13g2_fill_2 FILLER_20_65 ();
 sg13g2_fill_1 FILLER_20_71 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_123 ();
 sg13g2_fill_2 FILLER_20_163 ();
 sg13g2_fill_2 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_185 ();
 sg13g2_fill_1 FILLER_20_192 ();
 sg13g2_decap_8 FILLER_20_206 ();
 sg13g2_fill_2 FILLER_20_216 ();
 sg13g2_fill_2 FILLER_20_222 ();
 sg13g2_fill_1 FILLER_20_228 ();
 sg13g2_fill_2 FILLER_20_233 ();
 sg13g2_decap_4 FILLER_20_240 ();
 sg13g2_fill_2 FILLER_20_244 ();
 sg13g2_fill_1 FILLER_20_250 ();
 sg13g2_fill_2 FILLER_20_255 ();
 sg13g2_fill_2 FILLER_20_285 ();
 sg13g2_fill_1 FILLER_20_287 ();
 sg13g2_fill_2 FILLER_20_292 ();
 sg13g2_fill_1 FILLER_20_302 ();
 sg13g2_fill_2 FILLER_20_318 ();
 sg13g2_fill_2 FILLER_20_362 ();
 sg13g2_fill_1 FILLER_20_374 ();
 sg13g2_fill_2 FILLER_20_400 ();
 sg13g2_fill_2 FILLER_20_407 ();
 sg13g2_fill_1 FILLER_20_409 ();
 sg13g2_fill_2 FILLER_20_424 ();
 sg13g2_fill_1 FILLER_21_39 ();
 sg13g2_fill_1 FILLER_21_45 ();
 sg13g2_fill_1 FILLER_21_125 ();
 sg13g2_fill_1 FILLER_21_145 ();
 sg13g2_fill_1 FILLER_21_151 ();
 sg13g2_fill_1 FILLER_21_156 ();
 sg13g2_fill_2 FILLER_21_187 ();
 sg13g2_fill_2 FILLER_21_197 ();
 sg13g2_fill_2 FILLER_21_212 ();
 sg13g2_fill_1 FILLER_21_251 ();
 sg13g2_fill_1 FILLER_21_256 ();
 sg13g2_fill_2 FILLER_21_266 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_decap_4 FILLER_21_299 ();
 sg13g2_fill_1 FILLER_21_303 ();
 sg13g2_fill_1 FILLER_21_370 ();
 sg13g2_fill_2 FILLER_21_391 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_21_414 ();
 sg13g2_fill_1 FILLER_22_47 ();
 sg13g2_fill_1 FILLER_22_71 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_fill_1 FILLER_22_83 ();
 sg13g2_fill_1 FILLER_22_89 ();
 sg13g2_fill_2 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_122 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_154 ();
 sg13g2_fill_1 FILLER_22_178 ();
 sg13g2_fill_2 FILLER_22_209 ();
 sg13g2_fill_1 FILLER_22_211 ();
 sg13g2_fill_2 FILLER_22_242 ();
 sg13g2_fill_2 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_250 ();
 sg13g2_fill_1 FILLER_22_256 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_1 FILLER_22_325 ();
 sg13g2_fill_2 FILLER_22_337 ();
 sg13g2_fill_1 FILLER_22_348 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_2 FILLER_22_374 ();
 sg13g2_fill_2 FILLER_22_392 ();
 sg13g2_fill_1 FILLER_22_398 ();
 sg13g2_fill_2 FILLER_22_412 ();
 sg13g2_fill_2 FILLER_22_427 ();
 sg13g2_fill_1 FILLER_22_429 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_7 ();
 sg13g2_fill_1 FILLER_23_69 ();
 sg13g2_fill_1 FILLER_23_161 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_188 ();
 sg13g2_fill_2 FILLER_23_200 ();
 sg13g2_decap_8 FILLER_23_206 ();
 sg13g2_decap_8 FILLER_23_213 ();
 sg13g2_decap_4 FILLER_23_220 ();
 sg13g2_fill_1 FILLER_23_224 ();
 sg13g2_fill_1 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_266 ();
 sg13g2_fill_1 FILLER_23_276 ();
 sg13g2_fill_1 FILLER_23_324 ();
 sg13g2_fill_1 FILLER_23_329 ();
 sg13g2_decap_4 FILLER_23_343 ();
 sg13g2_fill_2 FILLER_23_347 ();
 sg13g2_fill_1 FILLER_23_357 ();
 sg13g2_fill_2 FILLER_23_367 ();
 sg13g2_fill_1 FILLER_23_369 ();
 sg13g2_fill_1 FILLER_23_374 ();
 sg13g2_fill_2 FILLER_23_381 ();
 sg13g2_fill_1 FILLER_23_383 ();
 sg13g2_fill_1 FILLER_23_394 ();
 sg13g2_fill_1 FILLER_23_415 ();
 sg13g2_fill_2 FILLER_23_424 ();
 sg13g2_fill_1 FILLER_24_36 ();
 sg13g2_fill_2 FILLER_24_42 ();
 sg13g2_fill_1 FILLER_24_74 ();
 sg13g2_fill_1 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_93 ();
 sg13g2_fill_2 FILLER_24_110 ();
 sg13g2_fill_2 FILLER_24_158 ();
 sg13g2_fill_1 FILLER_24_192 ();
 sg13g2_fill_1 FILLER_24_198 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_2 FILLER_24_211 ();
 sg13g2_fill_1 FILLER_24_231 ();
 sg13g2_fill_2 FILLER_24_241 ();
 sg13g2_fill_1 FILLER_24_243 ();
 sg13g2_fill_2 FILLER_24_249 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_fill_2 FILLER_24_261 ();
 sg13g2_decap_8 FILLER_24_267 ();
 sg13g2_fill_1 FILLER_24_274 ();
 sg13g2_fill_1 FILLER_24_279 ();
 sg13g2_fill_2 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_335 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_386 ();
 sg13g2_fill_2 FILLER_24_412 ();
 sg13g2_fill_2 FILLER_24_418 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_65 ();
 sg13g2_fill_2 FILLER_25_96 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_fill_1 FILLER_25_192 ();
 sg13g2_fill_1 FILLER_25_197 ();
 sg13g2_fill_1 FILLER_25_223 ();
 sg13g2_fill_1 FILLER_25_232 ();
 sg13g2_fill_1 FILLER_25_237 ();
 sg13g2_fill_1 FILLER_25_247 ();
 sg13g2_fill_2 FILLER_25_253 ();
 sg13g2_fill_1 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_266 ();
 sg13g2_fill_2 FILLER_25_289 ();
 sg13g2_fill_1 FILLER_25_377 ();
 sg13g2_fill_2 FILLER_25_388 ();
 sg13g2_fill_1 FILLER_25_411 ();
 sg13g2_decap_8 FILLER_25_419 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_27 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_155 ();
 sg13g2_fill_1 FILLER_26_162 ();
 sg13g2_fill_1 FILLER_26_171 ();
 sg13g2_fill_2 FILLER_26_180 ();
 sg13g2_fill_1 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_186 ();
 sg13g2_fill_1 FILLER_26_191 ();
 sg13g2_fill_1 FILLER_26_196 ();
 sg13g2_fill_1 FILLER_26_210 ();
 sg13g2_fill_2 FILLER_26_214 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_262 ();
 sg13g2_fill_1 FILLER_26_277 ();
 sg13g2_fill_1 FILLER_26_282 ();
 sg13g2_fill_1 FILLER_26_306 ();
 sg13g2_fill_1 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_321 ();
 sg13g2_fill_1 FILLER_26_327 ();
 sg13g2_fill_1 FILLER_26_333 ();
 sg13g2_fill_1 FILLER_26_338 ();
 sg13g2_fill_1 FILLER_26_365 ();
 sg13g2_fill_2 FILLER_26_403 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_2 FILLER_27_59 ();
 sg13g2_fill_1 FILLER_27_99 ();
 sg13g2_fill_2 FILLER_27_135 ();
 sg13g2_fill_1 FILLER_27_171 ();
 sg13g2_decap_4 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_218 ();
 sg13g2_fill_1 FILLER_27_225 ();
 sg13g2_fill_1 FILLER_27_231 ();
 sg13g2_fill_1 FILLER_27_242 ();
 sg13g2_fill_2 FILLER_27_247 ();
 sg13g2_fill_2 FILLER_27_257 ();
 sg13g2_fill_2 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_285 ();
 sg13g2_fill_2 FILLER_27_292 ();
 sg13g2_fill_1 FILLER_27_333 ();
 sg13g2_fill_2 FILLER_27_353 ();
 sg13g2_fill_2 FILLER_27_364 ();
 sg13g2_fill_2 FILLER_27_379 ();
 sg13g2_fill_2 FILLER_27_398 ();
 sg13g2_fill_1 FILLER_27_400 ();
 sg13g2_decap_8 FILLER_27_408 ();
 sg13g2_fill_1 FILLER_28_39 ();
 sg13g2_fill_2 FILLER_28_45 ();
 sg13g2_fill_1 FILLER_28_152 ();
 sg13g2_fill_1 FILLER_28_159 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_fill_1 FILLER_28_174 ();
 sg13g2_fill_2 FILLER_28_188 ();
 sg13g2_fill_1 FILLER_28_190 ();
 sg13g2_fill_2 FILLER_28_195 ();
 sg13g2_fill_2 FILLER_28_201 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_208 ();
 sg13g2_decap_4 FILLER_28_215 ();
 sg13g2_fill_1 FILLER_28_219 ();
 sg13g2_fill_1 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_249 ();
 sg13g2_fill_1 FILLER_28_254 ();
 sg13g2_fill_2 FILLER_28_263 ();
 sg13g2_fill_1 FILLER_28_265 ();
 sg13g2_fill_2 FILLER_28_271 ();
 sg13g2_fill_1 FILLER_28_327 ();
 sg13g2_fill_1 FILLER_28_347 ();
 sg13g2_fill_2 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_404 ();
 sg13g2_fill_1 FILLER_28_409 ();
 sg13g2_fill_1 FILLER_28_414 ();
 sg13g2_fill_2 FILLER_28_418 ();
 sg13g2_fill_2 FILLER_28_428 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_7 ();
 sg13g2_fill_2 FILLER_29_12 ();
 sg13g2_fill_2 FILLER_29_89 ();
 sg13g2_fill_1 FILLER_29_105 ();
 sg13g2_fill_2 FILLER_29_110 ();
 sg13g2_fill_2 FILLER_29_117 ();
 sg13g2_fill_1 FILLER_29_184 ();
 sg13g2_decap_8 FILLER_29_203 ();
 sg13g2_fill_2 FILLER_29_210 ();
 sg13g2_fill_2 FILLER_29_220 ();
 sg13g2_fill_1 FILLER_29_227 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_2 FILLER_29_247 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_257 ();
 sg13g2_fill_1 FILLER_29_281 ();
 sg13g2_fill_1 FILLER_29_295 ();
 sg13g2_fill_1 FILLER_29_300 ();
 sg13g2_fill_1 FILLER_29_327 ();
 sg13g2_fill_2 FILLER_29_355 ();
 sg13g2_fill_1 FILLER_29_357 ();
 sg13g2_fill_2 FILLER_29_382 ();
 sg13g2_fill_1 FILLER_29_397 ();
 sg13g2_fill_2 FILLER_29_410 ();
 sg13g2_fill_2 FILLER_29_428 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_fill_1 FILLER_30_162 ();
 sg13g2_fill_1 FILLER_30_168 ();
 sg13g2_fill_2 FILLER_30_179 ();
 sg13g2_fill_1 FILLER_30_186 ();
 sg13g2_fill_1 FILLER_30_233 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_fill_1 FILLER_30_251 ();
 sg13g2_fill_2 FILLER_30_323 ();
 sg13g2_fill_1 FILLER_30_329 ();
 sg13g2_fill_2 FILLER_30_364 ();
 sg13g2_fill_2 FILLER_30_405 ();
 sg13g2_fill_1 FILLER_30_422 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_fill_1 FILLER_31_88 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_2 FILLER_31_115 ();
 sg13g2_fill_1 FILLER_31_190 ();
 sg13g2_fill_2 FILLER_31_199 ();
 sg13g2_fill_1 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_208 ();
 sg13g2_decap_4 FILLER_31_220 ();
 sg13g2_fill_1 FILLER_31_281 ();
 sg13g2_fill_1 FILLER_31_300 ();
 sg13g2_fill_1 FILLER_31_329 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_415 ();
 sg13g2_fill_2 FILLER_32_6 ();
 sg13g2_fill_2 FILLER_32_62 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_fill_2 FILLER_32_80 ();
 sg13g2_fill_1 FILLER_32_100 ();
 sg13g2_fill_1 FILLER_32_164 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_fill_1 FILLER_32_210 ();
 sg13g2_fill_1 FILLER_32_215 ();
 sg13g2_fill_1 FILLER_32_219 ();
 sg13g2_fill_2 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_264 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_fill_2 FILLER_32_274 ();
 sg13g2_fill_2 FILLER_32_281 ();
 sg13g2_fill_2 FILLER_32_287 ();
 sg13g2_fill_1 FILLER_32_289 ();
 sg13g2_fill_2 FILLER_32_315 ();
 sg13g2_fill_1 FILLER_32_317 ();
 sg13g2_fill_1 FILLER_32_323 ();
 sg13g2_fill_2 FILLER_32_328 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_fill_1 FILLER_32_377 ();
 sg13g2_fill_1 FILLER_32_400 ();
 sg13g2_decap_4 FILLER_32_426 ();
 sg13g2_fill_1 FILLER_33_87 ();
 sg13g2_fill_1 FILLER_33_119 ();
 sg13g2_fill_2 FILLER_33_129 ();
 sg13g2_fill_2 FILLER_33_145 ();
 sg13g2_fill_1 FILLER_33_173 ();
 sg13g2_fill_1 FILLER_33_179 ();
 sg13g2_fill_2 FILLER_33_194 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_decap_4 FILLER_33_215 ();
 sg13g2_decap_4 FILLER_33_222 ();
 sg13g2_fill_1 FILLER_33_231 ();
 sg13g2_fill_2 FILLER_33_257 ();
 sg13g2_fill_1 FILLER_33_259 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_fill_1 FILLER_33_303 ();
 sg13g2_fill_2 FILLER_33_324 ();
 sg13g2_fill_1 FILLER_33_347 ();
 sg13g2_fill_1 FILLER_33_352 ();
 sg13g2_fill_1 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_367 ();
 sg13g2_fill_1 FILLER_33_406 ();
 sg13g2_fill_1 FILLER_33_411 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_34_83 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_2 FILLER_34_109 ();
 sg13g2_fill_1 FILLER_34_119 ();
 sg13g2_fill_1 FILLER_34_125 ();
 sg13g2_decap_4 FILLER_34_167 ();
 sg13g2_fill_1 FILLER_34_179 ();
 sg13g2_fill_1 FILLER_34_185 ();
 sg13g2_fill_1 FILLER_34_194 ();
 sg13g2_fill_2 FILLER_34_200 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_decap_4 FILLER_34_214 ();
 sg13g2_fill_1 FILLER_34_229 ();
 sg13g2_fill_2 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_246 ();
 sg13g2_fill_1 FILLER_34_263 ();
 sg13g2_fill_2 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_276 ();
 sg13g2_fill_2 FILLER_34_293 ();
 sg13g2_fill_2 FILLER_34_318 ();
 sg13g2_decap_4 FILLER_34_332 ();
 sg13g2_fill_1 FILLER_34_336 ();
 sg13g2_decap_4 FILLER_34_396 ();
 sg13g2_fill_1 FILLER_34_400 ();
 sg13g2_fill_1 FILLER_34_429 ();
 sg13g2_fill_1 FILLER_35_26 ();
 sg13g2_fill_2 FILLER_35_67 ();
 sg13g2_fill_1 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_158 ();
 sg13g2_fill_1 FILLER_35_164 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_fill_2 FILLER_35_199 ();
 sg13g2_decap_4 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_213 ();
 sg13g2_fill_1 FILLER_35_215 ();
 sg13g2_fill_2 FILLER_35_220 ();
 sg13g2_fill_1 FILLER_35_222 ();
 sg13g2_fill_1 FILLER_35_240 ();
 sg13g2_fill_2 FILLER_35_255 ();
 sg13g2_fill_1 FILLER_35_266 ();
 sg13g2_fill_1 FILLER_35_271 ();
 sg13g2_fill_1 FILLER_35_276 ();
 sg13g2_fill_2 FILLER_35_307 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_1 FILLER_35_351 ();
 sg13g2_fill_1 FILLER_35_373 ();
 sg13g2_fill_1 FILLER_35_377 ();
 sg13g2_fill_1 FILLER_35_391 ();
 sg13g2_fill_1 FILLER_35_397 ();
 sg13g2_fill_1 FILLER_35_416 ();
 sg13g2_fill_1 FILLER_36_6 ();
 sg13g2_fill_2 FILLER_36_36 ();
 sg13g2_fill_1 FILLER_36_133 ();
 sg13g2_fill_2 FILLER_36_205 ();
 sg13g2_fill_1 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_224 ();
 sg13g2_fill_1 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_240 ();
 sg13g2_decap_8 FILLER_36_246 ();
 sg13g2_fill_2 FILLER_36_253 ();
 sg13g2_fill_1 FILLER_36_255 ();
 sg13g2_fill_2 FILLER_36_265 ();
 sg13g2_fill_1 FILLER_36_284 ();
 sg13g2_fill_1 FILLER_36_293 ();
 sg13g2_fill_1 FILLER_36_307 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_317 ();
 sg13g2_fill_2 FILLER_36_340 ();
 sg13g2_fill_1 FILLER_36_386 ();
 sg13g2_fill_2 FILLER_36_402 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_36_414 ();
 sg13g2_fill_1 FILLER_36_423 ();
 sg13g2_fill_2 FILLER_36_428 ();
 sg13g2_fill_1 FILLER_37_34 ();
 sg13g2_fill_2 FILLER_37_84 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_2 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_148 ();
 sg13g2_fill_1 FILLER_37_171 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_fill_1 FILLER_37_234 ();
 sg13g2_decap_4 FILLER_37_255 ();
 sg13g2_fill_1 FILLER_37_259 ();
 sg13g2_fill_2 FILLER_37_286 ();
 sg13g2_fill_1 FILLER_37_292 ();
 sg13g2_fill_1 FILLER_37_299 ();
 sg13g2_fill_1 FILLER_37_328 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_2 FILLER_37_339 ();
 sg13g2_fill_1 FILLER_37_345 ();
 sg13g2_fill_2 FILLER_37_351 ();
 sg13g2_fill_1 FILLER_37_385 ();
 sg13g2_fill_1 FILLER_37_394 ();
 sg13g2_fill_2 FILLER_37_398 ();
 sg13g2_fill_2 FILLER_37_415 ();
 sg13g2_fill_2 FILLER_38_14 ();
 sg13g2_fill_1 FILLER_38_59 ();
 sg13g2_fill_1 FILLER_38_70 ();
 sg13g2_fill_1 FILLER_38_81 ();
 sg13g2_fill_1 FILLER_38_87 ();
 sg13g2_fill_2 FILLER_38_102 ();
 sg13g2_fill_2 FILLER_38_148 ();
 sg13g2_fill_1 FILLER_38_181 ();
 sg13g2_fill_2 FILLER_38_186 ();
 sg13g2_fill_1 FILLER_38_206 ();
 sg13g2_fill_2 FILLER_38_290 ();
 sg13g2_fill_1 FILLER_38_299 ();
 sg13g2_fill_1 FILLER_38_361 ();
 sg13g2_fill_2 FILLER_38_403 ();
 sg13g2_fill_2 FILLER_38_420 ();
 sg13g2_fill_2 FILLER_38_428 ();
 sg13g2_fill_1 FILLER_39_43 ();
 sg13g2_fill_2 FILLER_39_117 ();
 sg13g2_fill_1 FILLER_39_124 ();
 sg13g2_fill_1 FILLER_39_132 ();
 sg13g2_fill_2 FILLER_39_143 ();
 sg13g2_fill_1 FILLER_39_174 ();
 sg13g2_fill_2 FILLER_39_207 ();
 sg13g2_fill_1 FILLER_39_236 ();
 sg13g2_fill_1 FILLER_39_241 ();
 sg13g2_fill_2 FILLER_39_255 ();
 sg13g2_fill_1 FILLER_39_261 ();
 sg13g2_fill_1 FILLER_39_267 ();
 sg13g2_fill_2 FILLER_39_272 ();
 sg13g2_fill_1 FILLER_39_279 ();
 sg13g2_fill_2 FILLER_39_299 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_311 ();
 sg13g2_fill_1 FILLER_39_332 ();
 sg13g2_fill_2 FILLER_39_359 ();
 sg13g2_fill_2 FILLER_39_379 ();
 sg13g2_fill_1 FILLER_39_385 ();
 sg13g2_decap_4 FILLER_39_391 ();
 sg13g2_fill_1 FILLER_39_395 ();
 sg13g2_fill_1 FILLER_39_404 ();
 sg13g2_fill_2 FILLER_39_410 ();
 sg13g2_fill_2 FILLER_40_40 ();
 sg13g2_fill_1 FILLER_40_63 ();
 sg13g2_fill_2 FILLER_40_100 ();
 sg13g2_fill_2 FILLER_40_119 ();
 sg13g2_decap_4 FILLER_40_173 ();
 sg13g2_fill_2 FILLER_40_182 ();
 sg13g2_fill_2 FILLER_40_206 ();
 sg13g2_fill_2 FILLER_40_219 ();
 sg13g2_fill_1 FILLER_40_221 ();
 sg13g2_fill_2 FILLER_40_246 ();
 sg13g2_fill_1 FILLER_40_265 ();
 sg13g2_fill_2 FILLER_40_274 ();
 sg13g2_fill_1 FILLER_40_280 ();
 sg13g2_fill_2 FILLER_40_290 ();
 sg13g2_fill_1 FILLER_40_297 ();
 sg13g2_fill_2 FILLER_40_315 ();
 sg13g2_fill_1 FILLER_40_321 ();
 sg13g2_decap_4 FILLER_40_330 ();
 sg13g2_fill_1 FILLER_40_400 ();
 sg13g2_fill_1 FILLER_40_409 ();
 sg13g2_fill_2 FILLER_40_428 ();
 sg13g2_fill_1 FILLER_41_63 ();
 sg13g2_fill_2 FILLER_41_101 ();
 sg13g2_fill_1 FILLER_41_103 ();
 sg13g2_fill_1 FILLER_41_123 ();
 sg13g2_fill_2 FILLER_41_140 ();
 sg13g2_fill_1 FILLER_41_142 ();
 sg13g2_fill_1 FILLER_41_148 ();
 sg13g2_fill_1 FILLER_41_154 ();
 sg13g2_fill_2 FILLER_41_163 ();
 sg13g2_fill_1 FILLER_41_170 ();
 sg13g2_fill_1 FILLER_41_176 ();
 sg13g2_fill_1 FILLER_41_181 ();
 sg13g2_fill_2 FILLER_41_192 ();
 sg13g2_decap_4 FILLER_41_198 ();
 sg13g2_fill_2 FILLER_41_220 ();
 sg13g2_fill_2 FILLER_41_231 ();
 sg13g2_fill_2 FILLER_41_237 ();
 sg13g2_fill_1 FILLER_41_243 ();
 sg13g2_fill_2 FILLER_41_249 ();
 sg13g2_fill_1 FILLER_41_251 ();
 sg13g2_fill_2 FILLER_41_256 ();
 sg13g2_fill_1 FILLER_41_258 ();
 sg13g2_fill_1 FILLER_41_263 ();
 sg13g2_decap_4 FILLER_41_268 ();
 sg13g2_fill_1 FILLER_41_272 ();
 sg13g2_fill_2 FILLER_41_277 ();
 sg13g2_fill_2 FILLER_41_364 ();
 sg13g2_fill_1 FILLER_41_366 ();
 sg13g2_fill_2 FILLER_41_381 ();
 sg13g2_fill_1 FILLER_41_419 ();
 sg13g2_fill_2 FILLER_42_0 ();
 sg13g2_fill_1 FILLER_42_8 ();
 sg13g2_fill_2 FILLER_42_65 ();
 sg13g2_fill_2 FILLER_42_72 ();
 sg13g2_fill_1 FILLER_42_89 ();
 sg13g2_fill_1 FILLER_42_153 ();
 sg13g2_fill_1 FILLER_42_174 ();
 sg13g2_fill_1 FILLER_42_196 ();
 sg13g2_fill_1 FILLER_42_205 ();
 sg13g2_fill_1 FILLER_42_211 ();
 sg13g2_fill_2 FILLER_42_219 ();
 sg13g2_fill_1 FILLER_42_238 ();
 sg13g2_fill_1 FILLER_42_250 ();
 sg13g2_fill_2 FILLER_42_265 ();
 sg13g2_decap_4 FILLER_42_277 ();
 sg13g2_fill_1 FILLER_42_289 ();
 sg13g2_fill_1 FILLER_42_317 ();
 sg13g2_fill_1 FILLER_42_321 ();
 sg13g2_fill_2 FILLER_42_329 ();
 sg13g2_fill_2 FILLER_42_344 ();
 sg13g2_fill_2 FILLER_42_377 ();
 sg13g2_fill_2 FILLER_42_386 ();
 sg13g2_fill_1 FILLER_42_391 ();
 sg13g2_fill_1 FILLER_42_399 ();
 sg13g2_fill_2 FILLER_42_427 ();
 sg13g2_fill_1 FILLER_42_429 ();
 sg13g2_fill_2 FILLER_43_34 ();
 sg13g2_fill_1 FILLER_43_65 ();
 sg13g2_fill_2 FILLER_43_116 ();
 sg13g2_fill_1 FILLER_43_128 ();
 sg13g2_fill_1 FILLER_43_137 ();
 sg13g2_fill_1 FILLER_43_143 ();
 sg13g2_fill_2 FILLER_43_200 ();
 sg13g2_decap_4 FILLER_43_221 ();
 sg13g2_fill_2 FILLER_43_225 ();
 sg13g2_fill_1 FILLER_43_232 ();
 sg13g2_decap_8 FILLER_43_242 ();
 sg13g2_fill_2 FILLER_43_249 ();
 sg13g2_fill_1 FILLER_43_289 ();
 sg13g2_decap_8 FILLER_43_303 ();
 sg13g2_fill_2 FILLER_43_310 ();
 sg13g2_fill_1 FILLER_43_312 ();
 sg13g2_fill_2 FILLER_43_335 ();
 sg13g2_fill_2 FILLER_43_354 ();
 sg13g2_fill_2 FILLER_43_378 ();
 sg13g2_fill_2 FILLER_43_390 ();
 sg13g2_fill_2 FILLER_43_397 ();
 sg13g2_decap_4 FILLER_43_426 ();
 sg13g2_fill_2 FILLER_44_70 ();
 sg13g2_fill_2 FILLER_44_88 ();
 sg13g2_fill_1 FILLER_44_108 ();
 sg13g2_fill_1 FILLER_44_113 ();
 sg13g2_fill_2 FILLER_44_132 ();
 sg13g2_fill_2 FILLER_44_151 ();
 sg13g2_fill_1 FILLER_44_153 ();
 sg13g2_fill_1 FILLER_44_171 ();
 sg13g2_fill_1 FILLER_44_175 ();
 sg13g2_fill_1 FILLER_44_180 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_199 ();
 sg13g2_fill_2 FILLER_44_217 ();
 sg13g2_fill_2 FILLER_44_224 ();
 sg13g2_fill_1 FILLER_44_226 ();
 sg13g2_decap_8 FILLER_44_231 ();
 sg13g2_fill_2 FILLER_44_245 ();
 sg13g2_fill_1 FILLER_44_247 ();
 sg13g2_fill_2 FILLER_44_253 ();
 sg13g2_decap_8 FILLER_44_272 ();
 sg13g2_fill_1 FILLER_44_305 ();
 sg13g2_fill_2 FILLER_44_347 ();
 sg13g2_fill_2 FILLER_44_390 ();
 sg13g2_fill_1 FILLER_44_415 ();
 sg13g2_decap_4 FILLER_44_425 ();
 sg13g2_fill_1 FILLER_44_429 ();
 sg13g2_fill_1 FILLER_45_109 ();
 sg13g2_fill_1 FILLER_45_167 ();
 sg13g2_fill_1 FILLER_45_171 ();
 sg13g2_fill_2 FILLER_45_207 ();
 sg13g2_fill_1 FILLER_45_213 ();
 sg13g2_fill_2 FILLER_45_219 ();
 sg13g2_decap_4 FILLER_45_234 ();
 sg13g2_fill_2 FILLER_45_238 ();
 sg13g2_fill_2 FILLER_45_244 ();
 sg13g2_decap_4 FILLER_45_253 ();
 sg13g2_fill_2 FILLER_45_271 ();
 sg13g2_decap_4 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_290 ();
 sg13g2_decap_4 FILLER_45_297 ();
 sg13g2_fill_1 FILLER_45_321 ();
 sg13g2_fill_1 FILLER_45_325 ();
 sg13g2_fill_2 FILLER_45_330 ();
 sg13g2_fill_2 FILLER_45_336 ();
 sg13g2_fill_2 FILLER_45_341 ();
 sg13g2_fill_2 FILLER_45_356 ();
 sg13g2_fill_2 FILLER_45_393 ();
 sg13g2_decap_4 FILLER_45_399 ();
 sg13g2_fill_2 FILLER_45_403 ();
 sg13g2_fill_1 FILLER_45_413 ();
 sg13g2_fill_1 FILLER_45_429 ();
 sg13g2_fill_1 FILLER_46_4 ();
 sg13g2_fill_1 FILLER_46_31 ();
 sg13g2_fill_1 FILLER_46_66 ();
 sg13g2_fill_2 FILLER_46_155 ();
 sg13g2_fill_1 FILLER_46_157 ();
 sg13g2_fill_2 FILLER_46_164 ();
 sg13g2_fill_1 FILLER_46_187 ();
 sg13g2_decap_4 FILLER_46_217 ();
 sg13g2_fill_1 FILLER_46_221 ();
 sg13g2_decap_4 FILLER_46_231 ();
 sg13g2_fill_2 FILLER_46_247 ();
 sg13g2_fill_1 FILLER_46_253 ();
 sg13g2_fill_2 FILLER_46_271 ();
 sg13g2_fill_1 FILLER_46_277 ();
 sg13g2_decap_4 FILLER_46_287 ();
 sg13g2_fill_2 FILLER_46_311 ();
 sg13g2_fill_2 FILLER_46_322 ();
 sg13g2_fill_2 FILLER_46_331 ();
 sg13g2_fill_1 FILLER_46_333 ();
 sg13g2_fill_2 FILLER_46_341 ();
 sg13g2_fill_2 FILLER_46_357 ();
 sg13g2_fill_2 FILLER_46_373 ();
 sg13g2_decap_4 FILLER_46_384 ();
 sg13g2_fill_1 FILLER_46_388 ();
 sg13g2_fill_2 FILLER_46_397 ();
 sg13g2_fill_1 FILLER_46_399 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_2 FILLER_46_420 ();
 sg13g2_fill_1 FILLER_46_422 ();
 sg13g2_fill_2 FILLER_46_428 ();
 sg13g2_fill_2 FILLER_47_43 ();
 sg13g2_fill_2 FILLER_47_53 ();
 sg13g2_fill_1 FILLER_47_64 ();
 sg13g2_fill_1 FILLER_47_76 ();
 sg13g2_fill_1 FILLER_47_124 ();
 sg13g2_fill_1 FILLER_47_129 ();
 sg13g2_fill_1 FILLER_47_138 ();
 sg13g2_fill_1 FILLER_47_181 ();
 sg13g2_fill_2 FILLER_47_221 ();
 sg13g2_fill_2 FILLER_47_258 ();
 sg13g2_fill_1 FILLER_47_265 ();
 sg13g2_fill_2 FILLER_47_275 ();
 sg13g2_fill_2 FILLER_47_281 ();
 sg13g2_fill_1 FILLER_47_283 ();
 sg13g2_fill_2 FILLER_47_289 ();
 sg13g2_fill_1 FILLER_47_291 ();
 sg13g2_fill_2 FILLER_47_297 ();
 sg13g2_decap_4 FILLER_47_307 ();
 sg13g2_fill_1 FILLER_47_328 ();
 sg13g2_fill_2 FILLER_47_341 ();
 sg13g2_fill_1 FILLER_47_367 ();
 sg13g2_fill_1 FILLER_47_395 ();
 sg13g2_fill_2 FILLER_47_408 ();
 sg13g2_fill_2 FILLER_47_423 ();
 sg13g2_fill_1 FILLER_47_429 ();
 sg13g2_fill_1 FILLER_48_0 ();
 sg13g2_fill_2 FILLER_48_9 ();
 sg13g2_fill_1 FILLER_48_15 ();
 sg13g2_fill_1 FILLER_48_114 ();
 sg13g2_fill_1 FILLER_48_118 ();
 sg13g2_fill_2 FILLER_48_168 ();
 sg13g2_fill_1 FILLER_48_174 ();
 sg13g2_fill_1 FILLER_48_180 ();
 sg13g2_fill_2 FILLER_48_186 ();
 sg13g2_fill_1 FILLER_48_188 ();
 sg13g2_fill_1 FILLER_48_214 ();
 sg13g2_fill_2 FILLER_48_245 ();
 sg13g2_fill_1 FILLER_48_267 ();
 sg13g2_fill_1 FILLER_48_306 ();
 sg13g2_fill_1 FILLER_48_311 ();
 sg13g2_fill_2 FILLER_48_321 ();
 sg13g2_fill_2 FILLER_48_337 ();
 sg13g2_fill_1 FILLER_48_339 ();
 sg13g2_fill_1 FILLER_48_345 ();
 sg13g2_fill_1 FILLER_48_353 ();
 sg13g2_fill_2 FILLER_48_367 ();
 sg13g2_fill_2 FILLER_48_376 ();
 sg13g2_decap_4 FILLER_48_396 ();
 sg13g2_fill_2 FILLER_48_404 ();
 sg13g2_fill_2 FILLER_48_414 ();
 sg13g2_fill_1 FILLER_48_416 ();
 sg13g2_fill_1 FILLER_48_425 ();
 sg13g2_fill_2 FILLER_49_123 ();
 sg13g2_fill_2 FILLER_49_208 ();
 sg13g2_fill_1 FILLER_49_229 ();
 sg13g2_fill_2 FILLER_49_234 ();
 sg13g2_decap_4 FILLER_49_248 ();
 sg13g2_fill_2 FILLER_49_252 ();
 sg13g2_fill_1 FILLER_49_258 ();
 sg13g2_decap_4 FILLER_49_268 ();
 sg13g2_fill_2 FILLER_49_285 ();
 sg13g2_fill_1 FILLER_49_287 ();
 sg13g2_decap_8 FILLER_49_292 ();
 sg13g2_fill_1 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_321 ();
 sg13g2_fill_1 FILLER_49_323 ();
 sg13g2_fill_2 FILLER_49_346 ();
 sg13g2_fill_1 FILLER_49_348 ();
 sg13g2_fill_1 FILLER_49_368 ();
 sg13g2_fill_1 FILLER_49_385 ();
 sg13g2_decap_4 FILLER_49_389 ();
 sg13g2_fill_2 FILLER_49_393 ();
 sg13g2_decap_8 FILLER_49_399 ();
 sg13g2_fill_2 FILLER_49_406 ();
 sg13g2_fill_1 FILLER_49_408 ();
 sg13g2_fill_2 FILLER_49_422 ();
 sg13g2_fill_1 FILLER_49_429 ();
 sg13g2_fill_1 FILLER_50_42 ();
 sg13g2_fill_2 FILLER_50_52 ();
 sg13g2_fill_1 FILLER_50_105 ();
 sg13g2_fill_2 FILLER_50_142 ();
 sg13g2_fill_1 FILLER_50_148 ();
 sg13g2_fill_2 FILLER_50_160 ();
 sg13g2_fill_1 FILLER_50_168 ();
 sg13g2_fill_1 FILLER_50_174 ();
 sg13g2_fill_1 FILLER_50_187 ();
 sg13g2_fill_1 FILLER_50_192 ();
 sg13g2_fill_2 FILLER_50_216 ();
 sg13g2_decap_4 FILLER_50_248 ();
 sg13g2_fill_1 FILLER_50_302 ();
 sg13g2_fill_2 FILLER_50_307 ();
 sg13g2_fill_1 FILLER_50_309 ();
 sg13g2_fill_2 FILLER_50_317 ();
 sg13g2_fill_1 FILLER_50_336 ();
 sg13g2_fill_1 FILLER_50_340 ();
 sg13g2_fill_1 FILLER_50_345 ();
 sg13g2_fill_1 FILLER_50_369 ();
 sg13g2_decap_4 FILLER_50_416 ();
 sg13g2_decap_4 FILLER_50_425 ();
 sg13g2_fill_1 FILLER_50_429 ();
 sg13g2_fill_2 FILLER_51_28 ();
 sg13g2_fill_1 FILLER_51_75 ();
 sg13g2_fill_1 FILLER_51_92 ();
 sg13g2_fill_1 FILLER_51_110 ();
 sg13g2_fill_1 FILLER_51_157 ();
 sg13g2_fill_1 FILLER_51_167 ();
 sg13g2_fill_2 FILLER_51_206 ();
 sg13g2_fill_2 FILLER_51_224 ();
 sg13g2_fill_1 FILLER_51_239 ();
 sg13g2_fill_2 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_259 ();
 sg13g2_fill_1 FILLER_51_265 ();
 sg13g2_fill_1 FILLER_51_276 ();
 sg13g2_decap_4 FILLER_51_290 ();
 sg13g2_fill_1 FILLER_51_294 ();
 sg13g2_fill_1 FILLER_51_299 ();
 sg13g2_fill_2 FILLER_51_319 ();
 sg13g2_fill_2 FILLER_51_325 ();
 sg13g2_fill_1 FILLER_51_390 ();
 sg13g2_decap_8 FILLER_51_403 ();
 sg13g2_fill_2 FILLER_51_410 ();
 sg13g2_decap_4 FILLER_51_426 ();
 sg13g2_fill_2 FILLER_52_0 ();
 sg13g2_fill_2 FILLER_52_51 ();
 sg13g2_fill_2 FILLER_52_159 ();
 sg13g2_fill_2 FILLER_52_185 ();
 sg13g2_fill_1 FILLER_52_192 ();
 sg13g2_fill_1 FILLER_52_210 ();
 sg13g2_fill_1 FILLER_52_215 ();
 sg13g2_decap_4 FILLER_52_228 ();
 sg13g2_fill_1 FILLER_52_241 ();
 sg13g2_fill_1 FILLER_52_246 ();
 sg13g2_fill_1 FILLER_52_252 ();
 sg13g2_fill_1 FILLER_52_261 ();
 sg13g2_decap_4 FILLER_52_281 ();
 sg13g2_fill_1 FILLER_52_285 ();
 sg13g2_fill_2 FILLER_52_317 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_397 ();
 sg13g2_fill_2 FILLER_52_428 ();
 sg13g2_fill_2 FILLER_53_61 ();
 sg13g2_fill_1 FILLER_53_98 ();
 sg13g2_fill_2 FILLER_53_111 ();
 sg13g2_fill_2 FILLER_53_145 ();
 sg13g2_fill_1 FILLER_53_173 ();
 sg13g2_fill_1 FILLER_53_184 ();
 sg13g2_fill_1 FILLER_53_193 ();
 sg13g2_fill_1 FILLER_53_209 ();
 sg13g2_fill_1 FILLER_53_220 ();
 sg13g2_decap_4 FILLER_53_228 ();
 sg13g2_fill_2 FILLER_53_258 ();
 sg13g2_fill_1 FILLER_53_260 ();
 sg13g2_fill_1 FILLER_53_276 ();
 sg13g2_decap_4 FILLER_53_282 ();
 sg13g2_decap_4 FILLER_53_291 ();
 sg13g2_fill_1 FILLER_53_295 ();
 sg13g2_fill_2 FILLER_53_307 ();
 sg13g2_fill_1 FILLER_53_309 ();
 sg13g2_fill_2 FILLER_53_315 ();
 sg13g2_fill_1 FILLER_53_317 ();
 sg13g2_fill_1 FILLER_53_346 ();
 sg13g2_decap_8 FILLER_53_367 ();
 sg13g2_fill_2 FILLER_53_374 ();
 sg13g2_fill_1 FILLER_53_403 ();
 sg13g2_decap_4 FILLER_53_407 ();
 sg13g2_fill_2 FILLER_53_411 ();
 sg13g2_fill_1 FILLER_53_421 ();
 sg13g2_fill_2 FILLER_53_427 ();
 sg13g2_fill_1 FILLER_53_429 ();
 sg13g2_fill_1 FILLER_54_25 ();
 sg13g2_fill_2 FILLER_54_38 ();
 sg13g2_fill_1 FILLER_54_148 ();
 sg13g2_fill_1 FILLER_54_154 ();
 sg13g2_fill_1 FILLER_54_160 ();
 sg13g2_fill_1 FILLER_54_210 ();
 sg13g2_fill_2 FILLER_54_221 ();
 sg13g2_fill_2 FILLER_54_232 ();
 sg13g2_decap_4 FILLER_54_239 ();
 sg13g2_fill_1 FILLER_54_243 ();
 sg13g2_decap_4 FILLER_54_265 ();
 sg13g2_decap_4 FILLER_54_291 ();
 sg13g2_fill_2 FILLER_54_313 ();
 sg13g2_fill_2 FILLER_54_343 ();
 sg13g2_fill_1 FILLER_54_345 ();
 sg13g2_fill_1 FILLER_54_375 ();
 sg13g2_fill_1 FILLER_54_385 ();
 sg13g2_fill_1 FILLER_54_391 ();
 sg13g2_fill_1 FILLER_54_400 ();
 sg13g2_decap_4 FILLER_54_409 ();
 sg13g2_fill_2 FILLER_54_413 ();
 sg13g2_fill_1 FILLER_54_429 ();
 sg13g2_fill_2 FILLER_55_24 ();
 sg13g2_fill_2 FILLER_55_45 ();
 sg13g2_fill_1 FILLER_55_69 ();
 sg13g2_fill_1 FILLER_55_97 ();
 sg13g2_fill_1 FILLER_55_123 ();
 sg13g2_fill_2 FILLER_55_221 ();
 sg13g2_fill_2 FILLER_55_247 ();
 sg13g2_fill_2 FILLER_55_254 ();
 sg13g2_decap_4 FILLER_55_260 ();
 sg13g2_fill_2 FILLER_55_264 ();
 sg13g2_fill_1 FILLER_55_275 ();
 sg13g2_fill_1 FILLER_55_281 ();
 sg13g2_fill_1 FILLER_55_290 ();
 sg13g2_fill_1 FILLER_55_308 ();
 sg13g2_fill_1 FILLER_55_313 ();
 sg13g2_fill_1 FILLER_55_318 ();
 sg13g2_fill_2 FILLER_55_322 ();
 sg13g2_decap_4 FILLER_55_328 ();
 sg13g2_fill_1 FILLER_55_348 ();
 sg13g2_fill_1 FILLER_55_352 ();
 sg13g2_fill_1 FILLER_55_361 ();
 sg13g2_fill_1 FILLER_55_365 ();
 sg13g2_fill_1 FILLER_55_374 ();
 sg13g2_decap_8 FILLER_55_380 ();
 sg13g2_fill_2 FILLER_55_387 ();
 sg13g2_fill_1 FILLER_55_412 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_fill_1 FILLER_56_19 ();
 sg13g2_fill_1 FILLER_56_45 ();
 sg13g2_fill_2 FILLER_56_186 ();
 sg13g2_fill_1 FILLER_56_199 ();
 sg13g2_fill_1 FILLER_56_221 ();
 sg13g2_fill_1 FILLER_56_238 ();
 sg13g2_fill_2 FILLER_56_261 ();
 sg13g2_fill_2 FILLER_56_283 ();
 sg13g2_fill_2 FILLER_56_290 ();
 sg13g2_fill_1 FILLER_56_296 ();
 sg13g2_fill_2 FILLER_56_301 ();
 sg13g2_fill_2 FILLER_56_307 ();
 sg13g2_fill_2 FILLER_56_314 ();
 sg13g2_fill_1 FILLER_56_316 ();
 sg13g2_decap_8 FILLER_56_330 ();
 sg13g2_fill_1 FILLER_56_342 ();
 sg13g2_fill_1 FILLER_56_348 ();
 sg13g2_fill_2 FILLER_56_376 ();
 sg13g2_fill_1 FILLER_56_386 ();
 sg13g2_fill_1 FILLER_56_390 ();
 sg13g2_fill_1 FILLER_56_396 ();
 sg13g2_fill_2 FILLER_56_402 ();
 sg13g2_fill_1 FILLER_56_412 ();
 sg13g2_decap_4 FILLER_56_417 ();
 sg13g2_fill_1 FILLER_57_5 ();
 sg13g2_fill_1 FILLER_57_11 ();
 sg13g2_fill_2 FILLER_57_70 ();
 sg13g2_fill_1 FILLER_57_85 ();
 sg13g2_fill_2 FILLER_57_98 ();
 sg13g2_fill_1 FILLER_57_113 ();
 sg13g2_fill_2 FILLER_57_132 ();
 sg13g2_fill_1 FILLER_57_148 ();
 sg13g2_fill_2 FILLER_57_154 ();
 sg13g2_fill_1 FILLER_57_228 ();
 sg13g2_fill_1 FILLER_57_233 ();
 sg13g2_decap_4 FILLER_57_261 ();
 sg13g2_fill_1 FILLER_57_273 ();
 sg13g2_fill_1 FILLER_57_330 ();
 sg13g2_fill_2 FILLER_57_355 ();
 sg13g2_fill_1 FILLER_57_357 ();
 sg13g2_decap_4 FILLER_57_366 ();
 sg13g2_fill_1 FILLER_57_394 ();
 sg13g2_fill_1 FILLER_57_419 ();
 sg13g2_fill_1 FILLER_57_429 ();
 sg13g2_fill_2 FILLER_58_56 ();
 sg13g2_fill_2 FILLER_58_84 ();
 sg13g2_fill_2 FILLER_58_105 ();
 sg13g2_fill_2 FILLER_58_143 ();
 sg13g2_fill_1 FILLER_58_183 ();
 sg13g2_fill_1 FILLER_58_217 ();
 sg13g2_fill_2 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_241 ();
 sg13g2_fill_2 FILLER_58_246 ();
 sg13g2_fill_2 FILLER_58_257 ();
 sg13g2_fill_1 FILLER_58_263 ();
 sg13g2_fill_2 FILLER_58_269 ();
 sg13g2_fill_1 FILLER_58_279 ();
 sg13g2_fill_2 FILLER_58_289 ();
 sg13g2_fill_2 FILLER_58_310 ();
 sg13g2_fill_1 FILLER_58_312 ();
 sg13g2_fill_1 FILLER_58_317 ();
 sg13g2_fill_1 FILLER_58_337 ();
 sg13g2_fill_1 FILLER_58_347 ();
 sg13g2_fill_2 FILLER_58_351 ();
 sg13g2_fill_1 FILLER_58_353 ();
 sg13g2_fill_2 FILLER_58_363 ();
 sg13g2_fill_1 FILLER_58_365 ();
 sg13g2_fill_2 FILLER_58_379 ();
 sg13g2_fill_1 FILLER_58_411 ();
 sg13g2_fill_1 FILLER_58_429 ();
 sg13g2_fill_1 FILLER_59_0 ();
 sg13g2_fill_2 FILLER_59_9 ();
 sg13g2_fill_1 FILLER_59_41 ();
 sg13g2_fill_1 FILLER_59_60 ();
 sg13g2_fill_1 FILLER_59_66 ();
 sg13g2_fill_1 FILLER_59_76 ();
 sg13g2_fill_1 FILLER_59_99 ();
 sg13g2_fill_2 FILLER_59_105 ();
 sg13g2_fill_2 FILLER_59_210 ();
 sg13g2_fill_1 FILLER_59_219 ();
 sg13g2_fill_1 FILLER_59_224 ();
 sg13g2_fill_1 FILLER_59_234 ();
 sg13g2_fill_1 FILLER_59_251 ();
 sg13g2_fill_1 FILLER_59_260 ();
 sg13g2_fill_1 FILLER_59_270 ();
 sg13g2_fill_1 FILLER_59_275 ();
 sg13g2_fill_2 FILLER_59_293 ();
 sg13g2_decap_4 FILLER_59_308 ();
 sg13g2_fill_2 FILLER_59_312 ();
 sg13g2_fill_1 FILLER_59_335 ();
 sg13g2_fill_2 FILLER_59_353 ();
 sg13g2_fill_2 FILLER_59_373 ();
 sg13g2_fill_2 FILLER_59_398 ();
 sg13g2_fill_2 FILLER_59_404 ();
 sg13g2_fill_1 FILLER_59_406 ();
 sg13g2_fill_2 FILLER_59_415 ();
 sg13g2_fill_1 FILLER_59_417 ();
 sg13g2_fill_1 FILLER_60_63 ();
 sg13g2_fill_1 FILLER_60_87 ();
 sg13g2_fill_2 FILLER_60_97 ();
 sg13g2_fill_1 FILLER_60_133 ();
 sg13g2_fill_1 FILLER_60_143 ();
 sg13g2_fill_2 FILLER_60_148 ();
 sg13g2_fill_1 FILLER_60_159 ();
 sg13g2_fill_1 FILLER_60_165 ();
 sg13g2_fill_1 FILLER_60_212 ();
 sg13g2_fill_1 FILLER_60_220 ();
 sg13g2_fill_2 FILLER_60_263 ();
 sg13g2_fill_2 FILLER_60_296 ();
 sg13g2_fill_1 FILLER_60_311 ();
 sg13g2_decap_8 FILLER_60_351 ();
 sg13g2_fill_1 FILLER_60_389 ();
 sg13g2_fill_2 FILLER_60_394 ();
 sg13g2_fill_2 FILLER_60_400 ();
 sg13g2_fill_1 FILLER_60_419 ();
 sg13g2_decap_4 FILLER_60_425 ();
 sg13g2_fill_1 FILLER_60_429 ();
 sg13g2_fill_2 FILLER_61_38 ();
 sg13g2_fill_1 FILLER_61_52 ();
 sg13g2_fill_1 FILLER_61_81 ();
 sg13g2_fill_2 FILLER_61_105 ();
 sg13g2_fill_1 FILLER_61_115 ();
 sg13g2_fill_1 FILLER_61_122 ();
 sg13g2_fill_1 FILLER_61_127 ();
 sg13g2_fill_2 FILLER_61_132 ();
 sg13g2_fill_2 FILLER_61_165 ();
 sg13g2_fill_1 FILLER_61_174 ();
 sg13g2_fill_1 FILLER_61_199 ();
 sg13g2_fill_1 FILLER_61_203 ();
 sg13g2_fill_1 FILLER_61_217 ();
 sg13g2_fill_1 FILLER_61_226 ();
 sg13g2_fill_1 FILLER_61_243 ();
 sg13g2_fill_1 FILLER_61_260 ();
 sg13g2_fill_1 FILLER_61_272 ();
 sg13g2_fill_2 FILLER_61_303 ();
 sg13g2_fill_2 FILLER_61_309 ();
 sg13g2_fill_1 FILLER_61_311 ();
 sg13g2_fill_1 FILLER_61_317 ();
 sg13g2_fill_2 FILLER_61_334 ();
 sg13g2_fill_1 FILLER_61_336 ();
 sg13g2_fill_2 FILLER_61_358 ();
 sg13g2_fill_1 FILLER_61_360 ();
 sg13g2_decap_4 FILLER_61_382 ();
 sg13g2_decap_4 FILLER_61_393 ();
 sg13g2_fill_1 FILLER_61_400 ();
 sg13g2_fill_1 FILLER_61_404 ();
 sg13g2_fill_2 FILLER_61_414 ();
 sg13g2_decap_4 FILLER_61_426 ();
 sg13g2_fill_1 FILLER_62_57 ();
 sg13g2_fill_2 FILLER_62_104 ();
 sg13g2_fill_2 FILLER_62_130 ();
 sg13g2_fill_1 FILLER_62_164 ();
 sg13g2_fill_1 FILLER_62_182 ();
 sg13g2_fill_2 FILLER_62_188 ();
 sg13g2_fill_1 FILLER_62_204 ();
 sg13g2_fill_1 FILLER_62_208 ();
 sg13g2_fill_1 FILLER_62_213 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_fill_2 FILLER_62_261 ();
 sg13g2_fill_1 FILLER_62_275 ();
 sg13g2_fill_1 FILLER_62_289 ();
 sg13g2_fill_1 FILLER_62_326 ();
 sg13g2_fill_1 FILLER_62_339 ();
 sg13g2_fill_2 FILLER_62_345 ();
 sg13g2_fill_1 FILLER_62_347 ();
 sg13g2_fill_2 FILLER_62_366 ();
 sg13g2_fill_1 FILLER_62_376 ();
 sg13g2_fill_2 FILLER_62_380 ();
 sg13g2_fill_1 FILLER_62_404 ();
 sg13g2_fill_2 FILLER_62_409 ();
 sg13g2_fill_2 FILLER_62_428 ();
 sg13g2_fill_2 FILLER_63_32 ();
 sg13g2_fill_1 FILLER_63_91 ();
 sg13g2_fill_2 FILLER_63_180 ();
 sg13g2_fill_2 FILLER_63_228 ();
 sg13g2_fill_2 FILLER_63_245 ();
 sg13g2_fill_1 FILLER_63_252 ();
 sg13g2_fill_1 FILLER_63_268 ();
 sg13g2_fill_1 FILLER_63_272 ();
 sg13g2_fill_2 FILLER_63_284 ();
 sg13g2_fill_1 FILLER_63_294 ();
 sg13g2_fill_1 FILLER_63_306 ();
 sg13g2_fill_1 FILLER_63_311 ();
 sg13g2_fill_2 FILLER_63_320 ();
 sg13g2_fill_1 FILLER_63_322 ();
 sg13g2_fill_1 FILLER_63_328 ();
 sg13g2_fill_2 FILLER_63_358 ();
 sg13g2_fill_1 FILLER_63_360 ();
 sg13g2_fill_2 FILLER_63_402 ();
 sg13g2_fill_2 FILLER_63_409 ();
 sg13g2_fill_1 FILLER_63_424 ();
 sg13g2_fill_1 FILLER_63_429 ();
 sg13g2_fill_2 FILLER_64_0 ();
 sg13g2_fill_1 FILLER_64_39 ();
 sg13g2_fill_2 FILLER_64_56 ();
 sg13g2_fill_2 FILLER_64_79 ();
 sg13g2_fill_1 FILLER_64_136 ();
 sg13g2_fill_2 FILLER_64_142 ();
 sg13g2_fill_1 FILLER_64_171 ();
 sg13g2_fill_2 FILLER_64_199 ();
 sg13g2_fill_1 FILLER_64_270 ();
 sg13g2_fill_2 FILLER_64_275 ();
 sg13g2_fill_1 FILLER_64_285 ();
 sg13g2_fill_1 FILLER_64_298 ();
 sg13g2_fill_1 FILLER_64_307 ();
 sg13g2_fill_1 FILLER_64_317 ();
 sg13g2_fill_1 FILLER_64_326 ();
 sg13g2_fill_1 FILLER_64_331 ();
 sg13g2_fill_2 FILLER_64_374 ();
 sg13g2_fill_2 FILLER_64_380 ();
 sg13g2_fill_1 FILLER_64_395 ();
 sg13g2_fill_1 FILLER_64_399 ();
 sg13g2_fill_1 FILLER_64_404 ();
 sg13g2_fill_2 FILLER_64_408 ();
 sg13g2_decap_4 FILLER_64_421 ();
 sg13g2_fill_1 FILLER_65_0 ();
 sg13g2_fill_1 FILLER_65_14 ();
 sg13g2_fill_1 FILLER_65_41 ();
 sg13g2_fill_1 FILLER_65_68 ();
 sg13g2_fill_1 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_105 ();
 sg13g2_fill_1 FILLER_65_127 ();
 sg13g2_fill_2 FILLER_65_137 ();
 sg13g2_fill_1 FILLER_65_144 ();
 sg13g2_fill_2 FILLER_65_164 ();
 sg13g2_fill_1 FILLER_65_178 ();
 sg13g2_fill_1 FILLER_65_199 ();
 sg13g2_fill_2 FILLER_65_208 ();
 sg13g2_fill_1 FILLER_65_214 ();
 sg13g2_fill_1 FILLER_65_258 ();
 sg13g2_fill_2 FILLER_65_286 ();
 sg13g2_fill_2 FILLER_65_309 ();
 sg13g2_fill_2 FILLER_65_316 ();
 sg13g2_fill_2 FILLER_65_323 ();
 sg13g2_fill_2 FILLER_65_348 ();
 sg13g2_fill_1 FILLER_65_355 ();
 sg13g2_fill_1 FILLER_65_360 ();
 sg13g2_fill_1 FILLER_65_365 ();
 sg13g2_decap_4 FILLER_65_374 ();
 sg13g2_fill_1 FILLER_65_378 ();
 sg13g2_fill_2 FILLER_65_387 ();
 sg13g2_fill_1 FILLER_65_389 ();
 sg13g2_fill_1 FILLER_65_393 ();
 sg13g2_fill_1 FILLER_65_402 ();
 sg13g2_fill_1 FILLER_65_419 ();
 sg13g2_fill_1 FILLER_65_429 ();
 sg13g2_fill_1 FILLER_66_98 ();
 sg13g2_fill_2 FILLER_66_133 ();
 sg13g2_fill_1 FILLER_66_198 ();
 sg13g2_fill_2 FILLER_66_234 ();
 sg13g2_fill_1 FILLER_66_241 ();
 sg13g2_fill_1 FILLER_66_245 ();
 sg13g2_fill_1 FILLER_66_267 ();
 sg13g2_fill_1 FILLER_66_271 ();
 sg13g2_fill_1 FILLER_66_276 ();
 sg13g2_fill_2 FILLER_66_286 ();
 sg13g2_fill_1 FILLER_66_304 ();
 sg13g2_fill_1 FILLER_66_364 ();
 sg13g2_fill_1 FILLER_66_372 ();
 sg13g2_fill_1 FILLER_66_391 ();
 sg13g2_fill_2 FILLER_66_415 ();
 sg13g2_fill_2 FILLER_67_31 ();
 sg13g2_fill_1 FILLER_67_47 ();
 sg13g2_fill_1 FILLER_67_52 ();
 sg13g2_fill_1 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_230 ();
 sg13g2_fill_1 FILLER_67_235 ();
 sg13g2_fill_1 FILLER_67_240 ();
 sg13g2_fill_1 FILLER_67_244 ();
 sg13g2_fill_1 FILLER_67_250 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_276 ();
 sg13g2_fill_1 FILLER_67_281 ();
 sg13g2_fill_1 FILLER_67_301 ();
 sg13g2_fill_2 FILLER_67_319 ();
 sg13g2_fill_1 FILLER_67_334 ();
 sg13g2_fill_2 FILLER_67_356 ();
 sg13g2_fill_1 FILLER_67_358 ();
 sg13g2_decap_8 FILLER_67_395 ();
 sg13g2_fill_1 FILLER_68_20 ();
 sg13g2_fill_2 FILLER_68_55 ();
 sg13g2_fill_1 FILLER_68_88 ();
 sg13g2_fill_1 FILLER_68_143 ();
 sg13g2_fill_1 FILLER_68_164 ();
 sg13g2_fill_1 FILLER_68_169 ();
 sg13g2_fill_1 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_219 ();
 sg13g2_fill_2 FILLER_68_226 ();
 sg13g2_fill_2 FILLER_68_281 ();
 sg13g2_fill_1 FILLER_68_341 ();
 sg13g2_fill_1 FILLER_68_358 ();
 sg13g2_fill_2 FILLER_68_372 ();
 sg13g2_decap_8 FILLER_68_382 ();
 sg13g2_decap_4 FILLER_68_389 ();
 sg13g2_decap_4 FILLER_68_396 ();
 sg13g2_fill_2 FILLER_68_400 ();
 sg13g2_fill_1 FILLER_68_410 ();
 sg13g2_fill_1 FILLER_68_419 ();
 sg13g2_fill_1 FILLER_69_0 ();
 sg13g2_fill_2 FILLER_69_94 ();
 sg13g2_fill_1 FILLER_69_100 ();
 sg13g2_fill_1 FILLER_69_105 ();
 sg13g2_fill_1 FILLER_69_110 ();
 sg13g2_fill_1 FILLER_69_116 ();
 sg13g2_fill_1 FILLER_69_143 ();
 sg13g2_fill_1 FILLER_69_180 ();
 sg13g2_fill_1 FILLER_69_275 ();
 sg13g2_fill_2 FILLER_69_302 ();
 sg13g2_fill_1 FILLER_69_319 ();
 sg13g2_fill_2 FILLER_69_335 ();
 sg13g2_fill_1 FILLER_69_357 ();
 sg13g2_decap_4 FILLER_69_362 ();
 sg13g2_fill_2 FILLER_69_370 ();
 sg13g2_fill_1 FILLER_69_372 ();
 sg13g2_fill_2 FILLER_69_377 ();
 sg13g2_fill_1 FILLER_69_384 ();
 sg13g2_fill_1 FILLER_69_390 ();
 sg13g2_fill_1 FILLER_69_400 ();
 sg13g2_fill_1 FILLER_69_404 ();
 sg13g2_fill_1 FILLER_69_410 ();
 sg13g2_fill_2 FILLER_69_423 ();
 sg13g2_fill_1 FILLER_69_425 ();
 sg13g2_fill_1 FILLER_70_26 ();
 sg13g2_fill_2 FILLER_70_76 ();
 sg13g2_fill_1 FILLER_70_102 ();
 sg13g2_fill_2 FILLER_70_220 ();
 sg13g2_fill_1 FILLER_70_240 ();
 sg13g2_fill_1 FILLER_70_250 ();
 sg13g2_fill_1 FILLER_70_282 ();
 sg13g2_fill_1 FILLER_70_291 ();
 sg13g2_fill_1 FILLER_70_304 ();
 sg13g2_fill_1 FILLER_70_313 ();
 sg13g2_fill_1 FILLER_70_322 ();
 sg13g2_fill_2 FILLER_70_371 ();
 sg13g2_fill_1 FILLER_70_414 ();
 sg13g2_fill_2 FILLER_70_428 ();
 sg13g2_fill_2 FILLER_71_0 ();
 sg13g2_fill_1 FILLER_71_150 ();
 sg13g2_fill_2 FILLER_71_159 ();
 sg13g2_fill_1 FILLER_71_182 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_fill_2 FILLER_71_256 ();
 sg13g2_fill_1 FILLER_71_272 ();
 sg13g2_fill_2 FILLER_71_286 ();
 sg13g2_fill_2 FILLER_71_315 ();
 sg13g2_fill_1 FILLER_71_325 ();
 sg13g2_fill_2 FILLER_71_333 ();
 sg13g2_fill_1 FILLER_71_343 ();
 sg13g2_decap_4 FILLER_71_384 ();
 sg13g2_fill_2 FILLER_71_405 ();
 sg13g2_decap_4 FILLER_71_416 ();
 sg13g2_fill_1 FILLER_71_420 ();
 sg13g2_decap_4 FILLER_71_426 ();
 sg13g2_fill_2 FILLER_72_26 ();
 sg13g2_fill_1 FILLER_72_87 ();
 sg13g2_fill_2 FILLER_72_133 ();
 sg13g2_fill_2 FILLER_72_189 ();
 sg13g2_fill_2 FILLER_72_244 ();
 sg13g2_fill_2 FILLER_72_267 ();
 sg13g2_fill_2 FILLER_72_273 ();
 sg13g2_fill_2 FILLER_72_284 ();
 sg13g2_fill_1 FILLER_72_290 ();
 sg13g2_fill_1 FILLER_72_295 ();
 sg13g2_fill_2 FILLER_72_300 ();
 sg13g2_fill_1 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_388 ();
 sg13g2_fill_1 FILLER_72_397 ();
 sg13g2_fill_1 FILLER_73_48 ();
 sg13g2_fill_1 FILLER_73_154 ();
 sg13g2_fill_1 FILLER_73_186 ();
 sg13g2_fill_1 FILLER_73_191 ();
 sg13g2_fill_1 FILLER_73_206 ();
 sg13g2_fill_2 FILLER_73_239 ();
 sg13g2_fill_1 FILLER_73_246 ();
 sg13g2_fill_1 FILLER_73_253 ();
 sg13g2_fill_1 FILLER_73_272 ();
 sg13g2_fill_1 FILLER_73_293 ();
 sg13g2_fill_1 FILLER_73_360 ();
 sg13g2_fill_1 FILLER_73_371 ();
 sg13g2_fill_2 FILLER_73_402 ();
 sg13g2_fill_2 FILLER_73_417 ();
 sg13g2_fill_1 FILLER_73_424 ();
 sg13g2_fill_1 FILLER_73_429 ();
 sg13g2_fill_1 FILLER_74_8 ();
 sg13g2_fill_1 FILLER_74_35 ();
 sg13g2_fill_1 FILLER_74_44 ();
 sg13g2_fill_1 FILLER_74_75 ();
 sg13g2_fill_1 FILLER_74_158 ();
 sg13g2_fill_2 FILLER_74_186 ();
 sg13g2_fill_1 FILLER_74_193 ();
 sg13g2_fill_1 FILLER_74_207 ();
 sg13g2_fill_1 FILLER_74_310 ();
 sg13g2_fill_1 FILLER_74_319 ();
 sg13g2_fill_1 FILLER_74_328 ();
 sg13g2_fill_1 FILLER_74_346 ();
 sg13g2_fill_1 FILLER_74_352 ();
 sg13g2_fill_1 FILLER_74_357 ();
 sg13g2_fill_1 FILLER_74_362 ();
 sg13g2_fill_2 FILLER_74_424 ();
 sg13g2_fill_1 FILLER_75_39 ();
 sg13g2_fill_2 FILLER_75_81 ();
 sg13g2_fill_1 FILLER_75_155 ();
 sg13g2_fill_1 FILLER_75_169 ();
 sg13g2_fill_1 FILLER_75_210 ();
 sg13g2_fill_1 FILLER_75_279 ();
 sg13g2_fill_1 FILLER_75_284 ();
 sg13g2_fill_1 FILLER_75_301 ();
 sg13g2_fill_1 FILLER_75_311 ();
 sg13g2_fill_1 FILLER_75_338 ();
 sg13g2_fill_1 FILLER_75_372 ();
 sg13g2_fill_1 FILLER_75_377 ();
 sg13g2_fill_1 FILLER_75_386 ();
 sg13g2_fill_1 FILLER_75_411 ();
 sg13g2_fill_2 FILLER_76_207 ();
 sg13g2_fill_1 FILLER_76_213 ();
 sg13g2_fill_2 FILLER_76_262 ();
 sg13g2_fill_1 FILLER_76_281 ();
 sg13g2_fill_1 FILLER_76_337 ();
 sg13g2_fill_2 FILLER_76_346 ();
 sg13g2_fill_1 FILLER_76_356 ();
 sg13g2_fill_1 FILLER_76_365 ();
 sg13g2_fill_1 FILLER_76_370 ();
 sg13g2_fill_1 FILLER_76_378 ();
 sg13g2_fill_1 FILLER_76_403 ();
 sg13g2_fill_2 FILLER_76_425 ();
 sg13g2_fill_2 FILLER_77_0 ();
 sg13g2_fill_1 FILLER_77_32 ();
 sg13g2_fill_1 FILLER_77_156 ();
 sg13g2_fill_1 FILLER_77_161 ();
 sg13g2_fill_1 FILLER_77_175 ();
 sg13g2_fill_2 FILLER_77_184 ();
 sg13g2_fill_1 FILLER_77_220 ();
 sg13g2_fill_2 FILLER_77_233 ();
 sg13g2_fill_2 FILLER_77_269 ();
 sg13g2_fill_1 FILLER_77_279 ();
 sg13g2_fill_1 FILLER_77_293 ();
 sg13g2_fill_1 FILLER_77_300 ();
 sg13g2_fill_1 FILLER_77_372 ();
 sg13g2_fill_2 FILLER_77_408 ();
 sg13g2_fill_1 FILLER_77_429 ();
 sg13g2_fill_2 FILLER_78_0 ();
 sg13g2_fill_1 FILLER_78_54 ();
 sg13g2_fill_2 FILLER_78_161 ();
 sg13g2_fill_2 FILLER_78_167 ();
 sg13g2_fill_1 FILLER_78_226 ();
 sg13g2_fill_1 FILLER_78_232 ();
 sg13g2_fill_1 FILLER_78_243 ();
 sg13g2_fill_1 FILLER_78_270 ();
 sg13g2_fill_1 FILLER_78_285 ();
 sg13g2_fill_2 FILLER_78_346 ();
 sg13g2_fill_1 FILLER_78_391 ();
 sg13g2_fill_1 FILLER_78_400 ();
 sg13g2_fill_1 FILLER_78_405 ();
 sg13g2_fill_1 FILLER_78_411 ();
 sg13g2_fill_2 FILLER_78_424 ();
 sg13g2_fill_1 FILLER_78_429 ();
 sg13g2_fill_2 FILLER_79_0 ();
 sg13g2_fill_2 FILLER_79_60 ();
 sg13g2_fill_1 FILLER_79_175 ();
 sg13g2_fill_1 FILLER_79_180 ();
 sg13g2_fill_2 FILLER_79_271 ();
 sg13g2_fill_1 FILLER_79_343 ();
 sg13g2_fill_1 FILLER_79_383 ();
 sg13g2_fill_1 FILLER_80_86 ();
 sg13g2_fill_1 FILLER_80_132 ();
 sg13g2_fill_1 FILLER_80_141 ();
 sg13g2_fill_2 FILLER_80_172 ();
 sg13g2_fill_1 FILLER_80_204 ();
 sg13g2_fill_2 FILLER_80_309 ();
 sg13g2_fill_1 FILLER_80_318 ();
 sg13g2_fill_1 FILLER_80_384 ();
 sg13g2_fill_1 FILLER_80_402 ();
 sg13g2_fill_1 FILLER_80_416 ();
endmodule
