module tt_um_algofoogle_tinyvga_fun_wrapper (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire clknet_0_clk;
 wire net83;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[2] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;
 wire \depth[0] ;
 wire \depth[1] ;
 wire \depth[2] ;
 wire \dither_threshold[0] ;
 wire \dither_threshold[1] ;
 wire \dither_threshold[2] ;
 wire \dither_threshold[3] ;
 wire \dither_threshold[4] ;
 wire \dither_threshold[5] ;
 wire \dither_threshold[6] ;
 wire hsync;
 wire \i_project.controller_0.divider[0] ;
 wire \i_project.controller_0.divider[1] ;
 wire \i_project.controller_0.grey_pass[10] ;
 wire \i_project.controller_0.grey_pass[11] ;
 wire \i_project.controller_0.grey_pass[12] ;
 wire \i_project.controller_0.grey_pass[13] ;
 wire \i_project.controller_0.grey_pass[14] ;
 wire \i_project.controller_0.grey_pass[15] ;
 wire \i_project.controller_0.h[0] ;
 wire \i_project.controller_0.h[1] ;
 wire \i_project.controller_0.h[2] ;
 wire \i_project.controller_0.h[3] ;
 wire \i_project.controller_0.h[4] ;
 wire \i_project.controller_0.h[5] ;
 wire \i_project.controller_0.h[6] ;
 wire \i_project.controller_0.h[7] ;
 wire \i_project.controller_0.h[8] ;
 wire \i_project.controller_0.h[9] ;
 wire \i_project.controller_0.mode[0] ;
 wire \i_project.controller_0.mode[1] ;
 wire \i_project.controller_0.mode[2] ;
 wire \i_project.controller_0.mode_ramp_base[0] ;
 wire \i_project.controller_0.mode_ramp_base[1] ;
 wire \i_project.controller_0.mode_ramp_base[2] ;
 wire \i_project.controller_0.mode_ramp_base[3] ;
 wire \i_project.controller_0.mode_ramp_base[4] ;
 wire \i_project.controller_0.mode_ramp_base[5] ;
 wire \i_project.controller_0.mode_ramp_base[6] ;
 wire \i_project.controller_0.mode_ramp_base[7] ;
 wire \i_project.controller_0.rst_n ;
 wire \i_project.controller_0.t[10] ;
 wire \i_project.controller_0.t[11] ;
 wire \i_project.controller_0.t[8] ;
 wire \i_project.controller_0.t[9] ;
 wire \i_project.controller_0.v[0] ;
 wire \i_project.controller_0.v[1] ;
 wire \i_project.controller_0.v[2] ;
 wire \i_project.controller_0.v[3] ;
 wire \i_project.controller_0.v[4] ;
 wire \i_project.controller_0.v[5] ;
 wire \i_project.controller_0.v[6] ;
 wire \i_project.controller_0.v[7] ;
 wire \i_project.controller_0.v[8] ;
 wire \i_project.controller_0.v[9] ;
 wire \i_project.controller_0.vga_sync.hsync ;
 wire \i_project.controller_0.vga_sync.mode ;
 wire \i_project.controller_0.vga_sync.o_vsync ;
 wire \i_project.controller_0.vga_sync.vsync ;
 wire \i_project.controller_0.voffset[0] ;
 wire \i_project.controller_0.voffset[1] ;
 wire \i_project.controller_0.voffset[2] ;
 wire \i_project.controller_0.voffset[3] ;
 wire \i_project.controller_0.voffset[4] ;
 wire \i_project.controller_0.voffset[5] ;
 wire \i_project.controller_0.voffset[6] ;
 wire \i_project.controller_0.voffset[7] ;
 wire prev_vsync;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sg13g2_xnor2_1 _2295_ (.Y(_0292_),
    .A(_0212_),
    .B(_0211_));
 sg13g2_xnor2_1 _2296_ (.Y(_0293_),
    .A(_0292_),
    .B(_2197_));
 sg13g2_xnor2_1 _2297_ (.Y(_0294_),
    .A(_2040_),
    .B(net18));
 sg13g2_nand3_1 _2298_ (.B(_0294_),
    .C(_0172_),
    .A(_0167_),
    .Y(_0295_));
 sg13g2_nand2_1 _2299_ (.Y(_0296_),
    .A(_0295_),
    .B(_2155_));
 sg13g2_nand2b_1 _2300_ (.Y(_0297_),
    .B(_0296_),
    .A_N(_0293_));
 sg13g2_nand3_1 _2301_ (.B(_2155_),
    .C(_0293_),
    .A(_0295_),
    .Y(_0298_));
 sg13g2_buf_1 _2302_ (.A(net42),
    .X(_0299_));
 sg13g2_nand3_1 _2303_ (.B(_0298_),
    .C(_0299_),
    .A(_0297_),
    .Y(_0300_));
 sg13g2_xnor2_1 _2304_ (.Y(_0301_),
    .A(_1732_),
    .B(net19));
 sg13g2_inv_1 _2305_ (.Y(_0302_),
    .A(_0301_));
 sg13g2_a21oi_1 _2306_ (.A1(_0302_),
    .A2(_0228_),
    .Y(_0303_),
    .B1(_0224_));
 sg13g2_inv_1 _2307_ (.Y(_0304_),
    .A(_0303_));
 sg13g2_nand2_1 _2308_ (.Y(_0305_),
    .A(_0300_),
    .B(_0304_));
 sg13g2_xnor2_1 _2309_ (.Y(_0306_),
    .A(_1709_),
    .B(net18));
 sg13g2_inv_1 _2310_ (.Y(_0307_),
    .A(_0306_));
 sg13g2_buf_1 _2311_ (.A(_0233_),
    .X(_0308_));
 sg13g2_a21oi_1 _2312_ (.A1(_0307_),
    .A2(_0308_),
    .Y(_0309_),
    .B1(net34));
 sg13g2_nand2_1 _2313_ (.Y(_0310_),
    .A(_0305_),
    .B(_0309_));
 sg13g2_nor2b_1 _2314_ (.A(net52),
    .B_N(_0051_),
    .Y(_0311_));
 sg13g2_a21oi_1 _2315_ (.A1(net52),
    .A2(_0048_),
    .Y(_0312_),
    .B1(_0311_));
 sg13g2_nor2_1 _2316_ (.A(net50),
    .B(_0241_),
    .Y(_0313_));
 sg13g2_a21o_1 _2317_ (.A2(_0312_),
    .A1(net50),
    .B1(_0313_),
    .X(_0314_));
 sg13g2_buf_1 _2318_ (.A(_0314_),
    .X(_0315_));
 sg13g2_xnor2_1 _2319_ (.Y(_0316_),
    .A(_0315_),
    .B(_0254_));
 sg13g2_buf_1 _2320_ (.A(_0235_),
    .X(_0317_));
 sg13g2_a21oi_1 _2321_ (.A1(_0316_),
    .A2(_0317_),
    .Y(_0318_),
    .B1(net41));
 sg13g2_nand2_1 _2322_ (.Y(_0319_),
    .A(_0310_),
    .B(_0318_));
 sg13g2_buf_1 _2323_ (.A(net41),
    .X(_0320_));
 sg13g2_a21oi_1 _2324_ (.A1(_0315_),
    .A2(net38),
    .Y(_0321_),
    .B1(_0263_));
 sg13g2_nand2_1 _2325_ (.Y(_0322_),
    .A(_0319_),
    .B(_0321_));
 sg13g2_nand2_1 _2326_ (.Y(_0323_),
    .A(_0322_),
    .B(_0289_));
 sg13g2_nand2_1 _2327_ (.Y(_0324_),
    .A(_0323_),
    .B(net43));
 sg13g2_inv_1 _2328_ (.Y(_0325_),
    .A(_2106_));
 sg13g2_buf_1 _2329_ (.A(_0046_),
    .X(_0326_));
 sg13g2_inv_1 _2330_ (.Y(_0327_),
    .A(_0326_));
 sg13g2_nor3_1 _2331_ (.A(_2107_),
    .B(_0325_),
    .C(_0327_),
    .Y(_0328_));
 sg13g2_buf_1 _2332_ (.A(_0328_),
    .X(_0329_));
 sg13g2_nand2_1 _2333_ (.Y(_0330_),
    .A(_1807_),
    .B(_2099_));
 sg13g2_nand2_2 _2334_ (.Y(_0331_),
    .A(_0330_),
    .B(_2091_));
 sg13g2_inv_2 _2335_ (.Y(_0332_),
    .A(_0331_));
 sg13g2_nand2_1 _2336_ (.Y(_0333_),
    .A(_1815_),
    .B(_0050_));
 sg13g2_nor2b_1 _2337_ (.A(_0332_),
    .B_N(_0333_),
    .Y(_0334_));
 sg13g2_buf_1 _2338_ (.A(_0334_),
    .X(_0335_));
 sg13g2_nand3_1 _2339_ (.B(net46),
    .C(_0335_),
    .A(_0324_),
    .Y(_0336_));
 sg13g2_inv_1 _2340_ (.Y(_0337_),
    .A(net42));
 sg13g2_nor2b_1 _2341_ (.A(_0208_),
    .B_N(_0207_),
    .Y(_0338_));
 sg13g2_nor2b_1 _2342_ (.A(_0338_),
    .B_N(_0191_),
    .Y(_0339_));
 sg13g2_xor2_1 _2343_ (.B(_0339_),
    .A(_0192_),
    .X(_0340_));
 sg13g2_xnor2_1 _2344_ (.Y(_0341_),
    .A(_0162_),
    .B(_0153_));
 sg13g2_xnor2_1 _2345_ (.Y(_0342_),
    .A(_0340_),
    .B(_0341_));
 sg13g2_xnor2_1 _2346_ (.Y(_0343_),
    .A(net59),
    .B(net22));
 sg13g2_a21oi_1 _2347_ (.A1(_0343_),
    .A2(_0228_),
    .Y(_0344_),
    .B1(net42));
 sg13g2_inv_1 _2348_ (.Y(_0345_),
    .A(_0344_));
 sg13g2_o21ai_1 _2349_ (.B1(_0345_),
    .Y(_0346_),
    .A1(net37),
    .A2(_0342_));
 sg13g2_xnor2_1 _2350_ (.Y(_0347_),
    .A(_1720_),
    .B(_2229_));
 sg13g2_inv_1 _2351_ (.Y(_0348_),
    .A(_0347_));
 sg13g2_a21oi_1 _2352_ (.A1(_0348_),
    .A2(net51),
    .Y(_0349_),
    .B1(net34));
 sg13g2_nand2_1 _2353_ (.Y(_0350_),
    .A(_0346_),
    .B(_0349_));
 sg13g2_inv_1 _2354_ (.Y(_0351_),
    .A(net38));
 sg13g2_buf_1 _2355_ (.A(_0254_),
    .X(_0352_));
 sg13g2_nand2_1 _2356_ (.Y(_0353_),
    .A(net52),
    .B(_0051_));
 sg13g2_inv_1 _2357_ (.Y(_0354_),
    .A(_0353_));
 sg13g2_a21oi_1 _2358_ (.A1(_1687_),
    .A2(_0053_),
    .Y(_0355_),
    .B1(_0354_));
 sg13g2_inv_1 _2359_ (.Y(_0356_),
    .A(_0355_));
 sg13g2_nand2_1 _2360_ (.Y(_0357_),
    .A(_0250_),
    .B(net50));
 sg13g2_o21ai_1 _2361_ (.B1(_0357_),
    .Y(_0358_),
    .A1(net50),
    .A2(_0356_));
 sg13g2_inv_1 _2362_ (.Y(_0359_),
    .A(_0358_));
 sg13g2_inv_1 _2363_ (.Y(_0360_),
    .A(_0235_));
 sg13g2_a21oi_1 _2364_ (.A1(_0352_),
    .A2(_0359_),
    .Y(_0361_),
    .B1(_0360_));
 sg13g2_o21ai_1 _2365_ (.B1(_0361_),
    .Y(_0362_),
    .A1(net29),
    .A2(_0359_));
 sg13g2_nand3_1 _2366_ (.B(net33),
    .C(_0362_),
    .A(_0350_),
    .Y(_0363_));
 sg13g2_buf_1 _2367_ (.A(net41),
    .X(_0364_));
 sg13g2_buf_1 _2368_ (.A(net27),
    .X(_0365_));
 sg13g2_a21oi_1 _2369_ (.A1(_0358_),
    .A2(net36),
    .Y(_0366_),
    .B1(net25));
 sg13g2_nand2_1 _2370_ (.Y(_0367_),
    .A(_0363_),
    .B(_0366_));
 sg13g2_nand2_1 _2371_ (.Y(_0368_),
    .A(_0367_),
    .B(net17));
 sg13g2_nand2_1 _2372_ (.Y(_0369_),
    .A(_0368_),
    .B(net43));
 sg13g2_nand2_2 _2373_ (.Y(_0370_),
    .A(_2106_),
    .B(_2107_));
 sg13g2_nor2_1 _2374_ (.A(_0326_),
    .B(_0370_),
    .Y(_0371_));
 sg13g2_nor3_2 _2375_ (.A(_2107_),
    .B(_0325_),
    .C(_2108_),
    .Y(_0372_));
 sg13g2_inv_1 _2376_ (.Y(_0373_),
    .A(_2107_));
 sg13g2_nor3_1 _2377_ (.A(_2106_),
    .B(_0373_),
    .C(_2108_),
    .Y(_0374_));
 sg13g2_nor3_1 _2378_ (.A(_0371_),
    .B(_0372_),
    .C(_0374_),
    .Y(_0375_));
 sg13g2_nor2_1 _2379_ (.A(_0375_),
    .B(_0332_),
    .Y(_0376_));
 sg13g2_inv_1 _2380_ (.Y(_0377_),
    .A(_0376_));
 sg13g2_a21oi_1 _2381_ (.A1(_0018_),
    .A2(net49),
    .Y(_0378_),
    .B1(_0377_));
 sg13g2_a21oi_1 _2382_ (.A1(_0325_),
    .A2(_0373_),
    .Y(_0379_),
    .B1(_0327_));
 sg13g2_inv_1 _2383_ (.Y(_0380_),
    .A(_0370_));
 sg13g2_nor2_1 _2384_ (.A(\depth[2] ),
    .B(_0380_),
    .Y(_0381_));
 sg13g2_inv_1 _2385_ (.Y(_0382_),
    .A(_0381_));
 sg13g2_nor2_1 _2386_ (.A(_0379_),
    .B(_0382_),
    .Y(_0383_));
 sg13g2_buf_1 _2387_ (.A(_0383_),
    .X(_0384_));
 sg13g2_a21oi_1 _2388_ (.A1(_0369_),
    .A2(_0378_),
    .Y(_0385_),
    .B1(_0384_));
 sg13g2_nand2_1 _2389_ (.Y(_0386_),
    .A(_0336_),
    .B(_0385_));
 sg13g2_inv_1 _2390_ (.Y(_0387_),
    .A(_0153_));
 sg13g2_nand2_1 _2391_ (.Y(_0388_),
    .A(_0172_),
    .B(_0162_));
 sg13g2_nand2_1 _2392_ (.Y(_0389_),
    .A(_2197_),
    .B(_0294_));
 sg13g2_nor3_1 _2393_ (.A(_0387_),
    .B(_0388_),
    .C(_0389_),
    .Y(_0390_));
 sg13g2_a21oi_1 _2394_ (.A1(_0170_),
    .A2(_0165_),
    .Y(_0391_),
    .B1(_2134_));
 sg13g2_nand2_1 _2395_ (.Y(_0392_),
    .A(net19),
    .B(_2184_));
 sg13g2_a21oi_1 _2396_ (.A1(_2153_),
    .A2(_0392_),
    .Y(_0393_),
    .B1(_2201_));
 sg13g2_o21ai_1 _2397_ (.B1(_0393_),
    .Y(_0394_),
    .A1(_0391_),
    .A2(_0389_));
 sg13g2_nor2_1 _2398_ (.A(_0390_),
    .B(_0394_),
    .Y(_0395_));
 sg13g2_nor2b_1 _2399_ (.A(_0218_),
    .B_N(_0217_),
    .Y(_0396_));
 sg13g2_nand2_1 _2400_ (.Y(_0397_),
    .A(_2208_),
    .B(_0396_));
 sg13g2_inv_1 _2401_ (.Y(_0398_),
    .A(_0396_));
 sg13g2_nand2_1 _2402_ (.Y(_0399_),
    .A(_2183_),
    .B(_0398_));
 sg13g2_nand3_1 _2403_ (.B(_0399_),
    .C(_0215_),
    .A(_0397_),
    .Y(_0400_));
 sg13g2_nand2_1 _2404_ (.Y(_0401_),
    .A(_2183_),
    .B(_0396_));
 sg13g2_nand3_1 _2405_ (.B(_2182_),
    .C(_0398_),
    .A(_2181_),
    .Y(_0402_));
 sg13g2_nand3_1 _2406_ (.B(_0402_),
    .C(_0216_),
    .A(_0401_),
    .Y(_0403_));
 sg13g2_nand2_1 _2407_ (.Y(_0404_),
    .A(_0400_),
    .B(_0403_));
 sg13g2_nand2_1 _2408_ (.Y(_0405_),
    .A(_0395_),
    .B(_0404_));
 sg13g2_nand3_1 _2409_ (.B(_0399_),
    .C(_0216_),
    .A(_0397_),
    .Y(_0406_));
 sg13g2_nand3_1 _2410_ (.B(_0402_),
    .C(_0215_),
    .A(_0401_),
    .Y(_0407_));
 sg13g2_nand2_1 _2411_ (.Y(_0408_),
    .A(_0406_),
    .B(_0407_));
 sg13g2_nor2_1 _2412_ (.A(_0391_),
    .B(_0389_),
    .Y(_0409_));
 sg13g2_nor2b_1 _2413_ (.A(_0409_),
    .B_N(_0393_),
    .Y(_0410_));
 sg13g2_nor2_1 _2414_ (.A(_0388_),
    .B(_0389_),
    .Y(_0411_));
 sg13g2_nand2_1 _2415_ (.Y(_0412_),
    .A(_0411_),
    .B(_0153_));
 sg13g2_nand2_1 _2416_ (.Y(_0413_),
    .A(_0410_),
    .B(_0412_));
 sg13g2_nand2_1 _2417_ (.Y(_0414_),
    .A(_0408_),
    .B(_0413_));
 sg13g2_nand3_1 _2418_ (.B(_0414_),
    .C(_0225_),
    .A(_0405_),
    .Y(_0415_));
 sg13g2_a21o_1 _2419_ (.A2(_0228_),
    .A1(_0232_),
    .B1(_0224_),
    .X(_0416_));
 sg13g2_nand2_1 _2420_ (.Y(_0417_),
    .A(_0415_),
    .B(_0416_));
 sg13g2_a21oi_1 _2421_ (.A1(_0302_),
    .A2(net51),
    .Y(_0418_),
    .B1(net34));
 sg13g2_nand2_1 _2422_ (.Y(_0419_),
    .A(_0417_),
    .B(_0418_));
 sg13g2_inv_1 _2423_ (.Y(_0420_),
    .A(_0027_));
 sg13g2_a21oi_1 _2424_ (.A1(_0420_),
    .A2(_1687_),
    .Y(_0421_),
    .B1(net50));
 sg13g2_nand2b_1 _2425_ (.Y(_0422_),
    .B(_0238_),
    .A_N(_0049_));
 sg13g2_nand2_1 _2426_ (.Y(_0423_),
    .A(_0239_),
    .B(_1686_));
 sg13g2_o21ai_1 _2427_ (.B1(_0423_),
    .Y(_0424_),
    .A1(net52),
    .A2(_0048_));
 sg13g2_inv_1 _2428_ (.Y(_0425_),
    .A(_0424_));
 sg13g2_a22oi_1 _2429_ (.Y(_0426_),
    .B1(_1691_),
    .B2(_0425_),
    .A2(_0422_),
    .A1(_0421_));
 sg13g2_xnor2_1 _2430_ (.Y(_0427_),
    .A(_0426_),
    .B(_0254_));
 sg13g2_a21oi_1 _2431_ (.A1(_0427_),
    .A2(net34),
    .Y(_0428_),
    .B1(net41));
 sg13g2_nand2_1 _2432_ (.Y(_0429_),
    .A(_0419_),
    .B(_0428_));
 sg13g2_a21oi_1 _2433_ (.A1(_0426_),
    .A2(net38),
    .Y(_0430_),
    .B1(net27));
 sg13g2_nand2_1 _2434_ (.Y(_0431_),
    .A(_0429_),
    .B(_0430_));
 sg13g2_nor2_2 _2435_ (.A(_1815_),
    .B(_0287_),
    .Y(_0432_));
 sg13g2_nand2_1 _2436_ (.Y(_0433_),
    .A(_0431_),
    .B(_0432_));
 sg13g2_nor2_1 _2437_ (.A(_0047_),
    .B(_2092_),
    .Y(_0434_));
 sg13g2_inv_1 _2438_ (.Y(_0435_),
    .A(_0434_));
 sg13g2_nand2_1 _2439_ (.Y(_0436_),
    .A(_0433_),
    .B(_0435_));
 sg13g2_nor2_1 _2440_ (.A(_0327_),
    .B(_0370_),
    .Y(_0437_));
 sg13g2_inv_1 _2441_ (.Y(_0438_),
    .A(_0437_));
 sg13g2_nor2_1 _2442_ (.A(_0438_),
    .B(_0332_),
    .Y(_0439_));
 sg13g2_buf_2 _2443_ (.A(_0439_),
    .X(_0440_));
 sg13g2_nand2_1 _2444_ (.Y(_0441_),
    .A(_0436_),
    .B(_0440_));
 sg13g2_nor2b_1 _2445_ (.A(_0386_),
    .B_N(_0441_),
    .Y(_0442_));
 sg13g2_a21oi_1 _2446_ (.A1(_0433_),
    .A2(_0435_),
    .Y(_0443_),
    .B1(_0332_));
 sg13g2_nor3_1 _2447_ (.A(_2106_),
    .B(_0373_),
    .C(_0327_),
    .Y(_0444_));
 sg13g2_buf_2 _2448_ (.A(_0444_),
    .X(_0445_));
 sg13g2_nand2_1 _2449_ (.Y(_0446_),
    .A(_0443_),
    .B(_0445_));
 sg13g2_nand2_1 _2450_ (.Y(_0447_),
    .A(_0442_),
    .B(_0446_));
 sg13g2_nor2_1 _2451_ (.A(_0291_),
    .B(_0447_),
    .Y(_0448_));
 sg13g2_inv_1 _2452_ (.Y(_0449_),
    .A(_0372_));
 sg13g2_nand2_1 _2453_ (.Y(_0450_),
    .A(_0265_),
    .B(_0289_));
 sg13g2_nand2_1 _2454_ (.Y(_0451_),
    .A(_0450_),
    .B(net43));
 sg13g2_nand2_1 _2455_ (.Y(_0452_),
    .A(_0451_),
    .B(_2104_));
 sg13g2_buf_8 _2456_ (.A(_0452_),
    .X(_0453_));
 sg13g2_nor2_1 _2457_ (.A(_0449_),
    .B(_0453_),
    .Y(_0454_));
 sg13g2_inv_1 _2458_ (.Y(_0455_),
    .A(_0374_));
 sg13g2_nor2_1 _2459_ (.A(_0455_),
    .B(_0332_),
    .Y(_0456_));
 sg13g2_nand2_1 _2460_ (.Y(_0457_),
    .A(_0436_),
    .B(_0456_));
 sg13g2_a21oi_1 _2461_ (.A1(_0207_),
    .A2(_0209_),
    .Y(_0458_),
    .B1(_0194_));
 sg13g2_o21ai_1 _2462_ (.B1(_0199_),
    .Y(_0459_),
    .A1(_0197_),
    .A2(_0458_));
 sg13g2_xnor2_1 _2463_ (.Y(_0460_),
    .A(_0195_),
    .B(_0459_));
 sg13g2_nor2b_1 _2464_ (.A(_2153_),
    .B_N(_2154_),
    .Y(_0461_));
 sg13g2_xnor2_1 _2465_ (.Y(_0462_),
    .A(_0460_),
    .B(_0461_));
 sg13g2_a21oi_1 _2466_ (.A1(_0167_),
    .A2(_0172_),
    .Y(_0463_),
    .B1(_2134_));
 sg13g2_xnor2_1 _2467_ (.Y(_0464_),
    .A(_0462_),
    .B(_0463_));
 sg13g2_nand2_1 _2468_ (.Y(_0465_),
    .A(_0464_),
    .B(net40));
 sg13g2_a21oi_1 _2469_ (.A1(_0307_),
    .A2(_0228_),
    .Y(_0466_),
    .B1(_0224_));
 sg13g2_inv_1 _2470_ (.Y(_0467_),
    .A(_0466_));
 sg13g2_nand2_1 _2471_ (.Y(_0468_),
    .A(_0465_),
    .B(_0467_));
 sg13g2_xnor2_1 _2472_ (.Y(_0469_),
    .A(_1742_),
    .B(net20));
 sg13g2_inv_1 _2473_ (.Y(_0470_),
    .A(_0469_));
 sg13g2_a21oi_1 _2474_ (.A1(_0470_),
    .A2(net51),
    .Y(_0471_),
    .B1(net39));
 sg13g2_nand2_1 _2475_ (.Y(_0472_),
    .A(_0468_),
    .B(_0471_));
 sg13g2_nand2_1 _2476_ (.Y(_0473_),
    .A(_0355_),
    .B(net50));
 sg13g2_o21ai_1 _2477_ (.B1(_0473_),
    .Y(_0474_),
    .A1(net50),
    .A2(_0425_));
 sg13g2_xnor2_1 _2478_ (.Y(_0475_),
    .A(_0474_),
    .B(_0352_));
 sg13g2_a21oi_1 _2479_ (.A1(_0475_),
    .A2(net39),
    .Y(_0476_),
    .B1(net38));
 sg13g2_nand2_1 _2480_ (.Y(_0477_),
    .A(_0472_),
    .B(_0476_));
 sg13g2_a21oi_1 _2481_ (.A1(_0474_),
    .A2(net36),
    .Y(_0478_),
    .B1(net25));
 sg13g2_nand2_1 _2482_ (.Y(_0479_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_nand2_1 _2483_ (.Y(_0480_),
    .A(_0479_),
    .B(_0432_));
 sg13g2_nand2b_1 _2484_ (.Y(_0481_),
    .B(_1816_),
    .A_N(_0052_));
 sg13g2_nand2_1 _2485_ (.Y(_0482_),
    .A(_0480_),
    .B(_0481_));
 sg13g2_buf_1 _2486_ (.A(net36),
    .X(_0483_));
 sg13g2_inv_1 _2487_ (.Y(_0484_),
    .A(_0251_));
 sg13g2_xor2_1 _2488_ (.B(_0204_),
    .A(_0203_),
    .X(_0485_));
 sg13g2_nor2b_1 _2489_ (.A(_2219_),
    .B_N(_2214_),
    .Y(_0486_));
 sg13g2_xnor2_1 _2490_ (.Y(_0487_),
    .A(_2218_),
    .B(_0486_));
 sg13g2_xnor2_1 _2491_ (.Y(_0488_),
    .A(_0485_),
    .B(_0487_));
 sg13g2_xnor2_1 _2492_ (.Y(_0489_),
    .A(_1715_),
    .B(_0282_));
 sg13g2_o21ai_1 _2493_ (.B1(net37),
    .Y(_0490_),
    .A1(_0229_),
    .A2(_0489_));
 sg13g2_o21ai_1 _2494_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net37),
    .A2(_0488_));
 sg13g2_xnor2_1 _2495_ (.Y(_0492_),
    .A(net60),
    .B(net35));
 sg13g2_buf_1 _2496_ (.A(net34),
    .X(_0493_));
 sg13g2_a21oi_1 _2497_ (.A1(_0492_),
    .A2(net51),
    .Y(_0494_),
    .B1(net31));
 sg13g2_nand2_1 _2498_ (.Y(_0495_),
    .A(_0491_),
    .B(_0494_));
 sg13g2_xnor2_1 _2499_ (.Y(_0496_),
    .A(_0484_),
    .B(net29));
 sg13g2_a21oi_1 _2500_ (.A1(_0496_),
    .A2(net31),
    .Y(_0497_),
    .B1(net36));
 sg13g2_a221oi_1 _2501_ (.B2(_0497_),
    .C1(net25),
    .B1(_0495_),
    .A1(net32),
    .Y(_0498_),
    .A2(_0484_));
 sg13g2_nor4_1 _2502_ (.A(_0326_),
    .B(net49),
    .C(_0370_),
    .D(_0330_),
    .Y(_0499_));
 sg13g2_nand2_1 _2503_ (.Y(_0500_),
    .A(net17),
    .B(_0499_));
 sg13g2_inv_2 _2504_ (.Y(_0501_),
    .A(_0384_));
 sg13g2_o21ai_1 _2505_ (.B1(_0501_),
    .Y(_0502_),
    .A1(_0498_),
    .A2(_0500_));
 sg13g2_a21oi_1 _2506_ (.A1(_0482_),
    .A2(_0440_),
    .Y(_0503_),
    .B1(_0502_));
 sg13g2_nand2_1 _2507_ (.Y(_0504_),
    .A(_0457_),
    .B(_0503_));
 sg13g2_nand3_1 _2508_ (.B(net47),
    .C(_0335_),
    .A(_0324_),
    .Y(_0505_));
 sg13g2_nor2b_1 _2509_ (.A(_0504_),
    .B_N(_0505_),
    .Y(_0506_));
 sg13g2_o21ai_1 _2510_ (.B1(_0443_),
    .Y(_0507_),
    .A1(_0445_),
    .A2(net46));
 sg13g2_nand2_1 _2511_ (.Y(_0508_),
    .A(_0506_),
    .B(_0507_));
 sg13g2_nor2_1 _2512_ (.A(_0454_),
    .B(_0508_),
    .Y(_0509_));
 sg13g2_nor2_1 _2513_ (.A(_0448_),
    .B(_0509_),
    .Y(_0510_));
 sg13g2_buf_1 _2514_ (.A(_0384_),
    .X(_0511_));
 sg13g2_nand2_2 _2515_ (.Y(_0512_),
    .A(_0453_),
    .B(_0511_));
 sg13g2_nor2_1 _2516_ (.A(_0381_),
    .B(_0332_),
    .Y(_0513_));
 sg13g2_a21oi_1 _2517_ (.A1(_0482_),
    .A2(_0513_),
    .Y(_0514_),
    .B1(net24));
 sg13g2_nand2_1 _2518_ (.Y(_0515_),
    .A(_0446_),
    .B(_0514_));
 sg13g2_nand2_1 _2519_ (.Y(_0516_),
    .A(_0512_),
    .B(_0515_));
 sg13g2_inv_1 _2520_ (.Y(_0517_),
    .A(_0453_));
 sg13g2_nand2_1 _2521_ (.Y(_0518_),
    .A(_0517_),
    .B(net46));
 sg13g2_nand2_2 _2522_ (.Y(_0519_),
    .A(_0516_),
    .B(_0518_));
 sg13g2_nand2_1 _2523_ (.Y(_0520_),
    .A(_0510_),
    .B(_0519_));
 sg13g2_nand3_1 _2524_ (.B(_0331_),
    .C(net47),
    .A(_0436_),
    .Y(_0521_));
 sg13g2_nand2_1 _2525_ (.Y(_0522_),
    .A(_0521_),
    .B(_0501_));
 sg13g2_nor2_1 _2526_ (.A(_0440_),
    .B(_0376_),
    .Y(_0523_));
 sg13g2_inv_1 _2527_ (.Y(_0524_),
    .A(_0523_));
 sg13g2_nand2_1 _2528_ (.Y(_0525_),
    .A(_0436_),
    .B(_0524_));
 sg13g2_nand3b_1 _2529_ (.B(_0507_),
    .C(_0525_),
    .Y(_0526_),
    .A_N(_0522_));
 sg13g2_nand2_2 _2530_ (.Y(_0527_),
    .A(_0526_),
    .B(_0512_));
 sg13g2_inv_4 _2531_ (.A(_0527_),
    .Y(_0528_));
 sg13g2_nand2_1 _2532_ (.Y(_0529_),
    .A(_0520_),
    .B(_0528_));
 sg13g2_nor2_1 _2533_ (.A(_0445_),
    .B(net24),
    .Y(_0530_));
 sg13g2_nand2_1 _2534_ (.Y(_0531_),
    .A(_0324_),
    .B(_0335_));
 sg13g2_inv_1 _2535_ (.Y(_0532_),
    .A(_0531_));
 sg13g2_inv_1 _2536_ (.Y(_0533_),
    .A(_0329_));
 sg13g2_nand2_1 _2537_ (.Y(_0534_),
    .A(_0533_),
    .B(_0381_));
 sg13g2_nand2_1 _2538_ (.Y(_0535_),
    .A(_0532_),
    .B(_0534_));
 sg13g2_o21ai_1 _2539_ (.B1(_0535_),
    .Y(_0536_),
    .A1(_0530_),
    .A2(_0453_));
 sg13g2_nor2_1 _2540_ (.A(_0371_),
    .B(_0372_),
    .Y(_0537_));
 sg13g2_nor4_2 _2541_ (.A(net49),
    .B(_0330_),
    .C(_0537_),
    .Y(_0538_),
    .D(_0287_));
 sg13g2_inv_1 _2542_ (.Y(_0539_),
    .A(_0233_));
 sg13g2_buf_1 _2543_ (.A(_0539_),
    .X(_0540_));
 sg13g2_buf_1 _2544_ (.A(_0360_),
    .X(_0541_));
 sg13g2_o21ai_1 _2545_ (.B1(net30),
    .Y(_0542_),
    .A1(net45),
    .A2(_0489_));
 sg13g2_xnor2_1 _2546_ (.Y(_0543_),
    .A(_0208_),
    .B(_0207_));
 sg13g2_xnor2_1 _2547_ (.Y(_0544_),
    .A(_2220_),
    .B(_0148_));
 sg13g2_xnor2_1 _2548_ (.Y(_0545_),
    .A(_0543_),
    .B(_0544_));
 sg13g2_a21oi_1 _2549_ (.A1(_0348_),
    .A2(_0228_),
    .Y(_0546_),
    .B1(net42));
 sg13g2_a21oi_1 _2550_ (.A1(_0545_),
    .A2(net40),
    .Y(_0547_),
    .B1(_0546_));
 sg13g2_nand2_1 _2551_ (.Y(_0548_),
    .A(_1687_),
    .B(_0038_));
 sg13g2_a21oi_1 _2552_ (.A1(net52),
    .A2(_0037_),
    .Y(_0549_),
    .B1(_1689_));
 sg13g2_nand2_1 _2553_ (.Y(_0550_),
    .A(net52),
    .B(_0053_));
 sg13g2_o21ai_1 _2554_ (.B1(_0550_),
    .Y(_0551_),
    .A1(net52),
    .A2(_1800_));
 sg13g2_inv_1 _2555_ (.Y(_0552_),
    .A(_0551_));
 sg13g2_a22oi_1 _2556_ (.Y(_0553_),
    .B1(_1689_),
    .B2(_0552_),
    .A2(_0549_),
    .A1(_0548_));
 sg13g2_buf_1 _2557_ (.A(net29),
    .X(_0554_));
 sg13g2_xor2_1 _2558_ (.B(_0554_),
    .A(_0553_),
    .X(_0555_));
 sg13g2_a21oi_1 _2559_ (.A1(_0555_),
    .A2(net31),
    .Y(_0556_),
    .B1(net32));
 sg13g2_o21ai_1 _2560_ (.B1(_0556_),
    .Y(_0557_),
    .A1(_0542_),
    .A2(_0547_));
 sg13g2_nand2b_1 _2561_ (.Y(_0558_),
    .B(net32),
    .A_N(_0553_));
 sg13g2_nand3_1 _2562_ (.B(_0262_),
    .C(_0558_),
    .A(_0557_),
    .Y(_0559_));
 sg13g2_nand2_1 _2563_ (.Y(_0560_),
    .A(_0538_),
    .B(_0559_));
 sg13g2_o21ai_1 _2564_ (.B1(_0560_),
    .Y(_0561_),
    .A1(_0438_),
    .A2(_0531_));
 sg13g2_nor2_1 _2565_ (.A(_0561_),
    .B(_0522_),
    .Y(_0562_));
 sg13g2_a21oi_1 _2566_ (.A1(_0379_),
    .A2(_0370_),
    .Y(_0563_),
    .B1(_0374_));
 sg13g2_inv_1 _2567_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nand3_1 _2568_ (.B(_2104_),
    .C(_0564_),
    .A(_0451_),
    .Y(_0565_));
 sg13g2_nand2_1 _2569_ (.Y(_0566_),
    .A(_0562_),
    .B(_0565_));
 sg13g2_nand2_1 _2570_ (.Y(_0567_),
    .A(_2107_),
    .B(_0326_));
 sg13g2_nand2_1 _2571_ (.Y(_0568_),
    .A(_0501_),
    .B(_0567_));
 sg13g2_nand3_1 _2572_ (.B(_2104_),
    .C(_0568_),
    .A(_0451_),
    .Y(_0569_));
 sg13g2_a21o_1 _2573_ (.A2(net51),
    .A1(_0343_),
    .B1(net31),
    .X(_0570_));
 sg13g2_xnor2_1 _2574_ (.Y(_0571_),
    .A(_0197_),
    .B(_0458_));
 sg13g2_xnor2_1 _2575_ (.Y(_0572_),
    .A(_0172_),
    .B(_0167_));
 sg13g2_xnor2_1 _2576_ (.Y(_0573_),
    .A(_0571_),
    .B(_0572_));
 sg13g2_a21oi_1 _2577_ (.A1(_0470_),
    .A2(_0228_),
    .Y(_0574_),
    .B1(net42));
 sg13g2_a21oi_1 _2578_ (.A1(_0573_),
    .A2(_0299_),
    .Y(_0575_),
    .B1(_0574_));
 sg13g2_nor2_1 _2579_ (.A(_1689_),
    .B(_0551_),
    .Y(_0576_));
 sg13g2_a21o_1 _2580_ (.A2(_0312_),
    .A1(_1689_),
    .B1(_0576_),
    .X(_0577_));
 sg13g2_xnor2_1 _2581_ (.Y(_0578_),
    .A(_0577_),
    .B(_0554_));
 sg13g2_a21oi_1 _2582_ (.A1(_0578_),
    .A2(_0493_),
    .Y(_0579_),
    .B1(net32));
 sg13g2_o21ai_1 _2583_ (.B1(_0579_),
    .Y(_0580_),
    .A1(_0570_),
    .A2(_0575_));
 sg13g2_a21oi_1 _2584_ (.A1(_0577_),
    .A2(_0483_),
    .Y(_0581_),
    .B1(net25));
 sg13g2_a21oi_1 _2585_ (.A1(_0580_),
    .A2(_0581_),
    .Y(_0582_),
    .B1(_0287_));
 sg13g2_nand2b_1 _2586_ (.Y(_0583_),
    .B(_2092_),
    .A_N(_0582_));
 sg13g2_nand3_1 _2587_ (.B(_0438_),
    .C(_0382_),
    .A(_0331_),
    .Y(_0584_));
 sg13g2_a21oi_1 _2588_ (.A1(_0017_),
    .A2(net49),
    .Y(_0585_),
    .B1(_0584_));
 sg13g2_a22oi_1 _2589_ (.Y(_0586_),
    .B1(net46),
    .B2(_0443_),
    .A2(_0585_),
    .A1(_0583_));
 sg13g2_nand2_1 _2590_ (.Y(_0587_),
    .A(_0569_),
    .B(_0586_));
 sg13g2_nand3_1 _2591_ (.B(_0566_),
    .C(_0587_),
    .A(_0536_),
    .Y(_0588_));
 sg13g2_nand2_1 _2592_ (.Y(_0589_),
    .A(_0588_),
    .B(_0517_));
 sg13g2_nand2_1 _2593_ (.Y(_0590_),
    .A(_0529_),
    .B(_0589_));
 sg13g2_nor2_1 _2594_ (.A(_0453_),
    .B(_0519_),
    .Y(_0591_));
 sg13g2_nand3_1 _2595_ (.B(_0336_),
    .C(_0385_),
    .A(_0441_),
    .Y(_0592_));
 sg13g2_nor2b_1 _2596_ (.A(_0592_),
    .B_N(_0446_),
    .Y(_0593_));
 sg13g2_nand3_1 _2597_ (.B(_2104_),
    .C(net47),
    .A(_0451_),
    .Y(_0594_));
 sg13g2_nand2_1 _2598_ (.Y(_0595_),
    .A(_0593_),
    .B(_0594_));
 sg13g2_nand3_1 _2599_ (.B(_0587_),
    .C(_0512_),
    .A(_0595_),
    .Y(_0596_));
 sg13g2_nand2_1 _2600_ (.Y(_0597_),
    .A(_0591_),
    .B(_0596_));
 sg13g2_inv_1 _2601_ (.Y(_0598_),
    .A(_0536_));
 sg13g2_a21oi_1 _2602_ (.A1(_0526_),
    .A2(_0517_),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_nand2_1 _2603_ (.Y(_0600_),
    .A(_0597_),
    .B(_0599_));
 sg13g2_nand3_1 _2604_ (.B(_0566_),
    .C(_0512_),
    .A(_0595_),
    .Y(_0601_));
 sg13g2_inv_1 _2605_ (.Y(_0602_),
    .A(_0587_));
 sg13g2_nand2_1 _2606_ (.Y(_0603_),
    .A(_0601_),
    .B(_0602_));
 sg13g2_nor2_1 _2607_ (.A(_0517_),
    .B(_0516_),
    .Y(_0604_));
 sg13g2_nand2_1 _2608_ (.Y(_0605_),
    .A(_0603_),
    .B(_0604_));
 sg13g2_nand3_1 _2609_ (.B(_0600_),
    .C(_0605_),
    .A(_0590_),
    .Y(_0606_));
 sg13g2_buf_1 _2610_ (.A(_0606_),
    .X(_0607_));
 sg13g2_nand4_1 _2611_ (.B(_0600_),
    .C(_0605_),
    .A(_0590_),
    .Y(_0608_),
    .D(_0528_));
 sg13g2_nand2_1 _2612_ (.Y(_0609_),
    .A(_0607_),
    .B(_0527_));
 sg13g2_nand2_2 _2613_ (.Y(_0610_),
    .A(_0608_),
    .B(_0609_));
 sg13g2_nor2_1 _2614_ (.A(_0519_),
    .B(_0610_),
    .Y(_0611_));
 sg13g2_inv_1 _2615_ (.Y(_0612_),
    .A(_0519_));
 sg13g2_xnor2_1 _2616_ (.Y(_0613_),
    .A(_0528_),
    .B(_0607_));
 sg13g2_buf_2 _2617_ (.A(_0613_),
    .X(_0614_));
 sg13g2_nor2_1 _2618_ (.A(_0612_),
    .B(_0614_),
    .Y(_0615_));
 sg13g2_nor2_1 _2619_ (.A(_0611_),
    .B(_0615_),
    .Y(_0616_));
 sg13g2_xnor2_1 _2620_ (.Y(_0617_),
    .A(_0517_),
    .B(_0527_));
 sg13g2_nand4_1 _2621_ (.B(_0600_),
    .C(_0605_),
    .A(_0590_),
    .Y(_0618_),
    .D(_0617_));
 sg13g2_nand2_1 _2622_ (.Y(_0619_),
    .A(_0607_),
    .B(_0453_));
 sg13g2_nand2_2 _2623_ (.Y(_0620_),
    .A(_0618_),
    .B(_0619_));
 sg13g2_xnor2_1 _2624_ (.Y(_0621_),
    .A(_0598_),
    .B(_0620_));
 sg13g2_nand2_1 _2625_ (.Y(_0622_),
    .A(_0616_),
    .B(_0621_));
 sg13g2_inv_1 _2626_ (.Y(_0623_),
    .A(_0622_));
 sg13g2_inv_1 _2627_ (.Y(_0624_),
    .A(_0512_));
 sg13g2_nor2_1 _2628_ (.A(_0624_),
    .B(_0509_),
    .Y(_0625_));
 sg13g2_inv_1 _2629_ (.Y(_0626_),
    .A(_0625_));
 sg13g2_nand2_2 _2630_ (.Y(_0627_),
    .A(_0614_),
    .B(_0626_));
 sg13g2_nand2_1 _2631_ (.Y(_0628_),
    .A(_0566_),
    .B(_0512_));
 sg13g2_nand3_1 _2632_ (.B(_0619_),
    .C(_0628_),
    .A(_0618_),
    .Y(_0629_));
 sg13g2_inv_1 _2633_ (.Y(_0630_),
    .A(_0628_));
 sg13g2_nand2_1 _2634_ (.Y(_0631_),
    .A(_0620_),
    .B(_0630_));
 sg13g2_inv_1 _2635_ (.Y(_0632_),
    .A(_0631_));
 sg13g2_a21oi_1 _2636_ (.A1(_0627_),
    .A2(_0629_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_inv_2 _2637_ (.Y(_0634_),
    .A(_0633_));
 sg13g2_nor2_1 _2638_ (.A(_0624_),
    .B(_0448_),
    .Y(_0635_));
 sg13g2_nand2_1 _2639_ (.Y(_0636_),
    .A(_0610_),
    .B(_0635_));
 sg13g2_inv_1 _2640_ (.Y(_0637_),
    .A(_0635_));
 sg13g2_nand3_1 _2641_ (.B(_0609_),
    .C(_0637_),
    .A(_0608_),
    .Y(_0638_));
 sg13g2_nand2_1 _2642_ (.Y(_0639_),
    .A(_0636_),
    .B(_0638_));
 sg13g2_nand2_1 _2643_ (.Y(_0640_),
    .A(_0620_),
    .B(_0587_));
 sg13g2_nand3_1 _2644_ (.B(_0619_),
    .C(_0602_),
    .A(_0618_),
    .Y(_0641_));
 sg13g2_nand2_1 _2645_ (.Y(_0642_),
    .A(_0640_),
    .B(_0641_));
 sg13g2_nor2_1 _2646_ (.A(_0639_),
    .B(_0642_),
    .Y(_0643_));
 sg13g2_nand3_1 _2647_ (.B(_0634_),
    .C(_0643_),
    .A(_0623_),
    .Y(_0644_));
 sg13g2_nor2_1 _2648_ (.A(_0637_),
    .B(_0614_),
    .Y(_0645_));
 sg13g2_inv_1 _2649_ (.Y(_0646_),
    .A(_0640_));
 sg13g2_a21oi_1 _2650_ (.A1(_0645_),
    .A2(_0641_),
    .Y(_0647_),
    .B1(_0646_));
 sg13g2_nor2_1 _2651_ (.A(_0647_),
    .B(_0622_),
    .Y(_0648_));
 sg13g2_inv_1 _2652_ (.Y(_0649_),
    .A(_0620_));
 sg13g2_nand2_1 _2653_ (.Y(_0650_),
    .A(_0649_),
    .B(_0598_));
 sg13g2_nor2_1 _2654_ (.A(_0598_),
    .B(_0649_),
    .Y(_0651_));
 sg13g2_a21oi_1 _2655_ (.A1(_0650_),
    .A2(_0615_),
    .Y(_0652_),
    .B1(_0651_));
 sg13g2_nor2b_1 _2656_ (.A(_0648_),
    .B_N(_0652_),
    .Y(_0653_));
 sg13g2_nand2_1 _2657_ (.Y(_0654_),
    .A(_0644_),
    .B(_0653_));
 sg13g2_nand2b_1 _2658_ (.Y(_0655_),
    .B(_0654_),
    .A_N(_0607_));
 sg13g2_inv_1 _2659_ (.Y(_0656_),
    .A(\dither_threshold[6] ));
 sg13g2_nand2b_1 _2660_ (.Y(_0657_),
    .B(_0656_),
    .A_N(_0655_));
 sg13g2_nand2_1 _2661_ (.Y(_0658_),
    .A(_0655_),
    .B(\dither_threshold[6] ));
 sg13g2_nand2_1 _2662_ (.Y(_0659_),
    .A(_0657_),
    .B(_0658_));
 sg13g2_nor2_1 _2663_ (.A(_0635_),
    .B(_0610_),
    .Y(_0660_));
 sg13g2_o21ai_1 _2664_ (.B1(_0636_),
    .Y(_0661_),
    .A1(_0631_),
    .A2(_0660_));
 sg13g2_nand2_1 _2665_ (.Y(_0662_),
    .A(_0610_),
    .B(_0519_));
 sg13g2_nand3_1 _2666_ (.B(_0609_),
    .C(_0612_),
    .A(_0608_),
    .Y(_0663_));
 sg13g2_nand2_1 _2667_ (.Y(_0664_),
    .A(_0662_),
    .B(_0663_));
 sg13g2_nor2_1 _2668_ (.A(_0664_),
    .B(_0642_),
    .Y(_0665_));
 sg13g2_a21oi_1 _2669_ (.A1(_0662_),
    .A2(_0640_),
    .Y(_0666_),
    .B1(_0611_));
 sg13g2_a21oi_1 _2670_ (.A1(_0661_),
    .A2(_0665_),
    .Y(_0667_),
    .B1(_0666_));
 sg13g2_nand2_1 _2671_ (.Y(_0668_),
    .A(_0631_),
    .B(_0629_));
 sg13g2_nor2_1 _2672_ (.A(_0639_),
    .B(_0668_),
    .Y(_0669_));
 sg13g2_nand3_1 _2673_ (.B(_0665_),
    .C(_0627_),
    .A(_0669_),
    .Y(_0670_));
 sg13g2_nand2_1 _2674_ (.Y(_0671_),
    .A(_0667_),
    .B(_0670_));
 sg13g2_inv_1 _2675_ (.Y(_0672_),
    .A(_0621_));
 sg13g2_nand2_1 _2676_ (.Y(_0673_),
    .A(_0671_),
    .B(_0672_));
 sg13g2_nand3_1 _2677_ (.B(_0670_),
    .C(_0621_),
    .A(_0667_),
    .Y(_0674_));
 sg13g2_nand3_1 _2678_ (.B(_0674_),
    .C(_1895_),
    .A(_0673_),
    .Y(_0675_));
 sg13g2_nand2_1 _2679_ (.Y(_0676_),
    .A(_0671_),
    .B(_0621_));
 sg13g2_nand3_1 _2680_ (.B(_0670_),
    .C(_0672_),
    .A(_0667_),
    .Y(_0677_));
 sg13g2_nand3_1 _2681_ (.B(_0677_),
    .C(_1894_),
    .A(_0676_),
    .Y(_0678_));
 sg13g2_nand2_1 _2682_ (.Y(_0679_),
    .A(_0675_),
    .B(_0678_));
 sg13g2_nor2_1 _2683_ (.A(_0659_),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nand2_1 _2684_ (.Y(_0681_),
    .A(_0634_),
    .B(_0643_));
 sg13g2_nand2_1 _2685_ (.Y(_0682_),
    .A(_0681_),
    .B(_0647_));
 sg13g2_nand2_1 _2686_ (.Y(_0683_),
    .A(_0682_),
    .B(_0616_));
 sg13g2_nand3_1 _2687_ (.B(_0664_),
    .C(_0647_),
    .A(_0681_),
    .Y(_0684_));
 sg13g2_nand2_1 _2688_ (.Y(_0685_),
    .A(_0683_),
    .B(_0684_));
 sg13g2_nand2_1 _2689_ (.Y(_0686_),
    .A(_0685_),
    .B(_1886_));
 sg13g2_nand3_1 _2690_ (.B(_0684_),
    .C(_1885_),
    .A(_0683_),
    .Y(_0687_));
 sg13g2_nand2_1 _2691_ (.Y(_0688_),
    .A(_0669_),
    .B(_0627_));
 sg13g2_inv_1 _2692_ (.Y(_0689_),
    .A(_0661_));
 sg13g2_nand2_1 _2693_ (.Y(_0690_),
    .A(_0688_),
    .B(_0689_));
 sg13g2_inv_1 _2694_ (.Y(_0691_),
    .A(_0642_));
 sg13g2_nand2_1 _2695_ (.Y(_0692_),
    .A(_0690_),
    .B(_0691_));
 sg13g2_nand3_1 _2696_ (.B(_0642_),
    .C(_0689_),
    .A(_0688_),
    .Y(_0693_));
 sg13g2_nand2_1 _2697_ (.Y(_0694_),
    .A(_0692_),
    .B(_0693_));
 sg13g2_nor2_1 _2698_ (.A(\dither_threshold[3] ),
    .B(_0694_),
    .Y(_0695_));
 sg13g2_nand3_1 _2699_ (.B(_0687_),
    .C(_0695_),
    .A(_0686_),
    .Y(_0696_));
 sg13g2_nand3_1 _2700_ (.B(_0684_),
    .C(_1857_),
    .A(_0683_),
    .Y(_0697_));
 sg13g2_nand2_1 _2701_ (.Y(_0698_),
    .A(_0696_),
    .B(_0697_));
 sg13g2_nand2_1 _2702_ (.Y(_0699_),
    .A(_0673_),
    .B(_0674_));
 sg13g2_nand3_1 _2703_ (.B(_0699_),
    .C(_1856_),
    .A(_0658_),
    .Y(_0700_));
 sg13g2_nand2_1 _2704_ (.Y(_0701_),
    .A(_0700_),
    .B(_0657_));
 sg13g2_a21oi_1 _2705_ (.A1(_0680_),
    .A2(_0698_),
    .Y(_0702_),
    .B1(_0701_));
 sg13g2_xor2_1 _2706_ (.B(_0668_),
    .A(_0627_),
    .X(_0703_));
 sg13g2_xnor2_1 _2707_ (.Y(_0704_),
    .A(_1870_),
    .B(_0703_));
 sg13g2_xnor2_1 _2708_ (.Y(_0705_),
    .A(_0639_),
    .B(_0633_));
 sg13g2_nand2b_1 _2709_ (.Y(_0706_),
    .B(_1874_),
    .A_N(_0705_));
 sg13g2_nand2_1 _2710_ (.Y(_0707_),
    .A(_0705_),
    .B(_1854_));
 sg13g2_nand2_1 _2711_ (.Y(_0708_),
    .A(_0706_),
    .B(_0707_));
 sg13g2_nor2_1 _2712_ (.A(_0704_),
    .B(_0708_),
    .Y(_0709_));
 sg13g2_xnor2_1 _2713_ (.Y(_0710_),
    .A(_0626_),
    .B(_0610_));
 sg13g2_nand2_1 _2714_ (.Y(_0711_),
    .A(_0710_),
    .B(_1849_));
 sg13g2_nand2_1 _2715_ (.Y(_0712_),
    .A(_0709_),
    .B(_0711_));
 sg13g2_nor2_1 _2716_ (.A(_1851_),
    .B(_0703_),
    .Y(_0713_));
 sg13g2_inv_1 _2717_ (.Y(_0714_),
    .A(_0706_));
 sg13g2_a21oi_1 _2718_ (.A1(_0707_),
    .A2(_0713_),
    .Y(_0715_),
    .B1(_0714_));
 sg13g2_nand2_1 _2719_ (.Y(_0716_),
    .A(_0712_),
    .B(_0715_));
 sg13g2_xnor2_1 _2720_ (.Y(_0717_),
    .A(_1878_),
    .B(_0694_));
 sg13g2_nand2_1 _2721_ (.Y(_0718_),
    .A(_0686_),
    .B(_0687_));
 sg13g2_nor2_1 _2722_ (.A(_0717_),
    .B(_0718_),
    .Y(_0719_));
 sg13g2_nand3_1 _2723_ (.B(_0716_),
    .C(_0719_),
    .A(_0680_),
    .Y(_0720_));
 sg13g2_nand2_1 _2724_ (.Y(_0721_),
    .A(_0702_),
    .B(_0720_));
 sg13g2_xnor2_1 _2725_ (.Y(_0722_),
    .A(_1850_),
    .B(_0710_));
 sg13g2_nand2_1 _2726_ (.Y(_0723_),
    .A(_0709_),
    .B(_0722_));
 sg13g2_nor2_1 _2727_ (.A(_0717_),
    .B(_0723_),
    .Y(_0724_));
 sg13g2_nand3b_1 _2728_ (.B(_0680_),
    .C(_0724_),
    .Y(_0725_),
    .A_N(_0718_));
 sg13g2_nand3_1 _2729_ (.B(_0614_),
    .C(_0725_),
    .A(_0721_),
    .Y(_0726_));
 sg13g2_nand2_1 _2730_ (.Y(_0727_),
    .A(_0726_),
    .B(_0649_));
 sg13g2_nand4_1 _2731_ (.B(_0620_),
    .C(_0614_),
    .A(_0721_),
    .Y(_0728_),
    .D(_0725_));
 sg13g2_nand2_1 _2732_ (.Y(net8),
    .A(_0727_),
    .B(_0728_));
 sg13g2_inv_1 _2733_ (.Y(_0729_),
    .A(_0039_));
 sg13g2_xnor2_1 _2734_ (.Y(_0730_),
    .A(_0729_),
    .B(_2179_));
 sg13g2_xnor2_1 _2735_ (.Y(_0731_),
    .A(net70),
    .B(_2039_));
 sg13g2_nand2_1 _2736_ (.Y(_0732_),
    .A(net58),
    .B(net65));
 sg13g2_xor2_1 _2737_ (.B(net53),
    .A(net59),
    .X(_0733_));
 sg13g2_inv_1 _2738_ (.Y(_0734_),
    .A(_0733_));
 sg13g2_nand2_1 _2739_ (.Y(_0735_),
    .A(net59),
    .B(net53));
 sg13g2_o21ai_1 _2740_ (.B1(_0735_),
    .Y(_0736_),
    .A1(_0732_),
    .A2(_0734_));
 sg13g2_xnor2_1 _2741_ (.Y(_0737_),
    .A(net57),
    .B(net66));
 sg13g2_xor2_1 _2742_ (.B(_2042_),
    .A(net61),
    .X(_0738_));
 sg13g2_inv_1 _2743_ (.Y(_0739_),
    .A(_0738_));
 sg13g2_nor2_1 _2744_ (.A(_0737_),
    .B(_0739_),
    .Y(_0740_));
 sg13g2_nand2_1 _2745_ (.Y(_0741_),
    .A(net61),
    .B(net54));
 sg13g2_nand2_1 _2746_ (.Y(_0742_),
    .A(net57),
    .B(net66));
 sg13g2_o21ai_1 _2747_ (.B1(_0742_),
    .Y(_0743_),
    .A1(_0741_),
    .A2(_0737_));
 sg13g2_a21oi_1 _2748_ (.A1(_0736_),
    .A2(_0740_),
    .Y(_0744_),
    .B1(_0743_));
 sg13g2_nand2_1 _2749_ (.Y(_0745_),
    .A(_1712_),
    .B(_2052_));
 sg13g2_xnor2_1 _2750_ (.Y(_0746_),
    .A(net71),
    .B(net64));
 sg13g2_nand2_1 _2751_ (.Y(_0747_),
    .A(net71),
    .B(net64));
 sg13g2_o21ai_1 _2752_ (.B1(_0747_),
    .Y(_0748_),
    .A1(_0745_),
    .A2(_0746_));
 sg13g2_buf_1 _2753_ (.A(_0748_),
    .X(_0749_));
 sg13g2_xor2_1 _2754_ (.B(net65),
    .A(net58),
    .X(_0750_));
 sg13g2_inv_1 _2755_ (.Y(_0751_),
    .A(_0750_));
 sg13g2_nor2_1 _2756_ (.A(_0751_),
    .B(_0734_),
    .Y(_0752_));
 sg13g2_nand3_1 _2757_ (.B(_0752_),
    .C(_0740_),
    .A(_0749_),
    .Y(_0753_));
 sg13g2_nand2_1 _2758_ (.Y(_0754_),
    .A(_0744_),
    .B(_0753_));
 sg13g2_xor2_1 _2759_ (.B(_2040_),
    .A(net72),
    .X(_0755_));
 sg13g2_nand2_1 _2760_ (.Y(_0756_),
    .A(_0754_),
    .B(_0755_));
 sg13g2_o21ai_1 _2761_ (.B1(_0756_),
    .Y(_0757_),
    .A1(_1732_),
    .A2(_2058_));
 sg13g2_xnor2_1 _2762_ (.Y(_0758_),
    .A(_0731_),
    .B(_0757_));
 sg13g2_xnor2_1 _2763_ (.Y(_0759_),
    .A(_0730_),
    .B(_0758_));
 sg13g2_xnor2_1 _2764_ (.Y(_0760_),
    .A(_2047_),
    .B(net20));
 sg13g2_inv_1 _2765_ (.Y(_0761_),
    .A(_0044_));
 sg13g2_xnor2_1 _2766_ (.Y(_0762_),
    .A(_0761_),
    .B(_2229_));
 sg13g2_inv_2 _2767_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_xnor2_1 _2768_ (.Y(_0764_),
    .A(_2052_),
    .B(net26));
 sg13g2_nor2b_1 _2769_ (.A(_0763_),
    .B_N(_0764_),
    .Y(_0765_));
 sg13g2_nor2b_2 _2770_ (.A(net35),
    .B_N(net63),
    .Y(_0766_));
 sg13g2_nand2_1 _2771_ (.Y(_0767_),
    .A(_0765_),
    .B(_0766_));
 sg13g2_nor2_1 _2772_ (.A(_0045_),
    .B(net26),
    .Y(_0768_));
 sg13g2_nor2_1 _2773_ (.A(_0044_),
    .B(_2229_),
    .Y(_0769_));
 sg13g2_a21oi_1 _2774_ (.A1(_0762_),
    .A2(_0768_),
    .Y(_0770_),
    .B1(_0769_));
 sg13g2_nand2_1 _2775_ (.Y(_0771_),
    .A(_0767_),
    .B(_0770_));
 sg13g2_xnor2_1 _2776_ (.Y(_0772_),
    .A(_2049_),
    .B(net22));
 sg13g2_inv_1 _2777_ (.Y(_0773_),
    .A(_0772_));
 sg13g2_nand2_1 _2778_ (.Y(_0774_),
    .A(_0771_),
    .B(_0773_));
 sg13g2_xnor2_1 _2779_ (.Y(_0775_),
    .A(_2112_),
    .B(net19));
 sg13g2_xnor2_1 _2780_ (.Y(_0776_),
    .A(_0164_),
    .B(_2152_));
 sg13g2_inv_1 _2781_ (.Y(_0777_),
    .A(_0776_));
 sg13g2_nand2b_1 _2782_ (.Y(_0778_),
    .B(_0777_),
    .A_N(_0775_));
 sg13g2_nor3_1 _2783_ (.A(_0760_),
    .B(_0774_),
    .C(_0778_),
    .Y(_0779_));
 sg13g2_inv_1 _2784_ (.Y(_0780_),
    .A(_0778_));
 sg13g2_inv_1 _2785_ (.Y(_0781_),
    .A(net22));
 sg13g2_inv_1 _2786_ (.Y(_0782_),
    .A(_0043_));
 sg13g2_nand2_1 _2787_ (.Y(_0783_),
    .A(_0781_),
    .B(_0782_));
 sg13g2_nor2_1 _2788_ (.A(_0042_),
    .B(net20),
    .Y(_0784_));
 sg13g2_inv_1 _2789_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_o21ai_1 _2790_ (.B1(_0785_),
    .Y(_0786_),
    .A1(_0783_),
    .A2(_0760_));
 sg13g2_inv_1 _2791_ (.Y(_0787_),
    .A(_2112_));
 sg13g2_inv_1 _2792_ (.Y(_0788_),
    .A(net19));
 sg13g2_nor2_1 _2793_ (.A(_0164_),
    .B(net18),
    .Y(_0789_));
 sg13g2_o21ai_1 _2794_ (.B1(_0789_),
    .Y(_0790_),
    .A1(_0787_),
    .A2(_0788_));
 sg13g2_o21ai_1 _2795_ (.B1(_0790_),
    .Y(_0791_),
    .A1(_2112_),
    .A2(net19));
 sg13g2_a21oi_1 _2796_ (.A1(_0780_),
    .A2(_0786_),
    .Y(_0792_),
    .B1(_0791_));
 sg13g2_nand2b_1 _2797_ (.Y(_0793_),
    .B(_0792_),
    .A_N(_0779_));
 sg13g2_nor2_1 _2798_ (.A(_0759_),
    .B(_0793_),
    .Y(_0794_));
 sg13g2_a21oi_1 _2799_ (.A1(_0793_),
    .A2(_0759_),
    .Y(_0795_),
    .B1(_0337_));
 sg13g2_nand2b_1 _2800_ (.Y(_0796_),
    .B(_0795_),
    .A_N(_0794_));
 sg13g2_a21oi_1 _2801_ (.A1(_0229_),
    .A2(_0244_),
    .Y(_0797_),
    .B1(_0416_));
 sg13g2_nor2_1 _2802_ (.A(_0308_),
    .B(_0797_),
    .Y(_0798_));
 sg13g2_nand2_1 _2803_ (.Y(_0799_),
    .A(_0796_),
    .B(_0798_));
 sg13g2_inv_1 _2804_ (.Y(_0800_),
    .A(_2179_));
 sg13g2_nor2_1 _2805_ (.A(_0023_),
    .B(_0539_),
    .Y(_0801_));
 sg13g2_a21oi_1 _2806_ (.A1(_0800_),
    .A2(_0801_),
    .Y(_0802_),
    .B1(_0256_));
 sg13g2_nand2_1 _2807_ (.Y(_0803_),
    .A(_0799_),
    .B(_0802_));
 sg13g2_inv_1 _2808_ (.Y(_0804_),
    .A(_0254_));
 sg13g2_xnor2_1 _2809_ (.Y(_0805_),
    .A(net28),
    .B(_2179_));
 sg13g2_a21oi_1 _2810_ (.A1(_0805_),
    .A2(net39),
    .Y(_0806_),
    .B1(net38));
 sg13g2_nand2_1 _2811_ (.Y(_0807_),
    .A(_0803_),
    .B(_0806_));
 sg13g2_a21oi_1 _2812_ (.A1(_0800_),
    .A2(_0320_),
    .Y(_0808_),
    .B1(net27));
 sg13g2_nand2_1 _2813_ (.Y(_0809_),
    .A(_0807_),
    .B(_0808_));
 sg13g2_nor2_1 _2814_ (.A(_2100_),
    .B(_0287_),
    .Y(_0810_));
 sg13g2_a21oi_1 _2815_ (.A1(_0809_),
    .A2(_0810_),
    .Y(_0811_),
    .B1(_2101_));
 sg13g2_buf_2 _2816_ (.A(_0811_),
    .X(_0812_));
 sg13g2_nand2_1 _2817_ (.Y(_0813_),
    .A(_0812_),
    .B(net24));
 sg13g2_buf_2 _2818_ (.A(_0813_),
    .X(_0814_));
 sg13g2_inv_1 _2819_ (.Y(_0815_),
    .A(_0814_));
 sg13g2_nor2_1 _2820_ (.A(_0563_),
    .B(_0812_),
    .Y(_0816_));
 sg13g2_a21o_1 _2821_ (.A2(_0752_),
    .A1(_0749_),
    .B1(_0736_),
    .X(_0817_));
 sg13g2_nand2_1 _2822_ (.Y(_0818_),
    .A(_0817_),
    .B(_0738_));
 sg13g2_nand2_1 _2823_ (.Y(_0819_),
    .A(_0818_),
    .B(_0741_));
 sg13g2_xnor2_1 _2824_ (.Y(_0820_),
    .A(_0737_),
    .B(_0819_));
 sg13g2_nor3_1 _2825_ (.A(_0772_),
    .B(_0760_),
    .C(_0770_),
    .Y(_0821_));
 sg13g2_nor2_1 _2826_ (.A(_0821_),
    .B(_0786_),
    .Y(_0822_));
 sg13g2_inv_1 _2827_ (.Y(_0823_),
    .A(_0760_));
 sg13g2_nand4_1 _2828_ (.B(_0773_),
    .C(_0765_),
    .A(_0823_),
    .Y(_0824_),
    .D(_0766_));
 sg13g2_nand2_1 _2829_ (.Y(_0825_),
    .A(_0822_),
    .B(_0824_));
 sg13g2_nand2_1 _2830_ (.Y(_0826_),
    .A(_0825_),
    .B(_0777_));
 sg13g2_nand3_1 _2831_ (.B(_0776_),
    .C(_0824_),
    .A(_0822_),
    .Y(_0827_));
 sg13g2_nand3b_1 _2832_ (.B(_0826_),
    .C(_0827_),
    .Y(_0828_),
    .A_N(_0820_));
 sg13g2_nand2_1 _2833_ (.Y(_0829_),
    .A(_0826_),
    .B(_0827_));
 sg13g2_nand2_1 _2834_ (.Y(_0830_),
    .A(_0829_),
    .B(_0820_));
 sg13g2_nand3_1 _2835_ (.B(_0830_),
    .C(net40),
    .A(_0828_),
    .Y(_0831_));
 sg13g2_inv_1 _2836_ (.Y(_0832_),
    .A(_0315_));
 sg13g2_nand2_1 _2837_ (.Y(_0833_),
    .A(_0229_),
    .B(_0539_));
 sg13g2_buf_2 _2838_ (.A(_0833_),
    .X(_0834_));
 sg13g2_o21ai_1 _2839_ (.B1(_0466_),
    .Y(_0835_),
    .A1(_0832_),
    .A2(_0834_));
 sg13g2_nand2_1 _2840_ (.Y(_0836_),
    .A(_0831_),
    .B(_0835_));
 sg13g2_inv_1 _2841_ (.Y(_0837_),
    .A(_0168_));
 sg13g2_nor2_1 _2842_ (.A(_0051_),
    .B(net45),
    .Y(_0838_));
 sg13g2_a21oi_1 _2843_ (.A1(_0837_),
    .A2(_0838_),
    .Y(_0839_),
    .B1(net31));
 sg13g2_nand2_1 _2844_ (.Y(_0840_),
    .A(_0836_),
    .B(_0839_));
 sg13g2_xnor2_1 _2845_ (.Y(_0841_),
    .A(net28),
    .B(_0168_));
 sg13g2_a21oi_1 _2846_ (.A1(_0841_),
    .A2(net31),
    .Y(_0842_),
    .B1(net36));
 sg13g2_nand2_1 _2847_ (.Y(_0843_),
    .A(_0840_),
    .B(_0842_));
 sg13g2_a21oi_1 _2848_ (.A1(_0837_),
    .A2(_0483_),
    .Y(_0844_),
    .B1(net25));
 sg13g2_nand2_1 _2849_ (.Y(_0845_),
    .A(_0843_),
    .B(_0844_));
 sg13g2_a21oi_1 _2850_ (.A1(_0845_),
    .A2(net17),
    .Y(_0846_),
    .B1(net49));
 sg13g2_nor2b_1 _2851_ (.A(_0846_),
    .B_N(_0335_),
    .Y(_0847_));
 sg13g2_nand2_1 _2852_ (.Y(_0848_),
    .A(_0847_),
    .B(_0437_));
 sg13g2_xnor2_1 _2853_ (.Y(_0849_),
    .A(_0755_),
    .B(_0754_));
 sg13g2_xor2_1 _2854_ (.B(_0775_),
    .A(_0849_),
    .X(_0850_));
 sg13g2_nor2_1 _2855_ (.A(_0760_),
    .B(_0776_),
    .Y(_0851_));
 sg13g2_inv_1 _2856_ (.Y(_0852_),
    .A(_0769_));
 sg13g2_o21ai_1 _2857_ (.B1(_0783_),
    .Y(_0853_),
    .A1(_0852_),
    .A2(_0772_));
 sg13g2_nand2_1 _2858_ (.Y(_0854_),
    .A(net18),
    .B(_0164_));
 sg13g2_a21oi_1 _2859_ (.A1(_0854_),
    .A2(_0784_),
    .Y(_0855_),
    .B1(_0789_));
 sg13g2_inv_1 _2860_ (.Y(_0856_),
    .A(_0855_));
 sg13g2_a21oi_1 _2861_ (.A1(_0851_),
    .A2(_0853_),
    .Y(_0857_),
    .B1(_0856_));
 sg13g2_a21o_1 _2862_ (.A2(_0766_),
    .A1(_0764_),
    .B1(_0768_),
    .X(_0858_));
 sg13g2_nor2_1 _2863_ (.A(_0763_),
    .B(_0772_),
    .Y(_0859_));
 sg13g2_nand3_1 _2864_ (.B(_0858_),
    .C(_0859_),
    .A(_0851_),
    .Y(_0860_));
 sg13g2_nand2_1 _2865_ (.Y(_0861_),
    .A(_0857_),
    .B(_0860_));
 sg13g2_nand2b_1 _2866_ (.Y(_0862_),
    .B(_0861_),
    .A_N(_0850_));
 sg13g2_nand3_1 _2867_ (.B(_0860_),
    .C(_0850_),
    .A(_0857_),
    .Y(_0863_));
 sg13g2_nand3_1 _2868_ (.B(_0863_),
    .C(net42),
    .A(_0862_),
    .Y(_0864_));
 sg13g2_inv_1 _2869_ (.Y(_0865_),
    .A(_0426_));
 sg13g2_o21ai_1 _2870_ (.B1(_0303_),
    .Y(_0866_),
    .A1(_0865_),
    .A2(_0834_));
 sg13g2_nand2_1 _2871_ (.Y(_0867_),
    .A(_0864_),
    .B(_0866_));
 sg13g2_nor2_1 _2872_ (.A(_0048_),
    .B(_0539_),
    .Y(_0868_));
 sg13g2_a21oi_1 _2873_ (.A1(_0788_),
    .A2(_0868_),
    .Y(_0869_),
    .B1(net34));
 sg13g2_nand2_1 _2874_ (.Y(_0870_),
    .A(_0867_),
    .B(_0869_));
 sg13g2_xnor2_1 _2875_ (.Y(_0871_),
    .A(_0804_),
    .B(net19));
 sg13g2_a21oi_1 _2876_ (.A1(_0871_),
    .A2(net34),
    .Y(_0872_),
    .B1(net41));
 sg13g2_nand2_1 _2877_ (.Y(_0873_),
    .A(_0870_),
    .B(_0872_));
 sg13g2_a21oi_1 _2878_ (.A1(_0788_),
    .A2(_0320_),
    .Y(_0874_),
    .B1(net27));
 sg13g2_nand2_1 _2879_ (.Y(_0875_),
    .A(_0873_),
    .B(_0874_));
 sg13g2_nand2_1 _2880_ (.Y(_0876_),
    .A(_0875_),
    .B(_0432_));
 sg13g2_a21oi_2 _2881_ (.B1(_0332_),
    .Y(_0877_),
    .A2(_0435_),
    .A1(_0876_));
 sg13g2_a21oi_1 _2882_ (.A1(_0877_),
    .A2(net47),
    .Y(_0878_),
    .B1(_0511_));
 sg13g2_xor2_1 _2883_ (.B(_0746_),
    .A(_0745_),
    .X(_0879_));
 sg13g2_xor2_1 _2884_ (.B(_0764_),
    .A(_0766_),
    .X(_0880_));
 sg13g2_xor2_1 _2885_ (.B(_0880_),
    .A(_0879_),
    .X(_0881_));
 sg13g2_inv_1 _2886_ (.Y(_0882_),
    .A(_0490_));
 sg13g2_o21ai_1 _2887_ (.B1(_0882_),
    .Y(_0883_),
    .A1(_0553_),
    .A2(_0834_));
 sg13g2_o21ai_1 _2888_ (.B1(_0883_),
    .Y(_0884_),
    .A1(net37),
    .A2(_0881_));
 sg13g2_inv_1 _2889_ (.Y(_0885_),
    .A(net26));
 sg13g2_nor2_1 _2890_ (.A(_0038_),
    .B(net45),
    .Y(_0886_));
 sg13g2_a21oi_1 _2891_ (.A1(_0885_),
    .A2(_0886_),
    .Y(_0887_),
    .B1(net31));
 sg13g2_nand2_1 _2892_ (.Y(_0888_),
    .A(_0884_),
    .B(_0887_));
 sg13g2_a21oi_1 _2893_ (.A1(net23),
    .A2(net26),
    .Y(_0889_),
    .B1(net30));
 sg13g2_o21ai_1 _2894_ (.B1(_0889_),
    .Y(_0890_),
    .A1(net26),
    .A2(net23));
 sg13g2_nand3_1 _2895_ (.B(net33),
    .C(_0890_),
    .A(_0888_),
    .Y(_0891_));
 sg13g2_o21ai_1 _2896_ (.B1(_0891_),
    .Y(_0892_),
    .A1(net26),
    .A2(net33));
 sg13g2_o21ai_1 _2897_ (.B1(_0538_),
    .Y(_0893_),
    .A1(net25),
    .A2(_0892_));
 sg13g2_nand3_1 _2898_ (.B(_0878_),
    .C(_0893_),
    .A(_0848_),
    .Y(_0894_));
 sg13g2_nor2_1 _2899_ (.A(_0816_),
    .B(_0894_),
    .Y(_0895_));
 sg13g2_nor2_1 _2900_ (.A(_0815_),
    .B(_0895_),
    .Y(_0896_));
 sg13g2_nand2_1 _2901_ (.Y(_0897_),
    .A(_0876_),
    .B(_0435_));
 sg13g2_nand2_1 _2902_ (.Y(_0898_),
    .A(_0897_),
    .B(_0440_));
 sg13g2_xnor2_1 _2903_ (.Y(_0899_),
    .A(_0751_),
    .B(_0749_));
 sg13g2_xnor2_1 _2904_ (.Y(_0900_),
    .A(_0762_),
    .B(_0858_));
 sg13g2_xnor2_1 _2905_ (.Y(_0901_),
    .A(_0899_),
    .B(_0900_));
 sg13g2_o21ai_1 _2906_ (.B1(_0546_),
    .Y(_0902_),
    .A1(_0359_),
    .A2(_0834_));
 sg13g2_o21ai_1 _2907_ (.B1(_0902_),
    .Y(_0903_),
    .A1(net37),
    .A2(_0901_));
 sg13g2_nor2_1 _2908_ (.A(_0037_),
    .B(net45),
    .Y(_0904_));
 sg13g2_a21oi_1 _2909_ (.A1(_0150_),
    .A2(_0904_),
    .Y(_0905_),
    .B1(net39));
 sg13g2_nand2_1 _2910_ (.Y(_0906_),
    .A(_0903_),
    .B(_0905_));
 sg13g2_a21oi_1 _2911_ (.A1(net28),
    .A2(_0150_),
    .Y(_0907_),
    .B1(_0360_));
 sg13g2_o21ai_1 _2912_ (.B1(_0907_),
    .Y(_0908_),
    .A1(_0150_),
    .A2(net28));
 sg13g2_nand3_1 _2913_ (.B(net33),
    .C(_0908_),
    .A(_0906_),
    .Y(_0909_));
 sg13g2_a21oi_1 _2914_ (.A1(_0150_),
    .A2(_0364_),
    .Y(_0910_),
    .B1(_0365_));
 sg13g2_a21oi_1 _2915_ (.A1(_0909_),
    .A2(_0910_),
    .Y(_0911_),
    .B1(_0287_));
 sg13g2_nand2b_1 _2916_ (.Y(_0912_),
    .B(net43),
    .A_N(_0911_));
 sg13g2_a21oi_1 _2917_ (.A1(_0912_),
    .A2(_0378_),
    .Y(_0913_),
    .B1(_0384_));
 sg13g2_nand2_1 _2918_ (.Y(_0914_),
    .A(_0898_),
    .B(_0913_));
 sg13g2_a21oi_1 _2919_ (.A1(_0445_),
    .A2(_0877_),
    .Y(_0915_),
    .B1(_0914_));
 sg13g2_nand2_1 _2920_ (.Y(_0916_),
    .A(_0847_),
    .B(net46));
 sg13g2_inv_4 _2921_ (.A(_0812_),
    .Y(_0917_));
 sg13g2_nand2_1 _2922_ (.Y(_0918_),
    .A(_0917_),
    .B(net47));
 sg13g2_nand3_1 _2923_ (.B(_0916_),
    .C(_0918_),
    .A(_0915_),
    .Y(_0919_));
 sg13g2_buf_1 _2924_ (.A(_0919_),
    .X(_0920_));
 sg13g2_nand2_1 _2925_ (.Y(_0921_),
    .A(_0896_),
    .B(_0920_));
 sg13g2_nor2b_1 _2926_ (.A(_0834_),
    .B_N(_0577_),
    .Y(_0922_));
 sg13g2_nand2_1 _2927_ (.Y(_0923_),
    .A(_0749_),
    .B(_0750_));
 sg13g2_nand2_1 _2928_ (.Y(_0924_),
    .A(_0923_),
    .B(_0732_));
 sg13g2_xnor2_1 _2929_ (.Y(_0925_),
    .A(_0734_),
    .B(_0924_));
 sg13g2_xnor2_1 _2930_ (.Y(_0926_),
    .A(_0772_),
    .B(_0771_));
 sg13g2_xnor2_1 _2931_ (.Y(_0927_),
    .A(_0925_),
    .B(_0926_));
 sg13g2_nand2_1 _2932_ (.Y(_0928_),
    .A(_0927_),
    .B(net40));
 sg13g2_o21ai_1 _2933_ (.B1(_0928_),
    .Y(_0929_),
    .A1(_0345_),
    .A2(_0922_));
 sg13g2_nor2_1 _2934_ (.A(_0024_),
    .B(net45),
    .Y(_0930_));
 sg13g2_a21oi_1 _2935_ (.A1(_0781_),
    .A2(_0930_),
    .Y(_0931_),
    .B1(_0493_));
 sg13g2_nand2_1 _2936_ (.Y(_0932_),
    .A(_0929_),
    .B(_0931_));
 sg13g2_a21oi_1 _2937_ (.A1(net23),
    .A2(net22),
    .Y(_0933_),
    .B1(_0541_));
 sg13g2_o21ai_1 _2938_ (.B1(_0933_),
    .Y(_0934_),
    .A1(net22),
    .A2(net23));
 sg13g2_nand3_1 _2939_ (.B(_0351_),
    .C(_0934_),
    .A(_0932_),
    .Y(_0935_));
 sg13g2_a21oi_1 _2940_ (.A1(_0781_),
    .A2(net32),
    .Y(_0936_),
    .B1(net25));
 sg13g2_a21oi_1 _2941_ (.A1(_0935_),
    .A2(_0936_),
    .Y(_0937_),
    .B1(_0287_));
 sg13g2_nand2b_1 _2942_ (.Y(_0938_),
    .B(net43),
    .A_N(_0937_));
 sg13g2_a21oi_1 _2943_ (.A1(_0938_),
    .A2(_0585_),
    .Y(_0939_),
    .B1(net24));
 sg13g2_nand2b_1 _2944_ (.Y(_0940_),
    .B(_0917_),
    .A_N(_0567_));
 sg13g2_nand2_1 _2945_ (.Y(_0941_),
    .A(_0877_),
    .B(net46));
 sg13g2_nand3_1 _2946_ (.B(_0940_),
    .C(_0941_),
    .A(_0939_),
    .Y(_0942_));
 sg13g2_nand2_1 _2947_ (.Y(_0943_),
    .A(_0942_),
    .B(_0814_));
 sg13g2_nand2_1 _2948_ (.Y(_0944_),
    .A(_0877_),
    .B(_0445_));
 sg13g2_xnor2_1 _2949_ (.Y(_0945_),
    .A(_0739_),
    .B(_0817_));
 sg13g2_nand2_1 _2950_ (.Y(_0946_),
    .A(_0774_),
    .B(_0783_));
 sg13g2_nand2_1 _2951_ (.Y(_0947_),
    .A(_0946_),
    .B(_0823_));
 sg13g2_nand3_1 _2952_ (.B(_0760_),
    .C(_0783_),
    .A(_0774_),
    .Y(_0948_));
 sg13g2_nand2_1 _2953_ (.Y(_0949_),
    .A(_0947_),
    .B(_0948_));
 sg13g2_xnor2_1 _2954_ (.Y(_0950_),
    .A(_0945_),
    .B(_0949_));
 sg13g2_inv_1 _2955_ (.Y(_0951_),
    .A(_0474_));
 sg13g2_o21ai_1 _2956_ (.B1(_0574_),
    .Y(_0952_),
    .A1(_0951_),
    .A2(_0834_));
 sg13g2_o21ai_1 _2957_ (.B1(_0952_),
    .Y(_0953_),
    .A1(net37),
    .A2(_0950_));
 sg13g2_inv_1 _2958_ (.Y(_0954_),
    .A(net20));
 sg13g2_nor2_1 _2959_ (.A(_0053_),
    .B(_0540_),
    .Y(_0955_));
 sg13g2_a21oi_1 _2960_ (.A1(_0954_),
    .A2(_0955_),
    .Y(_0956_),
    .B1(_0317_));
 sg13g2_nand2_1 _2961_ (.Y(_0957_),
    .A(_0953_),
    .B(_0956_));
 sg13g2_xor2_1 _2962_ (.B(net29),
    .A(_2133_),
    .X(_0958_));
 sg13g2_a21oi_1 _2963_ (.A1(_0958_),
    .A2(net39),
    .Y(_0959_),
    .B1(net38));
 sg13g2_nand2_1 _2964_ (.Y(_0960_),
    .A(_0957_),
    .B(_0959_));
 sg13g2_a21oi_1 _2965_ (.A1(_0954_),
    .A2(_0364_),
    .Y(_0961_),
    .B1(_0365_));
 sg13g2_nand2_1 _2966_ (.Y(_0962_),
    .A(_0960_),
    .B(_0961_));
 sg13g2_nand2_1 _2967_ (.Y(_0963_),
    .A(_0962_),
    .B(_0432_));
 sg13g2_nand2_1 _2968_ (.Y(_0964_),
    .A(_0963_),
    .B(_0481_));
 sg13g2_nand2_1 _2969_ (.Y(_0965_),
    .A(_0964_),
    .B(_0513_));
 sg13g2_nand3_1 _2970_ (.B(_0965_),
    .C(_0501_),
    .A(_0944_),
    .Y(_0966_));
 sg13g2_nand3_1 _2971_ (.B(_0501_),
    .C(_0812_),
    .A(_0966_),
    .Y(_0967_));
 sg13g2_a21oi_1 _2972_ (.A1(_0921_),
    .A2(_0943_),
    .Y(_0968_),
    .B1(_0967_));
 sg13g2_nand2_1 _2973_ (.Y(_0969_),
    .A(_0897_),
    .B(_0524_));
 sg13g2_nand4_1 _2974_ (.B(_0944_),
    .C(_0941_),
    .A(_0878_),
    .Y(_0970_),
    .D(_0969_));
 sg13g2_nand2_1 _2975_ (.Y(_0971_),
    .A(_0970_),
    .B(_0814_));
 sg13g2_a21oi_1 _2976_ (.A1(_0847_),
    .A2(_2110_),
    .Y(_0972_),
    .B1(net24));
 sg13g2_a22oi_1 _2977_ (.Y(_0973_),
    .B1(_0440_),
    .B2(_0964_),
    .A2(_0456_),
    .A1(_0897_));
 sg13g2_nand2_1 _2978_ (.Y(_0974_),
    .A(_0972_),
    .B(_0973_));
 sg13g2_xor2_1 _2979_ (.B(net63),
    .A(net60),
    .X(_0975_));
 sg13g2_xnor2_1 _2980_ (.Y(_0976_),
    .A(_2053_),
    .B(_0975_));
 sg13g2_o21ai_1 _2981_ (.B1(net40),
    .Y(_0977_),
    .A1(net35),
    .A2(_0976_));
 sg13g2_a21oi_1 _2982_ (.A1(net35),
    .A2(_0976_),
    .Y(_0978_),
    .B1(_0977_));
 sg13g2_nor3_1 _2983_ (.A(_0251_),
    .B(_0834_),
    .C(_0978_),
    .Y(_0979_));
 sg13g2_a21oi_1 _2984_ (.A1(_0492_),
    .A2(_0228_),
    .Y(_0980_),
    .B1(net40));
 sg13g2_nor2_1 _2985_ (.A(_0980_),
    .B(_0978_),
    .Y(_0981_));
 sg13g2_nor2_1 _2986_ (.A(net31),
    .B(_0981_),
    .Y(_0982_));
 sg13g2_inv_1 _2987_ (.Y(_0983_),
    .A(net35));
 sg13g2_nand3_1 _2988_ (.B(net51),
    .C(_1905_),
    .A(_0983_),
    .Y(_0984_));
 sg13g2_nand3b_1 _2989_ (.B(_0982_),
    .C(_0984_),
    .Y(_0985_),
    .A_N(_0979_));
 sg13g2_a21oi_1 _2990_ (.A1(net28),
    .A2(_0983_),
    .Y(_0986_),
    .B1(net30));
 sg13g2_o21ai_1 _2991_ (.B1(_0986_),
    .Y(_0987_),
    .A1(_0983_),
    .A2(net28));
 sg13g2_nand3_1 _2992_ (.B(_0987_),
    .C(net33),
    .A(_0985_),
    .Y(_0988_));
 sg13g2_nand2_1 _2993_ (.Y(_0989_),
    .A(_0983_),
    .B(net32));
 sg13g2_nand3_1 _2994_ (.B(_0262_),
    .C(_0989_),
    .A(_0988_),
    .Y(_0990_));
 sg13g2_nor2b_1 _2995_ (.A(_0500_),
    .B_N(_0990_),
    .Y(_0991_));
 sg13g2_nor2_1 _2996_ (.A(_0449_),
    .B(_0812_),
    .Y(_0992_));
 sg13g2_nand2_1 _2997_ (.Y(_0993_),
    .A(_0941_),
    .B(_0944_));
 sg13g2_nor3_1 _2998_ (.A(_0991_),
    .B(_0992_),
    .C(_0993_),
    .Y(_0994_));
 sg13g2_nor2b_1 _2999_ (.A(_0974_),
    .B_N(_0994_),
    .Y(_0995_));
 sg13g2_nor2_1 _3000_ (.A(_0533_),
    .B(_0812_),
    .Y(_0996_));
 sg13g2_nand2_1 _3001_ (.Y(_0997_),
    .A(_0966_),
    .B(_0814_));
 sg13g2_nand2b_1 _3002_ (.Y(_0998_),
    .B(_0997_),
    .A_N(_0996_));
 sg13g2_nand2_1 _3003_ (.Y(_0999_),
    .A(_0998_),
    .B(_0920_));
 sg13g2_nor2_1 _3004_ (.A(_0995_),
    .B(_0999_),
    .Y(_1000_));
 sg13g2_nor2_1 _3005_ (.A(_0971_),
    .B(_1000_),
    .Y(_1001_));
 sg13g2_nand2_1 _3006_ (.Y(_1002_),
    .A(_0375_),
    .B(_0533_));
 sg13g2_o21ai_1 _3007_ (.B1(_0847_),
    .Y(_1003_),
    .A1(_0437_),
    .A2(_1002_));
 sg13g2_nand2_1 _3008_ (.Y(_1004_),
    .A(_0972_),
    .B(_1003_));
 sg13g2_nand2_1 _3009_ (.Y(_1005_),
    .A(_1004_),
    .B(_0814_));
 sg13g2_nand2_1 _3010_ (.Y(_1006_),
    .A(_0917_),
    .B(_0445_));
 sg13g2_nand2_1 _3011_ (.Y(_1007_),
    .A(_1005_),
    .B(_1006_));
 sg13g2_nor2b_1 _3012_ (.A(_0895_),
    .B_N(_0942_),
    .Y(_1008_));
 sg13g2_a21oi_1 _3013_ (.A1(_1007_),
    .A2(_1008_),
    .Y(_1009_),
    .B1(_0812_));
 sg13g2_nor2_1 _3014_ (.A(_1001_),
    .B(_1009_),
    .Y(_1010_));
 sg13g2_nor2_1 _3015_ (.A(_0968_),
    .B(_1010_),
    .Y(_1011_));
 sg13g2_nand3_1 _3016_ (.B(_0814_),
    .C(_0942_),
    .A(_0920_),
    .Y(_1012_));
 sg13g2_inv_2 _3017_ (.Y(_1013_),
    .A(_0998_));
 sg13g2_nand2_1 _3018_ (.Y(_1014_),
    .A(_1012_),
    .B(_1013_));
 sg13g2_nand2b_1 _3019_ (.Y(_1015_),
    .B(_1014_),
    .A_N(_0970_));
 sg13g2_nand2_1 _3020_ (.Y(_1016_),
    .A(_1015_),
    .B(_0917_));
 sg13g2_nand2_1 _3021_ (.Y(_1017_),
    .A(_1016_),
    .B(_1007_));
 sg13g2_nand3_1 _3022_ (.B(_1017_),
    .C(_0971_),
    .A(_1011_),
    .Y(_1018_));
 sg13g2_buf_1 _3023_ (.A(_1018_),
    .X(_1019_));
 sg13g2_nand2_1 _3024_ (.Y(_1020_),
    .A(_1019_),
    .B(_0917_));
 sg13g2_nand2_1 _3025_ (.Y(_1021_),
    .A(_1020_),
    .B(_0896_));
 sg13g2_inv_1 _3026_ (.Y(_1022_),
    .A(_0896_));
 sg13g2_nand3_1 _3027_ (.B(_0917_),
    .C(_1022_),
    .A(_1019_),
    .Y(_1023_));
 sg13g2_nand2_1 _3028_ (.Y(_1024_),
    .A(_1021_),
    .B(_1023_));
 sg13g2_nand2_1 _3029_ (.Y(_1025_),
    .A(_1011_),
    .B(_1017_));
 sg13g2_inv_1 _3030_ (.Y(_1026_),
    .A(_0971_));
 sg13g2_nand2_1 _3031_ (.Y(_1027_),
    .A(_1025_),
    .B(_1026_));
 sg13g2_nand2_1 _3032_ (.Y(_1028_),
    .A(_0920_),
    .B(_0814_));
 sg13g2_inv_1 _3033_ (.Y(_1029_),
    .A(_1028_));
 sg13g2_nand3_1 _3034_ (.B(_1019_),
    .C(_1029_),
    .A(_1027_),
    .Y(_1030_));
 sg13g2_nand2_1 _3035_ (.Y(_1031_),
    .A(_1025_),
    .B(_0971_));
 sg13g2_nand3_1 _3036_ (.B(_1017_),
    .C(_1026_),
    .A(_1011_),
    .Y(_1032_));
 sg13g2_nand3_1 _3037_ (.B(_1032_),
    .C(_1028_),
    .A(_1031_),
    .Y(_1033_));
 sg13g2_nand2_1 _3038_ (.Y(_1034_),
    .A(_1030_),
    .B(_1033_));
 sg13g2_nor2_1 _3039_ (.A(_1024_),
    .B(_1034_),
    .Y(_1035_));
 sg13g2_nor2_1 _3040_ (.A(_0815_),
    .B(_0995_),
    .Y(_1036_));
 sg13g2_inv_1 _3041_ (.Y(_1037_),
    .A(_1036_));
 sg13g2_nand3_1 _3042_ (.B(_1032_),
    .C(_1037_),
    .A(_1031_),
    .Y(_1038_));
 sg13g2_buf_1 _3043_ (.A(_1038_),
    .X(_1039_));
 sg13g2_nand2_1 _3044_ (.Y(_1040_),
    .A(_1035_),
    .B(_1039_));
 sg13g2_inv_1 _3045_ (.Y(_1041_),
    .A(_1021_));
 sg13g2_nand2_1 _3046_ (.Y(_1042_),
    .A(_1027_),
    .B(_1019_));
 sg13g2_buf_8 _3047_ (.A(_1042_),
    .X(_1043_));
 sg13g2_nor2_1 _3048_ (.A(_1028_),
    .B(_1043_),
    .Y(_1044_));
 sg13g2_a21oi_1 _3049_ (.A1(_1041_),
    .A2(_1033_),
    .Y(_1045_),
    .B1(_1044_));
 sg13g2_nand2_1 _3050_ (.Y(_1046_),
    .A(_1040_),
    .B(_1045_));
 sg13g2_inv_1 _3051_ (.Y(_1047_),
    .A(_0943_));
 sg13g2_nand2_1 _3052_ (.Y(_1048_),
    .A(_1020_),
    .B(_1047_));
 sg13g2_nand3_1 _3053_ (.B(_0917_),
    .C(_0943_),
    .A(_1019_),
    .Y(_1049_));
 sg13g2_nand2_1 _3054_ (.Y(_1050_),
    .A(_1048_),
    .B(_1049_));
 sg13g2_inv_1 _3055_ (.Y(_1051_),
    .A(_1050_));
 sg13g2_nand2_1 _3056_ (.Y(_1052_),
    .A(_1046_),
    .B(_1051_));
 sg13g2_nand3_1 _3057_ (.B(_1045_),
    .C(_1050_),
    .A(_1040_),
    .Y(_1053_));
 sg13g2_nand2_1 _3058_ (.Y(_1054_),
    .A(_1052_),
    .B(_1053_));
 sg13g2_xnor2_1 _3059_ (.Y(_1055_),
    .A(_1878_),
    .B(_1054_));
 sg13g2_a21oi_1 _3060_ (.A1(_1039_),
    .A2(_1023_),
    .Y(_1056_),
    .B1(_1041_));
 sg13g2_inv_1 _3061_ (.Y(_1057_),
    .A(_1056_));
 sg13g2_nor2_1 _3062_ (.A(_1050_),
    .B(_1034_),
    .Y(_1058_));
 sg13g2_nand2_1 _3063_ (.Y(_1059_),
    .A(_1057_),
    .B(_1058_));
 sg13g2_inv_1 _3064_ (.Y(_1060_),
    .A(_1048_));
 sg13g2_o21ai_1 _3065_ (.B1(_1049_),
    .Y(_1061_),
    .A1(_1044_),
    .A2(_1060_));
 sg13g2_nand2_1 _3066_ (.Y(_1062_),
    .A(_1059_),
    .B(_1061_));
 sg13g2_nor2_1 _3067_ (.A(_1013_),
    .B(_1043_),
    .Y(_1063_));
 sg13g2_nand2_1 _3068_ (.Y(_1064_),
    .A(_1043_),
    .B(_1013_));
 sg13g2_nor2b_1 _3069_ (.A(_1063_),
    .B_N(_1064_),
    .Y(_1065_));
 sg13g2_nand2_1 _3070_ (.Y(_1066_),
    .A(_1062_),
    .B(_1065_));
 sg13g2_nand2b_1 _3071_ (.Y(_1067_),
    .B(_1064_),
    .A_N(_1063_));
 sg13g2_nand3_1 _3072_ (.B(_1061_),
    .C(_1067_),
    .A(_1059_),
    .Y(_1068_));
 sg13g2_buf_1 _3073_ (.A(_1068_),
    .X(_1069_));
 sg13g2_nand2_1 _3074_ (.Y(_1070_),
    .A(_1066_),
    .B(_1069_));
 sg13g2_nand2_1 _3075_ (.Y(_1071_),
    .A(_1070_),
    .B(_1886_));
 sg13g2_nand3_1 _3076_ (.B(_1069_),
    .C(_1885_),
    .A(_1066_),
    .Y(_1072_));
 sg13g2_nand2_1 _3077_ (.Y(_1073_),
    .A(_1071_),
    .B(_1072_));
 sg13g2_nor2_1 _3078_ (.A(_1055_),
    .B(_1073_),
    .Y(_1074_));
 sg13g2_xor2_1 _3079_ (.B(_1056_),
    .A(_1034_),
    .X(_1075_));
 sg13g2_nor2_1 _3080_ (.A(_1874_),
    .B(_1075_),
    .Y(_1076_));
 sg13g2_inv_1 _3081_ (.Y(_1077_),
    .A(_1039_));
 sg13g2_xnor2_1 _3082_ (.Y(_1078_),
    .A(_1077_),
    .B(_1024_));
 sg13g2_xnor2_1 _3083_ (.Y(_1079_),
    .A(_1870_),
    .B(_1078_));
 sg13g2_nor2_1 _3084_ (.A(_1037_),
    .B(_1043_),
    .Y(_1080_));
 sg13g2_o21ai_1 _3085_ (.B1(_1850_),
    .Y(_1081_),
    .A1(_1080_),
    .A2(_1077_));
 sg13g2_nor2b_1 _3086_ (.A(_1079_),
    .B_N(_1081_),
    .Y(_1082_));
 sg13g2_nand2_1 _3087_ (.Y(_1083_),
    .A(_1075_),
    .B(_1874_));
 sg13g2_nand3b_1 _3088_ (.B(_1082_),
    .C(_1083_),
    .Y(_1084_),
    .A_N(_1076_));
 sg13g2_nor2b_1 _3089_ (.A(_1852_),
    .B_N(_1078_),
    .Y(_1085_));
 sg13g2_a21oi_1 _3090_ (.A1(_1083_),
    .A2(_1085_),
    .Y(_1086_),
    .B1(_1076_));
 sg13g2_nand2_1 _3091_ (.Y(_1087_),
    .A(_1084_),
    .B(_1086_));
 sg13g2_nand2_1 _3092_ (.Y(_1088_),
    .A(_1074_),
    .B(_1087_));
 sg13g2_nand2_1 _3093_ (.Y(_1089_),
    .A(_1070_),
    .B(_1885_));
 sg13g2_nand3_1 _3094_ (.B(_1069_),
    .C(_1886_),
    .A(_1066_),
    .Y(_1090_));
 sg13g2_nand2_1 _3095_ (.Y(_1091_),
    .A(_1089_),
    .B(_1090_));
 sg13g2_a21oi_1 _3096_ (.A1(_1052_),
    .A2(_1053_),
    .Y(_1092_),
    .B1(_0032_));
 sg13g2_a21oi_1 _3097_ (.A1(_1066_),
    .A2(_1069_),
    .Y(_1093_),
    .B1(_1857_));
 sg13g2_a21oi_1 _3098_ (.A1(_1091_),
    .A2(_1092_),
    .Y(_1094_),
    .B1(_1093_));
 sg13g2_nand2_1 _3099_ (.Y(_1095_),
    .A(_1088_),
    .B(_1094_));
 sg13g2_nor3_1 _3100_ (.A(_1050_),
    .B(_1067_),
    .C(_1045_),
    .Y(_1096_));
 sg13g2_a21oi_1 _3101_ (.A1(_1060_),
    .A2(_1064_),
    .Y(_1097_),
    .B1(_1063_));
 sg13g2_nor2b_1 _3102_ (.A(_1096_),
    .B_N(_1097_),
    .Y(_1098_));
 sg13g2_nand4_1 _3103_ (.B(_1065_),
    .C(_1039_),
    .A(_1035_),
    .Y(_1099_),
    .D(_1051_));
 sg13g2_nand2_1 _3104_ (.Y(_1100_),
    .A(_1098_),
    .B(_1099_));
 sg13g2_inv_1 _3105_ (.Y(_1101_),
    .A(_1007_));
 sg13g2_nor2_1 _3106_ (.A(_1026_),
    .B(_1025_),
    .Y(_1102_));
 sg13g2_nor2_1 _3107_ (.A(_0812_),
    .B(_1102_),
    .Y(_1103_));
 sg13g2_nor2_1 _3108_ (.A(_1101_),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_nand2_1 _3109_ (.Y(_1105_),
    .A(_1103_),
    .B(_1101_));
 sg13g2_nand2b_1 _3110_ (.Y(_1106_),
    .B(_1105_),
    .A_N(_1104_));
 sg13g2_inv_1 _3111_ (.Y(_1107_),
    .A(_1106_));
 sg13g2_nand2_1 _3112_ (.Y(_1108_),
    .A(_1100_),
    .B(_1107_));
 sg13g2_nand3_1 _3113_ (.B(_1099_),
    .C(_1106_),
    .A(_1098_),
    .Y(_1109_));
 sg13g2_nand2_1 _3114_ (.Y(_1110_),
    .A(_1108_),
    .B(_1109_));
 sg13g2_nand2_1 _3115_ (.Y(_1111_),
    .A(_1110_),
    .B(_1895_));
 sg13g2_nand3_1 _3116_ (.B(_1109_),
    .C(_1894_),
    .A(_1108_),
    .Y(_1112_));
 sg13g2_nand2_1 _3117_ (.Y(_1113_),
    .A(_1111_),
    .B(_1112_));
 sg13g2_nor3_1 _3118_ (.A(_1067_),
    .B(_1106_),
    .C(_1061_),
    .Y(_1114_));
 sg13g2_a21oi_1 _3119_ (.A1(_1105_),
    .A2(_1063_),
    .Y(_1115_),
    .B1(_1104_));
 sg13g2_nor2b_1 _3120_ (.A(_1114_),
    .B_N(_1115_),
    .Y(_1116_));
 sg13g2_nand4_1 _3121_ (.B(_1057_),
    .C(_1058_),
    .A(_1107_),
    .Y(_1117_),
    .D(_1065_));
 sg13g2_nand2_1 _3122_ (.Y(_1118_),
    .A(_1116_),
    .B(_1117_));
 sg13g2_inv_1 _3123_ (.Y(_1119_),
    .A(_1025_));
 sg13g2_nand2_1 _3124_ (.Y(_1120_),
    .A(_1118_),
    .B(_1119_));
 sg13g2_nand2_1 _3125_ (.Y(_1121_),
    .A(_1120_),
    .B(_1901_));
 sg13g2_inv_1 _3126_ (.Y(_1122_),
    .A(_1901_));
 sg13g2_nand3_1 _3127_ (.B(_1122_),
    .C(_1119_),
    .A(_1118_),
    .Y(_1123_));
 sg13g2_nand2_1 _3128_ (.Y(_1124_),
    .A(_1121_),
    .B(_1123_));
 sg13g2_nor2b_1 _3129_ (.A(_1113_),
    .B_N(_1124_),
    .Y(_1125_));
 sg13g2_nand2_1 _3130_ (.Y(_1126_),
    .A(_1095_),
    .B(_1125_));
 sg13g2_a21oi_1 _3131_ (.A1(_1108_),
    .A2(_1109_),
    .Y(_1127_),
    .B1(_1856_));
 sg13g2_a21oi_1 _3132_ (.A1(_1118_),
    .A2(_1119_),
    .Y(_1128_),
    .B1(_1901_));
 sg13g2_a21oi_1 _3133_ (.A1(_1124_),
    .A2(_1127_),
    .Y(_1129_),
    .B1(_1128_));
 sg13g2_nand3_1 _3134_ (.B(_1043_),
    .C(_1129_),
    .A(_1126_),
    .Y(_1130_));
 sg13g2_nand2_1 _3135_ (.Y(_1131_),
    .A(_1130_),
    .B(_1103_));
 sg13g2_nand4_1 _3136_ (.B(_1020_),
    .C(_1043_),
    .A(_1126_),
    .Y(_1132_),
    .D(_1129_));
 sg13g2_nand2_1 _3137_ (.Y(net9),
    .A(_1131_),
    .B(_1132_));
 sg13g2_nand2_1 _3138_ (.Y(_1133_),
    .A(_2127_),
    .B(_2128_));
 sg13g2_nand3_1 _3139_ (.B(_2129_),
    .C(_2126_),
    .A(_2122_),
    .Y(_1134_));
 sg13g2_nand2_1 _3140_ (.Y(_1135_),
    .A(_1742_),
    .B(_2049_));
 sg13g2_nand2_1 _3141_ (.Y(_1136_),
    .A(_1706_),
    .B(_2048_));
 sg13g2_nand2_1 _3142_ (.Y(_1137_),
    .A(_1135_),
    .B(_1136_));
 sg13g2_inv_1 _3143_ (.Y(_1138_),
    .A(_1137_));
 sg13g2_nand3_1 _3144_ (.B(_1134_),
    .C(_1138_),
    .A(_1133_),
    .Y(_1139_));
 sg13g2_nand3_1 _3145_ (.B(_2131_),
    .C(_1137_),
    .A(_2130_),
    .Y(_1140_));
 sg13g2_nand2_1 _3146_ (.Y(_1141_),
    .A(_1139_),
    .B(_1140_));
 sg13g2_nand2_1 _3147_ (.Y(_1142_),
    .A(_1718_),
    .B(_2051_));
 sg13g2_nand2_1 _3148_ (.Y(_1143_),
    .A(net59),
    .B(net64));
 sg13g2_inv_1 _3149_ (.Y(_1144_),
    .A(_1143_));
 sg13g2_a21oi_1 _3150_ (.A1(_0160_),
    .A2(_1142_),
    .Y(_1145_),
    .B1(_1144_));
 sg13g2_nand2_1 _3151_ (.Y(_1146_),
    .A(_1141_),
    .B(_1145_));
 sg13g2_xor2_1 _3152_ (.B(_2052_),
    .A(net58),
    .X(_1147_));
 sg13g2_nand2_1 _3153_ (.Y(_1148_),
    .A(_2229_),
    .B(_1147_));
 sg13g2_nand2_1 _3154_ (.Y(_1149_),
    .A(net58),
    .B(_2052_));
 sg13g2_nand2_1 _3155_ (.Y(_1150_),
    .A(_1148_),
    .B(_1149_));
 sg13g2_inv_1 _3156_ (.Y(_1151_),
    .A(_1150_));
 sg13g2_nand2_1 _3157_ (.Y(_1152_),
    .A(_1142_),
    .B(_1143_));
 sg13g2_nand2b_1 _3158_ (.Y(_1153_),
    .B(net22),
    .A_N(_1152_));
 sg13g2_nand3_1 _3159_ (.B(_0159_),
    .C(_1152_),
    .A(_0154_),
    .Y(_1154_));
 sg13g2_nand2_1 _3160_ (.Y(_1155_),
    .A(_1153_),
    .B(_1154_));
 sg13g2_nor2_2 _3161_ (.A(_1151_),
    .B(_1155_),
    .Y(_1156_));
 sg13g2_nor2_1 _3162_ (.A(_1145_),
    .B(_1141_),
    .Y(_1157_));
 sg13g2_a21oi_1 _3163_ (.A1(_1146_),
    .A2(_1156_),
    .Y(_1158_),
    .B1(_1157_));
 sg13g2_nand2_1 _3164_ (.Y(_1159_),
    .A(_1709_),
    .B(_2047_));
 sg13g2_nand2_1 _3165_ (.Y(_1160_),
    .A(_1708_),
    .B(_2046_));
 sg13g2_nand2_1 _3166_ (.Y(_1161_),
    .A(_1159_),
    .B(_1160_));
 sg13g2_nand2b_1 _3167_ (.Y(_1162_),
    .B(_2152_),
    .A_N(_1161_));
 sg13g2_nand3_1 _3168_ (.B(_2150_),
    .C(_1161_),
    .A(_2149_),
    .Y(_1163_));
 sg13g2_nand2_1 _3169_ (.Y(_1164_),
    .A(_1162_),
    .B(_1163_));
 sg13g2_nand2_1 _3170_ (.Y(_1165_),
    .A(_1139_),
    .B(_1136_));
 sg13g2_inv_1 _3171_ (.Y(_1166_),
    .A(_1165_));
 sg13g2_nand2_1 _3172_ (.Y(_1167_),
    .A(_1164_),
    .B(_1166_));
 sg13g2_nand3_1 _3173_ (.B(_1163_),
    .C(_1165_),
    .A(_1162_),
    .Y(_1168_));
 sg13g2_nand2_2 _3174_ (.Y(_1169_),
    .A(_1167_),
    .B(_1168_));
 sg13g2_xor2_1 _3175_ (.B(_2043_),
    .A(\i_project.controller_0.h[6] ),
    .X(_1170_));
 sg13g2_inv_1 _3176_ (.Y(_1171_),
    .A(_1170_));
 sg13g2_xnor2_1 _3177_ (.Y(_1172_),
    .A(_1171_),
    .B(_2206_));
 sg13g2_nand2_1 _3178_ (.Y(_1173_),
    .A(_1162_),
    .B(_1160_));
 sg13g2_nand2_1 _3179_ (.Y(_1174_),
    .A(_1172_),
    .B(_1173_));
 sg13g2_nand2_1 _3180_ (.Y(_1175_),
    .A(_2196_),
    .B(_1170_));
 sg13g2_nand3_1 _3181_ (.B(_2195_),
    .C(_1171_),
    .A(_2194_),
    .Y(_1176_));
 sg13g2_nand2_1 _3182_ (.Y(_1177_),
    .A(_1175_),
    .B(_1176_));
 sg13g2_inv_1 _3183_ (.Y(_1178_),
    .A(_1160_));
 sg13g2_a21oi_1 _3184_ (.A1(net18),
    .A2(_1159_),
    .Y(_1179_),
    .B1(_1178_));
 sg13g2_nand2_1 _3185_ (.Y(_1180_),
    .A(_1177_),
    .B(_1179_));
 sg13g2_nand2_1 _3186_ (.Y(_1181_),
    .A(_1174_),
    .B(_1180_));
 sg13g2_nor3_1 _3187_ (.A(_1158_),
    .B(_1169_),
    .C(_1181_),
    .Y(_1182_));
 sg13g2_inv_1 _3188_ (.Y(_1183_),
    .A(_1168_));
 sg13g2_inv_1 _3189_ (.Y(_1184_),
    .A(_1174_));
 sg13g2_a21oi_1 _3190_ (.A1(_1183_),
    .A2(_1180_),
    .Y(_1185_),
    .B1(_1184_));
 sg13g2_nor2b_1 _3191_ (.A(_1182_),
    .B_N(_1185_),
    .Y(_1186_));
 sg13g2_nor2_1 _3192_ (.A(_1169_),
    .B(_1181_),
    .Y(_1187_));
 sg13g2_inv_1 _3193_ (.Y(_1188_),
    .A(net63));
 sg13g2_xor2_1 _3194_ (.B(net63),
    .A(net71),
    .X(_1189_));
 sg13g2_nand2_1 _3195_ (.Y(_1190_),
    .A(net26),
    .B(_1189_));
 sg13g2_o21ai_1 _3196_ (.B1(_1190_),
    .Y(_1191_),
    .A1(_1715_),
    .A2(_1188_));
 sg13g2_xor2_1 _3197_ (.B(_2229_),
    .A(_1147_),
    .X(_1192_));
 sg13g2_nor2_1 _3198_ (.A(_1191_),
    .B(_1192_),
    .Y(_1193_));
 sg13g2_xnor2_1 _3199_ (.Y(_1194_),
    .A(_1189_),
    .B(net26));
 sg13g2_inv_1 _3200_ (.Y(_1195_),
    .A(_0056_));
 sg13g2_nor2_1 _3201_ (.A(_1195_),
    .B(net35),
    .Y(_1196_));
 sg13g2_nand2_1 _3202_ (.Y(_1197_),
    .A(_1194_),
    .B(_1196_));
 sg13g2_xnor2_1 _3203_ (.Y(_1198_),
    .A(_2035_),
    .B(net35));
 sg13g2_nor2_1 _3204_ (.A(_0269_),
    .B(_1198_),
    .Y(_1199_));
 sg13g2_nor2_1 _3205_ (.A(_1196_),
    .B(_1194_),
    .Y(_1200_));
 sg13g2_a21oi_2 _3206_ (.B1(_1200_),
    .Y(_1201_),
    .A2(_1199_),
    .A1(_1197_));
 sg13g2_nand2_1 _3207_ (.Y(_1202_),
    .A(_1192_),
    .B(_1191_));
 sg13g2_o21ai_1 _3208_ (.B1(_1202_),
    .Y(_1203_),
    .A1(_1193_),
    .A2(_1201_));
 sg13g2_buf_2 _3209_ (.A(_1203_),
    .X(_1204_));
 sg13g2_inv_1 _3210_ (.Y(_1205_),
    .A(_1157_));
 sg13g2_nand2_2 _3211_ (.Y(_1206_),
    .A(_1205_),
    .B(_1146_));
 sg13g2_nand2_1 _3212_ (.Y(_1207_),
    .A(_1155_),
    .B(_1151_));
 sg13g2_nand2b_1 _3213_ (.Y(_1208_),
    .B(_1207_),
    .A_N(_1156_));
 sg13g2_nor2_1 _3214_ (.A(_1206_),
    .B(_1208_),
    .Y(_1209_));
 sg13g2_nand3_1 _3215_ (.B(_1204_),
    .C(_1209_),
    .A(_1187_),
    .Y(_1210_));
 sg13g2_nand2_1 _3216_ (.Y(_1211_),
    .A(_1186_),
    .B(_1210_));
 sg13g2_o21ai_1 _3217_ (.B1(_1175_),
    .Y(_1212_),
    .A1(_1732_),
    .A2(_2059_));
 sg13g2_xnor2_1 _3218_ (.Y(_1213_),
    .A(net70),
    .B(net66));
 sg13g2_xnor2_1 _3219_ (.Y(_1214_),
    .A(_1213_),
    .B(_2179_));
 sg13g2_xor2_1 _3220_ (.B(_1214_),
    .A(_1212_),
    .X(_1215_));
 sg13g2_nand2_1 _3221_ (.Y(_1216_),
    .A(_1211_),
    .B(_1215_));
 sg13g2_inv_1 _3222_ (.Y(_1217_),
    .A(_1215_));
 sg13g2_nand3_1 _3223_ (.B(_1210_),
    .C(_1217_),
    .A(_1186_),
    .Y(_1218_));
 sg13g2_nand3_1 _3224_ (.B(_1218_),
    .C(_0233_),
    .A(_1216_),
    .Y(_1219_));
 sg13g2_xor2_1 _3225_ (.B(net66),
    .A(net72),
    .X(_1220_));
 sg13g2_nand2_1 _3226_ (.Y(_1221_),
    .A(net58),
    .B(net64));
 sg13g2_xnor2_1 _3227_ (.Y(_1222_),
    .A(net59),
    .B(net65));
 sg13g2_nand2_1 _3228_ (.Y(_1223_),
    .A(net59),
    .B(net65));
 sg13g2_o21ai_1 _3229_ (.B1(_1223_),
    .Y(_1224_),
    .A1(_1221_),
    .A2(_1222_));
 sg13g2_xnor2_1 _3230_ (.Y(_1225_),
    .A(net61),
    .B(net53));
 sg13g2_nor2_1 _3231_ (.A(net57),
    .B(net54),
    .Y(_1226_));
 sg13g2_nand2_1 _3232_ (.Y(_1227_),
    .A(net57),
    .B(net54));
 sg13g2_nor2b_1 _3233_ (.A(_1226_),
    .B_N(_1227_),
    .Y(_1228_));
 sg13g2_nor2b_1 _3234_ (.A(_1225_),
    .B_N(_1228_),
    .Y(_1229_));
 sg13g2_nand2_1 _3235_ (.Y(_1230_),
    .A(net61),
    .B(net53));
 sg13g2_o21ai_1 _3236_ (.B1(_1227_),
    .Y(_1231_),
    .A1(_1230_),
    .A2(_1226_));
 sg13g2_a21oi_1 _3237_ (.A1(_1224_),
    .A2(_1229_),
    .Y(_1232_),
    .B1(_1231_));
 sg13g2_nand2_1 _3238_ (.Y(_1233_),
    .A(_1712_),
    .B(\i_project.controller_0.mode_ramp_base[1] ));
 sg13g2_xnor2_1 _3239_ (.Y(_1234_),
    .A(net71),
    .B(_2052_));
 sg13g2_nor2_1 _3240_ (.A(_1233_),
    .B(_1234_),
    .Y(_1235_));
 sg13g2_nand2_1 _3241_ (.Y(_1236_),
    .A(net71),
    .B(_2052_));
 sg13g2_nor2b_1 _3242_ (.A(_1235_),
    .B_N(_1236_),
    .Y(_1237_));
 sg13g2_inv_1 _3243_ (.Y(_1238_),
    .A(_1237_));
 sg13g2_nand2_1 _3244_ (.Y(_1239_),
    .A(_1720_),
    .B(_2051_));
 sg13g2_nand2_1 _3245_ (.Y(_1240_),
    .A(_1239_),
    .B(_1221_));
 sg13g2_nor2_1 _3246_ (.A(_1222_),
    .B(_1240_),
    .Y(_1241_));
 sg13g2_nand3_1 _3247_ (.B(_1229_),
    .C(_1241_),
    .A(_1238_),
    .Y(_1242_));
 sg13g2_nand2_1 _3248_ (.Y(_1243_),
    .A(_1232_),
    .B(_1242_));
 sg13g2_xnor2_1 _3249_ (.Y(_1244_),
    .A(_1220_),
    .B(_1243_));
 sg13g2_xnor2_1 _3250_ (.Y(_1245_),
    .A(_0729_),
    .B(net19));
 sg13g2_xnor2_1 _3251_ (.Y(_1246_),
    .A(_1244_),
    .B(_1245_));
 sg13g2_nor2_1 _3252_ (.A(_0164_),
    .B(net20),
    .Y(_1247_));
 sg13g2_inv_1 _3253_ (.Y(_1248_),
    .A(_1247_));
 sg13g2_xnor2_1 _3254_ (.Y(_1249_),
    .A(_2112_),
    .B(net18));
 sg13g2_nor2_1 _3255_ (.A(_1248_),
    .B(_1249_),
    .Y(_1250_));
 sg13g2_a21oi_1 _3256_ (.A1(_0787_),
    .A2(_0837_),
    .Y(_1251_),
    .B1(_1250_));
 sg13g2_nor2_1 _3257_ (.A(_0044_),
    .B(_2213_),
    .Y(_1252_));
 sg13g2_xnor2_1 _3258_ (.Y(_1253_),
    .A(net64),
    .B(_2213_));
 sg13g2_nor2_1 _3259_ (.A(_2053_),
    .B(net35),
    .Y(_1254_));
 sg13g2_nand2_1 _3260_ (.Y(_1255_),
    .A(_1253_),
    .B(_1254_));
 sg13g2_nand2b_1 _3261_ (.Y(_1256_),
    .B(_1255_),
    .A_N(_1252_));
 sg13g2_xnor2_1 _3262_ (.Y(_1257_),
    .A(_2049_),
    .B(_2229_));
 sg13g2_inv_1 _3263_ (.Y(_1258_),
    .A(_1257_));
 sg13g2_nand2_1 _3264_ (.Y(_1259_),
    .A(_1256_),
    .B(_1258_));
 sg13g2_nand2_1 _3265_ (.Y(_1260_),
    .A(_0150_),
    .B(_0782_));
 sg13g2_nand2_1 _3266_ (.Y(_1261_),
    .A(_1259_),
    .B(_1260_));
 sg13g2_xnor2_1 _3267_ (.Y(_1262_),
    .A(net53),
    .B(net22));
 sg13g2_nand2_1 _3268_ (.Y(_1263_),
    .A(_1261_),
    .B(_1262_));
 sg13g2_nand2_1 _3269_ (.Y(_1264_),
    .A(_0781_),
    .B(_0151_));
 sg13g2_nand2_1 _3270_ (.Y(_1265_),
    .A(_1263_),
    .B(_1264_));
 sg13g2_xnor2_1 _3271_ (.Y(_1266_),
    .A(_2059_),
    .B(net20));
 sg13g2_nor2_1 _3272_ (.A(_1266_),
    .B(_1249_),
    .Y(_1267_));
 sg13g2_nand2_1 _3273_ (.Y(_1268_),
    .A(_1265_),
    .B(_1267_));
 sg13g2_nand2_1 _3274_ (.Y(_1269_),
    .A(_1251_),
    .B(_1268_));
 sg13g2_nand2b_1 _3275_ (.Y(_1270_),
    .B(_1269_),
    .A_N(_1246_));
 sg13g2_nand3_1 _3276_ (.B(_1268_),
    .C(_1246_),
    .A(_1251_),
    .Y(_1271_));
 sg13g2_nand3_1 _3277_ (.B(_1271_),
    .C(net42),
    .A(_1270_),
    .Y(_1272_));
 sg13g2_a21oi_1 _3278_ (.A1(_1272_),
    .A2(_0304_),
    .Y(_1273_),
    .B1(_0235_));
 sg13g2_nand2_1 _3279_ (.Y(_1274_),
    .A(_1219_),
    .B(_1273_));
 sg13g2_xnor2_1 _3280_ (.Y(_1275_),
    .A(net66),
    .B(_0254_));
 sg13g2_a21oi_1 _3281_ (.A1(_1275_),
    .A2(net34),
    .Y(_1276_),
    .B1(net41));
 sg13g2_nand2_1 _3282_ (.Y(_1277_),
    .A(_1274_),
    .B(_1276_));
 sg13g2_a21oi_1 _3283_ (.A1(_0787_),
    .A2(net41),
    .Y(_1278_),
    .B1(net27));
 sg13g2_nand2_1 _3284_ (.Y(_1279_),
    .A(_1277_),
    .B(_1278_));
 sg13g2_nand2_1 _3285_ (.Y(_1280_),
    .A(_1279_),
    .B(_0288_));
 sg13g2_nand2_1 _3286_ (.Y(_1281_),
    .A(_1280_),
    .B(net43));
 sg13g2_nand2_1 _3287_ (.Y(_1282_),
    .A(_1281_),
    .B(_2104_));
 sg13g2_buf_8 _3288_ (.A(_1282_),
    .X(_1283_));
 sg13g2_nor2_1 _3289_ (.A(_0530_),
    .B(_1283_),
    .Y(_1284_));
 sg13g2_xnor2_1 _3290_ (.Y(_1285_),
    .A(net54),
    .B(net20));
 sg13g2_nand2_1 _3291_ (.Y(_1286_),
    .A(_1265_),
    .B(_1285_));
 sg13g2_nand3_1 _3292_ (.B(_1266_),
    .C(_1264_),
    .A(_1263_),
    .Y(_1287_));
 sg13g2_nand2_1 _3293_ (.Y(_1288_),
    .A(_1286_),
    .B(_1287_));
 sg13g2_a21oi_1 _3294_ (.A1(_1238_),
    .A2(_1241_),
    .Y(_1289_),
    .B1(_1224_));
 sg13g2_xor2_1 _3295_ (.B(_1289_),
    .A(_1225_),
    .X(_1290_));
 sg13g2_nand2_1 _3296_ (.Y(_1291_),
    .A(_1288_),
    .B(_1290_));
 sg13g2_inv_1 _3297_ (.Y(_1292_),
    .A(_1290_));
 sg13g2_nand3_1 _3298_ (.B(_1287_),
    .C(_1292_),
    .A(_1286_),
    .Y(_1293_));
 sg13g2_nand3_1 _3299_ (.B(_1293_),
    .C(net40),
    .A(_1291_),
    .Y(_1294_));
 sg13g2_inv_1 _3300_ (.Y(_1295_),
    .A(_0574_));
 sg13g2_a21oi_1 _3301_ (.A1(_1294_),
    .A2(_1295_),
    .Y(_1296_),
    .B1(net39));
 sg13g2_nor2b_1 _3302_ (.A(_1156_),
    .B_N(_1207_),
    .Y(_1297_));
 sg13g2_nand2_1 _3303_ (.Y(_1298_),
    .A(_1297_),
    .B(_1204_));
 sg13g2_nand3b_1 _3304_ (.B(_1298_),
    .C(_1205_),
    .Y(_1299_),
    .A_N(_1156_));
 sg13g2_nand2_1 _3305_ (.Y(_1300_),
    .A(_1299_),
    .B(_1146_));
 sg13g2_nor2_1 _3306_ (.A(_1169_),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_a21oi_1 _3307_ (.A1(_1300_),
    .A2(_1169_),
    .Y(_1302_),
    .B1(net45));
 sg13g2_nand2b_1 _3308_ (.Y(_1303_),
    .B(_1302_),
    .A_N(_1301_));
 sg13g2_nand2_1 _3309_ (.Y(_1304_),
    .A(_1296_),
    .B(_1303_));
 sg13g2_xnor2_1 _3310_ (.Y(_1305_),
    .A(net53),
    .B(net29));
 sg13g2_a21oi_1 _3311_ (.A1(_1305_),
    .A2(net39),
    .Y(_1306_),
    .B1(net38));
 sg13g2_nand2_1 _3312_ (.Y(_1307_),
    .A(_1304_),
    .B(_1306_));
 sg13g2_a21oi_1 _3313_ (.A1(_0151_),
    .A2(net38),
    .Y(_1308_),
    .B1(net27));
 sg13g2_nand2_1 _3314_ (.Y(_1309_),
    .A(_1307_),
    .B(_1308_));
 sg13g2_nand2_1 _3315_ (.Y(_1310_),
    .A(_1309_),
    .B(net17));
 sg13g2_nand2_1 _3316_ (.Y(_1311_),
    .A(_1310_),
    .B(net43));
 sg13g2_nand3_1 _3317_ (.B(_0333_),
    .C(_0513_),
    .A(_1311_),
    .Y(_1312_));
 sg13g2_nand3_1 _3318_ (.B(net46),
    .C(_0335_),
    .A(_1311_),
    .Y(_1313_));
 sg13g2_nand2_1 _3319_ (.Y(_1314_),
    .A(_1312_),
    .B(_1313_));
 sg13g2_nor2_2 _3320_ (.A(_1284_),
    .B(_1314_),
    .Y(_1315_));
 sg13g2_inv_1 _3321_ (.Y(_1316_),
    .A(_0445_));
 sg13g2_inv_1 _3322_ (.Y(_1317_),
    .A(_1202_));
 sg13g2_a21oi_1 _3323_ (.A1(_1207_),
    .A2(_1317_),
    .Y(_1318_),
    .B1(_1156_));
 sg13g2_nor3_1 _3324_ (.A(_1206_),
    .B(_1318_),
    .C(_1169_),
    .Y(_1319_));
 sg13g2_a21oi_1 _3325_ (.A1(_1167_),
    .A2(_1157_),
    .Y(_1320_),
    .B1(_1183_));
 sg13g2_nor2b_1 _3326_ (.A(_1319_),
    .B_N(_1320_),
    .Y(_1321_));
 sg13g2_nor2_1 _3327_ (.A(_1206_),
    .B(_1169_),
    .Y(_1322_));
 sg13g2_inv_1 _3328_ (.Y(_1323_),
    .A(_1201_));
 sg13g2_nand2b_1 _3329_ (.Y(_1324_),
    .B(_1202_),
    .A_N(_1193_));
 sg13g2_nor2_1 _3330_ (.A(_1324_),
    .B(_1208_),
    .Y(_1325_));
 sg13g2_nand3_1 _3331_ (.B(_1323_),
    .C(_1325_),
    .A(_1322_),
    .Y(_1326_));
 sg13g2_nand2_1 _3332_ (.Y(_1327_),
    .A(_1321_),
    .B(_1326_));
 sg13g2_nand2b_1 _3333_ (.Y(_1328_),
    .B(_1327_),
    .A_N(_1181_));
 sg13g2_nand3_1 _3334_ (.B(_1326_),
    .C(_1181_),
    .A(_1321_),
    .Y(_1329_));
 sg13g2_nand3_1 _3335_ (.B(_1329_),
    .C(_0233_),
    .A(_1328_),
    .Y(_1330_));
 sg13g2_o21ai_1 _3336_ (.B1(_1230_),
    .Y(_1331_),
    .A1(_1225_),
    .A2(_1289_));
 sg13g2_xnor2_1 _3337_ (.Y(_1332_),
    .A(_1228_),
    .B(_1331_));
 sg13g2_xor2_1 _3338_ (.B(_1332_),
    .A(_1249_),
    .X(_1333_));
 sg13g2_a22oi_1 _3339_ (.Y(_1334_),
    .B1(_1252_),
    .B2(_1258_),
    .A2(_0150_),
    .A1(_0782_));
 sg13g2_nand2_1 _3340_ (.Y(_1335_),
    .A(_1285_),
    .B(_1262_));
 sg13g2_nor2_1 _3341_ (.A(_1334_),
    .B(_1335_),
    .Y(_1336_));
 sg13g2_o21ai_1 _3342_ (.B1(_1248_),
    .Y(_1337_),
    .A1(_1264_),
    .A2(_1266_));
 sg13g2_nor2_1 _3343_ (.A(_1336_),
    .B(_1337_),
    .Y(_1338_));
 sg13g2_nor2b_1 _3344_ (.A(_1257_),
    .B_N(_1253_),
    .Y(_1339_));
 sg13g2_nand4_1 _3345_ (.B(_1262_),
    .C(_1254_),
    .A(_1285_),
    .Y(_1340_),
    .D(_1339_));
 sg13g2_nand2_1 _3346_ (.Y(_1341_),
    .A(_1338_),
    .B(_1340_));
 sg13g2_xnor2_1 _3347_ (.Y(_1342_),
    .A(_1333_),
    .B(_1341_));
 sg13g2_nand2_1 _3348_ (.Y(_1343_),
    .A(_1342_),
    .B(net42));
 sg13g2_a21oi_1 _3349_ (.A1(_1343_),
    .A2(_0467_),
    .Y(_1344_),
    .B1(_0235_));
 sg13g2_nand2_1 _3350_ (.Y(_1345_),
    .A(_1330_),
    .B(_1344_));
 sg13g2_xnor2_1 _3351_ (.Y(_1346_),
    .A(net54),
    .B(_0254_));
 sg13g2_a21oi_1 _3352_ (.A1(_1346_),
    .A2(_0235_),
    .Y(_1347_),
    .B1(_0257_));
 sg13g2_nand2_1 _3353_ (.Y(_1348_),
    .A(_1345_),
    .B(_1347_));
 sg13g2_inv_1 _3354_ (.Y(_1349_),
    .A(_0164_));
 sg13g2_a21oi_1 _3355_ (.A1(_1349_),
    .A2(net41),
    .Y(_1350_),
    .B1(net27));
 sg13g2_nand2_1 _3356_ (.Y(_1351_),
    .A(_1348_),
    .B(_1350_));
 sg13g2_nand2_1 _3357_ (.Y(_1352_),
    .A(_1351_),
    .B(_0432_));
 sg13g2_nand2_1 _3358_ (.Y(_1353_),
    .A(_1352_),
    .B(_0435_));
 sg13g2_nand2_1 _3359_ (.Y(_1354_),
    .A(_1353_),
    .B(_0331_));
 sg13g2_a21oi_1 _3360_ (.A1(_1316_),
    .A2(_0533_),
    .Y(_1355_),
    .B1(_1354_));
 sg13g2_inv_1 _3361_ (.Y(_1356_),
    .A(_1239_));
 sg13g2_o21ai_1 _3362_ (.B1(_1221_),
    .Y(_1357_),
    .A1(_1356_),
    .A2(_1237_));
 sg13g2_xnor2_1 _3363_ (.Y(_1358_),
    .A(_1222_),
    .B(_1357_));
 sg13g2_xnor2_1 _3364_ (.Y(_1359_),
    .A(_1262_),
    .B(_1261_));
 sg13g2_xnor2_1 _3365_ (.Y(_1360_),
    .A(_1358_),
    .B(_1359_));
 sg13g2_o21ai_1 _3366_ (.B1(_0345_),
    .Y(_1361_),
    .A1(net37),
    .A2(_1360_));
 sg13g2_a21oi_1 _3367_ (.A1(_1204_),
    .A2(_1207_),
    .Y(_1362_),
    .B1(_1156_));
 sg13g2_xor2_1 _3368_ (.B(_1362_),
    .A(_1206_),
    .X(_1363_));
 sg13g2_nand2_1 _3369_ (.Y(_1364_),
    .A(_1363_),
    .B(net51));
 sg13g2_nand3_1 _3370_ (.B(_1364_),
    .C(_0541_),
    .A(_1361_),
    .Y(_1365_));
 sg13g2_a21oi_1 _3371_ (.A1(net29),
    .A2(_2049_),
    .Y(_1366_),
    .B1(_0360_));
 sg13g2_o21ai_1 _3372_ (.B1(_1366_),
    .Y(_1367_),
    .A1(_2049_),
    .A2(net23));
 sg13g2_nand3_1 _3373_ (.B(net33),
    .C(_1367_),
    .A(_1365_),
    .Y(_1368_));
 sg13g2_a21oi_1 _3374_ (.A1(_0782_),
    .A2(net36),
    .Y(_1369_),
    .B1(net25));
 sg13g2_nand2_1 _3375_ (.Y(_1370_),
    .A(_1368_),
    .B(_1369_));
 sg13g2_nand2_1 _3376_ (.Y(_1371_),
    .A(_1370_),
    .B(_0432_));
 sg13g2_nand2_1 _3377_ (.Y(_1372_),
    .A(_1371_),
    .B(_0481_));
 sg13g2_xnor2_1 _3378_ (.Y(_1373_),
    .A(_2035_),
    .B(net23));
 sg13g2_xnor2_1 _3379_ (.Y(_1374_),
    .A(_0054_),
    .B(_1198_));
 sg13g2_o21ai_1 _3380_ (.B1(net30),
    .Y(_1375_),
    .A1(net45),
    .A2(_1374_));
 sg13g2_o21ai_1 _3381_ (.B1(_1375_),
    .Y(_1376_),
    .A1(net30),
    .A2(_1373_));
 sg13g2_nand2_1 _3382_ (.Y(_1377_),
    .A(net32),
    .B(_1195_));
 sg13g2_nand3_1 _3383_ (.B(_0262_),
    .C(_1377_),
    .A(_1376_),
    .Y(_1378_));
 sg13g2_nand3_1 _3384_ (.B(_0499_),
    .C(_1378_),
    .A(net17),
    .Y(_1379_));
 sg13g2_nand2_1 _3385_ (.Y(_1380_),
    .A(_1379_),
    .B(_0501_));
 sg13g2_a21oi_1 _3386_ (.A1(_1372_),
    .A2(_0440_),
    .Y(_1381_),
    .B1(_1380_));
 sg13g2_nand2_1 _3387_ (.Y(_1382_),
    .A(_1353_),
    .B(_0456_));
 sg13g2_nand2_1 _3388_ (.Y(_1383_),
    .A(_1381_),
    .B(_1382_));
 sg13g2_nand3_1 _3389_ (.B(_2104_),
    .C(_0372_),
    .A(_1281_),
    .Y(_1384_));
 sg13g2_nand3_1 _3390_ (.B(net47),
    .C(_0335_),
    .A(_1311_),
    .Y(_1385_));
 sg13g2_nand2_1 _3391_ (.Y(_1386_),
    .A(_1384_),
    .B(_1385_));
 sg13g2_nor3_1 _3392_ (.A(_1355_),
    .B(_1383_),
    .C(_1386_),
    .Y(_1387_));
 sg13g2_nor2_1 _3393_ (.A(_1316_),
    .B(_1354_),
    .Y(_1388_));
 sg13g2_nand2_1 _3394_ (.Y(_1389_),
    .A(_1372_),
    .B(_0513_));
 sg13g2_nor2b_1 _3395_ (.A(_1388_),
    .B_N(_1389_),
    .Y(_1390_));
 sg13g2_inv_8 _3396_ (.Y(_1391_),
    .A(_1283_));
 sg13g2_nand2_1 _3397_ (.Y(_1392_),
    .A(_0501_),
    .B(_0533_));
 sg13g2_nand2_1 _3398_ (.Y(_1393_),
    .A(_1391_),
    .B(_1392_));
 sg13g2_nand2_2 _3399_ (.Y(_1394_),
    .A(_1390_),
    .B(_1393_));
 sg13g2_nor2b_1 _3400_ (.A(_1387_),
    .B_N(_1394_),
    .Y(_1395_));
 sg13g2_o21ai_1 _3401_ (.B1(net51),
    .Y(_1396_),
    .A1(_1201_),
    .A2(_1324_));
 sg13g2_a21oi_1 _3402_ (.A1(_1324_),
    .A2(_1201_),
    .Y(_1397_),
    .B1(_1396_));
 sg13g2_xor2_1 _3403_ (.B(_1234_),
    .A(_1233_),
    .X(_1398_));
 sg13g2_xor2_1 _3404_ (.B(_1253_),
    .A(_1254_),
    .X(_1399_));
 sg13g2_xor2_1 _3405_ (.B(_1399_),
    .A(_1398_),
    .X(_1400_));
 sg13g2_o21ai_1 _3406_ (.B1(_0490_),
    .Y(_1401_),
    .A1(net37),
    .A2(_1400_));
 sg13g2_nand3b_1 _3407_ (.B(net30),
    .C(_1401_),
    .Y(_1402_),
    .A_N(_1397_));
 sg13g2_a21oi_1 _3408_ (.A1(net29),
    .A2(_2053_),
    .Y(_1403_),
    .B1(net30));
 sg13g2_o21ai_1 _3409_ (.B1(_1403_),
    .Y(_1404_),
    .A1(_2053_),
    .A2(net23));
 sg13g2_nand3_1 _3410_ (.B(net33),
    .C(_1404_),
    .A(_1402_),
    .Y(_1405_));
 sg13g2_nand2b_1 _3411_ (.Y(_1406_),
    .B(net36),
    .A_N(_0045_));
 sg13g2_nand3_1 _3412_ (.B(_0262_),
    .C(_1406_),
    .A(_1405_),
    .Y(_1407_));
 sg13g2_a21oi_1 _3413_ (.A1(_1407_),
    .A2(net17),
    .Y(_1408_),
    .B1(net49));
 sg13g2_nand2b_1 _3414_ (.Y(_1409_),
    .B(_0378_),
    .A_N(_1408_));
 sg13g2_nand2_1 _3415_ (.Y(_1410_),
    .A(_1313_),
    .B(_1409_));
 sg13g2_nor2_1 _3416_ (.A(_1388_),
    .B(_1410_),
    .Y(_1411_));
 sg13g2_o21ai_1 _3417_ (.B1(_1391_),
    .Y(_1412_),
    .A1(net47),
    .A2(net24));
 sg13g2_nand2_1 _3418_ (.Y(_1413_),
    .A(_1353_),
    .B(_0440_));
 sg13g2_nand3_1 _3419_ (.B(_1412_),
    .C(_1413_),
    .A(_1411_),
    .Y(_1414_));
 sg13g2_buf_8 _3420_ (.A(_1414_),
    .X(_1415_));
 sg13g2_nand2_1 _3421_ (.Y(_1416_),
    .A(_1395_),
    .B(_1415_));
 sg13g2_a21oi_1 _3422_ (.A1(_0524_),
    .A2(_1353_),
    .Y(_1417_),
    .B1(_1355_));
 sg13g2_inv_2 _3423_ (.Y(_1418_),
    .A(_1354_));
 sg13g2_a21oi_1 _3424_ (.A1(_1418_),
    .A2(net47),
    .Y(_1419_),
    .B1(net24));
 sg13g2_nor2_1 _3425_ (.A(_0501_),
    .B(_1391_),
    .Y(_1420_));
 sg13g2_a21oi_1 _3426_ (.A1(_1417_),
    .A2(_1419_),
    .Y(_1421_),
    .B1(_1420_));
 sg13g2_nand2_1 _3427_ (.Y(_1422_),
    .A(_1416_),
    .B(_1421_));
 sg13g2_nor2_1 _3428_ (.A(_0567_),
    .B(_1283_),
    .Y(_1423_));
 sg13g2_nand2_1 _3429_ (.Y(_1424_),
    .A(_1418_),
    .B(net46));
 sg13g2_xnor2_1 _3430_ (.Y(_1425_),
    .A(_1204_),
    .B(_1297_));
 sg13g2_xnor2_1 _3431_ (.Y(_1426_),
    .A(_1240_),
    .B(_1237_));
 sg13g2_xnor2_1 _3432_ (.Y(_1427_),
    .A(_1258_),
    .B(_1256_));
 sg13g2_xnor2_1 _3433_ (.Y(_1428_),
    .A(_1426_),
    .B(_1427_));
 sg13g2_a21oi_1 _3434_ (.A1(_1428_),
    .A2(net40),
    .Y(_1429_),
    .B1(_0546_));
 sg13g2_nor2_1 _3435_ (.A(net39),
    .B(_1429_),
    .Y(_1430_));
 sg13g2_o21ai_1 _3436_ (.B1(_1430_),
    .Y(_1431_),
    .A1(_0540_),
    .A2(_1425_));
 sg13g2_a21oi_1 _3437_ (.A1(net29),
    .A2(_2051_),
    .Y(_1432_),
    .B1(_0360_));
 sg13g2_o21ai_1 _3438_ (.B1(_1432_),
    .Y(_1433_),
    .A1(_2051_),
    .A2(net23));
 sg13g2_nand3_1 _3439_ (.B(_0351_),
    .C(_1433_),
    .A(_1431_),
    .Y(_1434_));
 sg13g2_nand2_1 _3440_ (.Y(_1435_),
    .A(net36),
    .B(_0761_));
 sg13g2_nand3_1 _3441_ (.B(_0262_),
    .C(_1435_),
    .A(_1434_),
    .Y(_1436_));
 sg13g2_a21o_1 _3442_ (.A2(net17),
    .A1(_1436_),
    .B1(net49),
    .X(_1437_));
 sg13g2_a21oi_1 _3443_ (.A1(_1437_),
    .A2(_0585_),
    .Y(_1438_),
    .B1(net24));
 sg13g2_nand2_1 _3444_ (.Y(_1439_),
    .A(_1424_),
    .B(_1438_));
 sg13g2_nor2_1 _3445_ (.A(_1423_),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_nor2_1 _3446_ (.A(_1315_),
    .B(_1440_),
    .Y(_1441_));
 sg13g2_nand3_1 _3447_ (.B(_0440_),
    .C(_0333_),
    .A(_1311_),
    .Y(_1442_));
 sg13g2_nor2b_1 _3448_ (.A(_1200_),
    .B_N(_1197_),
    .Y(_1443_));
 sg13g2_xnor2_1 _3449_ (.Y(_1444_),
    .A(_1199_),
    .B(_1443_));
 sg13g2_o21ai_1 _3450_ (.B1(_0982_),
    .Y(_1445_),
    .A1(net45),
    .A2(_1444_));
 sg13g2_a21oi_1 _3451_ (.A1(net28),
    .A2(net63),
    .Y(_1446_),
    .B1(net30));
 sg13g2_o21ai_1 _3452_ (.B1(_1446_),
    .Y(_1447_),
    .A1(net63),
    .A2(net28));
 sg13g2_nand3_1 _3453_ (.B(net33),
    .C(_1447_),
    .A(_1445_),
    .Y(_1448_));
 sg13g2_nand2b_1 _3454_ (.Y(_1449_),
    .B(net32),
    .A_N(_0021_));
 sg13g2_nand3_1 _3455_ (.B(_0262_),
    .C(_1449_),
    .A(_1448_),
    .Y(_1450_));
 sg13g2_nand2_1 _3456_ (.Y(_1451_),
    .A(_0538_),
    .B(_1450_));
 sg13g2_nand2_1 _3457_ (.Y(_1452_),
    .A(_1442_),
    .B(_1451_));
 sg13g2_a21oi_1 _3458_ (.A1(_0564_),
    .A2(_1391_),
    .Y(_1453_),
    .B1(_1452_));
 sg13g2_nand2_1 _3459_ (.Y(_1454_),
    .A(_1453_),
    .B(_1419_));
 sg13g2_nand2_1 _3460_ (.Y(_1455_),
    .A(_1441_),
    .B(_1454_));
 sg13g2_nand2_1 _3461_ (.Y(_1456_),
    .A(_1455_),
    .B(_1391_));
 sg13g2_nand2_1 _3462_ (.Y(_1457_),
    .A(_1422_),
    .B(_1456_));
 sg13g2_nand2_1 _3463_ (.Y(_1458_),
    .A(_1415_),
    .B(_1454_));
 sg13g2_inv_2 _3464_ (.Y(_1459_),
    .A(_1440_));
 sg13g2_inv_1 _3465_ (.Y(_1460_),
    .A(_1420_));
 sg13g2_nand2_2 _3466_ (.Y(_1461_),
    .A(_1459_),
    .B(_1460_));
 sg13g2_nand2_1 _3467_ (.Y(_1462_),
    .A(_1458_),
    .B(_1461_));
 sg13g2_nor2_1 _3468_ (.A(_1391_),
    .B(_1390_),
    .Y(_1463_));
 sg13g2_nand2_1 _3469_ (.Y(_1464_),
    .A(_1462_),
    .B(_1463_));
 sg13g2_nand2_1 _3470_ (.Y(_1465_),
    .A(_1415_),
    .B(_1459_));
 sg13g2_nor2_1 _3471_ (.A(_1283_),
    .B(_1394_),
    .Y(_1466_));
 sg13g2_nand2_1 _3472_ (.Y(_1467_),
    .A(_1465_),
    .B(_1466_));
 sg13g2_nand2_1 _3473_ (.Y(_1468_),
    .A(_1417_),
    .B(_1419_));
 sg13g2_a21oi_1 _3474_ (.A1(_1468_),
    .A2(_1391_),
    .Y(_1469_),
    .B1(_1315_));
 sg13g2_nand2_1 _3475_ (.Y(_1470_),
    .A(_1467_),
    .B(_1469_));
 sg13g2_nand3_1 _3476_ (.B(_1464_),
    .C(_1470_),
    .A(_1457_),
    .Y(_1471_));
 sg13g2_nand2_1 _3477_ (.Y(_1472_),
    .A(_1471_),
    .B(_1283_));
 sg13g2_nand2_1 _3478_ (.Y(_1473_),
    .A(_1421_),
    .B(_1283_));
 sg13g2_nand2_1 _3479_ (.Y(_1474_),
    .A(_1468_),
    .B(_1460_));
 sg13g2_nand2_1 _3480_ (.Y(_1475_),
    .A(_1474_),
    .B(_1391_));
 sg13g2_nand2_1 _3481_ (.Y(_1476_),
    .A(_1473_),
    .B(_1475_));
 sg13g2_nand4_1 _3482_ (.B(_1464_),
    .C(_1470_),
    .A(_1457_),
    .Y(_1477_),
    .D(_1476_));
 sg13g2_nand2_1 _3483_ (.Y(_1478_),
    .A(_1472_),
    .B(_1477_));
 sg13g2_buf_8 _3484_ (.A(_1478_),
    .X(_1479_));
 sg13g2_xnor2_1 _3485_ (.Y(_1480_),
    .A(_1315_),
    .B(_1479_));
 sg13g2_xnor2_1 _3486_ (.Y(_1481_),
    .A(_1461_),
    .B(_1479_));
 sg13g2_nand2_1 _3487_ (.Y(_1482_),
    .A(_1471_),
    .B(_1421_));
 sg13g2_nand4_1 _3488_ (.B(_1464_),
    .C(_1470_),
    .A(_1457_),
    .Y(_1483_),
    .D(_1474_));
 sg13g2_buf_1 _3489_ (.A(_1483_),
    .X(_1484_));
 sg13g2_nand2_1 _3490_ (.Y(_1485_),
    .A(_1482_),
    .B(_1484_));
 sg13g2_buf_8 _3491_ (.A(_1485_),
    .X(_1486_));
 sg13g2_nand2_1 _3492_ (.Y(_1487_),
    .A(net16),
    .B(_1394_));
 sg13g2_inv_1 _3493_ (.Y(_1488_),
    .A(_1394_));
 sg13g2_nand3_1 _3494_ (.B(_1484_),
    .C(_1488_),
    .A(_1482_),
    .Y(_1489_));
 sg13g2_nand2_1 _3495_ (.Y(_1490_),
    .A(_1487_),
    .B(_1489_));
 sg13g2_nand2_1 _3496_ (.Y(_1491_),
    .A(_1481_),
    .B(_1490_));
 sg13g2_nand2_2 _3497_ (.Y(_1492_),
    .A(_1454_),
    .B(_1460_));
 sg13g2_a21oi_1 _3498_ (.A1(_1472_),
    .A2(_1477_),
    .Y(_1493_),
    .B1(_1492_));
 sg13g2_nand2b_1 _3499_ (.Y(_1494_),
    .B(net16),
    .A_N(_1415_));
 sg13g2_nand3_1 _3500_ (.B(_1484_),
    .C(_1415_),
    .A(_1482_),
    .Y(_1495_));
 sg13g2_inv_1 _3501_ (.Y(_1496_),
    .A(_1495_));
 sg13g2_a21oi_1 _3502_ (.A1(_1493_),
    .A2(_1494_),
    .Y(_1497_),
    .B1(_1496_));
 sg13g2_nor2_1 _3503_ (.A(_1491_),
    .B(_1497_),
    .Y(_1498_));
 sg13g2_inv_4 _3504_ (.A(_1479_),
    .Y(_1499_));
 sg13g2_nor2_1 _3505_ (.A(_1461_),
    .B(_1499_),
    .Y(_1500_));
 sg13g2_nand2_1 _3506_ (.Y(_1501_),
    .A(net16),
    .B(_1488_));
 sg13g2_nand3_1 _3507_ (.B(_1484_),
    .C(_1394_),
    .A(_1482_),
    .Y(_1502_));
 sg13g2_inv_1 _3508_ (.Y(_1503_),
    .A(_1502_));
 sg13g2_a21oi_1 _3509_ (.A1(_1500_),
    .A2(_1501_),
    .Y(_1504_),
    .B1(_1503_));
 sg13g2_nor2b_1 _3510_ (.A(_1498_),
    .B_N(_1504_),
    .Y(_1505_));
 sg13g2_nand2_1 _3511_ (.Y(_1506_),
    .A(_1494_),
    .B(_1495_));
 sg13g2_xor2_1 _3512_ (.B(_1479_),
    .A(_1492_),
    .X(_1507_));
 sg13g2_nor2_1 _3513_ (.A(_1506_),
    .B(_1507_),
    .Y(_1508_));
 sg13g2_nand2_1 _3514_ (.Y(_1509_),
    .A(_1501_),
    .B(_1502_));
 sg13g2_inv_1 _3515_ (.Y(_1510_),
    .A(_1461_));
 sg13g2_xnor2_1 _3516_ (.Y(_1511_),
    .A(_1510_),
    .B(_1479_));
 sg13g2_nor2_1 _3517_ (.A(_1509_),
    .B(_1511_),
    .Y(_1512_));
 sg13g2_nor2_1 _3518_ (.A(_1420_),
    .B(_1387_),
    .Y(_1513_));
 sg13g2_nand2b_2 _3519_ (.Y(_1514_),
    .B(net16),
    .A_N(_1513_));
 sg13g2_nand3_1 _3520_ (.B(_1512_),
    .C(_1514_),
    .A(_1508_),
    .Y(_1515_));
 sg13g2_nand2_1 _3521_ (.Y(_1516_),
    .A(_1505_),
    .B(_1515_));
 sg13g2_nand2b_1 _3522_ (.Y(_1517_),
    .B(_1516_),
    .A_N(_1480_));
 sg13g2_nand3_1 _3523_ (.B(_1515_),
    .C(_1480_),
    .A(_1505_),
    .Y(_1518_));
 sg13g2_nand2_1 _3524_ (.Y(_1519_),
    .A(_1517_),
    .B(_1518_));
 sg13g2_nand2_1 _3525_ (.Y(_1520_),
    .A(_1519_),
    .B(_1894_));
 sg13g2_nand3_1 _3526_ (.B(_1518_),
    .C(_1895_),
    .A(_1517_),
    .Y(_1521_));
 sg13g2_nand2_1 _3527_ (.Y(_1522_),
    .A(_1520_),
    .B(_1521_));
 sg13g2_nand2_1 _3528_ (.Y(_1523_),
    .A(_1480_),
    .B(_1490_));
 sg13g2_nand3_1 _3529_ (.B(_1477_),
    .C(_1492_),
    .A(_1472_),
    .Y(_1524_));
 sg13g2_a21oi_1 _3530_ (.A1(_1514_),
    .A2(_1524_),
    .Y(_1525_),
    .B1(_1493_));
 sg13g2_inv_1 _3531_ (.Y(_1526_),
    .A(_1525_));
 sg13g2_nor2_1 _3532_ (.A(_1506_),
    .B(_1511_),
    .Y(_1527_));
 sg13g2_nand3b_1 _3533_ (.B(_1526_),
    .C(_1527_),
    .Y(_1528_),
    .A_N(_1523_));
 sg13g2_nand2_1 _3534_ (.Y(_1529_),
    .A(_1499_),
    .B(_1461_));
 sg13g2_a21oi_1 _3535_ (.A1(_1529_),
    .A2(_1496_),
    .Y(_1530_),
    .B1(_1500_));
 sg13g2_nor2_1 _3536_ (.A(_1523_),
    .B(_1530_),
    .Y(_1531_));
 sg13g2_nand2_1 _3537_ (.Y(_1532_),
    .A(_1499_),
    .B(_1315_));
 sg13g2_nor2_1 _3538_ (.A(_1315_),
    .B(_1499_),
    .Y(_1533_));
 sg13g2_a21oi_1 _3539_ (.A1(_1532_),
    .A2(_1503_),
    .Y(_1534_),
    .B1(_1533_));
 sg13g2_nor2b_1 _3540_ (.A(_1531_),
    .B_N(_1534_),
    .Y(_1535_));
 sg13g2_nand2_1 _3541_ (.Y(_1536_),
    .A(_1528_),
    .B(_1535_));
 sg13g2_inv_1 _3542_ (.Y(_1537_),
    .A(_1471_));
 sg13g2_nand2_1 _3543_ (.Y(_1538_),
    .A(_1536_),
    .B(_1537_));
 sg13g2_nand2_1 _3544_ (.Y(_1539_),
    .A(_1538_),
    .B(_0656_));
 sg13g2_nand3_1 _3545_ (.B(\dither_threshold[6] ),
    .C(_1537_),
    .A(_1536_),
    .Y(_1540_));
 sg13g2_nand2_1 _3546_ (.Y(_1541_),
    .A(_1539_),
    .B(_1540_));
 sg13g2_nor2b_1 _3547_ (.A(_1522_),
    .B_N(_1541_),
    .Y(_1542_));
 sg13g2_nand2_1 _3548_ (.Y(_1543_),
    .A(_1526_),
    .B(_1527_));
 sg13g2_nand2_1 _3549_ (.Y(_1544_),
    .A(_1543_),
    .B(_1530_));
 sg13g2_nand2_1 _3550_ (.Y(_1545_),
    .A(_1544_),
    .B(_1490_));
 sg13g2_nand3_1 _3551_ (.B(_1530_),
    .C(_1509_),
    .A(_1543_),
    .Y(_1546_));
 sg13g2_nand2_1 _3552_ (.Y(_1547_),
    .A(_1545_),
    .B(_1546_));
 sg13g2_nand2_1 _3553_ (.Y(_1548_),
    .A(_1547_),
    .B(_1886_));
 sg13g2_nand3_1 _3554_ (.B(_1546_),
    .C(_1885_),
    .A(_1545_),
    .Y(_1549_));
 sg13g2_xnor2_1 _3555_ (.Y(_1550_),
    .A(_1415_),
    .B(_1486_));
 sg13g2_xnor2_1 _3556_ (.Y(_1551_),
    .A(_1492_),
    .B(_1479_));
 sg13g2_nand3_1 _3557_ (.B(_1551_),
    .C(_1514_),
    .A(_1550_),
    .Y(_1552_));
 sg13g2_nand2_1 _3558_ (.Y(_1553_),
    .A(_1552_),
    .B(_1497_));
 sg13g2_nand2_1 _3559_ (.Y(_1554_),
    .A(_1553_),
    .B(_1481_));
 sg13g2_nand3_1 _3560_ (.B(_1497_),
    .C(_1511_),
    .A(_1552_),
    .Y(_1555_));
 sg13g2_nand2_1 _3561_ (.Y(_1556_),
    .A(_1554_),
    .B(_1555_));
 sg13g2_nor2b_1 _3562_ (.A(_1556_),
    .B_N(_1887_),
    .Y(_1557_));
 sg13g2_nand3_1 _3563_ (.B(_1549_),
    .C(_1557_),
    .A(_1548_),
    .Y(_1558_));
 sg13g2_nand3_1 _3564_ (.B(_1546_),
    .C(_1857_),
    .A(_1545_),
    .Y(_1559_));
 sg13g2_nand2_1 _3565_ (.Y(_1560_),
    .A(_1558_),
    .B(_1559_));
 sg13g2_a21oi_1 _3566_ (.A1(_1517_),
    .A2(_1518_),
    .Y(_1561_),
    .B1(\dither_threshold[5] ));
 sg13g2_nand2_1 _3567_ (.Y(_1562_),
    .A(_1541_),
    .B(_1561_));
 sg13g2_nand3_1 _3568_ (.B(_0656_),
    .C(_1537_),
    .A(_1536_),
    .Y(_1563_));
 sg13g2_nand2_1 _3569_ (.Y(_1564_),
    .A(_1562_),
    .B(_1563_));
 sg13g2_a21oi_1 _3570_ (.A1(_1542_),
    .A2(_1560_),
    .Y(_1565_),
    .B1(_1564_));
 sg13g2_xor2_1 _3571_ (.B(net16),
    .A(_1513_),
    .X(_1566_));
 sg13g2_nor2_1 _3572_ (.A(_1867_),
    .B(_1566_),
    .Y(_1567_));
 sg13g2_xnor2_1 _3573_ (.Y(_1568_),
    .A(_1550_),
    .B(_1525_));
 sg13g2_nand2b_1 _3574_ (.Y(_1569_),
    .B(_1854_),
    .A_N(_1568_));
 sg13g2_xnor2_1 _3575_ (.Y(_1570_),
    .A(_1514_),
    .B(_1551_));
 sg13g2_xnor2_1 _3576_ (.Y(_1571_),
    .A(_0031_),
    .B(_1570_));
 sg13g2_nand2_1 _3577_ (.Y(_1572_),
    .A(_1568_),
    .B(_1874_));
 sg13g2_nand3_1 _3578_ (.B(_1571_),
    .C(_1572_),
    .A(_1569_),
    .Y(_1573_));
 sg13g2_o21ai_1 _3579_ (.B1(_1572_),
    .Y(_1574_),
    .A1(_1851_),
    .A2(_1570_));
 sg13g2_nand2_1 _3580_ (.Y(_1575_),
    .A(_1574_),
    .B(_1569_));
 sg13g2_o21ai_1 _3581_ (.B1(_1575_),
    .Y(_1576_),
    .A1(_1567_),
    .A2(_1573_));
 sg13g2_xnor2_1 _3582_ (.Y(_1577_),
    .A(_1878_),
    .B(_1556_));
 sg13g2_nand2_1 _3583_ (.Y(_1578_),
    .A(_1548_),
    .B(_1549_));
 sg13g2_nor2_1 _3584_ (.A(_1577_),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_nand3_1 _3585_ (.B(_1576_),
    .C(_1579_),
    .A(_1542_),
    .Y(_1580_));
 sg13g2_nand2_1 _3586_ (.Y(_1581_),
    .A(_1565_),
    .B(_1580_));
 sg13g2_nor2_1 _3587_ (.A(_1578_),
    .B(_1522_),
    .Y(_1582_));
 sg13g2_xnor2_1 _3588_ (.Y(_1583_),
    .A(_1850_),
    .B(_1566_));
 sg13g2_nor3_1 _3589_ (.A(_1573_),
    .B(_1583_),
    .C(_1577_),
    .Y(_1584_));
 sg13g2_nand3_1 _3590_ (.B(_1584_),
    .C(_1541_),
    .A(_1582_),
    .Y(_1585_));
 sg13g2_nand3_1 _3591_ (.B(net16),
    .C(_1585_),
    .A(_1581_),
    .Y(_1586_));
 sg13g2_nand2_1 _3592_ (.Y(_1587_),
    .A(_1586_),
    .B(_1499_));
 sg13g2_nand4_1 _3593_ (.B(_1479_),
    .C(net16),
    .A(_1581_),
    .Y(_1588_),
    .D(_1585_));
 sg13g2_nand2_1 _3594_ (.Y(net10),
    .A(_1587_),
    .B(_1588_));
 sg13g2_a21oi_1 _3595_ (.A1(_0721_),
    .A2(_0725_),
    .Y(_1589_),
    .B1(_0614_));
 sg13g2_nor2b_1 _3596_ (.A(_1589_),
    .B_N(_0726_),
    .Y(net12));
 sg13g2_a21oi_1 _3597_ (.A1(_1126_),
    .A2(_1129_),
    .Y(_1590_),
    .B1(_1043_));
 sg13g2_nor2b_1 _3598_ (.A(_1590_),
    .B_N(_1130_),
    .Y(net13));
 sg13g2_a21oi_1 _3599_ (.A1(_1581_),
    .A2(_1585_),
    .Y(_1591_),
    .B1(net16));
 sg13g2_nor2b_1 _3600_ (.A(_1591_),
    .B_N(_1586_),
    .Y(net14));
 sg13g2_buf_1 _3601_ (.A(\counter[10] ),
    .X(_1592_));
 sg13g2_inv_1 _3602_ (.Y(_1593_),
    .A(\counter[5] ));
 sg13g2_inv_1 _3603_ (.Y(_1594_),
    .A(\counter[4] ));
 sg13g2_inv_1 _3604_ (.Y(_1595_),
    .A(\counter[7] ));
 sg13g2_inv_1 _3605_ (.Y(_1596_),
    .A(\counter[6] ));
 sg13g2_nand4_1 _3606_ (.B(_1594_),
    .C(_1595_),
    .A(_1593_),
    .Y(_1597_),
    .D(_1596_));
 sg13g2_nor2_1 _3607_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1598_));
 sg13g2_inv_1 _3608_ (.Y(_1599_),
    .A(\counter[3] ));
 sg13g2_inv_1 _3609_ (.Y(_1600_),
    .A(\counter[2] ));
 sg13g2_nand3_1 _3610_ (.B(_1599_),
    .C(_1600_),
    .A(_1598_),
    .Y(_1601_));
 sg13g2_buf_1 _3611_ (.A(\counter[20] ),
    .X(_1602_));
 sg13g2_buf_1 _3612_ (.A(\counter[22] ),
    .X(_1603_));
 sg13g2_nor4_1 _3613_ (.A(\counter[21] ),
    .B(_1602_),
    .C(\counter[23] ),
    .D(_1603_),
    .Y(_1604_));
 sg13g2_buf_1 _3614_ (.A(\counter[16] ),
    .X(_1605_));
 sg13g2_buf_1 _3615_ (.A(\counter[19] ),
    .X(_1606_));
 sg13g2_buf_1 _3616_ (.A(\counter[18] ),
    .X(_1607_));
 sg13g2_nor4_1 _3617_ (.A(\counter[17] ),
    .B(_1605_),
    .C(_1606_),
    .D(_1607_),
    .Y(_1608_));
 sg13g2_buf_1 _3618_ (.A(\counter[24] ),
    .X(_1609_));
 sg13g2_nor3_1 _3619_ (.A(\counter[25] ),
    .B(_1609_),
    .C(\counter[26] ),
    .Y(_1610_));
 sg13g2_nand3_1 _3620_ (.B(_1608_),
    .C(_1610_),
    .A(_1604_),
    .Y(_1611_));
 sg13g2_nor4_1 _3621_ (.A(_1592_),
    .B(_1597_),
    .C(_1601_),
    .D(_1611_),
    .Y(_1612_));
 sg13g2_buf_1 _3622_ (.A(\counter[13] ),
    .X(_1613_));
 sg13g2_buf_1 _3623_ (.A(\counter[12] ),
    .X(_1614_));
 sg13g2_buf_1 _3624_ (.A(\counter[15] ),
    .X(_1615_));
 sg13g2_buf_1 _3625_ (.A(\counter[14] ),
    .X(_1616_));
 sg13g2_nor4_1 _3626_ (.A(_1613_),
    .B(_1614_),
    .C(_1615_),
    .D(_1616_),
    .Y(_1617_));
 sg13g2_buf_1 _3627_ (.A(\counter[11] ),
    .X(_1618_));
 sg13g2_nor3_1 _3628_ (.A(\counter[9] ),
    .B(\counter[8] ),
    .C(_1618_),
    .Y(_1619_));
 sg13g2_nand3_1 _3629_ (.B(_1617_),
    .C(_1619_),
    .A(_1612_),
    .Y(_0008_));
 sg13g2_buf_1 _3630_ (.A(rst_n),
    .X(_1620_));
 sg13g2_inv_2 _3631_ (.Y(_1621_),
    .A(_1620_));
 sg13g2_inv_1 _3632_ (.Y(_1622_),
    .A(\counter[28] ));
 sg13g2_nand2_1 _3633_ (.Y(_1623_),
    .A(\counter[26] ),
    .B(\counter[27] ));
 sg13g2_nand2_1 _3634_ (.Y(_1624_),
    .A(\counter[21] ),
    .B(_1602_));
 sg13g2_inv_1 _3635_ (.Y(_1625_),
    .A(\counter[17] ));
 sg13g2_inv_1 _3636_ (.Y(_1626_),
    .A(_1605_));
 sg13g2_nand2_1 _3637_ (.Y(_1627_),
    .A(_1606_),
    .B(_1607_));
 sg13g2_nor3_1 _3638_ (.A(_1625_),
    .B(_1626_),
    .C(_1627_),
    .Y(_1628_));
 sg13g2_inv_1 _3639_ (.Y(_1629_),
    .A(_1628_));
 sg13g2_inv_1 _3640_ (.Y(_1630_),
    .A(_1618_));
 sg13g2_inv_1 _3641_ (.Y(_1631_),
    .A(_1592_));
 sg13g2_inv_1 _3642_ (.Y(_1632_),
    .A(\counter[9] ));
 sg13g2_nand2_1 _3643_ (.Y(_1633_),
    .A(\counter[7] ),
    .B(\counter[6] ));
 sg13g2_nand2_1 _3644_ (.Y(_1634_),
    .A(\counter[1] ),
    .B(\counter[0] ));
 sg13g2_nor2_1 _3645_ (.A(_1600_),
    .B(_1634_),
    .Y(_1635_));
 sg13g2_inv_1 _3646_ (.Y(_1636_),
    .A(_1635_));
 sg13g2_nor2_1 _3647_ (.A(_1599_),
    .B(_1636_),
    .Y(_1637_));
 sg13g2_inv_1 _3648_ (.Y(_1638_),
    .A(_1637_));
 sg13g2_nor2_1 _3649_ (.A(_1594_),
    .B(_1638_),
    .Y(_1639_));
 sg13g2_inv_1 _3650_ (.Y(_1640_),
    .A(_1639_));
 sg13g2_nor2_1 _3651_ (.A(_1593_),
    .B(_1640_),
    .Y(_1641_));
 sg13g2_inv_1 _3652_ (.Y(_1642_),
    .A(_1641_));
 sg13g2_nor2_1 _3653_ (.A(_1633_),
    .B(_1642_),
    .Y(_1643_));
 sg13g2_nand2_1 _3654_ (.Y(_1644_),
    .A(_1643_),
    .B(\counter[8] ));
 sg13g2_nor2_1 _3655_ (.A(_1632_),
    .B(_1644_),
    .Y(_1645_));
 sg13g2_inv_1 _3656_ (.Y(_1646_),
    .A(_1645_));
 sg13g2_nor3_1 _3657_ (.A(_1630_),
    .B(_1631_),
    .C(_1646_),
    .Y(_1647_));
 sg13g2_nand2_1 _3658_ (.Y(_1648_),
    .A(_1647_),
    .B(_1614_));
 sg13g2_nor2b_1 _3659_ (.A(_1648_),
    .B_N(_1613_),
    .Y(_1649_));
 sg13g2_nand3_1 _3660_ (.B(_1615_),
    .C(_1616_),
    .A(_1649_),
    .Y(_1650_));
 sg13g2_nor3_2 _3661_ (.A(_1624_),
    .B(_1629_),
    .C(_1650_),
    .Y(_1651_));
 sg13g2_inv_1 _3662_ (.Y(_1652_),
    .A(\counter[25] ));
 sg13g2_inv_1 _3663_ (.Y(_1653_),
    .A(_1609_));
 sg13g2_nand2_1 _3664_ (.Y(_1654_),
    .A(\counter[23] ),
    .B(_1603_));
 sg13g2_nor3_2 _3665_ (.A(_1652_),
    .B(_1653_),
    .C(_1654_),
    .Y(_1655_));
 sg13g2_nand2_1 _3666_ (.Y(_1656_),
    .A(_1651_),
    .B(_1655_));
 sg13g2_nor3_1 _3667_ (.A(_1622_),
    .B(_1623_),
    .C(_1656_),
    .Y(_1657_));
 sg13g2_nor2_1 _3668_ (.A(\counter[29] ),
    .B(_1657_),
    .Y(_1658_));
 sg13g2_nand2_1 _3669_ (.Y(_1659_),
    .A(_1657_),
    .B(\counter[29] ));
 sg13g2_inv_1 _3670_ (.Y(_1660_),
    .A(_1659_));
 sg13g2_nor3_2 _3671_ (.A(_1621_),
    .B(_1658_),
    .C(_1660_),
    .Y(_0079_));
 sg13g2_inv_1 _3672_ (.Y(_1661_),
    .A(\counter[8] ));
 sg13g2_nand2_1 _3673_ (.Y(_1662_),
    .A(_1618_),
    .B(_1592_));
 sg13g2_nor4_1 _3674_ (.A(_1632_),
    .B(_1661_),
    .C(_1633_),
    .D(_1662_),
    .Y(_1663_));
 sg13g2_nand4_1 _3675_ (.B(_1663_),
    .C(_1613_),
    .A(_1641_),
    .Y(_1664_),
    .D(_1614_));
 sg13g2_nand3b_1 _3676_ (.B(_1615_),
    .C(_1616_),
    .Y(_1665_),
    .A_N(_1664_));
 sg13g2_nor4_1 _3677_ (.A(_1624_),
    .B(_1623_),
    .C(_1629_),
    .D(_1665_),
    .Y(_1666_));
 sg13g2_nand2_1 _3678_ (.Y(_1667_),
    .A(_1666_),
    .B(_1655_));
 sg13g2_nand3_1 _3679_ (.B(\counter[28] ),
    .C(_1655_),
    .A(_1666_),
    .Y(_1668_));
 sg13g2_buf_1 _3680_ (.A(_1620_),
    .X(_1669_));
 sg13g2_nand2_1 _3681_ (.Y(_1670_),
    .A(_1668_),
    .B(net73));
 sg13g2_a21oi_1 _3682_ (.A1(_1622_),
    .A2(_1667_),
    .Y(_0078_),
    .B1(_1670_));
 sg13g2_nand4_1 _3683_ (.B(\counter[25] ),
    .C(_1609_),
    .A(\counter[23] ),
    .Y(_1671_),
    .D(\counter[26] ));
 sg13g2_nand4_1 _3684_ (.B(_1613_),
    .C(_1614_),
    .A(_1618_),
    .Y(_1672_),
    .D(_1616_));
 sg13g2_nand4_1 _3685_ (.B(\counter[17] ),
    .C(_1605_),
    .A(_1615_),
    .Y(_1673_),
    .D(_1607_));
 sg13g2_nand4_1 _3686_ (.B(\counter[21] ),
    .C(_1602_),
    .A(_1606_),
    .Y(_1674_),
    .D(_1603_));
 sg13g2_nor4_1 _3687_ (.A(_1671_),
    .B(_1672_),
    .C(_1673_),
    .D(_1674_),
    .Y(_1675_));
 sg13g2_nor4_1 _3688_ (.A(_1599_),
    .B(_1593_),
    .C(_1594_),
    .D(_1596_),
    .Y(_1676_));
 sg13g2_nor4_1 _3689_ (.A(_1595_),
    .B(_1632_),
    .C(_1661_),
    .D(_1631_),
    .Y(_1677_));
 sg13g2_nand4_1 _3690_ (.B(_1635_),
    .C(_1676_),
    .A(_1675_),
    .Y(_1678_),
    .D(_1677_));
 sg13g2_xor2_1 _3691_ (.B(_1678_),
    .A(\counter[27] ),
    .X(_1679_));
 sg13g2_nor2_1 _3692_ (.A(_1621_),
    .B(_1679_),
    .Y(_0077_));
 sg13g2_inv_1 _3693_ (.Y(_1680_),
    .A(_0077_));
 sg13g2_nand2_1 _3694_ (.Y(_1681_),
    .A(_0078_),
    .B(_1680_));
 sg13g2_nor2_1 _3695_ (.A(_1680_),
    .B(_0078_),
    .Y(_1682_));
 sg13g2_a21oi_1 _3696_ (.A1(_0079_),
    .A2(_1681_),
    .Y(_0000_),
    .B1(_1682_));
 sg13g2_inv_1 _3697_ (.Y(_1683_),
    .A(_0079_));
 sg13g2_o21ai_1 _3698_ (.B1(_1681_),
    .Y(_0001_),
    .A1(_1682_),
    .A2(_1683_));
 sg13g2_a21o_1 _3699_ (.A2(_0078_),
    .A1(_0079_),
    .B1(_0077_),
    .X(_0002_));
 sg13g2_buf_1 _3700_ (.A(\i_project.controller_0.rst_n ),
    .X(_1684_));
 sg13g2_buf_1 _3701_ (.A(_1684_),
    .X(_1685_));
 sg13g2_buf_1 _3702_ (.A(\i_project.controller_0.divider[0] ),
    .X(_1686_));
 sg13g2_inv_1 _3703_ (.Y(_1687_),
    .A(_1686_));
 sg13g2_nor2_1 _3704_ (.A(net62),
    .B(\i_project.controller_0.grey_pass[10] ),
    .Y(_1688_));
 sg13g2_a21oi_1 _3705_ (.A1(net62),
    .A2(_1687_),
    .Y(_0003_),
    .B1(_1688_));
 sg13g2_buf_2 _3706_ (.A(\i_project.controller_0.divider[1] ),
    .X(_1689_));
 sg13g2_inv_1 _3707_ (.Y(_1690_),
    .A(_1689_));
 sg13g2_buf_1 _3708_ (.A(_1690_),
    .X(_1691_));
 sg13g2_nor2_1 _3709_ (.A(net62),
    .B(\i_project.controller_0.grey_pass[11] ),
    .Y(_1692_));
 sg13g2_a21oi_1 _3710_ (.A1(net62),
    .A2(_1691_),
    .Y(_0004_),
    .B1(_1692_));
 sg13g2_buf_1 _3711_ (.A(ui_in[7]),
    .X(_1693_));
 sg13g2_mux2_1 _3712_ (.A0(_0012_),
    .A1(net1),
    .S(net74),
    .X(_0009_));
 sg13g2_mux2_1 _3713_ (.A0(_0013_),
    .A1(net2),
    .S(net74),
    .X(_0010_));
 sg13g2_mux2_1 _3714_ (.A0(_0014_),
    .A1(net3),
    .S(net74),
    .X(_0011_));
 sg13g2_nand2_1 _3715_ (.Y(_1694_),
    .A(net74),
    .B(net5));
 sg13g2_o21ai_1 _3716_ (.B1(_1694_),
    .Y(_0005_),
    .A1(net74),
    .A2(_1653_));
 sg13g2_nand2_1 _3717_ (.Y(_1695_),
    .A(net74),
    .B(net6));
 sg13g2_o21ai_1 _3718_ (.B1(_1695_),
    .Y(_0006_),
    .A1(net74),
    .A2(_1652_));
 sg13g2_inv_1 _3719_ (.Y(_1696_),
    .A(\counter[26] ));
 sg13g2_nand2_1 _3720_ (.Y(_1697_),
    .A(_1693_),
    .B(net7));
 sg13g2_o21ai_1 _3721_ (.B1(_1697_),
    .Y(_0007_),
    .A1(_1693_),
    .A2(_1696_));
 sg13g2_buf_1 _3722_ (.A(\i_project.controller_0.h[9] ),
    .X(_1698_));
 sg13g2_buf_2 _3723_ (.A(\i_project.controller_0.h[8] ),
    .X(_1699_));
 sg13g2_inv_1 _3724_ (.Y(_1700_),
    .A(_1699_));
 sg13g2_nor2_1 _3725_ (.A(_1698_),
    .B(_1700_),
    .Y(_1701_));
 sg13g2_inv_1 _3726_ (.Y(_1702_),
    .A(_1701_));
 sg13g2_buf_1 _3727_ (.A(\i_project.controller_0.h[6] ),
    .X(_1703_));
 sg13g2_inv_1 _3728_ (.Y(_1704_),
    .A(\i_project.controller_0.h[7] ));
 sg13g2_nor2_1 _3729_ (.A(net72),
    .B(_1704_),
    .Y(_1705_));
 sg13g2_buf_1 _3730_ (.A(\i_project.controller_0.h[4] ),
    .X(_1706_));
 sg13g2_buf_1 _3731_ (.A(_1706_),
    .X(_1707_));
 sg13g2_buf_1 _3732_ (.A(\i_project.controller_0.h[5] ),
    .X(_1708_));
 sg13g2_inv_1 _3733_ (.Y(_1709_),
    .A(_1708_));
 sg13g2_nor2_1 _3734_ (.A(net61),
    .B(_1709_),
    .Y(_1710_));
 sg13g2_nand2_1 _3735_ (.Y(_1711_),
    .A(_1705_),
    .B(_1710_));
 sg13g2_buf_1 _3736_ (.A(\i_project.controller_0.h[0] ),
    .X(_1712_));
 sg13g2_buf_1 _3737_ (.A(_1712_),
    .X(_1713_));
 sg13g2_buf_1 _3738_ (.A(\i_project.controller_0.h[1] ),
    .X(_1714_));
 sg13g2_inv_1 _3739_ (.Y(_1715_),
    .A(net71));
 sg13g2_nor2_1 _3740_ (.A(net60),
    .B(_1715_),
    .Y(_1716_));
 sg13g2_buf_1 _3741_ (.A(\i_project.controller_0.h[3] ),
    .X(_1717_));
 sg13g2_inv_1 _3742_ (.Y(_1718_),
    .A(_1717_));
 sg13g2_buf_1 _3743_ (.A(\i_project.controller_0.h[2] ),
    .X(_1719_));
 sg13g2_inv_2 _3744_ (.Y(_1720_),
    .A(_1719_));
 sg13g2_nand3_1 _3745_ (.B(_1718_),
    .C(_1720_),
    .A(_1716_),
    .Y(_1721_));
 sg13g2_nor4_1 _3746_ (.A(_0022_),
    .B(_1702_),
    .C(_1711_),
    .D(_1721_),
    .Y(_1722_));
 sg13g2_nor2_2 _3747_ (.A(_1684_),
    .B(net73),
    .Y(_1723_));
 sg13g2_buf_1 _3748_ (.A(_1717_),
    .X(_1724_));
 sg13g2_buf_1 _3749_ (.A(_1719_),
    .X(_1725_));
 sg13g2_nor2_1 _3750_ (.A(_1714_),
    .B(net60),
    .Y(_1726_));
 sg13g2_inv_1 _3751_ (.Y(_1727_),
    .A(_1726_));
 sg13g2_nor3_1 _3752_ (.A(net59),
    .B(net58),
    .C(_1727_),
    .Y(_1728_));
 sg13g2_inv_1 _3753_ (.Y(_1729_),
    .A(_1698_));
 sg13g2_nor2_1 _3754_ (.A(_1699_),
    .B(_1729_),
    .Y(_1730_));
 sg13g2_and3_1 _3755_ (.X(_1731_),
    .A(_1728_),
    .B(_0022_),
    .C(_1730_));
 sg13g2_inv_2 _3756_ (.Y(_1732_),
    .A(net72));
 sg13g2_buf_1 _3757_ (.A(_1708_),
    .X(_1733_));
 sg13g2_nand2_1 _3758_ (.Y(_1734_),
    .A(net57),
    .B(net61));
 sg13g2_nor3_1 _3759_ (.A(_1732_),
    .B(_1704_),
    .C(_1734_),
    .Y(_1735_));
 sg13g2_and2_1 _3760_ (.A(_1731_),
    .B(_1735_),
    .X(_1736_));
 sg13g2_buf_1 _3761_ (.A(\i_project.controller_0.h[7] ),
    .X(_1737_));
 sg13g2_nor3_1 _3762_ (.A(_1732_),
    .B(net70),
    .C(_1734_),
    .Y(_1738_));
 sg13g2_nand2_1 _3763_ (.Y(_1739_),
    .A(_1724_),
    .B(net58));
 sg13g2_nor4_1 _3764_ (.A(_0022_),
    .B(_1739_),
    .C(_1727_),
    .D(_1702_),
    .Y(_1740_));
 sg13g2_inv_1 _3765_ (.Y(_1741_),
    .A(_1705_));
 sg13g2_inv_1 _3766_ (.Y(_1742_),
    .A(_1706_));
 sg13g2_nor2_1 _3767_ (.A(net57),
    .B(_1742_),
    .Y(_1743_));
 sg13g2_inv_1 _3768_ (.Y(_1744_),
    .A(_1743_));
 sg13g2_nor2_1 _3769_ (.A(_1741_),
    .B(_1744_),
    .Y(_1745_));
 sg13g2_a221oi_1 _3770_ (.B2(_1745_),
    .C1(\i_project.controller_0.vga_sync.hsync ),
    .B1(_1731_),
    .A1(_1738_),
    .Y(_1746_),
    .A2(_1740_));
 sg13g2_nor4_1 _3771_ (.A(_1722_),
    .B(_1723_),
    .C(_1736_),
    .D(_1746_),
    .Y(_0123_));
 sg13g2_buf_1 _3772_ (.A(\i_project.controller_0.v[7] ),
    .X(_1747_));
 sg13g2_buf_1 _3773_ (.A(\i_project.controller_0.v[6] ),
    .X(_1748_));
 sg13g2_nand2_1 _3774_ (.Y(_1749_),
    .A(_1747_),
    .B(net69));
 sg13g2_buf_8 _3775_ (.A(\i_project.controller_0.v[4] ),
    .X(_1750_));
 sg13g2_buf_2 _3776_ (.A(\i_project.controller_0.v[5] ),
    .X(_1751_));
 sg13g2_inv_1 _3777_ (.Y(_1752_),
    .A(_1751_));
 sg13g2_nor2_1 _3778_ (.A(_1750_),
    .B(_1752_),
    .Y(_1753_));
 sg13g2_buf_2 _3779_ (.A(\i_project.controller_0.v[8] ),
    .X(_1754_));
 sg13g2_buf_1 _3780_ (.A(\i_project.controller_0.v[9] ),
    .X(_1755_));
 sg13g2_inv_1 _3781_ (.Y(_1756_),
    .A(_1755_));
 sg13g2_nand3_1 _3782_ (.B(_1754_),
    .C(_1756_),
    .A(_1753_),
    .Y(_1757_));
 sg13g2_nor2_1 _3783_ (.A(_1749_),
    .B(_1757_),
    .Y(_1758_));
 sg13g2_inv_1 _3784_ (.Y(_1759_),
    .A(_1758_));
 sg13g2_buf_8 _3785_ (.A(\i_project.controller_0.v[2] ),
    .X(_1760_));
 sg13g2_buf_8 _3786_ (.A(\i_project.controller_0.v[3] ),
    .X(_1761_));
 sg13g2_inv_1 _3787_ (.Y(_1762_),
    .A(_1761_));
 sg13g2_nor2_1 _3788_ (.A(_1760_),
    .B(_1762_),
    .Y(_1763_));
 sg13g2_buf_1 _3789_ (.A(\i_project.controller_0.vga_sync.mode ),
    .X(_1764_));
 sg13g2_inv_1 _3790_ (.Y(_1765_),
    .A(net68));
 sg13g2_buf_8 _3791_ (.A(\i_project.controller_0.v[0] ),
    .X(_1766_));
 sg13g2_inv_1 _3792_ (.Y(_1767_),
    .A(_1766_));
 sg13g2_buf_8 _3793_ (.A(\i_project.controller_0.v[1] ),
    .X(_1768_));
 sg13g2_nand4_1 _3794_ (.B(_1765_),
    .C(_1767_),
    .A(_1763_),
    .Y(_1769_),
    .D(net67));
 sg13g2_inv_1 _3795_ (.Y(_1770_),
    .A(_1747_));
 sg13g2_nor2_1 _3796_ (.A(net69),
    .B(_1770_),
    .Y(_1771_));
 sg13g2_inv_1 _3797_ (.Y(_1772_),
    .A(_1771_));
 sg13g2_nor2_1 _3798_ (.A(_1750_),
    .B(_1751_),
    .Y(_1773_));
 sg13g2_inv_1 _3799_ (.Y(_1774_),
    .A(_1773_));
 sg13g2_inv_2 _3800_ (.Y(_1775_),
    .A(_1760_));
 sg13g2_nand2_1 _3801_ (.Y(_1776_),
    .A(_1754_),
    .B(_1755_));
 sg13g2_nor3_1 _3802_ (.A(_1775_),
    .B(_1761_),
    .C(_1776_),
    .Y(_1777_));
 sg13g2_inv_1 _3803_ (.Y(_1778_),
    .A(net67));
 sg13g2_nand4_1 _3804_ (.B(net68),
    .C(_1766_),
    .A(_1777_),
    .Y(_1779_),
    .D(_1778_));
 sg13g2_nor3_1 _3805_ (.A(_1772_),
    .B(_1774_),
    .C(_1779_),
    .Y(_1780_));
 sg13g2_nor2_1 _3806_ (.A(\i_project.controller_0.vga_sync.vsync ),
    .B(_1780_),
    .Y(_1781_));
 sg13g2_o21ai_1 _3807_ (.B1(_1781_),
    .Y(_1782_),
    .A1(_1759_),
    .A2(_1769_));
 sg13g2_nand2_1 _3808_ (.Y(_1783_),
    .A(net68),
    .B(_1754_));
 sg13g2_inv_1 _3809_ (.Y(_1784_),
    .A(_1763_));
 sg13g2_nor3_1 _3810_ (.A(_1756_),
    .B(_1783_),
    .C(_1784_),
    .Y(_1785_));
 sg13g2_nor2_1 _3811_ (.A(_1766_),
    .B(net67),
    .Y(_1786_));
 sg13g2_nand4_1 _3812_ (.B(_1786_),
    .C(_1771_),
    .A(_1785_),
    .Y(_1787_),
    .D(_1773_));
 sg13g2_nand2_1 _3813_ (.Y(_1788_),
    .A(_1760_),
    .B(_1761_));
 sg13g2_inv_1 _3814_ (.Y(_1789_),
    .A(_1786_));
 sg13g2_nor3_1 _3815_ (.A(net68),
    .B(_1788_),
    .C(_1789_),
    .Y(_1790_));
 sg13g2_a21oi_1 _3816_ (.A1(_1758_),
    .A2(_1790_),
    .Y(_1791_),
    .B1(_1723_));
 sg13g2_and3_1 _3817_ (.X(_0134_),
    .A(_1782_),
    .B(_1787_),
    .C(_1791_));
 sg13g2_inv_1 _3818_ (.Y(_1792_),
    .A(\i_project.controller_0.voffset[0] ));
 sg13g2_nor3_1 _3819_ (.A(net57),
    .B(net61),
    .C(_1741_),
    .Y(_1793_));
 sg13g2_nand2_1 _3820_ (.Y(_1794_),
    .A(_1700_),
    .B(_0023_));
 sg13g2_a21oi_1 _3821_ (.A1(_1793_),
    .A2(_1728_),
    .Y(_1795_),
    .B1(_1794_));
 sg13g2_inv_1 _3822_ (.Y(_1796_),
    .A(_1795_));
 sg13g2_nor2_1 _3823_ (.A(net68),
    .B(_1729_),
    .Y(_1797_));
 sg13g2_nor2_1 _3824_ (.A(net72),
    .B(net70),
    .Y(_1798_));
 sg13g2_nor3_1 _3825_ (.A(_1732_),
    .B(net70),
    .C(_1702_),
    .Y(_1799_));
 sg13g2_inv_1 _3826_ (.Y(_1800_),
    .A(_0024_));
 sg13g2_o21ai_1 _3827_ (.B1(_1733_),
    .Y(_1801_),
    .A1(_1707_),
    .A2(_1800_));
 sg13g2_nor2_1 _3828_ (.A(_1698_),
    .B(_1699_),
    .Y(_1802_));
 sg13g2_a221oi_1 _3829_ (.B2(_1801_),
    .C1(_1802_),
    .B1(_1799_),
    .A1(_1701_),
    .Y(_1803_),
    .A2(_1798_));
 sg13g2_nor2_1 _3830_ (.A(_1725_),
    .B(_1718_),
    .Y(_1804_));
 sg13g2_nand4_1 _3831_ (.B(_1710_),
    .C(_1726_),
    .A(_1799_),
    .Y(_1805_),
    .D(_1804_));
 sg13g2_nand2b_1 _3832_ (.Y(_1806_),
    .B(_1805_),
    .A_N(_1803_));
 sg13g2_a22oi_1 _3833_ (.Y(_1807_),
    .B1(net68),
    .B2(_1806_),
    .A2(_1797_),
    .A1(_1796_));
 sg13g2_xor2_1 _3834_ (.B(\i_project.controller_0.mode[2] ),
    .A(\i_project.controller_0.grey_pass[14] ),
    .X(_1808_));
 sg13g2_buf_2 _3835_ (.A(\i_project.controller_0.mode[1] ),
    .X(_1809_));
 sg13g2_xor2_1 _3836_ (.B(\i_project.controller_0.grey_pass[13] ),
    .A(_1809_),
    .X(_1810_));
 sg13g2_nor2_1 _3837_ (.A(_1808_),
    .B(_1810_),
    .Y(_1811_));
 sg13g2_buf_2 _3838_ (.A(\i_project.controller_0.mode[0] ),
    .X(_1812_));
 sg13g2_xnor2_1 _3839_ (.Y(_1813_),
    .A(_1812_),
    .B(\i_project.controller_0.grey_pass[12] ));
 sg13g2_inv_1 _3840_ (.Y(_1814_),
    .A(_0025_));
 sg13g2_nor3_2 _3841_ (.A(_1809_),
    .B(_1812_),
    .C(_1814_),
    .Y(_1815_));
 sg13g2_buf_1 _3842_ (.A(_1815_),
    .X(_1816_));
 sg13g2_a21oi_1 _3843_ (.A1(_1811_),
    .A2(_1813_),
    .Y(_1817_),
    .B1(_1816_));
 sg13g2_nand2b_1 _3844_ (.Y(_1818_),
    .B(_1817_),
    .A_N(_1807_));
 sg13g2_nand2_2 _3845_ (.Y(_1819_),
    .A(_1818_),
    .B(_1684_));
 sg13g2_inv_2 _3846_ (.Y(_1820_),
    .A(_1819_));
 sg13g2_nand2b_1 _3847_ (.Y(_1821_),
    .B(net62),
    .A_N(_1813_));
 sg13g2_inv_1 _3848_ (.Y(_1822_),
    .A(\i_project.controller_0.mode[2] ));
 sg13g2_nor3_1 _3849_ (.A(_1809_),
    .B(_1684_),
    .C(_1822_),
    .Y(_1823_));
 sg13g2_nand2_1 _3850_ (.Y(_1824_),
    .A(_1823_),
    .B(_0016_));
 sg13g2_nor2b_2 _3851_ (.A(_1820_),
    .B_N(_1824_),
    .Y(_1825_));
 sg13g2_a22oi_1 _3852_ (.Y(_0135_),
    .B1(_1821_),
    .B2(_1825_),
    .A2(_1820_),
    .A1(_1792_));
 sg13g2_a22oi_1 _3853_ (.Y(_1826_),
    .B1(_1685_),
    .B2(_1810_),
    .A2(_0015_),
    .A1(_1823_));
 sg13g2_buf_2 _3854_ (.A(\i_project.controller_0.voffset[1] ),
    .X(_1827_));
 sg13g2_nor2_1 _3855_ (.A(_1827_),
    .B(_1819_),
    .Y(_1828_));
 sg13g2_a21oi_1 _3856_ (.A1(_1819_),
    .A2(_1826_),
    .Y(_0136_),
    .B1(_1828_));
 sg13g2_buf_1 _3857_ (.A(\i_project.controller_0.voffset[2] ),
    .X(_1829_));
 sg13g2_inv_2 _3858_ (.Y(_1830_),
    .A(_1829_));
 sg13g2_nand2_1 _3859_ (.Y(_1831_),
    .A(_1808_),
    .B(net62));
 sg13g2_a22oi_1 _3860_ (.Y(_0137_),
    .B1(_1831_),
    .B2(_1825_),
    .A2(_1820_),
    .A1(_1830_));
 sg13g2_inv_1 _3861_ (.Y(_1832_),
    .A(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _3862_ (.Y(_1833_),
    .A(_1823_),
    .B(_0145_));
 sg13g2_o21ai_1 _3863_ (.B1(_1833_),
    .Y(_0138_),
    .A1(_1832_),
    .A2(_1819_));
 sg13g2_inv_1 _3864_ (.Y(_1834_),
    .A(\i_project.controller_0.voffset[4] ));
 sg13g2_o21ai_1 _3865_ (.B1(_1824_),
    .Y(_0139_),
    .A1(_1834_),
    .A2(_1819_));
 sg13g2_inv_1 _3866_ (.Y(_1835_),
    .A(\i_project.controller_0.voffset[5] ));
 sg13g2_buf_1 _3867_ (.A(net62),
    .X(_1836_));
 sg13g2_nand2_1 _3868_ (.Y(_1837_),
    .A(net48),
    .B(\i_project.controller_0.grey_pass[10] ));
 sg13g2_a22oi_1 _3869_ (.Y(_0140_),
    .B1(_1837_),
    .B2(_1825_),
    .A2(_1820_),
    .A1(_1835_));
 sg13g2_inv_1 _3870_ (.Y(_1838_),
    .A(\i_project.controller_0.voffset[6] ));
 sg13g2_nand2_1 _3871_ (.Y(_1839_),
    .A(net48),
    .B(\i_project.controller_0.grey_pass[11] ));
 sg13g2_a22oi_1 _3872_ (.Y(_0141_),
    .B1(_1839_),
    .B2(_1825_),
    .A2(_1820_),
    .A1(_1838_));
 sg13g2_inv_1 _3873_ (.Y(_1840_),
    .A(net62));
 sg13g2_inv_1 _3874_ (.Y(_1841_),
    .A(\i_project.controller_0.grey_pass[15] ));
 sg13g2_nor3_1 _3875_ (.A(_1840_),
    .B(_1841_),
    .C(_1818_),
    .Y(_1842_));
 sg13g2_a21o_1 _3876_ (.A2(_1820_),
    .A1(\i_project.controller_0.voffset[7] ),
    .B1(_1842_),
    .X(_0142_));
 sg13g2_inv_1 _3877_ (.Y(_1843_),
    .A(_1812_));
 sg13g2_nor2_1 _3878_ (.A(\i_project.controller_0.grey_pass[12] ),
    .B(net48),
    .Y(_1844_));
 sg13g2_a21oi_1 _3879_ (.A1(_1843_),
    .A2(net48),
    .Y(_0097_),
    .B1(_1844_));
 sg13g2_inv_1 _3880_ (.Y(_1845_),
    .A(_1809_));
 sg13g2_nor2_1 _3881_ (.A(\i_project.controller_0.grey_pass[13] ),
    .B(net48),
    .Y(_1846_));
 sg13g2_a21oi_1 _3882_ (.A1(_1845_),
    .A2(net48),
    .Y(_0098_),
    .B1(_1846_));
 sg13g2_nor2_1 _3883_ (.A(\i_project.controller_0.grey_pass[14] ),
    .B(_1836_),
    .Y(_1847_));
 sg13g2_a21oi_1 _3884_ (.A1(_1822_),
    .A2(_1836_),
    .Y(_0099_),
    .B1(_1847_));
 sg13g2_nand2_1 _3885_ (.Y(_1848_),
    .A(net68),
    .B(net48));
 sg13g2_o21ai_1 _3886_ (.B1(_1848_),
    .Y(_0100_),
    .A1(net48),
    .A2(_1841_));
 sg13g2_buf_1 _3887_ (.A(\dither_threshold[0] ),
    .X(_1849_));
 sg13g2_buf_2 _3888_ (.A(_0026_),
    .X(_1850_));
 sg13g2_buf_1 _3889_ (.A(\dither_threshold[1] ),
    .X(_1851_));
 sg13g2_inv_1 _3890_ (.Y(_1852_),
    .A(_1851_));
 sg13g2_a21oi_1 _3891_ (.A1(_1849_),
    .A2(_1850_),
    .Y(_1853_),
    .B1(_1852_));
 sg13g2_buf_1 _3892_ (.A(\dither_threshold[2] ),
    .X(_1854_));
 sg13g2_nor2_1 _3893_ (.A(\dither_threshold[3] ),
    .B(_1854_),
    .Y(_1855_));
 sg13g2_inv_1 _3894_ (.Y(_1856_),
    .A(\dither_threshold[5] ));
 sg13g2_inv_1 _3895_ (.Y(_1857_),
    .A(\dither_threshold[4] ));
 sg13g2_nand3_1 _3896_ (.B(_1856_),
    .C(_1857_),
    .A(_1855_),
    .Y(_1858_));
 sg13g2_o21ai_1 _3897_ (.B1(\dither_threshold[6] ),
    .Y(_1859_),
    .A1(_1853_),
    .A2(_1858_));
 sg13g2_buf_1 _3898_ (.A(_1859_),
    .X(_1860_));
 sg13g2_nor2_1 _3899_ (.A(_1849_),
    .B(_1860_),
    .Y(_1861_));
 sg13g2_xnor2_1 _3900_ (.Y(\i_project.controller_0.vga_sync.o_vsync ),
    .A(_1764_),
    .B(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_inv_1 _3901_ (.Y(_1862_),
    .A(\i_project.controller_0.vga_sync.o_vsync ));
 sg13g2_nand3_1 _3902_ (.B(_1841_),
    .C(prev_vsync),
    .A(_1862_),
    .Y(_1863_));
 sg13g2_nand3b_1 _3903_ (.B(\i_project.controller_0.vga_sync.o_vsync ),
    .C(\i_project.controller_0.grey_pass[15] ),
    .Y(_1864_),
    .A_N(prev_vsync));
 sg13g2_nand3_1 _3904_ (.B(_1864_),
    .C(_1669_),
    .A(_1863_),
    .Y(_1865_));
 sg13g2_buf_1 _3905_ (.A(_1865_),
    .X(_1866_));
 sg13g2_inv_1 _3906_ (.Y(_1867_),
    .A(_1849_));
 sg13g2_inv_2 _3907_ (.Y(_1868_),
    .A(_1860_));
 sg13g2_nor2_1 _3908_ (.A(_1867_),
    .B(_1868_),
    .Y(_1869_));
 sg13g2_nor3_1 _3909_ (.A(_1861_),
    .B(_1866_),
    .C(_1869_),
    .Y(_0090_));
 sg13g2_inv_1 _3910_ (.Y(_1870_),
    .A(_0031_));
 sg13g2_nor2_1 _3911_ (.A(_1851_),
    .B(_1849_),
    .Y(_1871_));
 sg13g2_nor2_1 _3912_ (.A(_1871_),
    .B(_1868_),
    .Y(_1872_));
 sg13g2_nand2_1 _3913_ (.Y(_1873_),
    .A(_1851_),
    .B(_1849_));
 sg13g2_a221oi_1 _3914_ (.B2(_1873_),
    .C1(_1866_),
    .B1(_1872_),
    .A1(_1870_),
    .Y(_0091_),
    .A2(_1868_));
 sg13g2_inv_2 _3915_ (.Y(_1874_),
    .A(_1854_));
 sg13g2_a21oi_1 _3916_ (.A1(_1852_),
    .A2(_1868_),
    .Y(_1875_),
    .B1(_1872_));
 sg13g2_inv_1 _3917_ (.Y(_1876_),
    .A(_1866_));
 sg13g2_o21ai_1 _3918_ (.B1(_1876_),
    .Y(_1877_),
    .A1(_1874_),
    .A2(_1875_));
 sg13g2_a21oi_1 _3919_ (.A1(_1874_),
    .A2(_1875_),
    .Y(_0092_),
    .B1(_1877_));
 sg13g2_inv_2 _3920_ (.Y(_1878_),
    .A(_0032_));
 sg13g2_a21oi_1 _3921_ (.A1(_1852_),
    .A2(_1850_),
    .Y(_1879_),
    .B1(_1874_));
 sg13g2_xnor2_1 _3922_ (.Y(_1880_),
    .A(_1878_),
    .B(_1879_));
 sg13g2_o21ai_1 _3923_ (.B1(\dither_threshold[3] ),
    .Y(_1881_),
    .A1(_1851_),
    .A2(_1854_));
 sg13g2_nand2_1 _3924_ (.Y(_1882_),
    .A(_1855_),
    .B(_1852_));
 sg13g2_nand2_1 _3925_ (.Y(_1883_),
    .A(_1881_),
    .B(_1882_));
 sg13g2_o21ai_1 _3926_ (.B1(_1876_),
    .Y(_1884_),
    .A1(_1860_),
    .A2(_1883_));
 sg13g2_a21oi_1 _3927_ (.A1(_1860_),
    .A2(_1880_),
    .Y(_0093_),
    .B1(_1884_));
 sg13g2_buf_1 _3928_ (.A(_0033_),
    .X(_1885_));
 sg13g2_inv_1 _3929_ (.Y(_1886_),
    .A(_1885_));
 sg13g2_inv_1 _3930_ (.Y(_1887_),
    .A(\dither_threshold[3] ));
 sg13g2_nor3_1 _3931_ (.A(_1887_),
    .B(_1874_),
    .C(_1871_),
    .Y(_1888_));
 sg13g2_xnor2_1 _3932_ (.Y(_1889_),
    .A(_1886_),
    .B(_1888_));
 sg13g2_nand3_1 _3933_ (.B(_1852_),
    .C(_1857_),
    .A(_1855_),
    .Y(_1890_));
 sg13g2_nand2_1 _3934_ (.Y(_1891_),
    .A(_1882_),
    .B(\dither_threshold[4] ));
 sg13g2_a21oi_1 _3935_ (.A1(_1890_),
    .A2(_1891_),
    .Y(_1892_),
    .B1(_1860_));
 sg13g2_a21oi_1 _3936_ (.A1(_1860_),
    .A2(_1889_),
    .Y(_1893_),
    .B1(_1892_));
 sg13g2_nor2_1 _3937_ (.A(_1866_),
    .B(_1893_),
    .Y(_0094_));
 sg13g2_buf_1 _3938_ (.A(_0034_),
    .X(_1894_));
 sg13g2_inv_1 _3939_ (.Y(_1895_),
    .A(_1894_));
 sg13g2_inv_1 _3940_ (.Y(_1896_),
    .A(_1888_));
 sg13g2_o21ai_1 _3941_ (.B1(_1885_),
    .Y(_1897_),
    .A1(\dither_threshold[4] ),
    .A2(_1896_));
 sg13g2_a21oi_1 _3942_ (.A1(_1897_),
    .A2(_1895_),
    .Y(_1898_),
    .B1(_1868_));
 sg13g2_o21ai_1 _3943_ (.B1(_1898_),
    .Y(_1899_),
    .A1(_1895_),
    .A2(_1897_));
 sg13g2_nand3_1 _3944_ (.B(\dither_threshold[5] ),
    .C(_1890_),
    .A(_1868_),
    .Y(_1900_));
 sg13g2_a21oi_1 _3945_ (.A1(_1899_),
    .A2(_1900_),
    .Y(_0095_),
    .B1(_1866_));
 sg13g2_buf_1 _3946_ (.A(_0035_),
    .X(_1901_));
 sg13g2_a21oi_1 _3947_ (.A1(_1896_),
    .A2(_1857_),
    .Y(_1902_),
    .B1(_1856_));
 sg13g2_nor2_1 _3948_ (.A(_1902_),
    .B(_1868_),
    .Y(_1903_));
 sg13g2_o21ai_1 _3949_ (.B1(_1876_),
    .Y(_1904_),
    .A1(_1901_),
    .A2(_1903_));
 sg13g2_a21oi_1 _3950_ (.A1(_1901_),
    .A2(_1903_),
    .Y(_0096_),
    .B1(_1904_));
 sg13g2_inv_1 _3951_ (.Y(_1905_),
    .A(_0054_));
 sg13g2_nand2_1 _3952_ (.Y(_1906_),
    .A(net71),
    .B(net60));
 sg13g2_nor4_1 _3953_ (.A(_0024_),
    .B(_0027_),
    .C(_1906_),
    .D(_1744_),
    .Y(_1907_));
 sg13g2_nand4_1 _3954_ (.B(net72),
    .C(net70),
    .A(_1729_),
    .Y(_1908_),
    .D(net68));
 sg13g2_nand2_1 _3955_ (.Y(_1909_),
    .A(_1908_),
    .B(_1720_));
 sg13g2_a21o_1 _3956_ (.A2(_1798_),
    .A1(_1797_),
    .B1(_1720_),
    .X(_1910_));
 sg13g2_nand3_1 _3957_ (.B(_1909_),
    .C(_1910_),
    .A(_1907_),
    .Y(_1911_));
 sg13g2_inv_1 _3958_ (.Y(_1912_),
    .A(_1911_));
 sg13g2_nor2_2 _3959_ (.A(_1723_),
    .B(_1912_),
    .Y(_1913_));
 sg13g2_inv_1 _3960_ (.Y(_1914_),
    .A(_1913_));
 sg13g2_nor2_1 _3961_ (.A(_1905_),
    .B(net21),
    .Y(_0113_));
 sg13g2_inv_1 _3962_ (.Y(_1915_),
    .A(_1906_));
 sg13g2_nor3_1 _3963_ (.A(_1726_),
    .B(_1915_),
    .C(net21),
    .Y(_0114_));
 sg13g2_nor2_1 _3964_ (.A(_1725_),
    .B(_1915_),
    .Y(_1916_));
 sg13g2_nor2_1 _3965_ (.A(_1720_),
    .B(_1906_),
    .Y(_1917_));
 sg13g2_nor3_1 _3966_ (.A(_1916_),
    .B(_1917_),
    .C(net21),
    .Y(_0115_));
 sg13g2_nor2_1 _3967_ (.A(_1724_),
    .B(_1917_),
    .Y(_1918_));
 sg13g2_nor2_1 _3968_ (.A(_1739_),
    .B(_1906_),
    .Y(_1919_));
 sg13g2_nor3_1 _3969_ (.A(_1918_),
    .B(_1919_),
    .C(net21),
    .Y(_0116_));
 sg13g2_nor2_1 _3970_ (.A(net61),
    .B(_1919_),
    .Y(_1920_));
 sg13g2_nand2_1 _3971_ (.Y(_1921_),
    .A(_1919_),
    .B(_1707_));
 sg13g2_inv_1 _3972_ (.Y(_1922_),
    .A(_1921_));
 sg13g2_nor3_1 _3973_ (.A(_1920_),
    .B(_1922_),
    .C(net21),
    .Y(_0117_));
 sg13g2_nor2_1 _3974_ (.A(_1733_),
    .B(_1922_),
    .Y(_1923_));
 sg13g2_nor2_1 _3975_ (.A(_1709_),
    .B(_1921_),
    .Y(_1924_));
 sg13g2_nor3_1 _3976_ (.A(_1923_),
    .B(_1924_),
    .C(net21),
    .Y(_0118_));
 sg13g2_nand2_1 _3977_ (.Y(_1925_),
    .A(_1924_),
    .B(_1703_));
 sg13g2_inv_1 _3978_ (.Y(_1926_),
    .A(_1925_));
 sg13g2_nor2_1 _3979_ (.A(net72),
    .B(_1924_),
    .Y(_1927_));
 sg13g2_nor3_1 _3980_ (.A(_1926_),
    .B(_1927_),
    .C(net21),
    .Y(_0119_));
 sg13g2_nor2_1 _3981_ (.A(net70),
    .B(_1926_),
    .Y(_1928_));
 sg13g2_nor2_1 _3982_ (.A(_1704_),
    .B(_1925_),
    .Y(_1929_));
 sg13g2_nor3_1 _3983_ (.A(_1928_),
    .B(_1929_),
    .C(net21),
    .Y(_0120_));
 sg13g2_nor2_1 _3984_ (.A(_1699_),
    .B(_1929_),
    .Y(_1930_));
 sg13g2_nand2_1 _3985_ (.Y(_1931_),
    .A(_1929_),
    .B(_1699_));
 sg13g2_inv_1 _3986_ (.Y(_1932_),
    .A(_1931_));
 sg13g2_nor3_1 _3987_ (.A(_1930_),
    .B(_1932_),
    .C(_1914_),
    .Y(_0121_));
 sg13g2_o21ai_1 _3988_ (.B1(_1913_),
    .Y(_1933_),
    .A1(_1729_),
    .A2(_1931_));
 sg13g2_a21oi_1 _3989_ (.A1(_1729_),
    .A2(_1931_),
    .Y(_0122_),
    .B1(_1933_));
 sg13g2_nand3_1 _3990_ (.B(_1909_),
    .C(_1910_),
    .A(_1907_),
    .Y(_1934_));
 sg13g2_nor2_1 _3991_ (.A(_1767_),
    .B(_1934_),
    .Y(_1935_));
 sg13g2_nor3_1 _3992_ (.A(_1747_),
    .B(net69),
    .C(_1774_),
    .Y(_1936_));
 sg13g2_inv_1 _3993_ (.Y(_1937_),
    .A(_1754_));
 sg13g2_nand3_1 _3994_ (.B(_1936_),
    .C(_1937_),
    .A(_1790_),
    .Y(_1938_));
 sg13g2_nand2_1 _3995_ (.Y(_1939_),
    .A(_1766_),
    .B(_1768_));
 sg13g2_nor2_1 _3996_ (.A(_1760_),
    .B(_1761_),
    .Y(_1940_));
 sg13g2_inv_1 _3997_ (.Y(_1941_),
    .A(_1940_));
 sg13g2_nor4_1 _3998_ (.A(_1750_),
    .B(net69),
    .C(_1939_),
    .D(_1941_),
    .Y(_1942_));
 sg13g2_nor4_1 _3999_ (.A(_1765_),
    .B(_1752_),
    .C(_1770_),
    .D(_1937_),
    .Y(_1943_));
 sg13g2_nand2_1 _4000_ (.Y(_1944_),
    .A(_1942_),
    .B(_1943_));
 sg13g2_a21o_1 _4001_ (.A2(_1944_),
    .A1(_1938_),
    .B1(_0028_),
    .X(_1945_));
 sg13g2_a21oi_1 _4002_ (.A1(_1945_),
    .A2(_1912_),
    .Y(_1946_),
    .B1(_1766_));
 sg13g2_nor3_1 _4003_ (.A(_1723_),
    .B(_1935_),
    .C(_1946_),
    .Y(_0124_));
 sg13g2_nor2_1 _4004_ (.A(_1768_),
    .B(_1935_),
    .Y(_1947_));
 sg13g2_nor2_1 _4005_ (.A(_1767_),
    .B(_1911_),
    .Y(_1948_));
 sg13g2_nand2_1 _4006_ (.Y(_1949_),
    .A(_1948_),
    .B(net67));
 sg13g2_inv_1 _4007_ (.Y(_1950_),
    .A(_1949_));
 sg13g2_nor3_1 _4008_ (.A(_1723_),
    .B(_1947_),
    .C(_1950_),
    .Y(_0125_));
 sg13g2_nor2_1 _4009_ (.A(_1775_),
    .B(_1949_),
    .Y(_1951_));
 sg13g2_nor2_1 _4010_ (.A(_1939_),
    .B(_1941_),
    .Y(_1952_));
 sg13g2_nand2_1 _4011_ (.Y(_1953_),
    .A(_1952_),
    .B(_1753_));
 sg13g2_nor3_1 _4012_ (.A(_1772_),
    .B(_1783_),
    .C(_1953_),
    .Y(_1954_));
 sg13g2_inv_1 _4013_ (.Y(_1955_),
    .A(_1954_));
 sg13g2_nor3_1 _4014_ (.A(_1754_),
    .B(_1788_),
    .C(_1789_),
    .Y(_1956_));
 sg13g2_nand3_1 _4015_ (.B(_1765_),
    .C(_1936_),
    .A(_1956_),
    .Y(_1957_));
 sg13g2_a21oi_1 _4016_ (.A1(_1955_),
    .A2(_1957_),
    .Y(_1958_),
    .B1(_0028_));
 sg13g2_inv_1 _4017_ (.Y(_1959_),
    .A(_1934_));
 sg13g2_nand2_2 _4018_ (.Y(_1960_),
    .A(_1958_),
    .B(_1959_));
 sg13g2_inv_1 _4019_ (.Y(_1961_),
    .A(_1723_));
 sg13g2_nand2_2 _4020_ (.Y(_1962_),
    .A(_1960_),
    .B(_1961_));
 sg13g2_nor2_1 _4021_ (.A(_1760_),
    .B(_1950_),
    .Y(_1963_));
 sg13g2_nor3_1 _4022_ (.A(_1951_),
    .B(_1962_),
    .C(_1963_),
    .Y(_0126_));
 sg13g2_nor2_1 _4023_ (.A(_1788_),
    .B(_1939_),
    .Y(_1964_));
 sg13g2_inv_1 _4024_ (.Y(_1965_),
    .A(_1964_));
 sg13g2_nor2_1 _4025_ (.A(_1965_),
    .B(_1934_),
    .Y(_1966_));
 sg13g2_nor2_1 _4026_ (.A(_1761_),
    .B(_1951_),
    .Y(_1967_));
 sg13g2_nor3_1 _4027_ (.A(_1966_),
    .B(_1962_),
    .C(_1967_),
    .Y(_0127_));
 sg13g2_nor2_1 _4028_ (.A(_1750_),
    .B(_1966_),
    .Y(_1968_));
 sg13g2_inv_1 _4029_ (.Y(_1969_),
    .A(_1750_));
 sg13g2_nor3_1 _4030_ (.A(_1969_),
    .B(_1788_),
    .C(_1949_),
    .Y(_1970_));
 sg13g2_nor3_1 _4031_ (.A(_1962_),
    .B(_1968_),
    .C(_1970_),
    .Y(_0128_));
 sg13g2_nor2_1 _4032_ (.A(_1969_),
    .B(_1965_),
    .Y(_1971_));
 sg13g2_xor2_1 _4033_ (.B(_1971_),
    .A(_0029_),
    .X(_1972_));
 sg13g2_nand3_1 _4034_ (.B(_1961_),
    .C(_1912_),
    .A(_1945_),
    .Y(_1973_));
 sg13g2_nand2_1 _4035_ (.Y(_1974_),
    .A(_1913_),
    .B(_1751_));
 sg13g2_o21ai_1 _4036_ (.B1(_1974_),
    .Y(_0129_),
    .A1(_1972_),
    .A2(_1973_));
 sg13g2_inv_1 _4037_ (.Y(_1975_),
    .A(_1748_));
 sg13g2_nand2_1 _4038_ (.Y(_1976_),
    .A(_1970_),
    .B(_1751_));
 sg13g2_nand3_1 _4039_ (.B(_1751_),
    .C(_1748_),
    .A(_1970_),
    .Y(_1977_));
 sg13g2_nand2b_1 _4040_ (.Y(_1978_),
    .B(_1977_),
    .A_N(_1962_));
 sg13g2_a21oi_1 _4041_ (.A1(_1975_),
    .A2(_1976_),
    .Y(_0130_),
    .B1(_1978_));
 sg13g2_xnor2_1 _4042_ (.Y(_1979_),
    .A(_1770_),
    .B(_1977_));
 sg13g2_nor2_1 _4043_ (.A(_1962_),
    .B(_1979_),
    .Y(_0131_));
 sg13g2_inv_1 _4044_ (.Y(_1980_),
    .A(_0030_));
 sg13g2_nor4_2 _4045_ (.A(_1969_),
    .B(_1752_),
    .C(_1749_),
    .Y(_1981_),
    .D(_1965_));
 sg13g2_xnor2_1 _4046_ (.Y(_1982_),
    .A(_1980_),
    .B(_1981_));
 sg13g2_nand2_1 _4047_ (.Y(_1983_),
    .A(_1913_),
    .B(_1754_));
 sg13g2_o21ai_1 _4048_ (.B1(_1983_),
    .Y(_0132_),
    .A1(_1982_),
    .A2(_1973_));
 sg13g2_nand2_1 _4049_ (.Y(_1984_),
    .A(_1981_),
    .B(_1754_));
 sg13g2_xnor2_1 _4050_ (.Y(_1985_),
    .A(_0028_),
    .B(_1984_));
 sg13g2_nand2_1 _4051_ (.Y(_1986_),
    .A(_1913_),
    .B(_1755_));
 sg13g2_o21ai_1 _4052_ (.B1(_1986_),
    .Y(_0133_),
    .A1(_1985_),
    .A2(_1973_));
 sg13g2_and2_1 _4053_ (.A(_0004_),
    .B(_0003_),
    .X(_0057_));
 sg13g2_nand2_1 _4054_ (.Y(_1987_),
    .A(net73),
    .B(_0055_));
 sg13g2_inv_1 _4055_ (.Y(_0058_),
    .A(_1987_));
 sg13g2_o21ai_1 _4056_ (.B1(net73),
    .Y(_1988_),
    .A1(_1631_),
    .A2(_1646_));
 sg13g2_a21oi_1 _4057_ (.A1(_1631_),
    .A2(_1646_),
    .Y(_0059_),
    .B1(_1988_));
 sg13g2_buf_1 _4058_ (.A(_1621_),
    .X(_1989_));
 sg13g2_a21oi_1 _4059_ (.A1(_1645_),
    .A2(_1592_),
    .Y(_1990_),
    .B1(_1618_));
 sg13g2_nor3_1 _4060_ (.A(net56),
    .B(_1990_),
    .C(_1647_),
    .Y(_0060_));
 sg13g2_nor2_1 _4061_ (.A(_1614_),
    .B(_1647_),
    .Y(_1991_));
 sg13g2_inv_1 _4062_ (.Y(_1992_),
    .A(_1648_));
 sg13g2_nor3_1 _4063_ (.A(net56),
    .B(_1991_),
    .C(_1992_),
    .Y(_0061_));
 sg13g2_nor2_1 _4064_ (.A(_1613_),
    .B(_1992_),
    .Y(_1993_));
 sg13g2_nor3_1 _4065_ (.A(_1989_),
    .B(_1649_),
    .C(_1993_),
    .Y(_0062_));
 sg13g2_nor2b_1 _4066_ (.A(_1664_),
    .B_N(_1616_),
    .Y(_1994_));
 sg13g2_nor2_1 _4067_ (.A(_1616_),
    .B(_1649_),
    .Y(_1995_));
 sg13g2_nor3_1 _4068_ (.A(_1989_),
    .B(_1994_),
    .C(_1995_),
    .Y(_0063_));
 sg13g2_a21oi_1 _4069_ (.A1(_1649_),
    .A2(_1616_),
    .Y(_1996_),
    .B1(_1615_));
 sg13g2_inv_1 _4070_ (.Y(_1997_),
    .A(_1650_));
 sg13g2_nor3_1 _4071_ (.A(net56),
    .B(_1996_),
    .C(_1997_),
    .Y(_0064_));
 sg13g2_o21ai_1 _4072_ (.B1(net73),
    .Y(_1998_),
    .A1(_1626_),
    .A2(_1665_));
 sg13g2_a21oi_1 _4073_ (.A1(_1626_),
    .A2(_1665_),
    .Y(_0065_),
    .B1(_1998_));
 sg13g2_nor3_1 _4074_ (.A(_1625_),
    .B(_1626_),
    .C(_1650_),
    .Y(_1999_));
 sg13g2_a21oi_1 _4075_ (.A1(_1997_),
    .A2(_1605_),
    .Y(_2000_),
    .B1(\counter[17] ));
 sg13g2_nor3_1 _4076_ (.A(net56),
    .B(_1999_),
    .C(_2000_),
    .Y(_0066_));
 sg13g2_nor2_1 _4077_ (.A(_1607_),
    .B(_1999_),
    .Y(_2001_));
 sg13g2_nand2_1 _4078_ (.Y(_2002_),
    .A(_1999_),
    .B(_1607_));
 sg13g2_inv_1 _4079_ (.Y(_2003_),
    .A(_2002_));
 sg13g2_nor3_1 _4080_ (.A(net56),
    .B(_2001_),
    .C(_2003_),
    .Y(_0067_));
 sg13g2_inv_1 _4081_ (.Y(_2004_),
    .A(_1606_));
 sg13g2_nor2_1 _4082_ (.A(_2004_),
    .B(_2002_),
    .Y(_2005_));
 sg13g2_nor2_1 _4083_ (.A(_1606_),
    .B(_2003_),
    .Y(_2006_));
 sg13g2_nor3_1 _4084_ (.A(net56),
    .B(_2005_),
    .C(_2006_),
    .Y(_0068_));
 sg13g2_buf_1 _4085_ (.A(_1621_),
    .X(_2007_));
 sg13g2_inv_1 _4086_ (.Y(_2008_),
    .A(_1634_));
 sg13g2_nor3_1 _4087_ (.A(net55),
    .B(_1598_),
    .C(_2008_),
    .Y(_0069_));
 sg13g2_nor2_1 _4088_ (.A(_1602_),
    .B(_2005_),
    .Y(_2009_));
 sg13g2_and2_1 _4089_ (.A(_2005_),
    .B(_1602_),
    .X(_2010_));
 sg13g2_nor3_1 _4090_ (.A(_2007_),
    .B(_2009_),
    .C(_2010_),
    .Y(_0070_));
 sg13g2_nor2_1 _4091_ (.A(\counter[21] ),
    .B(_2010_),
    .Y(_2011_));
 sg13g2_nor3_1 _4092_ (.A(net55),
    .B(_1651_),
    .C(_2011_),
    .Y(_0071_));
 sg13g2_inv_1 _4093_ (.Y(_2012_),
    .A(_1603_));
 sg13g2_inv_1 _4094_ (.Y(_2013_),
    .A(_1651_));
 sg13g2_o21ai_1 _4095_ (.B1(net73),
    .Y(_2014_),
    .A1(_2012_),
    .A2(_2013_));
 sg13g2_a21oi_1 _4096_ (.A1(_2012_),
    .A2(_2013_),
    .Y(_0072_),
    .B1(_2014_));
 sg13g2_nor2_1 _4097_ (.A(_1654_),
    .B(_2013_),
    .Y(_2015_));
 sg13g2_a21oi_1 _4098_ (.A1(_1651_),
    .A2(_1603_),
    .Y(_2016_),
    .B1(\counter[23] ));
 sg13g2_nor3_1 _4099_ (.A(_2007_),
    .B(_2015_),
    .C(_2016_),
    .Y(_0073_));
 sg13g2_o21ai_1 _4100_ (.B1(_1669_),
    .Y(_2017_),
    .A1(_1609_),
    .A2(_2015_));
 sg13g2_nand2_1 _4101_ (.Y(_2018_),
    .A(_2015_),
    .B(_1609_));
 sg13g2_nor2b_1 _4102_ (.A(_2017_),
    .B_N(_2018_),
    .Y(_0074_));
 sg13g2_a221oi_1 _4103_ (.B2(_1652_),
    .C1(net56),
    .B1(_2018_),
    .A1(_1655_),
    .Y(_0075_),
    .A2(_1651_));
 sg13g2_o21ai_1 _4104_ (.B1(net73),
    .Y(_2019_),
    .A1(_1696_),
    .A2(_1656_));
 sg13g2_a21oi_1 _4105_ (.A1(_1696_),
    .A2(_1656_),
    .Y(_0076_),
    .B1(_2019_));
 sg13g2_nor2_1 _4106_ (.A(\counter[2] ),
    .B(_2008_),
    .Y(_2020_));
 sg13g2_nor3_1 _4107_ (.A(net55),
    .B(_1635_),
    .C(_2020_),
    .Y(_0080_));
 sg13g2_nor2_1 _4108_ (.A(\counter[30] ),
    .B(_1660_),
    .Y(_2021_));
 sg13g2_nand2_1 _4109_ (.Y(_2022_),
    .A(_1660_),
    .B(\counter[30] ));
 sg13g2_inv_1 _4110_ (.Y(_2023_),
    .A(_2022_));
 sg13g2_nor3_1 _4111_ (.A(net55),
    .B(_2021_),
    .C(_2023_),
    .Y(_0081_));
 sg13g2_inv_1 _4112_ (.Y(_2024_),
    .A(\counter[31] ));
 sg13g2_o21ai_1 _4113_ (.B1(net73),
    .Y(_2025_),
    .A1(_2024_),
    .A2(_2022_));
 sg13g2_a21oi_1 _4114_ (.A1(_2024_),
    .A2(_2022_),
    .Y(_0082_),
    .B1(_2025_));
 sg13g2_nor2_1 _4115_ (.A(\counter[3] ),
    .B(_1635_),
    .Y(_2026_));
 sg13g2_nor3_1 _4116_ (.A(net55),
    .B(_2026_),
    .C(_1637_),
    .Y(_0083_));
 sg13g2_nor2_1 _4117_ (.A(\counter[4] ),
    .B(_1637_),
    .Y(_2027_));
 sg13g2_nor3_1 _4118_ (.A(net55),
    .B(_2027_),
    .C(_1639_),
    .Y(_0084_));
 sg13g2_nor2_1 _4119_ (.A(\counter[5] ),
    .B(_1639_),
    .Y(_2028_));
 sg13g2_nor3_1 _4120_ (.A(net55),
    .B(_2028_),
    .C(_1641_),
    .Y(_0085_));
 sg13g2_nor2_1 _4121_ (.A(\counter[6] ),
    .B(_1641_),
    .Y(_2029_));
 sg13g2_nor2_1 _4122_ (.A(_1596_),
    .B(_1642_),
    .Y(_2030_));
 sg13g2_nor3_1 _4123_ (.A(net55),
    .B(_2029_),
    .C(_2030_),
    .Y(_0086_));
 sg13g2_nor2_1 _4124_ (.A(\counter[7] ),
    .B(_2030_),
    .Y(_2031_));
 sg13g2_nor3_1 _4125_ (.A(_1621_),
    .B(_1643_),
    .C(_2031_),
    .Y(_0087_));
 sg13g2_nor2_1 _4126_ (.A(\counter[8] ),
    .B(_1643_),
    .Y(_2032_));
 sg13g2_inv_1 _4127_ (.Y(_2033_),
    .A(_1644_));
 sg13g2_nor3_1 _4128_ (.A(_1621_),
    .B(_2032_),
    .C(_2033_),
    .Y(_0088_));
 sg13g2_nor2_1 _4129_ (.A(\counter[9] ),
    .B(_2033_),
    .Y(_2034_));
 sg13g2_nor3_1 _4130_ (.A(_1621_),
    .B(_1645_),
    .C(_2034_),
    .Y(_0089_));
 sg13g2_inv_1 _4131_ (.Y(_2035_),
    .A(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_o21ai_1 _4132_ (.B1(_1685_),
    .Y(_2036_),
    .A1(_0056_),
    .A2(_1960_));
 sg13g2_a21oi_1 _4133_ (.A1(_2035_),
    .A2(_1960_),
    .Y(_0101_),
    .B1(_2036_));
 sg13g2_buf_1 _4134_ (.A(_1840_),
    .X(_2037_));
 sg13g2_inv_1 _4135_ (.Y(_2038_),
    .A(\i_project.controller_0.t[10] ));
 sg13g2_buf_2 _4136_ (.A(\i_project.controller_0.t[9] ),
    .X(_2039_));
 sg13g2_buf_2 _4137_ (.A(\i_project.controller_0.t[8] ),
    .X(_2040_));
 sg13g2_buf_1 _4138_ (.A(\i_project.controller_0.mode_ramp_base[7] ),
    .X(_2041_));
 sg13g2_buf_1 _4139_ (.A(\i_project.controller_0.mode_ramp_base[6] ),
    .X(_2042_));
 sg13g2_buf_1 _4140_ (.A(_2042_),
    .X(_2043_));
 sg13g2_nand4_1 _4141_ (.B(_2040_),
    .C(_2041_),
    .A(_2039_),
    .Y(_2044_),
    .D(_2043_));
 sg13g2_buf_1 _4142_ (.A(\i_project.controller_0.mode_ramp_base[5] ),
    .X(_2045_));
 sg13g2_buf_1 _4143_ (.A(_2045_),
    .X(_2046_));
 sg13g2_inv_2 _4144_ (.Y(_2047_),
    .A(_2046_));
 sg13g2_buf_1 _4145_ (.A(\i_project.controller_0.mode_ramp_base[4] ),
    .X(_2048_));
 sg13g2_inv_2 _4146_ (.Y(_2049_),
    .A(net65));
 sg13g2_buf_1 _4147_ (.A(\i_project.controller_0.mode_ramp_base[3] ),
    .X(_2050_));
 sg13g2_inv_1 _4148_ (.Y(_2051_),
    .A(_2050_));
 sg13g2_buf_2 _4149_ (.A(\i_project.controller_0.mode_ramp_base[2] ),
    .X(_2052_));
 sg13g2_inv_2 _4150_ (.Y(_2053_),
    .A(_2052_));
 sg13g2_nor4_1 _4151_ (.A(_2047_),
    .B(_2049_),
    .C(_2051_),
    .D(_2053_),
    .Y(_2054_));
 sg13g2_buf_1 _4152_ (.A(\i_project.controller_0.mode_ramp_base[1] ),
    .X(_2055_));
 sg13g2_nand3_1 _4153_ (.B(net63),
    .C(\i_project.controller_0.mode_ramp_base[0] ),
    .A(_2054_),
    .Y(_2056_));
 sg13g2_nor4_2 _4154_ (.A(_2038_),
    .B(_2044_),
    .C(_2056_),
    .Y(_2057_),
    .D(_1960_));
 sg13g2_inv_1 _4155_ (.Y(_2058_),
    .A(_2040_));
 sg13g2_inv_1 _4156_ (.Y(_2059_),
    .A(net54));
 sg13g2_nor2_1 _4157_ (.A(_1911_),
    .B(_1945_),
    .Y(_2060_));
 sg13g2_nand3_1 _4158_ (.B(net63),
    .C(\i_project.controller_0.mode_ramp_base[0] ),
    .A(_2060_),
    .Y(_2061_));
 sg13g2_nor2_1 _4159_ (.A(_2053_),
    .B(_2061_),
    .Y(_2062_));
 sg13g2_nand2_1 _4160_ (.Y(_2063_),
    .A(_2062_),
    .B(net64));
 sg13g2_nor2_1 _4161_ (.A(_2049_),
    .B(_2063_),
    .Y(_2064_));
 sg13g2_inv_1 _4162_ (.Y(_2065_),
    .A(_2064_));
 sg13g2_nor3_1 _4163_ (.A(_2059_),
    .B(_2047_),
    .C(_2065_),
    .Y(_2066_));
 sg13g2_nand2_1 _4164_ (.Y(_2067_),
    .A(_2066_),
    .B(net66));
 sg13g2_nor2_1 _4165_ (.A(_2058_),
    .B(_2067_),
    .Y(_2068_));
 sg13g2_nand2_1 _4166_ (.Y(_2069_),
    .A(_2068_),
    .B(_2039_));
 sg13g2_inv_1 _4167_ (.Y(_2070_),
    .A(_2069_));
 sg13g2_nor2_1 _4168_ (.A(\i_project.controller_0.t[10] ),
    .B(_2070_),
    .Y(_2071_));
 sg13g2_nor3_1 _4169_ (.A(_2037_),
    .B(_2057_),
    .C(_2071_),
    .Y(_0102_));
 sg13g2_buf_1 _4170_ (.A(\i_project.controller_0.t[11] ),
    .X(_2072_));
 sg13g2_xnor2_1 _4171_ (.Y(_2073_),
    .A(_2072_),
    .B(_2057_));
 sg13g2_nor2_1 _4172_ (.A(_2037_),
    .B(_2073_),
    .Y(_0103_));
 sg13g2_nor2_1 _4173_ (.A(_2035_),
    .B(_1960_),
    .Y(_2074_));
 sg13g2_nor2_1 _4174_ (.A(_2055_),
    .B(_2074_),
    .Y(_2075_));
 sg13g2_nand2_1 _4175_ (.Y(_2076_),
    .A(_2074_),
    .B(_2055_));
 sg13g2_inv_1 _4176_ (.Y(_2077_),
    .A(_2076_));
 sg13g2_nor3_1 _4177_ (.A(net44),
    .B(_2075_),
    .C(_2077_),
    .Y(_0104_));
 sg13g2_nor2_1 _4178_ (.A(_2053_),
    .B(_2076_),
    .Y(_2078_));
 sg13g2_nor2_1 _4179_ (.A(_2052_),
    .B(_2077_),
    .Y(_2079_));
 sg13g2_nor3_1 _4180_ (.A(net44),
    .B(_2078_),
    .C(_2079_),
    .Y(_0105_));
 sg13g2_nor2_1 _4181_ (.A(net64),
    .B(_2078_),
    .Y(_2080_));
 sg13g2_inv_1 _4182_ (.Y(_2081_),
    .A(_2063_));
 sg13g2_nor3_1 _4183_ (.A(net44),
    .B(_2080_),
    .C(_2081_),
    .Y(_0106_));
 sg13g2_nor2_1 _4184_ (.A(net65),
    .B(_2081_),
    .Y(_2082_));
 sg13g2_nor3_1 _4185_ (.A(net44),
    .B(_2064_),
    .C(_2082_),
    .Y(_0107_));
 sg13g2_nor2_1 _4186_ (.A(net53),
    .B(_2064_),
    .Y(_2083_));
 sg13g2_nor2_1 _4187_ (.A(_2047_),
    .B(_2065_),
    .Y(_2084_));
 sg13g2_nor3_1 _4188_ (.A(net44),
    .B(_2083_),
    .C(_2084_),
    .Y(_0108_));
 sg13g2_nor2_1 _4189_ (.A(net54),
    .B(_2084_),
    .Y(_2085_));
 sg13g2_nor3_1 _4190_ (.A(net44),
    .B(_2066_),
    .C(_2085_),
    .Y(_0109_));
 sg13g2_nor2_1 _4191_ (.A(net66),
    .B(_2066_),
    .Y(_2086_));
 sg13g2_inv_1 _4192_ (.Y(_2087_),
    .A(_2067_));
 sg13g2_nor3_1 _4193_ (.A(net44),
    .B(_2086_),
    .C(_2087_),
    .Y(_0110_));
 sg13g2_nor2_1 _4194_ (.A(_2040_),
    .B(_2087_),
    .Y(_2088_));
 sg13g2_nor3_1 _4195_ (.A(net44),
    .B(_2068_),
    .C(_2088_),
    .Y(_0111_));
 sg13g2_nor2_1 _4196_ (.A(_2039_),
    .B(_2068_),
    .Y(_2089_));
 sg13g2_nor3_1 _4197_ (.A(_1840_),
    .B(_2089_),
    .C(_2070_),
    .Y(_0112_));
 sg13g2_nor2_1 _4198_ (.A(net56),
    .B(_1862_),
    .Y(_0143_));
 sg13g2_nand2_1 _4199_ (.Y(_2090_),
    .A(net74),
    .B(net4));
 sg13g2_inv_1 _4200_ (.Y(_0144_),
    .A(_2090_));
 sg13g2_inv_1 _4201_ (.Y(_2091_),
    .A(_1815_));
 sg13g2_buf_1 _4202_ (.A(_2091_),
    .X(_2092_));
 sg13g2_nand2_1 _4203_ (.Y(_2093_),
    .A(_1786_),
    .B(_1940_));
 sg13g2_nor3_1 _4204_ (.A(_1937_),
    .B(_0029_),
    .C(_1749_),
    .Y(_2094_));
 sg13g2_nor2_1 _4205_ (.A(_1755_),
    .B(_2094_),
    .Y(_2095_));
 sg13g2_o21ai_1 _4206_ (.B1(_2095_),
    .Y(_2096_),
    .A1(_2093_),
    .A2(_1759_));
 sg13g2_nor3_1 _4207_ (.A(net69),
    .B(_1774_),
    .C(_1941_),
    .Y(_2097_));
 sg13g2_nor4_1 _4208_ (.A(_1765_),
    .B(_1770_),
    .C(_1776_),
    .D(_2097_),
    .Y(_2098_));
 sg13g2_a21oi_1 _4209_ (.A1(_2096_),
    .A2(_1765_),
    .Y(_2099_),
    .B1(_2098_));
 sg13g2_nand3_1 _4210_ (.B(net43),
    .C(_2099_),
    .A(_1807_),
    .Y(_2100_));
 sg13g2_nor2_1 _4211_ (.A(_0036_),
    .B(_2091_),
    .Y(_2101_));
 sg13g2_inv_1 _4212_ (.Y(_2102_),
    .A(_2101_));
 sg13g2_nand2_1 _4213_ (.Y(_2103_),
    .A(_2100_),
    .B(_2102_));
 sg13g2_buf_2 _4214_ (.A(_2103_),
    .X(_2104_));
 sg13g2_inv_1 _4215_ (.Y(_2105_),
    .A(_2104_));
 sg13g2_buf_1 _4216_ (.A(\depth[1] ),
    .X(_2106_));
 sg13g2_buf_2 _4217_ (.A(\depth[0] ),
    .X(_2107_));
 sg13g2_inv_1 _4218_ (.Y(_2108_),
    .A(\depth[2] ));
 sg13g2_nor3_1 _4219_ (.A(_2106_),
    .B(_2107_),
    .C(_2108_),
    .Y(_2109_));
 sg13g2_buf_1 _4220_ (.A(_2109_),
    .X(_2110_));
 sg13g2_inv_1 _4221_ (.Y(_2111_),
    .A(_2110_));
 sg13g2_buf_2 _4222_ (.A(_0040_),
    .X(_2112_));
 sg13g2_nand2_1 _4223_ (.Y(_2113_),
    .A(_1766_),
    .B(\i_project.controller_0.voffset[0] ));
 sg13g2_nor2_1 _4224_ (.A(net67),
    .B(_1827_),
    .Y(_2114_));
 sg13g2_nand2_1 _4225_ (.Y(_2115_),
    .A(net67),
    .B(_1827_));
 sg13g2_o21ai_1 _4226_ (.B1(_2115_),
    .Y(_2116_),
    .A1(_2113_),
    .A2(_2114_));
 sg13g2_xnor2_1 _4227_ (.Y(_2117_),
    .A(_1761_),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_nand2_1 _4228_ (.Y(_2118_),
    .A(_1775_),
    .B(_1830_));
 sg13g2_nand2_1 _4229_ (.Y(_2119_),
    .A(_1760_),
    .B(_1829_));
 sg13g2_nand2_1 _4230_ (.Y(_2120_),
    .A(_2118_),
    .B(_2119_));
 sg13g2_nor2_1 _4231_ (.A(_2117_),
    .B(_2120_),
    .Y(_2121_));
 sg13g2_nand2_1 _4232_ (.Y(_2122_),
    .A(_2116_),
    .B(_2121_));
 sg13g2_nor2_1 _4233_ (.A(_1761_),
    .B(\i_project.controller_0.voffset[3] ),
    .Y(_2123_));
 sg13g2_nand2_1 _4234_ (.Y(_2124_),
    .A(_1761_),
    .B(\i_project.controller_0.voffset[3] ));
 sg13g2_o21ai_1 _4235_ (.B1(_2124_),
    .Y(_2125_),
    .A1(_2119_),
    .A2(_2123_));
 sg13g2_inv_1 _4236_ (.Y(_2126_),
    .A(_2125_));
 sg13g2_nand2_1 _4237_ (.Y(_2127_),
    .A(_2122_),
    .B(_2126_));
 sg13g2_xnor2_1 _4238_ (.Y(_2128_),
    .A(_1750_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_inv_1 _4239_ (.Y(_2129_),
    .A(_2128_));
 sg13g2_nand2_1 _4240_ (.Y(_2130_),
    .A(_2127_),
    .B(_2129_));
 sg13g2_nand3_1 _4241_ (.B(_2128_),
    .C(_2126_),
    .A(_2122_),
    .Y(_2131_));
 sg13g2_nand2_1 _4242_ (.Y(_2132_),
    .A(_2130_),
    .B(_2131_));
 sg13g2_buf_8 _4243_ (.A(_2132_),
    .X(_2133_));
 sg13g2_nor2_1 _4244_ (.A(_2112_),
    .B(net20),
    .Y(_2134_));
 sg13g2_nor2_1 _4245_ (.A(_1760_),
    .B(_1829_),
    .Y(_2135_));
 sg13g2_o21ai_1 _4246_ (.B1(_2119_),
    .Y(_2136_),
    .A1(_2115_),
    .A2(_2135_));
 sg13g2_nor2_1 _4247_ (.A(_2128_),
    .B(_2117_),
    .Y(_2137_));
 sg13g2_nand2_1 _4248_ (.Y(_2138_),
    .A(_1750_),
    .B(\i_project.controller_0.voffset[4] ));
 sg13g2_nor2_1 _4249_ (.A(_1750_),
    .B(\i_project.controller_0.voffset[4] ),
    .Y(_2139_));
 sg13g2_a21oi_1 _4250_ (.A1(_2138_),
    .A2(_2124_),
    .Y(_2140_),
    .B1(_2139_));
 sg13g2_a21oi_1 _4251_ (.A1(_2136_),
    .A2(_2137_),
    .Y(_2141_),
    .B1(_2140_));
 sg13g2_xnor2_1 _4252_ (.Y(_2142_),
    .A(net67),
    .B(_1827_));
 sg13g2_nor2_1 _4253_ (.A(_2142_),
    .B(_2120_),
    .Y(_2143_));
 sg13g2_inv_1 _4254_ (.Y(_2144_),
    .A(_2113_));
 sg13g2_nand3_1 _4255_ (.B(_2143_),
    .C(_2144_),
    .A(_2137_),
    .Y(_2145_));
 sg13g2_nand2_1 _4256_ (.Y(_2146_),
    .A(_2141_),
    .B(_2145_));
 sg13g2_xnor2_1 _4257_ (.Y(_2147_),
    .A(_1751_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_inv_1 _4258_ (.Y(_2148_),
    .A(_2147_));
 sg13g2_nand2_1 _4259_ (.Y(_2149_),
    .A(_2146_),
    .B(_2148_));
 sg13g2_nand3_1 _4260_ (.B(_2145_),
    .C(_2147_),
    .A(_2141_),
    .Y(_2150_));
 sg13g2_nand2_1 _4261_ (.Y(_2151_),
    .A(_2149_),
    .B(_2150_));
 sg13g2_buf_8 _4262_ (.A(_2151_),
    .X(_2152_));
 sg13g2_nor2_1 _4263_ (.A(_0039_),
    .B(_2152_),
    .Y(_2153_));
 sg13g2_nand2_1 _4264_ (.Y(_2154_),
    .A(_2152_),
    .B(_0039_));
 sg13g2_o21ai_1 _4265_ (.B1(_2154_),
    .Y(_2155_),
    .A1(_2134_),
    .A2(_2153_));
 sg13g2_xor2_1 _4266_ (.B(_1827_),
    .A(net67),
    .X(_2156_));
 sg13g2_xor2_1 _4267_ (.B(_1829_),
    .A(_1760_),
    .X(_2157_));
 sg13g2_nand3_1 _4268_ (.B(_2157_),
    .C(_2144_),
    .A(_2156_),
    .Y(_2158_));
 sg13g2_inv_1 _4269_ (.Y(_2159_),
    .A(_2136_));
 sg13g2_nand2_1 _4270_ (.Y(_2160_),
    .A(_2158_),
    .B(_2159_));
 sg13g2_xnor2_1 _4271_ (.Y(_2161_),
    .A(net69),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_nor2_1 _4272_ (.A(_2161_),
    .B(_2147_),
    .Y(_2162_));
 sg13g2_and2_1 _4273_ (.A(_2162_),
    .B(_2137_),
    .X(_2163_));
 sg13g2_nand2_1 _4274_ (.Y(_2164_),
    .A(_2160_),
    .B(_2163_));
 sg13g2_nand2_1 _4275_ (.Y(_2165_),
    .A(_1751_),
    .B(\i_project.controller_0.voffset[5] ));
 sg13g2_nor2_1 _4276_ (.A(net69),
    .B(\i_project.controller_0.voffset[6] ),
    .Y(_2166_));
 sg13g2_nand2_1 _4277_ (.Y(_2167_),
    .A(net69),
    .B(\i_project.controller_0.voffset[6] ));
 sg13g2_o21ai_1 _4278_ (.B1(_2167_),
    .Y(_2168_),
    .A1(_2165_),
    .A2(_2166_));
 sg13g2_a21oi_1 _4279_ (.A1(_2162_),
    .A2(_2140_),
    .Y(_2169_),
    .B1(_2168_));
 sg13g2_nand2_1 _4280_ (.Y(_2170_),
    .A(_2164_),
    .B(_2169_));
 sg13g2_nor2_1 _4281_ (.A(_1747_),
    .B(\i_project.controller_0.voffset[7] ),
    .Y(_2171_));
 sg13g2_nand2_1 _4282_ (.Y(_2172_),
    .A(_1747_),
    .B(\i_project.controller_0.voffset[7] ));
 sg13g2_inv_1 _4283_ (.Y(_2173_),
    .A(_2172_));
 sg13g2_nor2_1 _4284_ (.A(_2171_),
    .B(_2173_),
    .Y(_2174_));
 sg13g2_nand2_1 _4285_ (.Y(_2175_),
    .A(_2170_),
    .B(_2174_));
 sg13g2_inv_1 _4286_ (.Y(_2176_),
    .A(_2174_));
 sg13g2_nand3_1 _4287_ (.B(_2176_),
    .C(_2169_),
    .A(_2164_),
    .Y(_2177_));
 sg13g2_nand2_1 _4288_ (.Y(_2178_),
    .A(_2175_),
    .B(_2177_));
 sg13g2_buf_8 _4289_ (.A(_2178_),
    .X(_2179_));
 sg13g2_inv_1 _4290_ (.Y(_2180_),
    .A(_0019_));
 sg13g2_nand2_1 _4291_ (.Y(_2181_),
    .A(_2179_),
    .B(_2180_));
 sg13g2_nand3_1 _4292_ (.B(_2177_),
    .C(_0019_),
    .A(_2175_),
    .Y(_2182_));
 sg13g2_nand2_1 _4293_ (.Y(_2183_),
    .A(_2181_),
    .B(_2182_));
 sg13g2_buf_1 _4294_ (.A(_0020_),
    .X(_2184_));
 sg13g2_inv_1 _4295_ (.Y(_2185_),
    .A(_2184_));
 sg13g2_nor2_1 _4296_ (.A(_2147_),
    .B(_2128_),
    .Y(_2186_));
 sg13g2_a21oi_1 _4297_ (.A1(_1752_),
    .A2(_1835_),
    .Y(_2187_),
    .B1(_2138_));
 sg13g2_nor2b_1 _4298_ (.A(_2187_),
    .B_N(_2165_),
    .Y(_2188_));
 sg13g2_inv_1 _4299_ (.Y(_2189_),
    .A(_2188_));
 sg13g2_a21oi_1 _4300_ (.A1(_2125_),
    .A2(_2186_),
    .Y(_2190_),
    .B1(_2189_));
 sg13g2_nand3_1 _4301_ (.B(_2121_),
    .C(_2186_),
    .A(_2116_),
    .Y(_2191_));
 sg13g2_nand2_1 _4302_ (.Y(_2192_),
    .A(_2190_),
    .B(_2191_));
 sg13g2_inv_1 _4303_ (.Y(_2193_),
    .A(_2161_));
 sg13g2_nand2_1 _4304_ (.Y(_2194_),
    .A(_2192_),
    .B(_2193_));
 sg13g2_nand3_1 _4305_ (.B(_2191_),
    .C(_2161_),
    .A(_2190_),
    .Y(_2195_));
 sg13g2_nand2_2 _4306_ (.Y(_2196_),
    .A(_2194_),
    .B(_2195_));
 sg13g2_xnor2_1 _4307_ (.Y(_2197_),
    .A(_2185_),
    .B(_2196_));
 sg13g2_nand2_1 _4308_ (.Y(_2198_),
    .A(_2183_),
    .B(_2197_));
 sg13g2_nor2_1 _4309_ (.A(_2155_),
    .B(_2198_),
    .Y(_2199_));
 sg13g2_nand2_1 _4310_ (.Y(_2200_),
    .A(_2179_),
    .B(_0019_));
 sg13g2_nor2_1 _4311_ (.A(_2184_),
    .B(_2196_),
    .Y(_2201_));
 sg13g2_nand3_1 _4312_ (.B(_2177_),
    .C(_2180_),
    .A(_2175_),
    .Y(_2202_));
 sg13g2_inv_1 _4313_ (.Y(_2203_),
    .A(_2202_));
 sg13g2_a21oi_1 _4314_ (.A1(_2200_),
    .A2(_2201_),
    .Y(_2204_),
    .B1(_2203_));
 sg13g2_nor2b_1 _4315_ (.A(_2199_),
    .B_N(_2204_),
    .Y(_2205_));
 sg13g2_buf_8 _4316_ (.A(_2196_),
    .X(_2206_));
 sg13g2_xnor2_1 _4317_ (.Y(_2207_),
    .A(_2184_),
    .B(_2206_));
 sg13g2_nand2_1 _4318_ (.Y(_2208_),
    .A(_2200_),
    .B(_2202_));
 sg13g2_nor2_1 _4319_ (.A(_2207_),
    .B(_2208_),
    .Y(_2209_));
 sg13g2_nand2_1 _4320_ (.Y(_2210_),
    .A(_2156_),
    .B(_2144_));
 sg13g2_nand2_1 _4321_ (.Y(_2211_),
    .A(_2142_),
    .B(_2113_));
 sg13g2_nand2_1 _4322_ (.Y(_2212_),
    .A(_2210_),
    .B(_2211_));
 sg13g2_buf_2 _4323_ (.A(_2212_),
    .X(_2213_));
 sg13g2_nand2_1 _4324_ (.Y(_2214_),
    .A(_2213_),
    .B(_0043_));
 sg13g2_nand2_1 _4325_ (.Y(_2215_),
    .A(_1767_),
    .B(_1792_));
 sg13g2_nand2_1 _4326_ (.Y(_2216_),
    .A(_2215_),
    .B(_2113_));
 sg13g2_buf_1 _4327_ (.A(_2216_),
    .X(_2217_));
 sg13g2_nor2_1 _4328_ (.A(_2051_),
    .B(_2217_),
    .Y(_2218_));
 sg13g2_nor2_1 _4329_ (.A(_0043_),
    .B(_2213_),
    .Y(_2219_));
 sg13g2_a21oi_1 _4330_ (.A1(_2214_),
    .A2(_2218_),
    .Y(_2220_),
    .B1(_2219_));
 sg13g2_inv_1 _4331_ (.Y(_2221_),
    .A(_2220_));
 sg13g2_inv_1 _4332_ (.Y(_2222_),
    .A(_1827_));
 sg13g2_nand2_1 _4333_ (.Y(_2223_),
    .A(_1778_),
    .B(_2222_));
 sg13g2_inv_1 _4334_ (.Y(_2224_),
    .A(_2115_));
 sg13g2_a21oi_1 _4335_ (.A1(_2144_),
    .A2(_2223_),
    .Y(_2225_),
    .B1(_2224_));
 sg13g2_nand2_1 _4336_ (.Y(_2226_),
    .A(_2225_),
    .B(_2120_));
 sg13g2_nand2_1 _4337_ (.Y(_2227_),
    .A(_2116_),
    .B(_2157_));
 sg13g2_nand2_1 _4338_ (.Y(_2228_),
    .A(_2226_),
    .B(_2227_));
 sg13g2_buf_8 _4339_ (.A(_2228_),
    .X(_2229_));
 sg13g2_nand2_1 _4340_ (.Y(_0146_),
    .A(_2229_),
    .B(net53));
 sg13g2_nand3_1 _4341_ (.B(_2227_),
    .C(_2047_),
    .A(_2226_),
    .Y(_0147_));
 sg13g2_nand2_1 _4342_ (.Y(_0148_),
    .A(_0146_),
    .B(_0147_));
 sg13g2_nand2_1 _4343_ (.Y(_0149_),
    .A(_2221_),
    .B(_0148_));
 sg13g2_inv_2 _4344_ (.Y(_0150_),
    .A(_2229_));
 sg13g2_inv_1 _4345_ (.Y(_0151_),
    .A(_0042_));
 sg13g2_nand2_1 _4346_ (.Y(_0152_),
    .A(_0150_),
    .B(_0151_));
 sg13g2_nand2_2 _4347_ (.Y(_0153_),
    .A(_0149_),
    .B(_0152_));
 sg13g2_nand3_1 _4348_ (.B(_2117_),
    .C(_2159_),
    .A(_2158_),
    .Y(_0154_));
 sg13g2_nand2_1 _4349_ (.Y(_0155_),
    .A(_2115_),
    .B(_2119_));
 sg13g2_inv_1 _4350_ (.Y(_0156_),
    .A(_0155_));
 sg13g2_nand2_1 _4351_ (.Y(_0157_),
    .A(_2210_),
    .B(_0156_));
 sg13g2_inv_1 _4352_ (.Y(_0158_),
    .A(_2117_));
 sg13g2_nand3_1 _4353_ (.B(_0158_),
    .C(_2118_),
    .A(_0157_),
    .Y(_0159_));
 sg13g2_nand2_1 _4354_ (.Y(_0160_),
    .A(_0154_),
    .B(_0159_));
 sg13g2_buf_8 _4355_ (.A(_0160_),
    .X(_0161_));
 sg13g2_xnor2_1 _4356_ (.Y(_0162_),
    .A(net54),
    .B(_0161_));
 sg13g2_nand2_1 _4357_ (.Y(_0163_),
    .A(_0153_),
    .B(_0162_));
 sg13g2_buf_2 _4358_ (.A(_0041_),
    .X(_0164_));
 sg13g2_nor2_1 _4359_ (.A(_0164_),
    .B(_0161_),
    .Y(_0165_));
 sg13g2_inv_1 _4360_ (.Y(_0166_),
    .A(_0165_));
 sg13g2_nand2_1 _4361_ (.Y(_0167_),
    .A(_0163_),
    .B(_0166_));
 sg13g2_buf_8 _4362_ (.A(_2152_),
    .X(_0168_));
 sg13g2_xnor2_1 _4363_ (.Y(_0169_),
    .A(_2058_),
    .B(net18));
 sg13g2_nand2_1 _4364_ (.Y(_0170_),
    .A(_2132_),
    .B(_2112_));
 sg13g2_nor2b_1 _4365_ (.A(_2134_),
    .B_N(_0170_),
    .Y(_0171_));
 sg13g2_buf_8 _4366_ (.A(_0171_),
    .X(_0172_));
 sg13g2_nor2b_1 _4367_ (.A(_0169_),
    .B_N(_0172_),
    .Y(_0173_));
 sg13g2_nand3_1 _4368_ (.B(_0167_),
    .C(_0173_),
    .A(_2209_),
    .Y(_0174_));
 sg13g2_nand2_1 _4369_ (.Y(_0175_),
    .A(_2205_),
    .B(_0174_));
 sg13g2_nor2_1 _4370_ (.A(_2161_),
    .B(_2176_),
    .Y(_0176_));
 sg13g2_nand3_1 _4371_ (.B(_2186_),
    .C(_0176_),
    .A(_2127_),
    .Y(_0177_));
 sg13g2_o21ai_1 _4372_ (.B1(_2172_),
    .Y(_0178_),
    .A1(_2167_),
    .A2(_2171_));
 sg13g2_a21oi_1 _4373_ (.A1(_2189_),
    .A2(_0176_),
    .Y(_0179_),
    .B1(_0178_));
 sg13g2_a21o_1 _4374_ (.A2(_0179_),
    .A1(_0177_),
    .B1(_1937_),
    .X(_0180_));
 sg13g2_nand3_1 _4375_ (.B(_1937_),
    .C(_0179_),
    .A(_0177_),
    .Y(_0181_));
 sg13g2_nand2_1 _4376_ (.Y(_0182_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_nand2b_1 _4377_ (.Y(_0183_),
    .B(_0182_),
    .A_N(_2072_));
 sg13g2_nand3_1 _4378_ (.B(_0181_),
    .C(_2072_),
    .A(_0180_),
    .Y(_0184_));
 sg13g2_nand2_1 _4379_ (.Y(_0185_),
    .A(_0183_),
    .B(_0184_));
 sg13g2_inv_1 _4380_ (.Y(_0186_),
    .A(_0185_));
 sg13g2_nand2_1 _4381_ (.Y(_0187_),
    .A(_0175_),
    .B(_0186_));
 sg13g2_nand3_1 _4382_ (.B(_0174_),
    .C(_0185_),
    .A(_2205_),
    .Y(_0188_));
 sg13g2_nand2_1 _4383_ (.Y(_0189_),
    .A(_0187_),
    .B(_0188_));
 sg13g2_xor2_1 _4384_ (.B(_2072_),
    .A(_1699_),
    .X(_0190_));
 sg13g2_nand2_1 _4385_ (.Y(_0191_),
    .A(net58),
    .B(_2045_));
 sg13g2_xnor2_1 _4386_ (.Y(_0192_),
    .A(_1717_),
    .B(_2042_));
 sg13g2_nand2_1 _4387_ (.Y(_0193_),
    .A(net59),
    .B(_2042_));
 sg13g2_o21ai_1 _4388_ (.B1(_0193_),
    .Y(_0194_),
    .A1(_0191_),
    .A2(_0192_));
 sg13g2_xnor2_1 _4389_ (.Y(_0195_),
    .A(_1708_),
    .B(_2040_));
 sg13g2_xor2_1 _4390_ (.B(_2041_),
    .A(_1706_),
    .X(_0196_));
 sg13g2_inv_1 _4391_ (.Y(_0197_),
    .A(_0196_));
 sg13g2_nor2_1 _4392_ (.A(_0195_),
    .B(_0197_),
    .Y(_0198_));
 sg13g2_nand2_1 _4393_ (.Y(_0199_),
    .A(_1706_),
    .B(net66));
 sg13g2_nand2_1 _4394_ (.Y(_0200_),
    .A(net57),
    .B(_2040_));
 sg13g2_o21ai_1 _4395_ (.B1(_0200_),
    .Y(_0201_),
    .A1(_0199_),
    .A2(_0195_));
 sg13g2_a21oi_1 _4396_ (.A1(_0194_),
    .A2(_0198_),
    .Y(_0202_),
    .B1(_0201_));
 sg13g2_nand2_1 _4397_ (.Y(_0203_),
    .A(_1712_),
    .B(net64));
 sg13g2_xnor2_1 _4398_ (.Y(_0204_),
    .A(\i_project.controller_0.h[1] ),
    .B(net65));
 sg13g2_nand2_1 _4399_ (.Y(_0205_),
    .A(net71),
    .B(net65));
 sg13g2_o21ai_1 _4400_ (.B1(_0205_),
    .Y(_0206_),
    .A1(_0203_),
    .A2(_0204_));
 sg13g2_buf_1 _4401_ (.A(_0206_),
    .X(_0207_));
 sg13g2_xnor2_1 _4402_ (.Y(_0208_),
    .A(_1719_),
    .B(_2045_));
 sg13g2_nor2_1 _4403_ (.A(_0192_),
    .B(_0208_),
    .Y(_0209_));
 sg13g2_nand3_1 _4404_ (.B(_0209_),
    .C(_0198_),
    .A(_0207_),
    .Y(_0210_));
 sg13g2_nand2_1 _4405_ (.Y(_0211_),
    .A(_0202_),
    .B(_0210_));
 sg13g2_xor2_1 _4406_ (.B(_2039_),
    .A(_1703_),
    .X(_0212_));
 sg13g2_nand2_1 _4407_ (.Y(_0213_),
    .A(_0211_),
    .B(_0212_));
 sg13g2_nand2_1 _4408_ (.Y(_0214_),
    .A(net72),
    .B(_2039_));
 sg13g2_nand2_1 _4409_ (.Y(_0215_),
    .A(_0213_),
    .B(_0214_));
 sg13g2_inv_1 _4410_ (.Y(_0216_),
    .A(_0215_));
 sg13g2_nand2_1 _4411_ (.Y(_0217_),
    .A(_1737_),
    .B(\i_project.controller_0.t[10] ));
 sg13g2_nor2_1 _4412_ (.A(_1737_),
    .B(\i_project.controller_0.t[10] ),
    .Y(_0218_));
 sg13g2_a21oi_1 _4413_ (.A1(_0216_),
    .A2(_0217_),
    .Y(_0219_),
    .B1(_0218_));
 sg13g2_xnor2_1 _4414_ (.Y(_0220_),
    .A(_0190_),
    .B(_0219_));
 sg13g2_nand2_1 _4415_ (.Y(_0221_),
    .A(_0189_),
    .B(_0220_));
 sg13g2_inv_1 _4416_ (.Y(_0222_),
    .A(_0220_));
 sg13g2_nand3_1 _4417_ (.B(_0188_),
    .C(_0222_),
    .A(_0187_),
    .Y(_0223_));
 sg13g2_nor3_2 _4418_ (.A(_1809_),
    .B(_1843_),
    .C(_1822_),
    .Y(_0224_));
 sg13g2_buf_1 _4419_ (.A(_0224_),
    .X(_0225_));
 sg13g2_nand3_1 _4420_ (.B(_0223_),
    .C(_0225_),
    .A(_0221_),
    .Y(_0226_));
 sg13g2_nor3_1 _4421_ (.A(_1812_),
    .B(_0025_),
    .C(_1845_),
    .Y(_0227_));
 sg13g2_buf_2 _4422_ (.A(_0227_),
    .X(_0228_));
 sg13g2_inv_1 _4423_ (.Y(_0229_),
    .A(_0228_));
 sg13g2_a21oi_1 _4424_ (.A1(_0182_),
    .A2(_1700_),
    .Y(_0230_),
    .B1(_0229_));
 sg13g2_o21ai_1 _4425_ (.B1(_0230_),
    .Y(_0231_),
    .A1(_1700_),
    .A2(_0182_));
 sg13g2_xnor2_1 _4426_ (.Y(_0232_),
    .A(net70),
    .B(_2179_));
 sg13g2_nor3_2 _4427_ (.A(_1809_),
    .B(_1812_),
    .C(_1822_),
    .Y(_0233_));
 sg13g2_nor3_1 _4428_ (.A(_1812_),
    .B(_1845_),
    .C(_1814_),
    .Y(_0234_));
 sg13g2_buf_1 _4429_ (.A(_0234_),
    .X(_0235_));
 sg13g2_a21oi_1 _4430_ (.A1(_0232_),
    .A2(_0233_),
    .Y(_0236_),
    .B1(_0235_));
 sg13g2_nand3_1 _4431_ (.B(_0231_),
    .C(_0236_),
    .A(_0226_),
    .Y(_0237_));
 sg13g2_buf_1 _4432_ (.A(_1686_),
    .X(_0238_));
 sg13g2_inv_1 _4433_ (.Y(_0239_),
    .A(_0023_));
 sg13g2_nand2_1 _4434_ (.Y(_0240_),
    .A(_0027_),
    .B(_0238_));
 sg13g2_o21ai_1 _4435_ (.B1(_0240_),
    .Y(_0241_),
    .A1(net52),
    .A2(_0239_));
 sg13g2_a21oi_1 _4436_ (.A1(_1687_),
    .A2(_1698_),
    .Y(_0242_),
    .B1(_1690_));
 sg13g2_a21o_1 _4437_ (.A2(net50),
    .A1(_0241_),
    .B1(_0242_),
    .X(_0243_));
 sg13g2_inv_1 _4438_ (.Y(_0244_),
    .A(_0243_));
 sg13g2_nor2_1 _4439_ (.A(_1754_),
    .B(_1755_),
    .Y(_0245_));
 sg13g2_inv_1 _4440_ (.Y(_0246_),
    .A(_0245_));
 sg13g2_nand2_1 _4441_ (.Y(_0247_),
    .A(_1687_),
    .B(_0054_));
 sg13g2_a21oi_1 _4442_ (.A1(_1686_),
    .A2(_0038_),
    .Y(_0248_),
    .B1(_1689_));
 sg13g2_nand2_1 _4443_ (.Y(_0249_),
    .A(_1800_),
    .B(_1686_));
 sg13g2_o21ai_1 _4444_ (.B1(_0249_),
    .Y(_0250_),
    .A1(_1686_),
    .A2(_0037_));
 sg13g2_a22oi_1 _4445_ (.Y(_0251_),
    .B1(_1689_),
    .B2(_0250_),
    .A2(_0248_),
    .A1(_0247_));
 sg13g2_nand2_1 _4446_ (.Y(_0252_),
    .A(_0246_),
    .B(_1905_));
 sg13g2_o21ai_1 _4447_ (.B1(_0252_),
    .Y(_0253_),
    .A1(_0246_),
    .A2(_0251_));
 sg13g2_buf_2 _4448_ (.A(_0253_),
    .X(_0254_));
 sg13g2_xnor2_1 _4449_ (.Y(_0255_),
    .A(_0244_),
    .B(_0254_));
 sg13g2_buf_1 _4450_ (.A(_0235_),
    .X(_0256_));
 sg13g2_nor3_1 _4451_ (.A(_1809_),
    .B(_1843_),
    .C(_1814_),
    .Y(_0257_));
 sg13g2_buf_1 _4452_ (.A(_0257_),
    .X(_0258_));
 sg13g2_a21oi_1 _4453_ (.A1(_0255_),
    .A2(_0256_),
    .Y(_0259_),
    .B1(_0258_));
 sg13g2_nand2_1 _4454_ (.Y(_0260_),
    .A(_0237_),
    .B(_0259_));
 sg13g2_nand2_1 _4455_ (.Y(_0261_),
    .A(_1738_),
    .B(_1730_));
 sg13g2_buf_2 _4456_ (.A(_0261_),
    .X(_0262_));
 sg13g2_inv_1 _4457_ (.Y(_0263_),
    .A(_0262_));
 sg13g2_a21oi_1 _4458_ (.A1(_0244_),
    .A2(_0258_),
    .Y(_0264_),
    .B1(net27));
 sg13g2_nand2_1 _4459_ (.Y(_0265_),
    .A(_0260_),
    .B(_0264_));
 sg13g2_nand2_1 _4460_ (.Y(_0266_),
    .A(_2173_),
    .B(_1980_));
 sg13g2_o21ai_1 _4461_ (.B1(_0266_),
    .Y(_0267_),
    .A1(_1937_),
    .A2(_2175_));
 sg13g2_nand2b_1 _4462_ (.Y(_0268_),
    .B(_1755_),
    .A_N(_0267_));
 sg13g2_inv_1 _4463_ (.Y(_0269_),
    .A(net60));
 sg13g2_nand2_1 _4464_ (.Y(_0270_),
    .A(_0267_),
    .B(_1756_));
 sg13g2_nand3_1 _4465_ (.B(_0269_),
    .C(_0270_),
    .A(_0268_),
    .Y(_0271_));
 sg13g2_nand2_1 _4466_ (.Y(_0272_),
    .A(_0182_),
    .B(_1713_));
 sg13g2_nor2_1 _4467_ (.A(_0038_),
    .B(_0037_),
    .Y(_0273_));
 sg13g2_nand3_1 _4468_ (.B(_0272_),
    .C(_0273_),
    .A(_0271_),
    .Y(_0274_));
 sg13g2_nand2_1 _4469_ (.Y(_0275_),
    .A(_0274_),
    .B(_1718_));
 sg13g2_a22oi_1 _4470_ (.Y(_0276_),
    .B1(_1716_),
    .B2(net18),
    .A2(_2133_),
    .A1(_1915_));
 sg13g2_nand2_1 _4471_ (.Y(_0277_),
    .A(_2179_),
    .B(_1726_));
 sg13g2_nand3_1 _4472_ (.B(_1715_),
    .C(net60),
    .A(net19),
    .Y(_0278_));
 sg13g2_nand3_1 _4473_ (.B(_0277_),
    .C(_0278_),
    .A(_0276_),
    .Y(_0279_));
 sg13g2_a21oi_1 _4474_ (.A1(_0150_),
    .A2(net60),
    .Y(_0280_),
    .B1(_1714_));
 sg13g2_o21ai_1 _4475_ (.B1(_0280_),
    .Y(_0281_),
    .A1(_1713_),
    .A2(net22));
 sg13g2_buf_8 _4476_ (.A(_2213_),
    .X(_0282_));
 sg13g2_a22oi_1 _4477_ (.Y(_0283_),
    .B1(_1716_),
    .B2(_0282_),
    .A2(_2217_),
    .A1(_1915_));
 sg13g2_a21oi_1 _4478_ (.A1(_0281_),
    .A2(_0283_),
    .Y(_0284_),
    .B1(_1739_));
 sg13g2_a21oi_1 _4479_ (.A1(_0279_),
    .A2(_1804_),
    .Y(_0285_),
    .B1(_0284_));
 sg13g2_a21oi_1 _4480_ (.A1(_0275_),
    .A2(_0285_),
    .Y(_0286_),
    .B1(_0262_));
 sg13g2_buf_2 _4481_ (.A(_0286_),
    .X(_0287_));
 sg13g2_inv_1 _4482_ (.Y(_0288_),
    .A(_0287_));
 sg13g2_buf_1 _4483_ (.A(_0288_),
    .X(_0289_));
 sg13g2_a21oi_1 _4484_ (.A1(_0265_),
    .A2(net17),
    .Y(_0290_),
    .B1(net49));
 sg13g2_nor3_1 _4485_ (.A(_2105_),
    .B(_2111_),
    .C(_0290_),
    .Y(_0291_));
 sg13g2_dfrbp_1 _4486_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net83),
    .D(_0000_),
    .Q_N(_2285_),
    .Q(_0012_));
 sg13g2_dfrbp_1 _4487_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net84),
    .D(_0001_),
    .Q_N(_2286_),
    .Q(_0013_));
 sg13g2_dfrbp_1 _4488_ (.CLK(clknet_4_7_0_clk),
    .RESET_B(net85),
    .D(_0002_),
    .Q_N(_2284_),
    .Q(_0014_));
 sg13g2_dfrbp_1 _4489_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net86),
    .D(_0057_),
    .Q_N(_2287_),
    .Q(_0016_));
 sg13g2_dfrbp_1 _4490_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net87),
    .D(_0003_),
    .Q_N(_2283_),
    .Q(_0015_));
 sg13g2_dfrbp_1 _4491_ (.CLK(clknet_4_12_0_clk),
    .RESET_B(net88),
    .D(_0004_),
    .Q_N(_2282_),
    .Q(_0145_));
 sg13g2_buf_1 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tiehi _4486__83 (.L_HI(net83));
 sg13g2_buf_1 _4494_ (.A(net89),
    .X(uio_oe[0]));
 sg13g2_buf_1 _4495_ (.A(net90),
    .X(uio_oe[1]));
 sg13g2_buf_1 _4496_ (.A(net91),
    .X(uio_oe[2]));
 sg13g2_buf_1 _4497_ (.A(net92),
    .X(uio_oe[3]));
 sg13g2_buf_1 _4498_ (.A(net93),
    .X(uio_oe[4]));
 sg13g2_buf_1 _4499_ (.A(net94),
    .X(uio_oe[5]));
 sg13g2_buf_1 _4500_ (.A(net95),
    .X(uio_oe[6]));
 sg13g2_buf_1 _4501_ (.A(net96),
    .X(uio_oe[7]));
 sg13g2_buf_1 _4502_ (.A(net75),
    .X(uio_out[0]));
 sg13g2_buf_1 _4503_ (.A(net76),
    .X(uio_out[1]));
 sg13g2_buf_1 _4504_ (.A(net77),
    .X(uio_out[2]));
 sg13g2_buf_1 _4505_ (.A(net78),
    .X(uio_out[3]));
 sg13g2_buf_1 _4506_ (.A(net79),
    .X(uio_out[4]));
 sg13g2_buf_1 _4507_ (.A(net80),
    .X(uio_out[5]));
 sg13g2_buf_1 _4508_ (.A(net81),
    .X(uio_out[6]));
 sg13g2_buf_1 _4509_ (.A(net82),
    .X(uio_out[7]));
 sg13g2_buf_1 _4510_ (.A(\i_project.controller_0.vga_sync.o_vsync ),
    .X(net11));
 sg13g2_buf_1 _4511_ (.A(hsync),
    .X(net15));
 sg13g2_dfrbp_1 \counter[0]$_SDFF_PN0_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net97),
    .D(_0058_),
    .Q_N(_0055_),
    .Q(\counter[0] ));
 sg13g2_dfrbp_1 \counter[10]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net98),
    .D(_0059_),
    .Q_N(_2281_),
    .Q(\counter[10] ));
 sg13g2_dfrbp_1 \counter[11]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net99),
    .D(_0060_),
    .Q_N(_2280_),
    .Q(\counter[11] ));
 sg13g2_dfrbp_1 \counter[12]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net100),
    .D(_0061_),
    .Q_N(_2279_),
    .Q(\counter[12] ));
 sg13g2_dfrbp_1 \counter[13]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net101),
    .D(_0062_),
    .Q_N(_2278_),
    .Q(\counter[13] ));
 sg13g2_dfrbp_1 \counter[14]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net102),
    .D(_0063_),
    .Q_N(_2277_),
    .Q(\counter[14] ));
 sg13g2_dfrbp_1 \counter[15]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net103),
    .D(_0064_),
    .Q_N(_2276_),
    .Q(\counter[15] ));
 sg13g2_dfrbp_1 \counter[16]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net104),
    .D(_0065_),
    .Q_N(_2275_),
    .Q(\counter[16] ));
 sg13g2_dfrbp_1 \counter[17]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net105),
    .D(_0066_),
    .Q_N(_2274_),
    .Q(\counter[17] ));
 sg13g2_dfrbp_1 \counter[18]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net106),
    .D(_0067_),
    .Q_N(_2273_),
    .Q(\counter[18] ));
 sg13g2_dfrbp_1 \counter[19]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net107),
    .D(_0068_),
    .Q_N(_2272_),
    .Q(\counter[19] ));
 sg13g2_dfrbp_1 \counter[1]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net108),
    .D(_0069_),
    .Q_N(_2271_),
    .Q(\counter[1] ));
 sg13g2_dfrbp_1 \counter[20]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net109),
    .D(_0070_),
    .Q_N(_2270_),
    .Q(\counter[20] ));
 sg13g2_dfrbp_1 \counter[21]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net110),
    .D(_0071_),
    .Q_N(_2269_),
    .Q(\counter[21] ));
 sg13g2_dfrbp_1 \counter[22]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net111),
    .D(_0072_),
    .Q_N(_2268_),
    .Q(\counter[22] ));
 sg13g2_dfrbp_1 \counter[23]$_SDFF_PN0_  (.CLK(clknet_4_3_0_clk),
    .RESET_B(net112),
    .D(_0073_),
    .Q_N(_2267_),
    .Q(\counter[23] ));
 sg13g2_dfrbp_1 \counter[24]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net113),
    .D(_0074_),
    .Q_N(_2266_),
    .Q(\counter[24] ));
 sg13g2_dfrbp_1 \counter[25]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net114),
    .D(_0075_),
    .Q_N(_2265_),
    .Q(\counter[25] ));
 sg13g2_dfrbp_1 \counter[26]$_SDFF_PN0_  (.CLK(clknet_4_2_0_clk),
    .RESET_B(net115),
    .D(_0076_),
    .Q_N(_2264_),
    .Q(\counter[26] ));
 sg13g2_dfrbp_1 \counter[27]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net116),
    .D(_0077_),
    .Q_N(_2263_),
    .Q(\counter[27] ));
 sg13g2_dfrbp_1 \counter[28]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net117),
    .D(_0078_),
    .Q_N(_2262_),
    .Q(\counter[28] ));
 sg13g2_dfrbp_1 \counter[29]$_SDFF_PN0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net118),
    .D(_0079_),
    .Q_N(_2261_),
    .Q(\counter[29] ));
 sg13g2_dfrbp_1 \counter[2]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net119),
    .D(_0080_),
    .Q_N(_2260_),
    .Q(\counter[2] ));
 sg13g2_dfrbp_1 \counter[30]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net120),
    .D(_0081_),
    .Q_N(_2259_),
    .Q(\counter[30] ));
 sg13g2_dfrbp_1 \counter[31]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net121),
    .D(_0082_),
    .Q_N(_2258_),
    .Q(\counter[31] ));
 sg13g2_dfrbp_1 \counter[3]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net122),
    .D(_0083_),
    .Q_N(_2257_),
    .Q(\counter[3] ));
 sg13g2_dfrbp_1 \counter[4]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net123),
    .D(_0084_),
    .Q_N(_2256_),
    .Q(\counter[4] ));
 sg13g2_dfrbp_1 \counter[5]$_SDFF_PN0_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net124),
    .D(_0085_),
    .Q_N(_2255_),
    .Q(\counter[5] ));
 sg13g2_dfrbp_1 \counter[6]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net125),
    .D(_0086_),
    .Q_N(_2254_),
    .Q(\counter[6] ));
 sg13g2_dfrbp_1 \counter[7]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net126),
    .D(_0087_),
    .Q_N(_2253_),
    .Q(\counter[7] ));
 sg13g2_dfrbp_1 \counter[8]$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net127),
    .D(_0088_),
    .Q_N(_2252_),
    .Q(\counter[8] ));
 sg13g2_dfrbp_1 \counter[9]$_SDFF_PN0_  (.CLK(clknet_4_1_0_clk),
    .RESET_B(net128),
    .D(_0089_),
    .Q_N(_2288_),
    .Q(\counter[9] ));
 sg13g2_dfrbp_1 \depth[0]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net129),
    .D(_0005_),
    .Q_N(_2289_),
    .Q(\depth[0] ));
 sg13g2_dfrbp_1 \depth[1]$_DFF_P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net130),
    .D(_0006_),
    .Q_N(_2290_),
    .Q(\depth[1] ));
 sg13g2_dfrbp_1 \depth[2]$_DFF_P_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net131),
    .D(_0007_),
    .Q_N(_0046_),
    .Q(\depth[2] ));
 sg13g2_dfrbp_1 \dither_threshold[0]$_SDFFE_PP0P_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net132),
    .D(_0090_),
    .Q_N(_0026_),
    .Q(\dither_threshold[0] ));
 sg13g2_dfrbp_1 \dither_threshold[1]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net133),
    .D(_0091_),
    .Q_N(_0031_),
    .Q(\dither_threshold[1] ));
 sg13g2_dfrbp_1 \dither_threshold[2]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net134),
    .D(_0092_),
    .Q_N(_2251_),
    .Q(\dither_threshold[2] ));
 sg13g2_dfrbp_1 \dither_threshold[3]$_SDFF_PP0_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net135),
    .D(_0093_),
    .Q_N(_0032_),
    .Q(\dither_threshold[3] ));
 sg13g2_dfrbp_1 \dither_threshold[4]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net136),
    .D(_0094_),
    .Q_N(_0033_),
    .Q(\dither_threshold[4] ));
 sg13g2_dfrbp_1 \dither_threshold[5]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net137),
    .D(_0095_),
    .Q_N(_0034_),
    .Q(\dither_threshold[5] ));
 sg13g2_dfrbp_1 \dither_threshold[6]$_SDFF_PP0_  (.CLK(clknet_4_5_0_clk),
    .RESET_B(net138),
    .D(_0096_),
    .Q_N(_0035_),
    .Q(\dither_threshold[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[2]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net139),
    .D(_0003_),
    .Q_N(_2250_),
    .Q(\i_project.controller_0.divider[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[3]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net140),
    .D(_0004_),
    .Q_N(_2249_),
    .Q(\i_project.controller_0.divider[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[4]$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net141),
    .D(_0097_),
    .Q_N(_2248_),
    .Q(\i_project.controller_0.mode[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[5]$_DFFE_PN_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net142),
    .D(_0098_),
    .Q_N(_2247_),
    .Q(\i_project.controller_0.mode[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[6]$_DFFE_PN_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net143),
    .D(_0099_),
    .Q_N(_0025_),
    .Q(\i_project.controller_0.mode[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.mode_params[7]$_DFFE_PN_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net144),
    .D(_0100_),
    .Q_N(_0022_),
    .Q(\i_project.controller_0.vga_sync.mode ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[0]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net145),
    .D(_0101_),
    .Q_N(_0056_),
    .Q(\i_project.controller_0.mode_ramp_base[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[10]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net146),
    .D(_0102_),
    .Q_N(_0019_),
    .Q(\i_project.controller_0.t[10] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[11]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net147),
    .D(_0103_),
    .Q_N(_2246_),
    .Q(\i_project.controller_0.t[11] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[1]$_SDFFE_PN0P_  (.CLK(clknet_4_4_0_clk),
    .RESET_B(net148),
    .D(_0104_),
    .Q_N(_0021_),
    .Q(\i_project.controller_0.mode_ramp_base[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[2]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net149),
    .D(_0105_),
    .Q_N(_0045_),
    .Q(\i_project.controller_0.mode_ramp_base[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[3]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net150),
    .D(_0106_),
    .Q_N(_0044_),
    .Q(\i_project.controller_0.mode_ramp_base[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[4]$_SDFFE_PN0P_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net151),
    .D(_0107_),
    .Q_N(_0043_),
    .Q(\i_project.controller_0.mode_ramp_base[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[5]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net152),
    .D(_0108_),
    .Q_N(_0042_),
    .Q(\i_project.controller_0.mode_ramp_base[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[6]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net153),
    .D(_0109_),
    .Q_N(_0041_),
    .Q(\i_project.controller_0.mode_ramp_base[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[7]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net154),
    .D(_0110_),
    .Q_N(_0040_),
    .Q(\i_project.controller_0.mode_ramp_base[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[8]$_SDFFE_PN0P_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net155),
    .D(_0111_),
    .Q_N(_0039_),
    .Q(\i_project.controller_0.t[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.t[9]$_SDFFE_PN0P_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net156),
    .D(_0112_),
    .Q_N(_0020_),
    .Q(\i_project.controller_0.t[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net157),
    .D(_0113_),
    .Q_N(_0054_),
    .Q(\i_project.controller_0.h[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net158),
    .D(_0114_),
    .Q_N(_0038_),
    .Q(\i_project.controller_0.h[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net159),
    .D(_0115_),
    .Q_N(_0037_),
    .Q(\i_project.controller_0.h[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0_  (.CLK(clknet_4_9_0_clk),
    .RESET_B(net160),
    .D(_0116_),
    .Q_N(_0024_),
    .Q(\i_project.controller_0.h[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net161),
    .D(_0117_),
    .Q_N(_0053_),
    .Q(\i_project.controller_0.h[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0_  (.CLK(clknet_4_8_0_clk),
    .RESET_B(net162),
    .D(_0118_),
    .Q_N(_0051_),
    .Q(\i_project.controller_0.h[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net163),
    .D(_0119_),
    .Q_N(_0048_),
    .Q(\i_project.controller_0.h[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net164),
    .D(_0120_),
    .Q_N(_0023_),
    .Q(\i_project.controller_0.h[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net165),
    .D(_0121_),
    .Q_N(_0027_),
    .Q(\i_project.controller_0.h[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net166),
    .D(_0122_),
    .Q_N(_0049_),
    .Q(\i_project.controller_0.h[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.hsync$_DFFE_PP_  (.CLK(clknet_4_10_0_clk),
    .RESET_B(net167),
    .D(_0123_),
    .Q_N(hsync),
    .Q(\i_project.controller_0.vga_sync.hsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net168),
    .D(_0124_),
    .Q_N(_2245_),
    .Q(\i_project.controller_0.v[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net169),
    .D(_0125_),
    .Q_N(_2244_),
    .Q(\i_project.controller_0.v[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net170),
    .D(_0126_),
    .Q_N(_2243_),
    .Q(\i_project.controller_0.v[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net171),
    .D(_0127_),
    .Q_N(_2242_),
    .Q(\i_project.controller_0.v[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net172),
    .D(_0128_),
    .Q_N(_2241_),
    .Q(\i_project.controller_0.v[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net173),
    .D(_0129_),
    .Q_N(_0029_),
    .Q(\i_project.controller_0.v[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net174),
    .D(_0130_),
    .Q_N(_2240_),
    .Q(\i_project.controller_0.v[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net175),
    .D(_0131_),
    .Q_N(_2239_),
    .Q(\i_project.controller_0.v[7] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P_  (.CLK(clknet_4_14_0_clk),
    .RESET_B(net176),
    .D(_0132_),
    .Q_N(_0030_),
    .Q(\i_project.controller_0.v[8] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net177),
    .D(_0133_),
    .Q_N(_0028_),
    .Q(\i_project.controller_0.v[9] ));
 sg13g2_dfrbp_1 \i_project.controller_0.vga_sync.vsync$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net178),
    .D(_0134_),
    .Q_N(_2238_),
    .Q(\i_project.controller_0.vga_sync.vsync ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[0]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net179),
    .D(_0135_),
    .Q_N(_2237_),
    .Q(\i_project.controller_0.voffset[0] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[1]$_DFFE_PP_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net180),
    .D(_0136_),
    .Q_N(_2236_),
    .Q(\i_project.controller_0.voffset[1] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[2]$_DFFE_PP_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net181),
    .D(_0137_),
    .Q_N(_2235_),
    .Q(\i_project.controller_0.voffset[2] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[3]$_SDFFCE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net182),
    .D(_0138_),
    .Q_N(_2234_),
    .Q(\i_project.controller_0.voffset[3] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[4]$_SDFFCE_PP0P_  (.CLK(clknet_4_12_0_clk),
    .RESET_B(net183),
    .D(_0139_),
    .Q_N(_2233_),
    .Q(\i_project.controller_0.voffset[4] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[5]$_DFFE_PP_  (.CLK(clknet_4_15_0_clk),
    .RESET_B(net184),
    .D(_0140_),
    .Q_N(_2232_),
    .Q(\i_project.controller_0.voffset[5] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[6]$_DFFE_PP_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net185),
    .D(_0141_),
    .Q_N(_2231_),
    .Q(\i_project.controller_0.voffset[6] ));
 sg13g2_dfrbp_1 \i_project.controller_0.voffset[7]$_SDFFCE_PN0P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net186),
    .D(_0142_),
    .Q_N(_2230_),
    .Q(\i_project.controller_0.voffset[7] ));
 sg13g2_dfrbp_1 \prev_vsync$_SDFF_PN0_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net187),
    .D(_0143_),
    .Q_N(_2291_),
    .Q(prev_vsync));
 sg13g2_dfrbp_1 \project_rst_n$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net188),
    .D(_0008_),
    .Q_N(_2292_),
    .Q(\i_project.controller_0.rst_n ));
 sg13g2_dfrbp_1 \project_ui_in[2]$_DFF_P_  (.CLK(clknet_4_0_0_clk),
    .RESET_B(net189),
    .D(\counter[30] ),
    .Q_N(_0018_),
    .Q(\i_project.controller_0.grey_pass[10] ));
 sg13g2_dfrbp_1 \project_ui_in[3]$_DFF_P_  (.CLK(clknet_4_6_0_clk),
    .RESET_B(net190),
    .D(\counter[31] ),
    .Q_N(_0017_),
    .Q(\i_project.controller_0.grey_pass[11] ));
 sg13g2_dfrbp_1 \project_ui_in[4]$_DFF_P_  (.CLK(clknet_4_11_0_clk),
    .RESET_B(net191),
    .D(_0009_),
    .Q_N(_0052_),
    .Q(\i_project.controller_0.grey_pass[12] ));
 sg13g2_dfrbp_1 \project_ui_in[5]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net192),
    .D(_0010_),
    .Q_N(_0050_),
    .Q(\i_project.controller_0.grey_pass[13] ));
 sg13g2_dfrbp_1 \project_ui_in[6]$_DFF_P_  (.CLK(clknet_4_13_0_clk),
    .RESET_B(net193),
    .D(_0011_),
    .Q_N(_0047_),
    .Q(\i_project.controller_0.grey_pass[14] ));
 sg13g2_dfrbp_1 \project_ui_in[7]$_SDFF_PN0_  (.CLK(clknet_4_7_0_clk),
    .RESET_B(net194),
    .D(_0144_),
    .Q_N(_0036_),
    .Q(\i_project.controller_0.grey_pass[15] ));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 output8 (.A(net8),
    .X(uo_out[0]));
 sg13g2_buf_1 output9 (.A(net9),
    .X(uo_out[1]));
 sg13g2_buf_1 output10 (.A(net10),
    .X(uo_out[2]));
 sg13g2_buf_1 output11 (.A(net11),
    .X(uo_out[3]));
 sg13g2_buf_1 output12 (.A(net12),
    .X(uo_out[4]));
 sg13g2_buf_1 output13 (.A(net13),
    .X(uo_out[5]));
 sg13g2_buf_1 output14 (.A(net14),
    .X(uo_out[6]));
 sg13g2_buf_1 output15 (.A(net15),
    .X(uo_out[7]));
 sg13g2_buf_2 fanout16 (.A(_1486_),
    .X(net16));
 sg13g2_buf_2 fanout17 (.A(_0289_),
    .X(net17));
 sg13g2_buf_2 fanout18 (.A(_0168_),
    .X(net18));
 sg13g2_buf_2 fanout19 (.A(_2206_),
    .X(net19));
 sg13g2_buf_2 fanout20 (.A(_2133_),
    .X(net20));
 sg13g2_buf_2 fanout21 (.A(_1914_),
    .X(net21));
 sg13g2_buf_2 fanout22 (.A(_0161_),
    .X(net22));
 sg13g2_buf_2 fanout23 (.A(_0554_),
    .X(net23));
 sg13g2_buf_2 fanout24 (.A(_0511_),
    .X(net24));
 sg13g2_buf_2 fanout25 (.A(_0365_),
    .X(net25));
 sg13g2_buf_2 fanout26 (.A(_0282_),
    .X(net26));
 sg13g2_buf_2 fanout27 (.A(_0263_),
    .X(net27));
 sg13g2_buf_2 fanout28 (.A(_0804_),
    .X(net28));
 sg13g2_buf_2 fanout29 (.A(_0352_),
    .X(net29));
 sg13g2_buf_2 fanout30 (.A(_0541_),
    .X(net30));
 sg13g2_buf_2 fanout31 (.A(_0493_),
    .X(net31));
 sg13g2_buf_2 fanout32 (.A(_0483_),
    .X(net32));
 sg13g2_buf_2 fanout33 (.A(_0351_),
    .X(net33));
 sg13g2_buf_2 fanout34 (.A(_0256_),
    .X(net34));
 sg13g2_buf_2 fanout35 (.A(_2217_),
    .X(net35));
 sg13g2_buf_2 fanout36 (.A(_0364_),
    .X(net36));
 sg13g2_buf_2 fanout37 (.A(_0337_),
    .X(net37));
 sg13g2_buf_2 fanout38 (.A(_0320_),
    .X(net38));
 sg13g2_buf_2 fanout39 (.A(_0317_),
    .X(net39));
 sg13g2_buf_2 fanout40 (.A(_0299_),
    .X(net40));
 sg13g2_buf_2 fanout41 (.A(_0258_),
    .X(net41));
 sg13g2_buf_2 fanout42 (.A(_0225_),
    .X(net42));
 sg13g2_buf_2 fanout43 (.A(_2092_),
    .X(net43));
 sg13g2_buf_2 fanout44 (.A(_2037_),
    .X(net44));
 sg13g2_buf_2 fanout45 (.A(_0540_),
    .X(net45));
 sg13g2_buf_2 fanout46 (.A(_0329_),
    .X(net46));
 sg13g2_buf_2 fanout47 (.A(_2110_),
    .X(net47));
 sg13g2_buf_2 fanout48 (.A(_1836_),
    .X(net48));
 sg13g2_buf_2 fanout49 (.A(_1816_),
    .X(net49));
 sg13g2_buf_2 fanout50 (.A(_1691_),
    .X(net50));
 sg13g2_buf_2 fanout51 (.A(_0308_),
    .X(net51));
 sg13g2_buf_2 fanout52 (.A(_0238_),
    .X(net52));
 sg13g2_buf_2 fanout53 (.A(_2046_),
    .X(net53));
 sg13g2_buf_2 fanout54 (.A(_2043_),
    .X(net54));
 sg13g2_buf_2 fanout55 (.A(_2007_),
    .X(net55));
 sg13g2_buf_2 fanout56 (.A(_1989_),
    .X(net56));
 sg13g2_buf_2 fanout57 (.A(_1733_),
    .X(net57));
 sg13g2_buf_2 fanout58 (.A(_1725_),
    .X(net58));
 sg13g2_buf_2 fanout59 (.A(_1724_),
    .X(net59));
 sg13g2_buf_2 fanout60 (.A(_1713_),
    .X(net60));
 sg13g2_buf_2 fanout61 (.A(_1707_),
    .X(net61));
 sg13g2_buf_2 fanout62 (.A(_1685_),
    .X(net62));
 sg13g2_buf_2 fanout63 (.A(_2055_),
    .X(net63));
 sg13g2_buf_2 fanout64 (.A(_2050_),
    .X(net64));
 sg13g2_buf_2 fanout65 (.A(_2048_),
    .X(net65));
 sg13g2_buf_2 fanout66 (.A(_2041_),
    .X(net66));
 sg13g2_buf_2 fanout67 (.A(_1768_),
    .X(net67));
 sg13g2_buf_2 fanout68 (.A(_1764_),
    .X(net68));
 sg13g2_buf_2 fanout69 (.A(_1748_),
    .X(net69));
 sg13g2_buf_2 fanout70 (.A(_1737_),
    .X(net70));
 sg13g2_buf_2 fanout71 (.A(_1714_),
    .X(net71));
 sg13g2_buf_2 fanout72 (.A(_1703_),
    .X(net72));
 sg13g2_buf_2 fanout73 (.A(_1669_),
    .X(net73));
 sg13g2_buf_2 fanout74 (.A(_1693_),
    .X(net74));
 sg13g2_tielo _4502__75 (.L_LO(net75));
 sg13g2_tielo _4503__76 (.L_LO(net76));
 sg13g2_tielo _4504__77 (.L_LO(net77));
 sg13g2_tielo _4505__78 (.L_LO(net78));
 sg13g2_tielo _4506__79 (.L_LO(net79));
 sg13g2_tielo _4507__80 (.L_LO(net80));
 sg13g2_tielo _4508__81 (.L_LO(net81));
 sg13g2_tielo _4509__82 (.L_LO(net82));
 sg13g2_tiehi _4487__84 (.L_HI(net84));
 sg13g2_tiehi _4488__85 (.L_HI(net85));
 sg13g2_tiehi _4489__86 (.L_HI(net86));
 sg13g2_tiehi _4490__87 (.L_HI(net87));
 sg13g2_tiehi _4491__88 (.L_HI(net88));
 sg13g2_tiehi _4494__89 (.L_HI(net89));
 sg13g2_tiehi _4495__90 (.L_HI(net90));
 sg13g2_tiehi _4496__91 (.L_HI(net91));
 sg13g2_tiehi _4497__92 (.L_HI(net92));
 sg13g2_tiehi _4498__93 (.L_HI(net93));
 sg13g2_tiehi _4499__94 (.L_HI(net94));
 sg13g2_tiehi _4500__95 (.L_HI(net95));
 sg13g2_tiehi _4501__96 (.L_HI(net96));
 sg13g2_tiehi \counter[0]$_SDFF_PN0__97  (.L_HI(net97));
 sg13g2_tiehi \counter[10]$_SDFF_PN0__98  (.L_HI(net98));
 sg13g2_tiehi \counter[11]$_SDFF_PN0__99  (.L_HI(net99));
 sg13g2_tiehi \counter[12]$_SDFF_PN0__100  (.L_HI(net100));
 sg13g2_tiehi \counter[13]$_SDFF_PN0__101  (.L_HI(net101));
 sg13g2_tiehi \counter[14]$_SDFF_PN0__102  (.L_HI(net102));
 sg13g2_tiehi \counter[15]$_SDFF_PN0__103  (.L_HI(net103));
 sg13g2_tiehi \counter[16]$_SDFF_PN0__104  (.L_HI(net104));
 sg13g2_tiehi \counter[17]$_SDFF_PN0__105  (.L_HI(net105));
 sg13g2_tiehi \counter[18]$_SDFF_PN0__106  (.L_HI(net106));
 sg13g2_tiehi \counter[19]$_SDFF_PN0__107  (.L_HI(net107));
 sg13g2_tiehi \counter[1]$_SDFF_PN0__108  (.L_HI(net108));
 sg13g2_tiehi \counter[20]$_SDFF_PN0__109  (.L_HI(net109));
 sg13g2_tiehi \counter[21]$_SDFF_PN0__110  (.L_HI(net110));
 sg13g2_tiehi \counter[22]$_SDFF_PN0__111  (.L_HI(net111));
 sg13g2_tiehi \counter[23]$_SDFF_PN0__112  (.L_HI(net112));
 sg13g2_tiehi \counter[24]$_SDFF_PN0__113  (.L_HI(net113));
 sg13g2_tiehi \counter[25]$_SDFF_PN0__114  (.L_HI(net114));
 sg13g2_tiehi \counter[26]$_SDFF_PN0__115  (.L_HI(net115));
 sg13g2_tiehi \counter[27]$_SDFF_PN0__116  (.L_HI(net116));
 sg13g2_tiehi \counter[28]$_SDFF_PN0__117  (.L_HI(net117));
 sg13g2_tiehi \counter[29]$_SDFF_PN0__118  (.L_HI(net118));
 sg13g2_tiehi \counter[2]$_SDFF_PN0__119  (.L_HI(net119));
 sg13g2_tiehi \counter[30]$_SDFF_PN0__120  (.L_HI(net120));
 sg13g2_tiehi \counter[31]$_SDFF_PN0__121  (.L_HI(net121));
 sg13g2_tiehi \counter[3]$_SDFF_PN0__122  (.L_HI(net122));
 sg13g2_tiehi \counter[4]$_SDFF_PN0__123  (.L_HI(net123));
 sg13g2_tiehi \counter[5]$_SDFF_PN0__124  (.L_HI(net124));
 sg13g2_tiehi \counter[6]$_SDFF_PN0__125  (.L_HI(net125));
 sg13g2_tiehi \counter[7]$_SDFF_PN0__126  (.L_HI(net126));
 sg13g2_tiehi \counter[8]$_SDFF_PN0__127  (.L_HI(net127));
 sg13g2_tiehi \counter[9]$_SDFF_PN0__128  (.L_HI(net128));
 sg13g2_tiehi \depth[0]$_DFF_P__129  (.L_HI(net129));
 sg13g2_tiehi \depth[1]$_DFF_P__130  (.L_HI(net130));
 sg13g2_tiehi \depth[2]$_DFF_P__131  (.L_HI(net131));
 sg13g2_tiehi \dither_threshold[0]$_SDFFE_PP0P__132  (.L_HI(net132));
 sg13g2_tiehi \dither_threshold[1]$_SDFF_PP0__133  (.L_HI(net133));
 sg13g2_tiehi \dither_threshold[2]$_SDFF_PP0__134  (.L_HI(net134));
 sg13g2_tiehi \dither_threshold[3]$_SDFF_PP0__135  (.L_HI(net135));
 sg13g2_tiehi \dither_threshold[4]$_SDFF_PP0__136  (.L_HI(net136));
 sg13g2_tiehi \dither_threshold[5]$_SDFF_PP0__137  (.L_HI(net137));
 sg13g2_tiehi \dither_threshold[6]$_SDFF_PP0__138  (.L_HI(net138));
 sg13g2_tiehi \i_project.controller_0.mode_params[2]$_DFFE_PN__139  (.L_HI(net139));
 sg13g2_tiehi \i_project.controller_0.mode_params[3]$_DFFE_PN__140  (.L_HI(net140));
 sg13g2_tiehi \i_project.controller_0.mode_params[4]$_DFFE_PN__141  (.L_HI(net141));
 sg13g2_tiehi \i_project.controller_0.mode_params[5]$_DFFE_PN__142  (.L_HI(net142));
 sg13g2_tiehi \i_project.controller_0.mode_params[6]$_DFFE_PN__143  (.L_HI(net143));
 sg13g2_tiehi \i_project.controller_0.mode_params[7]$_DFFE_PN__144  (.L_HI(net144));
 sg13g2_tiehi \i_project.controller_0.t[0]$_SDFFE_PN0P__145  (.L_HI(net145));
 sg13g2_tiehi \i_project.controller_0.t[10]$_SDFFE_PN0P__146  (.L_HI(net146));
 sg13g2_tiehi \i_project.controller_0.t[11]$_SDFFE_PN0P__147  (.L_HI(net147));
 sg13g2_tiehi \i_project.controller_0.t[1]$_SDFFE_PN0P__148  (.L_HI(net148));
 sg13g2_tiehi \i_project.controller_0.t[2]$_SDFFE_PN0P__149  (.L_HI(net149));
 sg13g2_tiehi \i_project.controller_0.t[3]$_SDFFE_PN0P__150  (.L_HI(net150));
 sg13g2_tiehi \i_project.controller_0.t[4]$_SDFFE_PN0P__151  (.L_HI(net151));
 sg13g2_tiehi \i_project.controller_0.t[5]$_SDFFE_PN0P__152  (.L_HI(net152));
 sg13g2_tiehi \i_project.controller_0.t[6]$_SDFFE_PN0P__153  (.L_HI(net153));
 sg13g2_tiehi \i_project.controller_0.t[7]$_SDFFE_PN0P__154  (.L_HI(net154));
 sg13g2_tiehi \i_project.controller_0.t[8]$_SDFFE_PN0P__155  (.L_HI(net155));
 sg13g2_tiehi \i_project.controller_0.t[9]$_SDFFE_PN0P__156  (.L_HI(net156));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[0]$_SDFF_PP0__157  (.L_HI(net157));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[1]$_SDFF_PP0__158  (.L_HI(net158));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[2]$_SDFF_PP0__159  (.L_HI(net159));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[3]$_SDFF_PP0__160  (.L_HI(net160));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[4]$_SDFF_PP0__161  (.L_HI(net161));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[5]$_SDFF_PP0__162  (.L_HI(net162));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[6]$_SDFF_PP0__163  (.L_HI(net163));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[7]$_SDFF_PP0__164  (.L_HI(net164));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[8]$_SDFF_PP0__165  (.L_HI(net165));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hpos[9]$_SDFF_PP0__166  (.L_HI(net166));
 sg13g2_tiehi \i_project.controller_0.vga_sync.hsync$_DFFE_PP__167  (.L_HI(net167));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[0]$_SDFFE_PP0P__168  (.L_HI(net168));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[1]$_SDFFE_PP0P__169  (.L_HI(net169));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[2]$_SDFFE_PP0P__170  (.L_HI(net170));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[3]$_SDFFE_PP0P__171  (.L_HI(net171));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[4]$_SDFFE_PP0P__172  (.L_HI(net172));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[5]$_SDFFE_PP0P__173  (.L_HI(net173));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[6]$_SDFFE_PP0P__174  (.L_HI(net174));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[7]$_SDFFE_PP0P__175  (.L_HI(net175));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[8]$_SDFFE_PP0P__176  (.L_HI(net176));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vpos[9]$_SDFFE_PP0P__177  (.L_HI(net177));
 sg13g2_tiehi \i_project.controller_0.vga_sync.vsync$_DFFE_PP__178  (.L_HI(net178));
 sg13g2_tiehi \i_project.controller_0.voffset[0]$_DFFE_PP__179  (.L_HI(net179));
 sg13g2_tiehi \i_project.controller_0.voffset[1]$_DFFE_PP__180  (.L_HI(net180));
 sg13g2_tiehi \i_project.controller_0.voffset[2]$_DFFE_PP__181  (.L_HI(net181));
 sg13g2_tiehi \i_project.controller_0.voffset[3]$_SDFFCE_PP0P__182  (.L_HI(net182));
 sg13g2_tiehi \i_project.controller_0.voffset[4]$_SDFFCE_PP0P__183  (.L_HI(net183));
 sg13g2_tiehi \i_project.controller_0.voffset[5]$_DFFE_PP__184  (.L_HI(net184));
 sg13g2_tiehi \i_project.controller_0.voffset[6]$_DFFE_PP__185  (.L_HI(net185));
 sg13g2_tiehi \i_project.controller_0.voffset[7]$_SDFFCE_PN0P__186  (.L_HI(net186));
 sg13g2_tiehi \prev_vsync$_SDFF_PN0__187  (.L_HI(net187));
 sg13g2_tiehi \project_rst_n$_DFF_P__188  (.L_HI(net188));
 sg13g2_tiehi \project_ui_in[2]$_DFF_P__189  (.L_HI(net189));
 sg13g2_tiehi \project_ui_in[3]$_DFF_P__190  (.L_HI(net190));
 sg13g2_tiehi \project_ui_in[4]$_DFF_P__191  (.L_HI(net191));
 sg13g2_tiehi \project_ui_in[5]$_DFF_P__192  (.L_HI(net192));
 sg13g2_tiehi \project_ui_in[6]$_DFF_P__193  (.L_HI(net193));
 sg13g2_tiehi \project_ui_in[7]$_SDFF_PN0__194  (.L_HI(net194));
 sg13g2_buf_2 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_2 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_2 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_2 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_2 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_2 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_2 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_2 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_2 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_2 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_2 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_2 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_2 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_2 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_2 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_2 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_inv_1 clkload0 (.A(clknet_4_1_0_clk));
 sg13g2_inv_1 clkload1 (.A(clknet_4_3_0_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_4_5_0_clk));
 sg13g2_inv_1 clkload3 (.A(clknet_4_7_0_clk));
 sg13g2_inv_1 clkload4 (.A(clknet_4_9_0_clk));
 sg13g2_inv_1 clkload5 (.A(clknet_4_11_0_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_4_13_0_clk));
 sg13g2_inv_1 clkload7 (.A(clknet_4_15_0_clk));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_54 ();
 sg13g2_decap_8 FILLER_0_61 ();
 sg13g2_decap_4 FILLER_0_68 ();
 sg13g2_fill_1 FILLER_0_72 ();
 sg13g2_fill_1 FILLER_0_104 ();
 sg13g2_fill_1 FILLER_0_131 ();
 sg13g2_fill_1 FILLER_0_198 ();
 sg13g2_decap_4 FILLER_0_210 ();
 sg13g2_fill_2 FILLER_0_214 ();
 sg13g2_fill_2 FILLER_0_228 ();
 sg13g2_fill_1 FILLER_0_230 ();
 sg13g2_fill_2 FILLER_0_247 ();
 sg13g2_fill_2 FILLER_0_253 ();
 sg13g2_fill_1 FILLER_0_255 ();
 sg13g2_fill_1 FILLER_0_261 ();
 sg13g2_decap_4 FILLER_0_267 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_fill_2 FILLER_0_280 ();
 sg13g2_fill_1 FILLER_0_282 ();
 sg13g2_fill_1 FILLER_0_295 ();
 sg13g2_fill_2 FILLER_0_326 ();
 sg13g2_decap_8 FILLER_0_358 ();
 sg13g2_decap_4 FILLER_0_365 ();
 sg13g2_fill_2 FILLER_0_369 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_4 FILLER_0_392 ();
 sg13g2_fill_1 FILLER_0_396 ();
 sg13g2_decap_8 FILLER_0_401 ();
 sg13g2_decap_8 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_0_415 ();
 sg13g2_decap_8 FILLER_0_422 ();
 sg13g2_fill_1 FILLER_0_429 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_fill_1 FILLER_1_28 ();
 sg13g2_fill_1 FILLER_1_34 ();
 sg13g2_decap_4 FILLER_1_40 ();
 sg13g2_fill_1 FILLER_1_44 ();
 sg13g2_fill_1 FILLER_1_54 ();
 sg13g2_fill_1 FILLER_1_116 ();
 sg13g2_fill_1 FILLER_1_121 ();
 sg13g2_fill_2 FILLER_1_134 ();
 sg13g2_fill_1 FILLER_1_136 ();
 sg13g2_fill_2 FILLER_1_146 ();
 sg13g2_fill_1 FILLER_1_187 ();
 sg13g2_fill_1 FILLER_1_193 ();
 sg13g2_fill_1 FILLER_1_202 ();
 sg13g2_fill_1 FILLER_1_209 ();
 sg13g2_fill_1 FILLER_1_222 ();
 sg13g2_fill_2 FILLER_1_231 ();
 sg13g2_fill_1 FILLER_1_263 ();
 sg13g2_decap_4 FILLER_1_294 ();
 sg13g2_fill_2 FILLER_1_298 ();
 sg13g2_fill_2 FILLER_1_307 ();
 sg13g2_fill_2 FILLER_1_313 ();
 sg13g2_fill_1 FILLER_1_315 ();
 sg13g2_fill_2 FILLER_1_320 ();
 sg13g2_fill_1 FILLER_1_322 ();
 sg13g2_fill_2 FILLER_1_336 ();
 sg13g2_fill_1 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_fill_1 FILLER_1_350 ();
 sg13g2_fill_1 FILLER_1_429 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_fill_2 FILLER_2_7 ();
 sg13g2_fill_1 FILLER_2_17 ();
 sg13g2_fill_1 FILLER_2_21 ();
 sg13g2_fill_1 FILLER_2_33 ();
 sg13g2_fill_1 FILLER_2_38 ();
 sg13g2_fill_2 FILLER_2_55 ();
 sg13g2_fill_1 FILLER_2_65 ();
 sg13g2_fill_2 FILLER_2_95 ();
 sg13g2_fill_2 FILLER_2_101 ();
 sg13g2_decap_4 FILLER_2_116 ();
 sg13g2_fill_2 FILLER_2_131 ();
 sg13g2_decap_8 FILLER_2_153 ();
 sg13g2_fill_2 FILLER_2_160 ();
 sg13g2_decap_4 FILLER_2_178 ();
 sg13g2_fill_2 FILLER_2_182 ();
 sg13g2_fill_2 FILLER_2_200 ();
 sg13g2_decap_4 FILLER_2_210 ();
 sg13g2_fill_1 FILLER_2_214 ();
 sg13g2_fill_1 FILLER_2_220 ();
 sg13g2_fill_1 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_234 ();
 sg13g2_fill_1 FILLER_2_243 ();
 sg13g2_fill_1 FILLER_2_255 ();
 sg13g2_fill_2 FILLER_2_260 ();
 sg13g2_fill_1 FILLER_2_266 ();
 sg13g2_decap_4 FILLER_2_278 ();
 sg13g2_fill_1 FILLER_2_282 ();
 sg13g2_fill_2 FILLER_2_329 ();
 sg13g2_fill_1 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_fill_1 FILLER_3_7 ();
 sg13g2_fill_1 FILLER_3_12 ();
 sg13g2_fill_1 FILLER_3_20 ();
 sg13g2_fill_2 FILLER_3_26 ();
 sg13g2_decap_4 FILLER_3_40 ();
 sg13g2_fill_1 FILLER_3_44 ();
 sg13g2_fill_1 FILLER_3_59 ();
 sg13g2_decap_4 FILLER_3_68 ();
 sg13g2_fill_1 FILLER_3_72 ();
 sg13g2_fill_2 FILLER_3_92 ();
 sg13g2_fill_1 FILLER_3_97 ();
 sg13g2_decap_4 FILLER_3_119 ();
 sg13g2_fill_2 FILLER_3_123 ();
 sg13g2_fill_1 FILLER_3_137 ();
 sg13g2_fill_2 FILLER_3_143 ();
 sg13g2_fill_2 FILLER_3_153 ();
 sg13g2_fill_2 FILLER_3_181 ();
 sg13g2_fill_1 FILLER_3_183 ();
 sg13g2_decap_4 FILLER_3_197 ();
 sg13g2_fill_1 FILLER_3_201 ();
 sg13g2_fill_2 FILLER_3_210 ();
 sg13g2_fill_1 FILLER_3_212 ();
 sg13g2_fill_1 FILLER_3_228 ();
 sg13g2_fill_2 FILLER_3_254 ();
 sg13g2_fill_1 FILLER_3_268 ();
 sg13g2_decap_4 FILLER_3_283 ();
 sg13g2_fill_1 FILLER_3_287 ();
 sg13g2_fill_2 FILLER_3_316 ();
 sg13g2_fill_1 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_324 ();
 sg13g2_decap_8 FILLER_3_331 ();
 sg13g2_decap_4 FILLER_3_338 ();
 sg13g2_fill_2 FILLER_3_342 ();
 sg13g2_decap_4 FILLER_3_351 ();
 sg13g2_fill_1 FILLER_3_368 ();
 sg13g2_fill_1 FILLER_3_382 ();
 sg13g2_fill_2 FILLER_3_409 ();
 sg13g2_fill_1 FILLER_3_415 ();
 sg13g2_decap_4 FILLER_3_424 ();
 sg13g2_fill_2 FILLER_3_428 ();
 sg13g2_decap_4 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_4 ();
 sg13g2_fill_1 FILLER_4_25 ();
 sg13g2_fill_1 FILLER_4_30 ();
 sg13g2_fill_1 FILLER_4_47 ();
 sg13g2_fill_2 FILLER_4_74 ();
 sg13g2_fill_2 FILLER_4_85 ();
 sg13g2_fill_1 FILLER_4_87 ();
 sg13g2_fill_2 FILLER_4_93 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_101 ();
 sg13g2_fill_2 FILLER_4_116 ();
 sg13g2_fill_1 FILLER_4_130 ();
 sg13g2_fill_2 FILLER_4_135 ();
 sg13g2_fill_1 FILLER_4_150 ();
 sg13g2_fill_2 FILLER_4_159 ();
 sg13g2_fill_1 FILLER_4_164 ();
 sg13g2_fill_2 FILLER_4_173 ();
 sg13g2_fill_1 FILLER_4_175 ();
 sg13g2_fill_2 FILLER_4_200 ();
 sg13g2_fill_1 FILLER_4_207 ();
 sg13g2_fill_2 FILLER_4_213 ();
 sg13g2_decap_4 FILLER_4_224 ();
 sg13g2_fill_2 FILLER_4_228 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_244 ();
 sg13g2_decap_4 FILLER_4_253 ();
 sg13g2_fill_2 FILLER_4_262 ();
 sg13g2_decap_4 FILLER_4_280 ();
 sg13g2_fill_2 FILLER_4_284 ();
 sg13g2_fill_1 FILLER_4_302 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_fill_1 FILLER_4_338 ();
 sg13g2_fill_2 FILLER_4_356 ();
 sg13g2_fill_1 FILLER_4_366 ();
 sg13g2_fill_1 FILLER_4_373 ();
 sg13g2_fill_1 FILLER_4_378 ();
 sg13g2_fill_1 FILLER_4_382 ();
 sg13g2_fill_1 FILLER_4_392 ();
 sg13g2_fill_2 FILLER_4_404 ();
 sg13g2_decap_8 FILLER_4_419 ();
 sg13g2_decap_4 FILLER_4_426 ();
 sg13g2_fill_2 FILLER_5_0 ();
 sg13g2_fill_1 FILLER_5_38 ();
 sg13g2_fill_2 FILLER_5_59 ();
 sg13g2_fill_1 FILLER_5_66 ();
 sg13g2_fill_2 FILLER_5_72 ();
 sg13g2_fill_1 FILLER_5_78 ();
 sg13g2_fill_2 FILLER_5_83 ();
 sg13g2_fill_2 FILLER_5_88 ();
 sg13g2_fill_2 FILLER_5_116 ();
 sg13g2_fill_1 FILLER_5_123 ();
 sg13g2_fill_1 FILLER_5_129 ();
 sg13g2_fill_1 FILLER_5_186 ();
 sg13g2_decap_4 FILLER_5_191 ();
 sg13g2_fill_2 FILLER_5_195 ();
 sg13g2_fill_1 FILLER_5_213 ();
 sg13g2_decap_4 FILLER_5_222 ();
 sg13g2_fill_1 FILLER_5_226 ();
 sg13g2_decap_4 FILLER_5_248 ();
 sg13g2_fill_1 FILLER_5_279 ();
 sg13g2_fill_2 FILLER_5_308 ();
 sg13g2_fill_1 FILLER_5_326 ();
 sg13g2_fill_1 FILLER_5_340 ();
 sg13g2_fill_1 FILLER_5_345 ();
 sg13g2_fill_1 FILLER_5_351 ();
 sg13g2_fill_1 FILLER_5_356 ();
 sg13g2_fill_1 FILLER_5_380 ();
 sg13g2_fill_1 FILLER_5_398 ();
 sg13g2_decap_4 FILLER_6_0 ();
 sg13g2_fill_2 FILLER_6_4 ();
 sg13g2_fill_1 FILLER_6_14 ();
 sg13g2_fill_1 FILLER_6_23 ();
 sg13g2_fill_1 FILLER_6_42 ();
 sg13g2_fill_1 FILLER_6_55 ();
 sg13g2_fill_1 FILLER_6_64 ();
 sg13g2_decap_4 FILLER_6_70 ();
 sg13g2_fill_1 FILLER_6_83 ();
 sg13g2_fill_1 FILLER_6_101 ();
 sg13g2_fill_2 FILLER_6_107 ();
 sg13g2_fill_2 FILLER_6_116 ();
 sg13g2_fill_1 FILLER_6_118 ();
 sg13g2_decap_8 FILLER_6_143 ();
 sg13g2_fill_2 FILLER_6_150 ();
 sg13g2_fill_1 FILLER_6_152 ();
 sg13g2_fill_2 FILLER_6_165 ();
 sg13g2_fill_1 FILLER_6_172 ();
 sg13g2_fill_1 FILLER_6_221 ();
 sg13g2_fill_2 FILLER_6_226 ();
 sg13g2_fill_1 FILLER_6_232 ();
 sg13g2_fill_2 FILLER_6_237 ();
 sg13g2_fill_2 FILLER_6_243 ();
 sg13g2_fill_2 FILLER_6_250 ();
 sg13g2_fill_1 FILLER_6_252 ();
 sg13g2_fill_2 FILLER_6_259 ();
 sg13g2_fill_1 FILLER_6_261 ();
 sg13g2_fill_2 FILLER_6_266 ();
 sg13g2_fill_1 FILLER_6_275 ();
 sg13g2_decap_4 FILLER_6_280 ();
 sg13g2_fill_1 FILLER_6_284 ();
 sg13g2_fill_1 FILLER_6_301 ();
 sg13g2_decap_4 FILLER_6_316 ();
 sg13g2_fill_2 FILLER_6_324 ();
 sg13g2_fill_1 FILLER_6_326 ();
 sg13g2_decap_4 FILLER_6_332 ();
 sg13g2_fill_2 FILLER_6_336 ();
 sg13g2_fill_2 FILLER_6_355 ();
 sg13g2_fill_2 FILLER_6_369 ();
 sg13g2_fill_1 FILLER_6_371 ();
 sg13g2_fill_1 FILLER_6_409 ();
 sg13g2_decap_8 FILLER_6_423 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_37 ();
 sg13g2_fill_2 FILLER_7_41 ();
 sg13g2_fill_1 FILLER_7_47 ();
 sg13g2_fill_2 FILLER_7_60 ();
 sg13g2_fill_1 FILLER_7_62 ();
 sg13g2_fill_1 FILLER_7_78 ();
 sg13g2_fill_1 FILLER_7_87 ();
 sg13g2_fill_2 FILLER_7_120 ();
 sg13g2_fill_2 FILLER_7_138 ();
 sg13g2_fill_1 FILLER_7_140 ();
 sg13g2_fill_1 FILLER_7_152 ();
 sg13g2_fill_1 FILLER_7_178 ();
 sg13g2_decap_4 FILLER_7_199 ();
 sg13g2_fill_2 FILLER_7_203 ();
 sg13g2_fill_1 FILLER_7_232 ();
 sg13g2_decap_8 FILLER_7_249 ();
 sg13g2_fill_1 FILLER_7_256 ();
 sg13g2_fill_1 FILLER_7_260 ();
 sg13g2_fill_1 FILLER_7_271 ();
 sg13g2_fill_2 FILLER_7_286 ();
 sg13g2_fill_1 FILLER_7_321 ();
 sg13g2_decap_4 FILLER_7_331 ();
 sg13g2_decap_4 FILLER_7_343 ();
 sg13g2_fill_2 FILLER_7_365 ();
 sg13g2_fill_1 FILLER_7_367 ();
 sg13g2_fill_2 FILLER_7_371 ();
 sg13g2_fill_1 FILLER_7_380 ();
 sg13g2_decap_4 FILLER_7_426 ();
 sg13g2_fill_1 FILLER_8_0 ();
 sg13g2_decap_4 FILLER_8_9 ();
 sg13g2_fill_2 FILLER_8_36 ();
 sg13g2_fill_2 FILLER_8_58 ();
 sg13g2_fill_1 FILLER_8_74 ();
 sg13g2_fill_1 FILLER_8_79 ();
 sg13g2_fill_1 FILLER_8_88 ();
 sg13g2_fill_1 FILLER_8_97 ();
 sg13g2_fill_1 FILLER_8_106 ();
 sg13g2_fill_1 FILLER_8_124 ();
 sg13g2_decap_4 FILLER_8_129 ();
 sg13g2_fill_2 FILLER_8_133 ();
 sg13g2_decap_4 FILLER_8_148 ();
 sg13g2_fill_2 FILLER_8_167 ();
 sg13g2_fill_1 FILLER_8_169 ();
 sg13g2_fill_2 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_189 ();
 sg13g2_fill_2 FILLER_8_225 ();
 sg13g2_fill_1 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_244 ();
 sg13g2_fill_2 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_decap_8 FILLER_8_262 ();
 sg13g2_decap_4 FILLER_8_269 ();
 sg13g2_fill_2 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_279 ();
 sg13g2_decap_8 FILLER_8_286 ();
 sg13g2_fill_1 FILLER_8_293 ();
 sg13g2_decap_4 FILLER_8_298 ();
 sg13g2_fill_1 FILLER_8_302 ();
 sg13g2_fill_2 FILLER_8_307 ();
 sg13g2_fill_1 FILLER_8_309 ();
 sg13g2_decap_4 FILLER_8_315 ();
 sg13g2_fill_1 FILLER_8_319 ();
 sg13g2_fill_2 FILLER_8_323 ();
 sg13g2_fill_2 FILLER_8_334 ();
 sg13g2_fill_1 FILLER_8_336 ();
 sg13g2_fill_2 FILLER_8_346 ();
 sg13g2_fill_2 FILLER_8_352 ();
 sg13g2_decap_4 FILLER_8_358 ();
 sg13g2_fill_1 FILLER_8_362 ();
 sg13g2_fill_2 FILLER_8_402 ();
 sg13g2_fill_2 FILLER_9_34 ();
 sg13g2_fill_1 FILLER_9_40 ();
 sg13g2_fill_2 FILLER_9_45 ();
 sg13g2_decap_4 FILLER_9_68 ();
 sg13g2_fill_2 FILLER_9_72 ();
 sg13g2_fill_1 FILLER_9_88 ();
 sg13g2_fill_1 FILLER_9_121 ();
 sg13g2_decap_4 FILLER_9_125 ();
 sg13g2_fill_2 FILLER_9_134 ();
 sg13g2_fill_2 FILLER_9_145 ();
 sg13g2_fill_1 FILLER_9_147 ();
 sg13g2_fill_2 FILLER_9_152 ();
 sg13g2_fill_1 FILLER_9_158 ();
 sg13g2_fill_2 FILLER_9_162 ();
 sg13g2_fill_1 FILLER_9_164 ();
 sg13g2_fill_2 FILLER_9_194 ();
 sg13g2_decap_4 FILLER_9_215 ();
 sg13g2_fill_1 FILLER_9_223 ();
 sg13g2_fill_2 FILLER_9_254 ();
 sg13g2_fill_1 FILLER_9_256 ();
 sg13g2_fill_2 FILLER_9_287 ();
 sg13g2_fill_2 FILLER_9_300 ();
 sg13g2_fill_1 FILLER_9_309 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_fill_2 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_366 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_59 ();
 sg13g2_decap_4 FILLER_10_68 ();
 sg13g2_fill_1 FILLER_10_72 ();
 sg13g2_decap_4 FILLER_10_94 ();
 sg13g2_fill_2 FILLER_10_98 ();
 sg13g2_decap_4 FILLER_10_104 ();
 sg13g2_fill_2 FILLER_10_113 ();
 sg13g2_fill_2 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_177 ();
 sg13g2_fill_1 FILLER_10_183 ();
 sg13g2_fill_2 FILLER_10_196 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_1 FILLER_10_203 ();
 sg13g2_fill_2 FILLER_10_209 ();
 sg13g2_fill_2 FILLER_10_215 ();
 sg13g2_fill_1 FILLER_10_217 ();
 sg13g2_fill_1 FILLER_10_261 ();
 sg13g2_fill_2 FILLER_10_276 ();
 sg13g2_decap_4 FILLER_10_287 ();
 sg13g2_fill_1 FILLER_10_337 ();
 sg13g2_fill_1 FILLER_10_356 ();
 sg13g2_fill_1 FILLER_10_367 ();
 sg13g2_fill_2 FILLER_10_415 ();
 sg13g2_fill_2 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_2 ();
 sg13g2_fill_1 FILLER_11_7 ();
 sg13g2_fill_1 FILLER_11_13 ();
 sg13g2_fill_1 FILLER_11_18 ();
 sg13g2_fill_1 FILLER_11_22 ();
 sg13g2_fill_1 FILLER_11_27 ();
 sg13g2_fill_1 FILLER_11_36 ();
 sg13g2_decap_4 FILLER_11_41 ();
 sg13g2_fill_1 FILLER_11_45 ();
 sg13g2_fill_2 FILLER_11_50 ();
 sg13g2_fill_1 FILLER_11_52 ();
 sg13g2_fill_1 FILLER_11_92 ();
 sg13g2_fill_2 FILLER_11_97 ();
 sg13g2_fill_2 FILLER_11_102 ();
 sg13g2_fill_1 FILLER_11_121 ();
 sg13g2_fill_2 FILLER_11_126 ();
 sg13g2_decap_4 FILLER_11_131 ();
 sg13g2_fill_2 FILLER_11_135 ();
 sg13g2_fill_2 FILLER_11_160 ();
 sg13g2_fill_2 FILLER_11_170 ();
 sg13g2_fill_1 FILLER_11_172 ();
 sg13g2_fill_2 FILLER_11_249 ();
 sg13g2_fill_1 FILLER_11_290 ();
 sg13g2_fill_2 FILLER_11_301 ();
 sg13g2_fill_2 FILLER_11_307 ();
 sg13g2_decap_4 FILLER_11_332 ();
 sg13g2_fill_2 FILLER_11_336 ();
 sg13g2_fill_2 FILLER_11_351 ();
 sg13g2_fill_2 FILLER_11_359 ();
 sg13g2_fill_1 FILLER_11_376 ();
 sg13g2_fill_1 FILLER_11_403 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_5 ();
 sg13g2_fill_2 FILLER_12_12 ();
 sg13g2_fill_2 FILLER_12_22 ();
 sg13g2_fill_1 FILLER_12_24 ();
 sg13g2_fill_2 FILLER_12_53 ();
 sg13g2_fill_1 FILLER_12_68 ();
 sg13g2_fill_2 FILLER_12_122 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_136 ();
 sg13g2_fill_1 FILLER_12_140 ();
 sg13g2_fill_1 FILLER_12_146 ();
 sg13g2_fill_1 FILLER_12_152 ();
 sg13g2_fill_1 FILLER_12_169 ();
 sg13g2_decap_4 FILLER_12_174 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_decap_4 FILLER_12_194 ();
 sg13g2_fill_1 FILLER_12_198 ();
 sg13g2_fill_2 FILLER_12_203 ();
 sg13g2_fill_2 FILLER_12_214 ();
 sg13g2_fill_1 FILLER_12_220 ();
 sg13g2_fill_2 FILLER_12_225 ();
 sg13g2_fill_2 FILLER_12_231 ();
 sg13g2_fill_1 FILLER_12_233 ();
 sg13g2_fill_2 FILLER_12_259 ();
 sg13g2_fill_2 FILLER_12_293 ();
 sg13g2_fill_1 FILLER_12_310 ();
 sg13g2_decap_4 FILLER_12_316 ();
 sg13g2_fill_1 FILLER_12_320 ();
 sg13g2_fill_2 FILLER_12_325 ();
 sg13g2_fill_1 FILLER_12_327 ();
 sg13g2_fill_1 FILLER_12_337 ();
 sg13g2_decap_4 FILLER_12_350 ();
 sg13g2_fill_2 FILLER_12_358 ();
 sg13g2_fill_1 FILLER_12_360 ();
 sg13g2_fill_1 FILLER_12_387 ();
 sg13g2_fill_2 FILLER_12_427 ();
 sg13g2_fill_1 FILLER_12_429 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_10 ();
 sg13g2_fill_1 FILLER_13_12 ();
 sg13g2_fill_2 FILLER_13_17 ();
 sg13g2_fill_1 FILLER_13_19 ();
 sg13g2_fill_2 FILLER_13_48 ();
 sg13g2_fill_1 FILLER_13_54 ();
 sg13g2_fill_1 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_173 ();
 sg13g2_fill_1 FILLER_13_179 ();
 sg13g2_fill_2 FILLER_13_185 ();
 sg13g2_fill_2 FILLER_13_212 ();
 sg13g2_decap_4 FILLER_13_221 ();
 sg13g2_fill_2 FILLER_13_225 ();
 sg13g2_fill_1 FILLER_13_273 ();
 sg13g2_fill_1 FILLER_13_281 ();
 sg13g2_fill_1 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_299 ();
 sg13g2_fill_2 FILLER_13_339 ();
 sg13g2_fill_1 FILLER_13_345 ();
 sg13g2_fill_1 FILLER_13_350 ();
 sg13g2_fill_1 FILLER_13_358 ();
 sg13g2_fill_2 FILLER_13_363 ();
 sg13g2_fill_1 FILLER_13_368 ();
 sg13g2_fill_2 FILLER_13_376 ();
 sg13g2_fill_2 FILLER_13_387 ();
 sg13g2_decap_8 FILLER_13_423 ();
 sg13g2_decap_4 FILLER_14_25 ();
 sg13g2_fill_1 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_50 ();
 sg13g2_fill_1 FILLER_14_60 ();
 sg13g2_fill_1 FILLER_14_66 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_fill_1 FILLER_14_84 ();
 sg13g2_fill_1 FILLER_14_92 ();
 sg13g2_fill_1 FILLER_14_97 ();
 sg13g2_fill_1 FILLER_14_101 ();
 sg13g2_fill_2 FILLER_14_110 ();
 sg13g2_fill_1 FILLER_14_120 ();
 sg13g2_decap_8 FILLER_14_125 ();
 sg13g2_fill_1 FILLER_14_149 ();
 sg13g2_fill_1 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_177 ();
 sg13g2_fill_1 FILLER_14_212 ();
 sg13g2_decap_4 FILLER_14_218 ();
 sg13g2_fill_1 FILLER_14_222 ();
 sg13g2_fill_1 FILLER_14_229 ();
 sg13g2_fill_2 FILLER_14_235 ();
 sg13g2_fill_2 FILLER_14_241 ();
 sg13g2_fill_1 FILLER_14_306 ();
 sg13g2_fill_2 FILLER_14_310 ();
 sg13g2_fill_1 FILLER_14_312 ();
 sg13g2_decap_4 FILLER_14_391 ();
 sg13g2_fill_2 FILLER_14_395 ();
 sg13g2_fill_1 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_6 ();
 sg13g2_fill_1 FILLER_15_16 ();
 sg13g2_fill_2 FILLER_15_21 ();
 sg13g2_fill_1 FILLER_15_39 ();
 sg13g2_fill_2 FILLER_15_48 ();
 sg13g2_fill_1 FILLER_15_50 ();
 sg13g2_fill_1 FILLER_15_54 ();
 sg13g2_fill_2 FILLER_15_91 ();
 sg13g2_fill_1 FILLER_15_111 ();
 sg13g2_fill_1 FILLER_15_130 ();
 sg13g2_fill_1 FILLER_15_136 ();
 sg13g2_fill_1 FILLER_15_147 ();
 sg13g2_fill_1 FILLER_15_152 ();
 sg13g2_fill_1 FILLER_15_167 ();
 sg13g2_fill_1 FILLER_15_198 ();
 sg13g2_fill_1 FILLER_15_211 ();
 sg13g2_fill_1 FILLER_15_220 ();
 sg13g2_fill_2 FILLER_15_282 ();
 sg13g2_fill_1 FILLER_15_322 ();
 sg13g2_fill_2 FILLER_15_327 ();
 sg13g2_fill_2 FILLER_15_336 ();
 sg13g2_fill_2 FILLER_15_344 ();
 sg13g2_fill_1 FILLER_15_352 ();
 sg13g2_fill_1 FILLER_15_359 ();
 sg13g2_fill_2 FILLER_15_373 ();
 sg13g2_fill_1 FILLER_15_375 ();
 sg13g2_fill_2 FILLER_15_402 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_fill_1 FILLER_16_47 ();
 sg13g2_fill_2 FILLER_16_65 ();
 sg13g2_fill_1 FILLER_16_82 ();
 sg13g2_fill_2 FILLER_16_93 ();
 sg13g2_fill_1 FILLER_16_95 ();
 sg13g2_fill_2 FILLER_16_101 ();
 sg13g2_fill_1 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_113 ();
 sg13g2_fill_1 FILLER_16_142 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_decap_8 FILLER_16_176 ();
 sg13g2_fill_1 FILLER_16_205 ();
 sg13g2_fill_2 FILLER_16_210 ();
 sg13g2_fill_1 FILLER_16_220 ();
 sg13g2_fill_1 FILLER_16_226 ();
 sg13g2_fill_1 FILLER_16_231 ();
 sg13g2_fill_2 FILLER_16_236 ();
 sg13g2_fill_1 FILLER_16_238 ();
 sg13g2_fill_2 FILLER_16_246 ();
 sg13g2_decap_4 FILLER_16_252 ();
 sg13g2_fill_2 FILLER_16_263 ();
 sg13g2_fill_1 FILLER_16_265 ();
 sg13g2_decap_8 FILLER_16_269 ();
 sg13g2_decap_8 FILLER_16_276 ();
 sg13g2_decap_4 FILLER_16_283 ();
 sg13g2_fill_1 FILLER_16_320 ();
 sg13g2_fill_2 FILLER_16_360 ();
 sg13g2_fill_1 FILLER_16_362 ();
 sg13g2_fill_1 FILLER_16_380 ();
 sg13g2_fill_2 FILLER_16_427 ();
 sg13g2_fill_1 FILLER_16_429 ();
 sg13g2_decap_4 FILLER_17_16 ();
 sg13g2_fill_1 FILLER_17_20 ();
 sg13g2_fill_1 FILLER_17_25 ();
 sg13g2_fill_1 FILLER_17_35 ();
 sg13g2_decap_4 FILLER_17_40 ();
 sg13g2_decap_4 FILLER_17_84 ();
 sg13g2_fill_1 FILLER_17_98 ();
 sg13g2_fill_1 FILLER_17_109 ();
 sg13g2_fill_2 FILLER_17_115 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_130 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_fill_1 FILLER_17_146 ();
 sg13g2_fill_1 FILLER_17_189 ();
 sg13g2_fill_1 FILLER_17_199 ();
 sg13g2_fill_2 FILLER_17_218 ();
 sg13g2_fill_1 FILLER_17_220 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_fill_2 FILLER_17_243 ();
 sg13g2_fill_1 FILLER_17_245 ();
 sg13g2_fill_2 FILLER_17_251 ();
 sg13g2_fill_1 FILLER_17_317 ();
 sg13g2_fill_1 FILLER_17_323 ();
 sg13g2_fill_1 FILLER_17_328 ();
 sg13g2_fill_1 FILLER_17_333 ();
 sg13g2_fill_2 FILLER_17_338 ();
 sg13g2_fill_2 FILLER_17_369 ();
 sg13g2_fill_1 FILLER_17_371 ();
 sg13g2_fill_2 FILLER_17_419 ();
 sg13g2_decap_4 FILLER_17_426 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_14 ();
 sg13g2_fill_2 FILLER_18_20 ();
 sg13g2_fill_1 FILLER_18_22 ();
 sg13g2_decap_4 FILLER_18_48 ();
 sg13g2_fill_2 FILLER_18_52 ();
 sg13g2_fill_2 FILLER_18_63 ();
 sg13g2_fill_1 FILLER_18_65 ();
 sg13g2_fill_1 FILLER_18_74 ();
 sg13g2_fill_1 FILLER_18_104 ();
 sg13g2_fill_1 FILLER_18_115 ();
 sg13g2_fill_2 FILLER_18_143 ();
 sg13g2_fill_1 FILLER_18_149 ();
 sg13g2_fill_2 FILLER_18_168 ();
 sg13g2_fill_1 FILLER_18_208 ();
 sg13g2_fill_1 FILLER_18_214 ();
 sg13g2_fill_1 FILLER_18_220 ();
 sg13g2_fill_1 FILLER_18_225 ();
 sg13g2_fill_2 FILLER_18_233 ();
 sg13g2_decap_8 FILLER_18_240 ();
 sg13g2_fill_2 FILLER_18_247 ();
 sg13g2_fill_2 FILLER_18_290 ();
 sg13g2_fill_2 FILLER_18_311 ();
 sg13g2_fill_1 FILLER_18_313 ();
 sg13g2_fill_1 FILLER_18_328 ();
 sg13g2_fill_2 FILLER_18_336 ();
 sg13g2_fill_2 FILLER_18_364 ();
 sg13g2_fill_2 FILLER_18_381 ();
 sg13g2_fill_2 FILLER_18_387 ();
 sg13g2_fill_1 FILLER_18_389 ();
 sg13g2_fill_1 FILLER_18_394 ();
 sg13g2_fill_2 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_403 ();
 sg13g2_fill_1 FILLER_19_34 ();
 sg13g2_fill_1 FILLER_19_43 ();
 sg13g2_fill_1 FILLER_19_49 ();
 sg13g2_fill_1 FILLER_19_55 ();
 sg13g2_fill_2 FILLER_19_62 ();
 sg13g2_fill_2 FILLER_19_88 ();
 sg13g2_fill_1 FILLER_19_99 ();
 sg13g2_fill_1 FILLER_19_105 ();
 sg13g2_fill_2 FILLER_19_113 ();
 sg13g2_fill_1 FILLER_19_124 ();
 sg13g2_fill_2 FILLER_19_134 ();
 sg13g2_fill_1 FILLER_19_136 ();
 sg13g2_fill_1 FILLER_19_157 ();
 sg13g2_fill_2 FILLER_19_168 ();
 sg13g2_fill_2 FILLER_19_174 ();
 sg13g2_fill_2 FILLER_19_180 ();
 sg13g2_fill_1 FILLER_19_190 ();
 sg13g2_fill_1 FILLER_19_199 ();
 sg13g2_fill_2 FILLER_19_213 ();
 sg13g2_fill_1 FILLER_19_227 ();
 sg13g2_fill_1 FILLER_19_300 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_fill_1 FILLER_19_314 ();
 sg13g2_fill_2 FILLER_19_351 ();
 sg13g2_fill_1 FILLER_19_410 ();
 sg13g2_decap_8 FILLER_19_415 ();
 sg13g2_decap_8 FILLER_19_422 ();
 sg13g2_fill_1 FILLER_19_429 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_11 ();
 sg13g2_fill_1 FILLER_20_31 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_fill_1 FILLER_20_52 ();
 sg13g2_fill_1 FILLER_20_58 ();
 sg13g2_fill_1 FILLER_20_72 ();
 sg13g2_fill_1 FILLER_20_77 ();
 sg13g2_fill_1 FILLER_20_81 ();
 sg13g2_fill_1 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_101 ();
 sg13g2_fill_2 FILLER_20_116 ();
 sg13g2_fill_2 FILLER_20_132 ();
 sg13g2_fill_1 FILLER_20_154 ();
 sg13g2_fill_1 FILLER_20_168 ();
 sg13g2_fill_1 FILLER_20_178 ();
 sg13g2_fill_1 FILLER_20_187 ();
 sg13g2_fill_1 FILLER_20_193 ();
 sg13g2_fill_1 FILLER_20_199 ();
 sg13g2_fill_1 FILLER_20_205 ();
 sg13g2_fill_1 FILLER_20_210 ();
 sg13g2_fill_2 FILLER_20_249 ();
 sg13g2_fill_1 FILLER_20_259 ();
 sg13g2_decap_4 FILLER_20_271 ();
 sg13g2_fill_2 FILLER_20_275 ();
 sg13g2_fill_2 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_297 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_321 ();
 sg13g2_fill_2 FILLER_20_338 ();
 sg13g2_fill_1 FILLER_20_359 ();
 sg13g2_fill_2 FILLER_20_364 ();
 sg13g2_fill_1 FILLER_20_371 ();
 sg13g2_fill_2 FILLER_20_378 ();
 sg13g2_fill_2 FILLER_20_384 ();
 sg13g2_fill_2 FILLER_20_390 ();
 sg13g2_fill_1 FILLER_20_396 ();
 sg13g2_fill_2 FILLER_21_31 ();
 sg13g2_fill_1 FILLER_21_33 ();
 sg13g2_fill_1 FILLER_21_42 ();
 sg13g2_fill_1 FILLER_21_53 ();
 sg13g2_fill_2 FILLER_21_79 ();
 sg13g2_fill_2 FILLER_21_89 ();
 sg13g2_fill_1 FILLER_21_91 ();
 sg13g2_fill_1 FILLER_21_97 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_109 ();
 sg13g2_fill_1 FILLER_21_115 ();
 sg13g2_fill_1 FILLER_21_121 ();
 sg13g2_decap_4 FILLER_21_127 ();
 sg13g2_decap_4 FILLER_21_136 ();
 sg13g2_fill_1 FILLER_21_140 ();
 sg13g2_decap_4 FILLER_21_153 ();
 sg13g2_fill_1 FILLER_21_157 ();
 sg13g2_decap_4 FILLER_21_167 ();
 sg13g2_fill_2 FILLER_21_171 ();
 sg13g2_decap_8 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_184 ();
 sg13g2_fill_1 FILLER_21_188 ();
 sg13g2_fill_2 FILLER_21_205 ();
 sg13g2_decap_4 FILLER_21_220 ();
 sg13g2_fill_2 FILLER_21_271 ();
 sg13g2_fill_1 FILLER_21_273 ();
 sg13g2_fill_1 FILLER_21_293 ();
 sg13g2_fill_2 FILLER_21_364 ();
 sg13g2_fill_2 FILLER_21_408 ();
 sg13g2_fill_1 FILLER_21_410 ();
 sg13g2_decap_8 FILLER_21_415 ();
 sg13g2_fill_1 FILLER_21_422 ();
 sg13g2_fill_2 FILLER_21_427 ();
 sg13g2_fill_1 FILLER_21_429 ();
 sg13g2_fill_1 FILLER_22_26 ();
 sg13g2_fill_1 FILLER_22_31 ();
 sg13g2_fill_2 FILLER_22_36 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_1 FILLER_22_49 ();
 sg13g2_decap_4 FILLER_22_55 ();
 sg13g2_fill_2 FILLER_22_68 ();
 sg13g2_decap_8 FILLER_22_75 ();
 sg13g2_fill_1 FILLER_22_82 ();
 sg13g2_decap_4 FILLER_22_88 ();
 sg13g2_fill_2 FILLER_22_92 ();
 sg13g2_fill_2 FILLER_22_99 ();
 sg13g2_fill_1 FILLER_22_106 ();
 sg13g2_fill_2 FILLER_22_114 ();
 sg13g2_fill_2 FILLER_22_121 ();
 sg13g2_fill_1 FILLER_22_128 ();
 sg13g2_fill_1 FILLER_22_134 ();
 sg13g2_fill_1 FILLER_22_139 ();
 sg13g2_fill_2 FILLER_22_149 ();
 sg13g2_fill_2 FILLER_22_155 ();
 sg13g2_fill_1 FILLER_22_157 ();
 sg13g2_fill_2 FILLER_22_182 ();
 sg13g2_fill_2 FILLER_22_192 ();
 sg13g2_fill_2 FILLER_22_198 ();
 sg13g2_fill_2 FILLER_22_204 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_222 ();
 sg13g2_decap_8 FILLER_22_227 ();
 sg13g2_decap_4 FILLER_22_238 ();
 sg13g2_fill_1 FILLER_22_258 ();
 sg13g2_fill_1 FILLER_22_290 ();
 sg13g2_fill_1 FILLER_22_294 ();
 sg13g2_fill_2 FILLER_22_300 ();
 sg13g2_fill_2 FILLER_22_306 ();
 sg13g2_fill_2 FILLER_22_313 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_2 FILLER_22_402 ();
 sg13g2_decap_4 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_4 ();
 sg13g2_decap_8 FILLER_23_10 ();
 sg13g2_decap_8 FILLER_23_17 ();
 sg13g2_decap_8 FILLER_23_24 ();
 sg13g2_decap_4 FILLER_23_31 ();
 sg13g2_decap_8 FILLER_23_39 ();
 sg13g2_decap_4 FILLER_23_46 ();
 sg13g2_decap_8 FILLER_23_54 ();
 sg13g2_fill_2 FILLER_23_61 ();
 sg13g2_fill_1 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_74 ();
 sg13g2_fill_2 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_83 ();
 sg13g2_fill_2 FILLER_23_102 ();
 sg13g2_fill_1 FILLER_23_117 ();
 sg13g2_fill_2 FILLER_23_133 ();
 sg13g2_fill_1 FILLER_23_143 ();
 sg13g2_decap_4 FILLER_23_153 ();
 sg13g2_fill_2 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_171 ();
 sg13g2_decap_8 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_2 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_231 ();
 sg13g2_fill_2 FILLER_23_237 ();
 sg13g2_fill_2 FILLER_23_244 ();
 sg13g2_fill_2 FILLER_23_251 ();
 sg13g2_fill_2 FILLER_23_272 ();
 sg13g2_fill_2 FILLER_23_282 ();
 sg13g2_decap_8 FILLER_23_340 ();
 sg13g2_decap_8 FILLER_23_347 ();
 sg13g2_decap_4 FILLER_23_406 ();
 sg13g2_fill_1 FILLER_23_410 ();
 sg13g2_decap_4 FILLER_23_419 ();
 sg13g2_fill_2 FILLER_23_427 ();
 sg13g2_fill_1 FILLER_23_429 ();
 sg13g2_decap_4 FILLER_24_0 ();
 sg13g2_fill_1 FILLER_24_4 ();
 sg13g2_fill_2 FILLER_24_29 ();
 sg13g2_fill_2 FILLER_24_56 ();
 sg13g2_fill_1 FILLER_24_91 ();
 sg13g2_fill_1 FILLER_24_96 ();
 sg13g2_fill_2 FILLER_24_101 ();
 sg13g2_fill_1 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_126 ();
 sg13g2_fill_1 FILLER_24_128 ();
 sg13g2_fill_2 FILLER_24_139 ();
 sg13g2_fill_1 FILLER_24_141 ();
 sg13g2_fill_2 FILLER_24_146 ();
 sg13g2_fill_1 FILLER_24_166 ();
 sg13g2_fill_2 FILLER_24_171 ();
 sg13g2_fill_1 FILLER_24_173 ();
 sg13g2_fill_1 FILLER_24_182 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_1 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_203 ();
 sg13g2_fill_1 FILLER_24_205 ();
 sg13g2_fill_1 FILLER_24_220 ();
 sg13g2_decap_4 FILLER_24_225 ();
 sg13g2_fill_2 FILLER_24_229 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_261 ();
 sg13g2_fill_1 FILLER_24_268 ();
 sg13g2_fill_1 FILLER_24_275 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_decap_4 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_303 ();
 sg13g2_fill_2 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_316 ();
 sg13g2_fill_2 FILLER_24_325 ();
 sg13g2_fill_2 FILLER_24_353 ();
 sg13g2_decap_4 FILLER_24_359 ();
 sg13g2_fill_2 FILLER_24_368 ();
 sg13g2_fill_2 FILLER_24_374 ();
 sg13g2_fill_2 FILLER_24_391 ();
 sg13g2_fill_2 FILLER_24_402 ();
 sg13g2_fill_2 FILLER_25_0 ();
 sg13g2_fill_1 FILLER_25_2 ();
 sg13g2_fill_1 FILLER_25_16 ();
 sg13g2_fill_1 FILLER_25_26 ();
 sg13g2_fill_1 FILLER_25_32 ();
 sg13g2_fill_1 FILLER_25_53 ();
 sg13g2_fill_1 FILLER_25_58 ();
 sg13g2_fill_1 FILLER_25_67 ();
 sg13g2_fill_2 FILLER_25_80 ();
 sg13g2_decap_8 FILLER_25_115 ();
 sg13g2_fill_2 FILLER_25_122 ();
 sg13g2_fill_1 FILLER_25_124 ();
 sg13g2_fill_2 FILLER_25_143 ();
 sg13g2_fill_2 FILLER_25_149 ();
 sg13g2_decap_4 FILLER_25_155 ();
 sg13g2_fill_1 FILLER_25_163 ();
 sg13g2_fill_1 FILLER_25_187 ();
 sg13g2_fill_1 FILLER_25_196 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_fill_1 FILLER_25_207 ();
 sg13g2_fill_1 FILLER_25_213 ();
 sg13g2_fill_1 FILLER_25_219 ();
 sg13g2_fill_1 FILLER_25_245 ();
 sg13g2_fill_2 FILLER_25_259 ();
 sg13g2_fill_1 FILLER_25_266 ();
 sg13g2_fill_1 FILLER_25_272 ();
 sg13g2_decap_4 FILLER_25_329 ();
 sg13g2_fill_1 FILLER_25_333 ();
 sg13g2_decap_4 FILLER_25_338 ();
 sg13g2_fill_1 FILLER_25_375 ();
 sg13g2_fill_2 FILLER_25_402 ();
 sg13g2_decap_4 FILLER_26_0 ();
 sg13g2_fill_2 FILLER_26_26 ();
 sg13g2_fill_1 FILLER_26_46 ();
 sg13g2_fill_2 FILLER_26_51 ();
 sg13g2_fill_2 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_84 ();
 sg13g2_fill_1 FILLER_26_86 ();
 sg13g2_fill_2 FILLER_26_92 ();
 sg13g2_fill_1 FILLER_26_94 ();
 sg13g2_fill_2 FILLER_26_129 ();
 sg13g2_fill_1 FILLER_26_131 ();
 sg13g2_fill_2 FILLER_26_140 ();
 sg13g2_fill_2 FILLER_26_164 ();
 sg13g2_fill_1 FILLER_26_166 ();
 sg13g2_fill_1 FILLER_26_172 ();
 sg13g2_fill_1 FILLER_26_218 ();
 sg13g2_fill_1 FILLER_26_225 ();
 sg13g2_fill_1 FILLER_26_235 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_249 ();
 sg13g2_fill_1 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_280 ();
 sg13g2_fill_1 FILLER_26_285 ();
 sg13g2_fill_2 FILLER_26_290 ();
 sg13g2_fill_2 FILLER_26_296 ();
 sg13g2_fill_1 FILLER_26_301 ();
 sg13g2_fill_2 FILLER_26_307 ();
 sg13g2_fill_1 FILLER_26_382 ();
 sg13g2_fill_1 FILLER_26_389 ();
 sg13g2_fill_1 FILLER_26_412 ();
 sg13g2_fill_2 FILLER_26_420 ();
 sg13g2_decap_4 FILLER_26_426 ();
 sg13g2_fill_1 FILLER_27_17 ();
 sg13g2_fill_2 FILLER_27_43 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_decap_4 FILLER_27_62 ();
 sg13g2_fill_2 FILLER_27_72 ();
 sg13g2_fill_1 FILLER_27_74 ();
 sg13g2_decap_8 FILLER_27_83 ();
 sg13g2_decap_8 FILLER_27_90 ();
 sg13g2_fill_2 FILLER_27_97 ();
 sg13g2_fill_1 FILLER_27_130 ();
 sg13g2_fill_2 FILLER_27_145 ();
 sg13g2_decap_4 FILLER_27_152 ();
 sg13g2_fill_1 FILLER_27_186 ();
 sg13g2_fill_1 FILLER_27_199 ();
 sg13g2_fill_1 FILLER_27_204 ();
 sg13g2_decap_4 FILLER_27_248 ();
 sg13g2_fill_2 FILLER_27_252 ();
 sg13g2_fill_1 FILLER_27_277 ();
 sg13g2_fill_2 FILLER_27_304 ();
 sg13g2_fill_1 FILLER_27_327 ();
 sg13g2_fill_1 FILLER_27_363 ();
 sg13g2_fill_2 FILLER_27_368 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_1 FILLER_28_4 ();
 sg13g2_fill_1 FILLER_28_23 ();
 sg13g2_fill_2 FILLER_28_28 ();
 sg13g2_decap_4 FILLER_28_47 ();
 sg13g2_fill_1 FILLER_28_51 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_88 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_fill_2 FILLER_28_112 ();
 sg13g2_fill_1 FILLER_28_114 ();
 sg13g2_decap_4 FILLER_28_124 ();
 sg13g2_fill_1 FILLER_28_132 ();
 sg13g2_fill_1 FILLER_28_138 ();
 sg13g2_decap_8 FILLER_28_148 ();
 sg13g2_fill_1 FILLER_28_165 ();
 sg13g2_fill_1 FILLER_28_170 ();
 sg13g2_fill_2 FILLER_28_179 ();
 sg13g2_decap_8 FILLER_28_185 ();
 sg13g2_decap_4 FILLER_28_192 ();
 sg13g2_fill_2 FILLER_28_210 ();
 sg13g2_fill_2 FILLER_28_220 ();
 sg13g2_fill_1 FILLER_28_222 ();
 sg13g2_fill_2 FILLER_28_227 ();
 sg13g2_fill_2 FILLER_28_233 ();
 sg13g2_fill_2 FILLER_28_253 ();
 sg13g2_fill_1 FILLER_28_255 ();
 sg13g2_fill_1 FILLER_28_284 ();
 sg13g2_decap_8 FILLER_28_289 ();
 sg13g2_fill_1 FILLER_28_353 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_380 ();
 sg13g2_fill_1 FILLER_28_385 ();
 sg13g2_fill_2 FILLER_28_420 ();
 sg13g2_fill_1 FILLER_28_429 ();
 sg13g2_decap_8 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_48 ();
 sg13g2_fill_2 FILLER_29_76 ();
 sg13g2_decap_8 FILLER_29_86 ();
 sg13g2_decap_8 FILLER_29_93 ();
 sg13g2_decap_8 FILLER_29_100 ();
 sg13g2_decap_4 FILLER_29_107 ();
 sg13g2_fill_1 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_119 ();
 sg13g2_fill_2 FILLER_29_125 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_fill_2 FILLER_29_132 ();
 sg13g2_fill_1 FILLER_29_134 ();
 sg13g2_fill_2 FILLER_29_139 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_fill_1 FILLER_29_160 ();
 sg13g2_fill_1 FILLER_29_170 ();
 sg13g2_fill_2 FILLER_29_180 ();
 sg13g2_fill_1 FILLER_29_182 ();
 sg13g2_decap_4 FILLER_29_194 ();
 sg13g2_fill_2 FILLER_29_198 ();
 sg13g2_decap_8 FILLER_29_204 ();
 sg13g2_fill_1 FILLER_29_211 ();
 sg13g2_decap_8 FILLER_29_216 ();
 sg13g2_fill_1 FILLER_29_233 ();
 sg13g2_fill_1 FILLER_29_239 ();
 sg13g2_fill_1 FILLER_29_249 ();
 sg13g2_fill_1 FILLER_29_264 ();
 sg13g2_fill_1 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_282 ();
 sg13g2_decap_4 FILLER_29_298 ();
 sg13g2_fill_1 FILLER_29_302 ();
 sg13g2_fill_1 FILLER_29_368 ();
 sg13g2_fill_1 FILLER_29_387 ();
 sg13g2_fill_2 FILLER_29_401 ();
 sg13g2_fill_1 FILLER_29_429 ();
 sg13g2_fill_2 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_2 ();
 sg13g2_decap_4 FILLER_30_26 ();
 sg13g2_fill_2 FILLER_30_30 ();
 sg13g2_fill_1 FILLER_30_36 ();
 sg13g2_decap_4 FILLER_30_41 ();
 sg13g2_fill_2 FILLER_30_45 ();
 sg13g2_decap_8 FILLER_30_60 ();
 sg13g2_fill_1 FILLER_30_67 ();
 sg13g2_decap_8 FILLER_30_96 ();
 sg13g2_decap_8 FILLER_30_103 ();
 sg13g2_fill_1 FILLER_30_110 ();
 sg13g2_decap_4 FILLER_30_114 ();
 sg13g2_fill_1 FILLER_30_118 ();
 sg13g2_decap_4 FILLER_30_141 ();
 sg13g2_decap_4 FILLER_30_149 ();
 sg13g2_fill_1 FILLER_30_153 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_fill_2 FILLER_30_210 ();
 sg13g2_fill_1 FILLER_30_234 ();
 sg13g2_fill_2 FILLER_30_250 ();
 sg13g2_fill_2 FILLER_30_270 ();
 sg13g2_fill_2 FILLER_30_335 ();
 sg13g2_fill_1 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_427 ();
 sg13g2_fill_1 FILLER_30_429 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_4 FILLER_31_7 ();
 sg13g2_fill_1 FILLER_31_19 ();
 sg13g2_fill_1 FILLER_31_33 ();
 sg13g2_decap_4 FILLER_31_41 ();
 sg13g2_fill_1 FILLER_31_45 ();
 sg13g2_fill_1 FILLER_31_59 ();
 sg13g2_fill_1 FILLER_31_65 ();
 sg13g2_fill_1 FILLER_31_71 ();
 sg13g2_fill_1 FILLER_31_77 ();
 sg13g2_fill_1 FILLER_31_89 ();
 sg13g2_fill_2 FILLER_31_95 ();
 sg13g2_fill_1 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_fill_1 FILLER_31_109 ();
 sg13g2_fill_1 FILLER_31_118 ();
 sg13g2_fill_1 FILLER_31_128 ();
 sg13g2_decap_8 FILLER_31_194 ();
 sg13g2_decap_8 FILLER_31_201 ();
 sg13g2_decap_4 FILLER_31_208 ();
 sg13g2_fill_2 FILLER_31_212 ();
 sg13g2_decap_4 FILLER_31_217 ();
 sg13g2_fill_1 FILLER_31_221 ();
 sg13g2_fill_1 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_250 ();
 sg13g2_fill_1 FILLER_31_261 ();
 sg13g2_fill_2 FILLER_31_296 ();
 sg13g2_fill_1 FILLER_31_328 ();
 sg13g2_fill_2 FILLER_31_337 ();
 sg13g2_fill_2 FILLER_31_343 ();
 sg13g2_fill_1 FILLER_31_345 ();
 sg13g2_fill_2 FILLER_31_350 ();
 sg13g2_fill_2 FILLER_31_369 ();
 sg13g2_fill_1 FILLER_31_378 ();
 sg13g2_fill_2 FILLER_31_428 ();
 sg13g2_fill_1 FILLER_32_40 ();
 sg13g2_fill_2 FILLER_32_55 ();
 sg13g2_fill_2 FILLER_32_61 ();
 sg13g2_fill_1 FILLER_32_63 ();
 sg13g2_fill_1 FILLER_32_72 ();
 sg13g2_fill_1 FILLER_32_78 ();
 sg13g2_fill_1 FILLER_32_83 ();
 sg13g2_fill_1 FILLER_32_89 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_116 ();
 sg13g2_fill_2 FILLER_32_138 ();
 sg13g2_decap_4 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_172 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_decap_8 FILLER_32_199 ();
 sg13g2_fill_2 FILLER_32_223 ();
 sg13g2_fill_1 FILLER_32_280 ();
 sg13g2_fill_1 FILLER_32_307 ();
 sg13g2_fill_1 FILLER_32_311 ();
 sg13g2_fill_2 FILLER_32_332 ();
 sg13g2_fill_1 FILLER_32_334 ();
 sg13g2_fill_2 FILLER_32_396 ();
 sg13g2_fill_1 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_16 ();
 sg13g2_fill_1 FILLER_33_18 ();
 sg13g2_fill_1 FILLER_33_24 ();
 sg13g2_fill_1 FILLER_33_30 ();
 sg13g2_fill_1 FILLER_33_35 ();
 sg13g2_fill_2 FILLER_33_45 ();
 sg13g2_decap_4 FILLER_33_51 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_decap_8 FILLER_33_65 ();
 sg13g2_fill_1 FILLER_33_72 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_decap_4 FILLER_33_105 ();
 sg13g2_fill_1 FILLER_33_109 ();
 sg13g2_fill_1 FILLER_33_126 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_183 ();
 sg13g2_fill_1 FILLER_33_185 ();
 sg13g2_decap_4 FILLER_33_191 ();
 sg13g2_fill_1 FILLER_33_195 ();
 sg13g2_fill_1 FILLER_33_200 ();
 sg13g2_decap_8 FILLER_33_206 ();
 sg13g2_fill_2 FILLER_33_226 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_234 ();
 sg13g2_fill_2 FILLER_33_239 ();
 sg13g2_fill_1 FILLER_33_241 ();
 sg13g2_fill_1 FILLER_33_246 ();
 sg13g2_fill_1 FILLER_33_251 ();
 sg13g2_fill_1 FILLER_33_261 ();
 sg13g2_fill_2 FILLER_33_265 ();
 sg13g2_decap_8 FILLER_33_277 ();
 sg13g2_decap_4 FILLER_33_284 ();
 sg13g2_fill_2 FILLER_33_288 ();
 sg13g2_decap_8 FILLER_33_298 ();
 sg13g2_fill_1 FILLER_33_305 ();
 sg13g2_fill_2 FILLER_33_310 ();
 sg13g2_decap_4 FILLER_33_316 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_fill_1 FILLER_33_396 ();
 sg13g2_fill_1 FILLER_33_405 ();
 sg13g2_fill_1 FILLER_33_410 ();
 sg13g2_fill_2 FILLER_33_427 ();
 sg13g2_fill_1 FILLER_33_429 ();
 sg13g2_fill_1 FILLER_34_34 ();
 sg13g2_fill_1 FILLER_34_99 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_fill_1 FILLER_34_109 ();
 sg13g2_decap_4 FILLER_34_117 ();
 sg13g2_fill_2 FILLER_34_121 ();
 sg13g2_fill_2 FILLER_34_136 ();
 sg13g2_fill_1 FILLER_34_207 ();
 sg13g2_decap_4 FILLER_34_212 ();
 sg13g2_fill_1 FILLER_34_221 ();
 sg13g2_fill_1 FILLER_34_226 ();
 sg13g2_fill_1 FILLER_34_232 ();
 sg13g2_fill_1 FILLER_34_239 ();
 sg13g2_decap_4 FILLER_34_244 ();
 sg13g2_fill_1 FILLER_34_253 ();
 sg13g2_fill_1 FILLER_34_265 ();
 sg13g2_decap_4 FILLER_34_270 ();
 sg13g2_fill_1 FILLER_34_274 ();
 sg13g2_fill_1 FILLER_34_311 ();
 sg13g2_fill_2 FILLER_34_315 ();
 sg13g2_fill_2 FILLER_34_347 ();
 sg13g2_fill_2 FILLER_34_387 ();
 sg13g2_fill_1 FILLER_34_394 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_7 ();
 sg13g2_fill_1 FILLER_35_99 ();
 sg13g2_fill_1 FILLER_35_104 ();
 sg13g2_fill_1 FILLER_35_115 ();
 sg13g2_fill_2 FILLER_35_120 ();
 sg13g2_fill_1 FILLER_35_126 ();
 sg13g2_fill_2 FILLER_35_132 ();
 sg13g2_decap_4 FILLER_35_151 ();
 sg13g2_fill_2 FILLER_35_155 ();
 sg13g2_fill_1 FILLER_35_161 ();
 sg13g2_decap_4 FILLER_35_176 ();
 sg13g2_fill_1 FILLER_35_184 ();
 sg13g2_fill_2 FILLER_35_194 ();
 sg13g2_decap_8 FILLER_35_200 ();
 sg13g2_decap_8 FILLER_35_207 ();
 sg13g2_decap_4 FILLER_35_214 ();
 sg13g2_fill_2 FILLER_35_226 ();
 sg13g2_fill_1 FILLER_35_228 ();
 sg13g2_decap_4 FILLER_35_271 ();
 sg13g2_fill_2 FILLER_35_283 ();
 sg13g2_fill_1 FILLER_35_285 ();
 sg13g2_fill_2 FILLER_35_321 ();
 sg13g2_fill_1 FILLER_35_323 ();
 sg13g2_fill_1 FILLER_35_368 ();
 sg13g2_fill_1 FILLER_35_393 ();
 sg13g2_fill_1 FILLER_35_425 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_fill_2 FILLER_36_7 ();
 sg13g2_fill_1 FILLER_36_9 ();
 sg13g2_fill_1 FILLER_36_57 ();
 sg13g2_fill_1 FILLER_36_62 ();
 sg13g2_fill_1 FILLER_36_85 ();
 sg13g2_fill_2 FILLER_36_99 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_1 FILLER_36_158 ();
 sg13g2_fill_1 FILLER_36_163 ();
 sg13g2_fill_2 FILLER_36_173 ();
 sg13g2_fill_2 FILLER_36_179 ();
 sg13g2_fill_2 FILLER_36_185 ();
 sg13g2_fill_1 FILLER_36_187 ();
 sg13g2_fill_1 FILLER_36_200 ();
 sg13g2_fill_2 FILLER_36_219 ();
 sg13g2_decap_8 FILLER_36_225 ();
 sg13g2_decap_4 FILLER_36_247 ();
 sg13g2_fill_2 FILLER_36_263 ();
 sg13g2_fill_2 FILLER_36_270 ();
 sg13g2_decap_4 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_1 FILLER_36_290 ();
 sg13g2_fill_2 FILLER_36_303 ();
 sg13g2_fill_1 FILLER_36_305 ();
 sg13g2_decap_4 FILLER_36_316 ();
 sg13g2_fill_1 FILLER_36_320 ();
 sg13g2_fill_2 FILLER_36_392 ();
 sg13g2_fill_1 FILLER_36_398 ();
 sg13g2_decap_4 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_13 ();
 sg13g2_fill_2 FILLER_37_53 ();
 sg13g2_fill_1 FILLER_37_96 ();
 sg13g2_fill_1 FILLER_37_105 ();
 sg13g2_fill_1 FILLER_37_110 ();
 sg13g2_fill_1 FILLER_37_131 ();
 sg13g2_fill_1 FILLER_37_148 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_fill_2 FILLER_37_193 ();
 sg13g2_fill_2 FILLER_37_221 ();
 sg13g2_fill_1 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_257 ();
 sg13g2_fill_1 FILLER_37_263 ();
 sg13g2_fill_1 FILLER_37_268 ();
 sg13g2_fill_2 FILLER_37_273 ();
 sg13g2_fill_1 FILLER_37_279 ();
 sg13g2_fill_2 FILLER_37_422 ();
 sg13g2_fill_1 FILLER_37_424 ();
 sg13g2_fill_1 FILLER_37_429 ();
 sg13g2_fill_1 FILLER_38_26 ();
 sg13g2_fill_1 FILLER_38_127 ();
 sg13g2_fill_1 FILLER_38_189 ();
 sg13g2_fill_1 FILLER_38_194 ();
 sg13g2_fill_1 FILLER_38_203 ();
 sg13g2_fill_2 FILLER_38_240 ();
 sg13g2_fill_1 FILLER_38_250 ();
 sg13g2_fill_1 FILLER_38_255 ();
 sg13g2_fill_1 FILLER_38_322 ();
 sg13g2_fill_1 FILLER_38_403 ();
endmodule
